`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GDjtpDLpTrwkCs+z3GE2+tDGSflarkIAnykdM550kGjK1Ce9i+ZWjfw4T0F8ie55+FB7xQomgSdP
exOo2LwyCw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ocrLj4slMX6IYCvT3Fxx3/1E+5RmtWeM7qcwVqFhppBkzzAYD3iexASL1kaNWcSJF3WVR85kixpm
jXw/hyccrXeqNjm/Qwo2acNXY0TvCBer6k1RqvM6LGGyehdf0jC6mn+0B/NBtPCuqqLFMd+Svr4k
zif+YnkNSeuPyix9swg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hd1O828ijlSZFj1eICielJkqOVqejY8vv1LyPQLkhD+ZIE7WXRzdUCvyBIrMkl7htlU9Tk0Aa9GI
UwqJ87HhLVvY4G0SzEleV3Z3ENcK8ueq8dA451VsSwwhlsRGCijmpiLlMAbKv8jTPaLS4uaQMfDw
tB+it8q/NtCOYH1tT93dn7V4McBE+Pptxw6DkZ8DpnaMqaM3WwmH800grXkoi1+vXi8+Zq/NTRLZ
WDFa5mGG0jbvTgxBhsNMy+qRftruFCJrSLrJa3XbSyCLvqqAf9MIR1ib8wXLxtOEXIJ4ec0dq4Cp
tQik68r/U9f1cRlcnGR6iRhvMLjplBWLqgqLnQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hd3fG8RdamuhXsfhLnMUhAnc0JijaAVPWK1C7gb+WbgLgu4o8EbZqG436+ymVWVaWUaYBoUQdqA6
pPnFEqGMU9i3MJ6jd6yWSZ5l91FyFstDzohHvNLsF/GyG0WVlbfrLiv3k5jvKMfuxts74XoOchKJ
HeJKmvAvD8jByx2Z4HrS2HXbHIwH2P68BcMy1r9pxm8Apa6STwyRamArTecy6KHKFGBYAnFs1ZKw
5epBuemssW2HJJ6XylDBG1hWHITipvj7+2FPUx/qMnNsY7aspBT+eNrDaPzv+k5fZ6o6BRhrx2p1
b0Dh7P+9KnF4PEGMgry+icQBmbaqO2+60QKkGA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HlKh+RG3201qhrHVxfwND3GCWQoi3/DiMmPI/Stx9v065LQ+yp8AlemtS+2TOT8cSKaAX1Gm/n4u
xHvqhz6G6WAKnMbFWs0M8uODhuJPxJmGgyUu8pqeGAUOu43aHTIEKd/nn+TX/ZnKwuk6m6n1IMiZ
tmDdcbCIqh3dxnO4+yiqdkltjm4QQhy4EoqMgylVJN27cAnaIpFg9H52wkdZR1wVUEQa8z/zZHke
io2PQhuHL/pIJ18ZThx0Os1eprgzF140cf6IFWWTpcekmTXHuUFHlKMicpxg5eTYNQNAnSZ/PijN
0Qvq8X5aavtHvKK0O7IuZzAagBKr3jKP6rI9gQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KD7FUY09rWLZruDGbmrJOXaDBraBxna2jboaVV/Qqxyjrby/ElxlNVTK0zj95OEJTsbJV4XL/9Jq
NgggzubaaCguemde7bL4KylHEXpX3G07ZtQwsi190p6nNYNnXpx5XZQtw6Ng08CDy+7acmhU6NB+
Dxf/RWARG92LDOdhMvo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cg2tVcuYYrV98PCK+rclTkZCoF+9HQytUf0yy1tFMAH0Zis5rEmDKTEc8EthWsDo6rRRqSD7GNSD
vrDOkoSGhni9EUzH2Lmb2We8YTELLp/C56B58wFCtFn9OseFZTXUyg2VTvS+eMeyzaddfG65JTTy
lxkif7uUdpdfqcNLwf0bt65bzLUo33DSeQma2qBH/+W2rdRkAFSD7n0JaVxN2O8pe2XOXzrFAVKH
su54BVqD4YaKNcyfD35oZlNkCLTm9oz3xw/aeF6fLf0KAfA9CkM+8RzoBfz+mZPgQLkREtrRHfMi
gNtkA1QUdbwqZp9n3G3OILNOPLk6lK55dySggA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
DXYxWFfHnnOsn20kNX1vymSvzNqGRrbSkMI1Acq/v+wqreEXKxZLv7R6rRgbgmxFK+8FG0TtB7+r
pcyyGqLmk0uVgDVsswfyc7tsns2Bm7VQHQK7W2PaotYXCtzKOEXmbYkLfodUpPlMRBX6A3JYGcBz
vQtYtRF6cZPx/NveYWTPkbEg7jZn7CZ5k7E3BaPGQhVW1kobXHXnj4qvO0wfVyYT6wNoqrxf3eF1
ZDPvlHAW0FIx1szxC/Cvo+v6RLfw1qzaX0xihI0GyrtQDam1xCBoHv/aAPxeOSUICIyDVfVq6/JD
G6Uoh6SZQIAOXga9nLB0puevWCWsRKRLqmo5gPFZYv4sjWADrHTfrUS0K5pZkolmKPYtgNVfg4sC
f02uccpF2a4q/SDIJ5MDidmcwQlUSQVl7r8vcTnRlKbXrASz65tFgJubW+3EhrkVMlo4l+c5sJdK
A/N6aG8ozw1i9lMauihSZ9Ykyt2mcLpobiOmiOn1Z+mv5Jdjl20EL4q+gxig7Gw9OYodk5yd/Oq9
uTlWHXoRUg7XAgDk7PduyZfghkeF7lpXaBQXt3f9FCQQLIzM7uPN9TSaRJhDbNEJ1D4kn9oK6p1P
ACE9BSZ9nPqCr+osGkXT99SGK/JVzDqbDNYO4gLAzK7/gKZqCx6rs7SNZhjq+jRVytgahxZ9W3cU
KruzA/Hwabm/FLze89DtCKzMIiUoGFG7FOGcyt4Br2/cZBvBvyoIfVbuGrI0NOrlF/LM6HD9iAFO
7nbaupUrsvCMI8tv6ZH/yEK+cVUufnSfrFhNeVRn1nqTukIs3IqroPNJObNnx3W1T5awB9gJQ4uz
Ya9MpL1JzZUahZuX9m4dP37gyLdztcXr3j+4asKHqvlv6xlgyefJijb2sK55R/jgKLnpXZP5zzmt
bA9sFlas+lDQFmNttTs70ohATrtI8MD95+rpHhGHYLhc6Ld/iIXswkG/8SAuw2IqGZalmhEC9FQI
dFSR0cNMT0g82d+1/Rq1S0s4taSiU11zW9nYC+mGRe4PY8S4LCvNFF/ikjTppMKDTJRzkx0xgmAA
LZC17kypKncdsFGujYjnJTaBYY0VG2L+6A4yJToqP8FvZrqWm6LwiOB2fi/CsAHfd4en9kPBVXOr
7IiTnOzvUR8MCZojTpGEUuxTOZ2qSR2wgBouwynqiDSUgw4YzMQc3nbWHVnT6E/+qN2UzcdsBdwx
YO/XQgdtRPY+7Pqw1dVNGFF1ItQZEAE7K9JjajBONV+3Cul0G2mjEju3PZB9lDNVL3KBP5KG+xsq
H8K/E3oFxvr/Y0qMbdBeBIR5zMLrzpHpK+Bc7Jwn1GaNGYOwvQAqxj18yNJJj80h/QFKyorE7fad
ppy6Gz0xaqhG9KTZHYxhMeTHMlOw/FDVxGieiU+lVGfKexA56e3wrXG5rOdDsbsFSOeaANuxwOpY
SgSNk9frP1fMGST8H3pFeFGPYmKWb88qZeEawcDeNmlLoIWzalRNsdRZz8qbQmr4VtZJwGoc2VzH
P75odFRhJz+3sztffYo90JaBzvJuczu88R2a1TDeNSXOdfoYB7ef6HGFk4dHiwCu2hPsnJVPQli3
+6qCpSkbylPVg5WVtS5VJuR0Pm2KuA1UWc+SywYJgdTuuKcOMVlfszG9AlXrpe1QDAASMltoqJK0
GBgJ5sMIoG63sO53uOQS5nwMocgJekHA8wkEWlAzGm2hx5Vqbv6leDpUbYT5U2s0rYisVyQpm9p5
fS9xZ01SQbc8FNFGVR+jXPj3+FZMjYPlUNlHFj+wXu/Gzo9Z42YbnTM1IDbRcoE/TiWuzgSzo/39
AZ/wPEmVQmjzR7vaPs6opMVLrOF8TBgJ3DnecOOCgpVUx1aGLUyRY58MawhtPOq3VkgrsbLC3KOo
OaojxwuboI5/EBJ4SDeLQ1NT0Az9ImlRod1zoxW9W/VvMclJB3s0kMINlcC7wTYW1UBOg8Epxihc
y4bIOWCdWuneOfbBCEBleBxEwZXIo4/XaVG/quo94gQOehngHy9fP1QbuS6svezrP1B1Qq1m3hvV
aijqA0s6jKcfGzAHTGGOOx+eYxwvLfzFNOqvFa+w+zS8KdCIkLq433sbuzpPgtTILWj3kHScfis3
pLIhUXab+cBJcjAJLR+FHFgj27E4lCj6VAlLcQmvb0+STFqt0c9WWFDsmHijqo6UbUX8smCEsduF
izPkhMRDmbvOpMbpIs9JUiI0lQBRO2fiUKTrWtLJXgnpDEnVhPer3jSJ2/eCLUXLoa4W0095I1Xz
3/lpSibfK+IeL7hkzVCoZYcxsaqZZKks/z1MLGYTDVDETkPPMHqu5ufAE25GM096kwUpp24RKAoh
h9dluID418WE8NKZaX5SN1T+Z6QgDvy3uQ+Q6eBQexm5XoLa45Ov6dhrYbCOjFWSbdbP3jPOC2lt
6vbUv4/+V56taL8I4CML3aoUc/VS+MSwUu/EpI5Y0GqoYBRq3YE6drzUqE6S3uWf98GIX6AZizf9
q4uS6rBLFCZncM5dMb0sFuqvIvbr1UAQgKs9kf1IFehD6ay3U81mkfEK3p3D+cclE/HVjspA4MZW
o6QVKZ1QqFpVIPnPMuItBgIS6mLwb37ElNK7G/tsLcxRxhhWHx5FVYx/7AfSwyYMb4OoQC1tZkow
tr1agKkKEiETYRnWiCPlWYl9Ba9EZDW0Fa3ZUyy6UmZ3Mx2yRiK3qhyHVda8r57nlHfjSXUA4TlR
6TVrouoHzHFiL8v3NXsZaCa26Cku5oGoZmwcusQ8Vt3a7m7H8tX4GTEBORhU7amnJ5iMDeOUcnfW
QaR4OMinLuweOs6c1KomqpMmpuAlFo/mivUbVi9HrMMIpoqJQ9SEVcPHYLrik/sQ76uq+X47IdCu
kfiAYMEf5tj1H09Wgc3zcUutg7+uBxiGHWSOd8t2CtXvaRht39Papfp71gLSI2wViv9COBAywKTn
MS72veSkCvX9IC9s/P4y8hzdUgEKDt4So+8msgUv/UCO4XXrqK6dAlgUWI8C+HvR1L4h/wBdeaoE
YRikbq4torYb0jTu0IsQ9jYaq/jYmBsBYspkkI1BcyB0dODQXLr8lYBkoHX3nXtTpo2fhtM0GNt6
38fPzYRn0e8GftVj3o4j8+OYQk+zYZGZub4SDkPkFc3POz5/54ciIE4XzIfMphR1rPmmY6zeOYAb
5fpBMtwzwfO12xAWkzY1//thsrAJEueUwxXkCSeJdOHiElB8GYzqfR+JD6pTnt1zy84Jfd2rtMAJ
T+GCx1SeSmjldsVhi+hw1w5/AAgOm37hTe1i/WPU8mL6BkkgwUkxMH3GpcnylF4oCUy8DXaJ/oj7
VpUBhNP/pP0/vkc3V7NZv+qKFlaLwFOvKgvlb5jD4FePoGU49K+IGFn3SVGLSGqJBm1OGGuWeo5s
g9lk7bOS7FVVxhU+EbHLDRYHjqm3IG0y1Sndle+pfTKI22q3F2V0ycskRt7u8bgRIB46C+nddBvv
y86ofHw++j+bc/c3lSlBxuroUuqrgczzogrc9aqJANK14bicmpFOwgL3pb89Kmhlvqh7Dmy7z8xG
r4R3YzoeskLp5qpEU0+sOWavKuVYGnn1GxLa/sjodnSYoVNp99SHyUa5lepFA8hFTfhcrJ5Rj0aW
OaNQh2Na/YUbRM4Z867LQwV3F2xZlsbNbGAFqUAbXfYsukH1KAkmjmYxmqNSnsE+9NnL34dMiyqG
ihmwFN7GXrKPEvYWez8HxFHARQHI8eeSoPn+nah1ng8tDR0gshdGcwmL+aL5G4NICaqLVSoiW1tr
xX+AW2yeWZ6JJdL7ZU4hrCwT1pjVv0CUfh5YWx/5NEIj2W5UtJmy7JgOAH4fl+sgy5WtfqPBPBVT
EuRnXl6AdT8fLJ//uS4hLZ9bIaYF/GAGUh3P6CFc/KGsEkIBKYFjvgiKxSKa9MA9lIA9LdNhbtNT
IS29fjpUWldOdFrRns3gpJ050oleAOI55WsvjtX//CgDUft6QNpq2BVz1jfZqzjgTI/fIYyBuj1T
aqngnxGRCD6BSiZmgaQOiDtT2bE5y2WKHRZR2yycRdODdXcypCak/2WMEKU/aQU2x5w1Zv1X2dTT
HNrBAgH2uKSyo5fGHXD9Wp+dxmkkMDHGdus9r1Jr3hT0P0qPDWFV12cQWP9Kt7aNmR/WtSLDg/aD
0JJzRcXMIAfcxE8d36C2Q+ebF2Q1W6QxXuNqUtD573TWcKAIHvOhG3oisaOTsfVu/Uc4IOgyxQPA
1NmrSySFPXgwpQpOeSFyQfBT38AP+faKbZVW+oVKfnpjyynSIW1etHYePIeiQztzSrv+hj0IIh/i
rwLfqsw/EQhFxECcyA4rcTevfkfHm7IXK4VfNMzAU8KYvBXg51YVL45scNiyH7TEP1s47zbXvavZ
tIJonV/0RWkyt7hxtNbaKjm0gEIERRMWqNzd1NrkxXx27IdqmMCTmW5VOycf/aeHF0Pk5KatzuA/
KGQF3ykEHpg1jgfzskNcEnXgXbxZk8UMFotGEhrkIBEuBcHS9p4yL225+hp0Nq6hkOl7dMgzKqXk
+v1tCwPVW4NlPdcw4BP8DSaMLkL5QYhBV67uwERVyfq4fvtyLgGVQJ1t6mKMCVbIyBE85WIynJ9p
7htG6nLk3gywx0W2aSW8nAtdtVUO1EOXaFkgJ7wvFZMmAZlhtaoil7SovloApH9kv4O3ZLCD7Kbp
pLrnSkYjIHK9naraAdgx5xauOGPtnapiiEsJetAn430iHgErwGsUUfe0H9UIPsT8P6BtwtU8P1cB
R9RBAmrcIwGcAGY81jUWN/MLY1Z2ajxJ6mjf5D+gPz54Zne849uQ6gitbqK3oPydAK42RJ31zCdr
nFadRbsgHB9grRr9MHOLbTe6vhGdYH3ZwWqC3TTwrAhOh2ksEdod5Os+XHSg53I9m0EX+B7r1Nph
3VsbxkeC39QbKioRyRviKvCohUdUJrN/cZTyIJOkUgtJgvA8SyFdsYYn+ayC7/IoYlVzg3D/kCdX
hv3qqpVixDuUPmivefBveDQBdXKydAMwPZrRl32cVL3bq6gmL03SJ7Gr5NPy4NzYa73HhOULO7Q/
izXamKpGfHHEzO9L6lS2x0AlJRStIpq+sY8x+qdEL5Ca/DbMBEWXIljsEswbXrm+uAol/4AA2mb5
YKNRNx2dILWhFb/Dm4mLuif+6XIUlrq4CGwRgVE1cq9N5pyJgExiEgRmEmcCiqejsKZV42Sv895G
cG1FvOjSV+zTPDVbk/ggZqzYbM9AQ0HBTKFw2WhdRrveKqbN0rjoebQpSH2arVEgAzfYULJ/b7py
yo1/0cSSOS9ZKcdWX3+XCi5XNUi0zr7rr2v9wF4MPb0EqSQAfNBLB2cnhwz2lA+WQ6E2Gz2uTH3X
4vdKh+inb2n7/TOojC0o3h/QRq8W5YyGYcA8LlOwtqi4Gl3yDzxoHMREaRQ61y3vzpHSGUEDaHA7
isPTScEsfmsBldeJgfnVM/xVWdqN7/+2TqE+C2Bao50t5ih85UWxvkhxmQbidumbn4FykVniagoA
LDznQI87sniS7dxP1eZtQo7fmQJpssPuhezBfgEJXFaXDJJj04iClDkeEZH3Z2Hg67RywAjPQHpJ
rSKIYISghNMMiRUfxzV5ljFUt79HTCv0qOwsrdIjiuGTrq38/Bdh13vcGeHvSIho7JdKa2r5Rr0Z
GYW7C8bIxGssIeHzv0i6OD7Fv6BSUiXaBcfslunRhx4d9+FyJlcfS8KH/OvzOitZoTSl7npbCxWM
W8/BkD198+4iXPmHHEMIeNLknXT2AbVmNtV9Cxb/UQn1R7+12IWAIMaWOkqIRBFiZ1r1KaBp+LNW
i55JkULkRRtEpDC20H6dXV0j8zo4DPncL5nmZ1ep0RQ0Q2qF0NcarULRxDz3pjOMzzmvCL0hHoUZ
ep8sCYGq9tqILJLT6Hu9ww33ZlKlJkI+Z7jLg7EmE+dUtf9W4si8EqVDVhmZvo71xWzC/iT3OTRm
RJQZ1uvO8GckEu23oiqz1PgxmrUFiQ0sqqwJ5K4pi6WM9XkiIzW3X4OzUvVsgOiCAarmrjZfDTrW
3VL5BRQTQCt6usBECm+kEJnLJXA/RvA7s8+1BCvoeRmrJH5qQXgQscnZuMpzyVNlWGoihtb9Vf0w
maDmbZB1pV8QFKbqGzvcr0qAPlYpJ/RTs1wxGv9AVrvkRSR65jbbaClTK8/Dux+4vPkHXRKdhwIn
/tIe2C3+9tX7B//KxVCoHTwJ0iG3num2Wa7FUlkQkCPwI/T/qQnwNHqzXVhXFwkYIO6H0PaITP7j
N3jMhiIs3VvVAE2umk29Q3cBu93MVzC9APitlw4bdWi0g5mGAsEtpX/Cxn+gjENoN+NhaVIBe1wK
JHm7PQGh5Jz6/Ef+2Km2gAUp3gdiaEJB8Y1S3BNlcClBnZtBvxV6OpRX8ljF5vCZ1332wSg5f1nJ
YS2OgR+OdCj05UgdFrPpPxHXHpCZqNNuuLpYl34xX6EtVY+V7/bv6ewUOJMK8h7N1C/bAZlLUkvD
CJqqQeHZPi80C/JyOAou0XjhOWyYYBMUwuJzFa5Sp8c/miVJW3okTAMzuermdwZU7PxPMj/WZPxI
S8Nesnk2vF2IPCQg2LEbJQ4KFynBhBBkbupQXPc8KXNnE/66zFU3K08+RhTt8W1EqsQlXNQgO7oE
nihcwZC3PSZkpF/08VBVPULvEMYuMMD/u+iOKNgOoo/zZkhiwqhAeQGXOMv1g/M8JoR7CtJ3h5o1
occsKLmWLSx6xftOhJKV8bBHzfMQ3023UR4gkMyvHWwJs55C10xz4DTPi7B3iIovepH2Y8EGG3cL
X+egdCu/ZHAcfogjLVyZL7OEmnaRngPjjqGXjJQ7GQecIMq0TTEvu8+gqoyoYSHYAWow2Koh36D2
1y4DPZl9FcBg+6Q4auySqsw5MFwJ016HcLz4dIL2hz0HvLK9fDW1Fj2MiucRSmvqYMZ7qophZO2B
waSDcT8cAB+1x//vUSe0TidkXtfjPBU2ts/hVal2EC1ohE5ms7e07rt9P8aQXF6ekGv6fqSRwVM/
7llkur1K6BQa4Q3zarN9Sgd64plBlnArJKuIKW98/cTGyyyqs0ZxSoHlQovlhFaXNS1R1hgUllRj
nSksHxM+r3FAjSXk8NISXTdhPcLu38vwZqfAMQN5odcy8xuWOqeXFVYNV5w+8vGPCtdgDxApIqoZ
xz9TETWtCvC/8LBFFda0HzhnZir3ctxVr2HBR0XxHivifmf+mPf+YQ6mX5CP11Jbwwu0BePEai8I
Yfifzou9MZQJVHUhrPi5jnvm6n9Bwohv1JPya4vj4axVKeh7YXPz4eQWNB9Heehspag3HRsE/jrN
v92J6Xr/PxemdwBxo79NkVH+HBvpvOeOdwpQCEQYATVVL2DEyiEKFB8UCcMMY1q4XBGBTZjZNG9F
QKpZ5grdDJYQH11yH4Qs51G1YnHGjdCMS4biDcdBxtnmaZZWp+Q47VlU3s3+HRMjgQt513b+ZoSU
cVdbQACmMON+FMdlC1oVzscyLSMLLC/LHV1rSTyYURsZG3qmV96F/zgB8wL//mY2mFqzj094hYoc
9hLwQfU9a5MvBTkmC/nZDIBC7S7kkQ4i4tzjk/PBukuENC/AQxnP12GTAMtzeILfx8FBLwDCFDjI
+bOPxzmJTIOWaRSE3cAlDZR1rs9yUA/Iz8ydhXM/N+pLsG9S5pDHlw0r+s1HAs8qYdgFhB9oT6yY
QcS3wA8+OK2esl+o+YL9yhAYBdWS69b5w6N0ingquHgxVlFeULYqM9cG6F+hrJXF2T12KvDtOYOZ
I1CJ+qsKWPbrvH/9rJ3K01EonVEAPXlhXnNws69J4VMi/s02PoxacwxEquEy+OJJ9bubtikY7NeT
yccYjtQ37wNFDnjhX6dZsvFSlApsVb5ezuKXFB0SrW2bWg1PuZQ6xSieXbahRtx7nZAmMk+Djuw6
EQL+edBZIt+KQklyy3vxMjkvRSlIu9NfqeCobUNaASVtizLNDDf+SMH0XLKXAOZhYeSYDjt0FjD8
o3ep1hPk03txi4I6NQgkt60k9yt3MsLgshxCR7VFah8TU0Ah1Ne+1m4V6kowoJtyOvCpxL4q9cxl
2l4Cm4WPvGIGaZYltizu7YFnRjbXhjVgUU73gaVYpSQDHRyWyYO3HUr6Z6JHlZi4O5r9PNhvd0RB
QDP0/SHN9QC42HNFGfUFn3aoV9mEES21KT5UkimLap5ZaE95kI5p2fYWhB+sNsJibZTq81mbvadB
hSN7QUwFYCI/yEUCsY4LtcA3m2yF1iG2zidTLd4vSeIb03+5iNRYzVjcYUCgsgfB7f+Fv7gLjhEg
4L4it+uTNwz11JZYihGxYIeHTD4jem63wHC3SmjoeLvf+MANB6bgfoWwxAGzOMXyjgI/PyY1BVOG
ULTEzxXY0M3Qh/Aq7LGV4eFx9YyR173SvI4ba8T7LlsyCccOnCbRnoOE43PY/bXJrJ93okY1zvro
P21gKC22Tdz0pwHQmafst1oFi7ZST/by0C6vrrcnR6f9zqXp3XL7eia/nQlyWLMtmVtpuiZ2dmhC
XXaiodIa6+s9hPMzezscLy44XbGrRfSmotZUuTxvU++Q4SGS3uKkHpc3UIE9kA5g/HV2UHrro4md
CvIOp/VSAwA5vIx+kx58XTqNwSo6jFBSDHlI+gVYTrpyfx8H4ZO2GlviwxRZq5A55CBUGr5mQUFb
T4cUHKl9D5nymLKQAWFbp7yasOeWHE+chKiAYEf6lLspky+jAVwBu/f4/CHHAjepbznhOi3i2ZiM
bnz2LS4VQZjwuRLAimtNK4z2ntmEzdkFjg8f/BdfJTaYfYf+RwkB9nMfsb2uz4ZLc9sUykx9gKlw
KIXtsgxzw15jCmvJxiVnLx7bmpDaUOP/J3tO7uaFrtCGzDQMu3sFjh3qgUbFJXWIclOTj/f/OgNN
8gCEVaoGYketfsBc9f7t0TBF/cUs84Bs9oUof0l2py6RphAxcVWOrJ6dZedjqsf1Eepz5ncQaRTd
rZbv+Qy6LD+92pn07N8clMfz8+vAl7/wvivcg1kk+HMZUPy8XWPrqBrZQb+t0kL5imS/JAixFlli
c9BbZP+eXRhaXHsfatozN+jniEKQU7t8a+0duKMdtklnqbAiAHqq+TxEZQ2/rtzB1UTts/6Gh1YN
v4SruNwsby8jZJO06hmFlqhK/O7nYq70MlI5mJQDi8UrubkhohYd517WxW2QPulJ/juTQy963wD0
mnSv5VO+5StToe4YlpsfC88H1cTup+r++gsg+SPBUHsIhoE71bdpdgkXriP5dQf1JGU9gghrkYeZ
WSNaXXu3Yyen9MlpK5h4BfbyU92Arv8IavCDYJhbNtvDUgHaca9RIHxScYlHr441tUyR6VB4FI90
gZ97/H/Tp2WL5KAnIsM5m81+4mhP0KkJM+kdP7AG98LcUlmfkv9K9fEMe+hihRr4F0qIJtWpEoCD
R/eM9nPf7QPNN2/jUXojQEg6Up6gWvwdBAhQ0ogjssHeeOXq7GSJiROrS3zQmJq91vkcR1j6x9d0
FGj1kHSCBLFngwbKIaIccVeTz+Eb123hFfZ0q6uyKsEkzWXrmB/5n+fCjng4qEtqz0I9Yb2Y18wr
ZNNyiR3nxzrGiIY4Ti5u4pbZ2ZxWaUVbXYyTxMWIDUBWDxt8VC2eAh15bZNT+EoLvevqhIwDDGno
W0uvKd5Jrkw7A8ueObOGCmUGLFlFEE0El9c+4Q/1Op6vym7VfXcWwY3CX3AihWoD/1TPN/8SpeS1
JGzWqGW8ogdGEydyuJHuRODN63IQWVI6zS5fffy0lk5rCUEvRJewOyfMAqKG1Gj+jOJ0r3Bmhu1M
2GHbJWTJCXvAhO6sBvyjdjemjnclFoKHpKxOVp4+p1z3vSWKZiJP2h7HJ5NumAyWzq6T+iw0alDN
cXGQn3k8JS3ixJ/6drubCd5EuLj2U1WlngVFvfVCthIWM45ezJLWR2ejIf4Bl5tbqxYrMJFCPGZN
lzH5ZydGnzA3DfNHO9IFtqqfOQrDAuGmmQ5AvEX52K0fCAPeliYQOWL6Q4sbKfuuTKt2npvnYTFd
v4E9vO9g4WQ6MqrVkVLR1Uyzkg/I7aovSH39+R7iXqlYVnO6UTEcxjENbVywHXjvsQ17wfh1/YEJ
yDY9alUM7S/YV0e4Htx42IsvVhkCnKDfKodylnkcO+rEV/9FanT2TcrX/b0cq/c9hC/L4Xqa6lP5
HQImIV4BVQNlWKTI4IBVrzuUQbRwrUygtV0sGHO9nXa2g2+nTFwCjm3JkNnlX1mhTP0HybB2bInl
QHAsBmQhGoX8ID7nh2RMT3f0GOHhbSn0gSzxZ8PDG2ebKOdowBXDwBeo0dmd/gPjQMdAcW5kTerU
NZmv2vVEfycRHR1/F86XEL5dRtWF/c5McCqcKq3x3jCHe5J/8hHmDy5tZV+X2guRY8L4wGtw0hTZ
ZV9ahxA0ZrcQUCLDHW4sVY24d/qrtBpTrG8DS1h2/Ri008BXMAbTnUbidmv8llbR3wdoSITtSM+/
tQ95BxeM/BsCK6ObTOiZ39JeaukjMyAyfA7VQ7Y8QWIiPiQf3rrjyIRLb9gXK5iPP82vFdfu7vCF
gN6xrcHHTzAfe4aqfqh8Mg7R+GuphhoMcc4mSemyQkNJfEQe1cO1QBUm6+CyXDsaFP1nDScBzmMp
KScMmTVH3jRF18eTAfatpNkCg2HmeQqajjSXScZPv4IQropaSAa6MZYxSE1VDvvO4GqCp6gmJNKH
sVK+e41C2YmaNZE72dGoIdnh/o8cE8wH7p0C/cdwCsWhSKzHwvidUSy3jFFvKUiy7F9UAO7KddXu
QWsjU5eZ5RDjfj1ATzjBMTEuGwUFtCWYW8NyUhCA8S3T58RtMYcyJw9qbhAZCvswTKbBolDvZmjg
awRCuKo9ddwVuy0X0IfqPOJXjTxWraPBX5Jjlauh/n6QSdYy2RLEsU4KVzOIMyd5zs/xKJ/2OF1S
XRKMt9Bj5XDMwE+Y0olf4DJlIC9HD/RWXiCP33HjtcvaAlRXrNGIB/jfeQZDToVQ4KwR+8aVW+jY
W9U/C23cay6azd23ihW1+4wFKbl+R36v2MWqtHmv5oGjwQAty5JuMP3RMh+8l+Sh4lrOTSGsbYL4
MZkgrU8PyQOUyXqxZjJ61U2EtsGUAIfrd0Ye2m4u0n53JGOyGwW+dJQm77bsvEsIf/jYI3dlsESq
yjJv9+8F6dRlMoA7Kxk5Rgfq2aXXifqQ/JBVkTwwlY6kKRUOPU55vTsn6MHVbJQ+FCT/rnxcbFBo
/j0KVTeyuqR5qIiMnh/xFz6nHItA3OXTQ6Ph2UalOL6KFGG6GDwYYzeqwxRWwauGCyxnTRFdZciz
ZqxiI9+M6ZQsL1NrhdkCJXi18WR0Z0s+10kmlKeF5FGhvKpnaMqKV1mr3/RQCP8QR2EUmR2NJorL
sza/mAGW/NVgbxiQpEhNiLL/Q/dO423NIvM8z4GRM+JZQ3y9DMh8iS6EJLtqpCBl+YvKG4nyFuIZ
mt7uKz1kthtGS9UzEU+BnyL9DZY9rxAR469UqY3oTSGcI6jYu55rqbJOaxrgJtxbkvdNC99quEnI
YMnSyLLTa+zn6Fn7j+6svuoMwRyaBtpOw3I3nUZVa6irOA/uJ8Y8ej5hVxkfqjsYzHSpVcTXz7OK
doYdPEAUw8hytZ0/5zIiJ9u7GksLdfdJj+SqRs9Gro+jriz3Wq07Llw/XmEHdAOKN+7DSh5r3EEm
Lc4G6FdxirP6JYrC7GRBwGnD6pr4tdN6a9Pom75CHpocYRHxFnctOPk40toPW6H2sUm8rKjDfQod
g/x3sfhjhS5c54qJ/l0RxfvUJRIe1L53gWJPM1ErE8Zx3OqmLWD0mJ/kg7194/WAK4GkupBhue24
fdWp28QQobTImlcerNBGndq4P+rIlFK1frG7+i1eEpEwwzRKN9F5YlAT08wmqnEgWgc/KfYQ/eL5
0dW4oUv+H3Yr0clg7pVHtPkawKrW3u1f/jvwCWFBahh2A+mpv8nTiFSH34dq02yqhKMub3ehiA9A
3JwWIHCkX98e/CAa+4mBLxtu1/z4o3vg5v8hh83EYAg3hdNgi5+V0zps0UGngDA5lzyxQkyplnpc
VmNpu8dEZT7Rjm/Fm8CVxnZI4//pfjn4ox3FjQFuOrRdxgI3bXHn4tMA9W3fomSNFqxTZ2LE/4u0
cjNUbph0q+Ia7I9evSXrYAU7TM8NqPHYCvtILgx/RwMKMtRKGiMAqP3MIiSialOoUic637MLuDCY
tipSH8XGNxDjhsJhT94qfzxyOdRcWzsoQY574Hxg7tRFPue37vQbj8ujtYtamZAmvAUaSXtwEHRm
hQnx+ze9BtfBdrW4s+4JK3lViPaqdAlS/Y/iPAG6OL1bDg6IbAC/xeJWzZOqna2Lk1FSq94fqbnC
P19NYGU+2CGScl8P6Srwf5cPqOJmbLR8oAbDrM0J+/E1bupEmNie67W1fYslSfdiNlSgG1R7spKE
yy65aOZsIZFX5Hbv94d+YTpzIe2og32h2mHglN9/VIH8So3IatwJjAkgk42m6XYNSb6mDaerbiy3
su1xj+xF7knyY3cXwiWm8xv96LeWowGL9A2mSPwQUiQ2PbJb2GiPyOgOOxI0iNC+sa4G7x5i2e2k
5MuWq2mGbtQ1NCmwopXrxM0koZBHzL9ZjzlrNeZ8yS9CKCDPUx6G2b9SBBkw1rqfYxlRlFGSF22S
whY1rKYwQTX2oQ6/rzposeV2jVo7YBbZQVrIO4Xh8KZ1ApWRC23SQLKO2EsHE7b/ksN3snXzlTQX
belcFHhYZU1YcBI2/gFoXNrxGcUy5IEBOXclxaHzqt5m/ds43eaNphvBk//nwwqZqwxs322P7XCP
IfmPIREbILG1IWN2doCma8pUx40qyXr9j9LEsT3PLrQ32702IaCQvFqyUYH2pfGvykMojgKv650Y
OyqESJ0WHB77mJG+5E3NihgK3G9yiG5XhI1W5bzm71TzaphswkmD/CoVDBKv3hcz4yvpYysLXwot
/k72GPtxEOoaB//R1GOCy6d1CDRtmYeduHZe8FGHg4tszT+20yKUId+A4X718eLtLjhMaV7WBGDo
wTJyaJcNGS6PRJT7Nd7i9V1eTGznTf2LPG9G/pJtxBXtNhWxTkHueWUgwjB969h19diIuWEJKqd7
alIwVbyMNeQ2JcFuJxdOhHPlLCI5zr9kysA6HfbYren4+Cg7vT1+Nq2n0HktHEG+LKDGSBw0svpw
ZNDy9hfVojMNix2cicXTogfSreYh1267XekLOj73zg4TdQRVNkGFUnRGdGweEA4fWGfGuqSZsERb
HbVauowy8sw9R2kdFIkYcETsRu/NMfyCxhIqitCgC3JONYXanOR6WY/1dSyDyT0F+JTEAGftRmTs
PjPQVAfvxhMPBMPSY3HNpvrw1+lXnx92BKU5OiDML3BHmzW16eyVHIdEH8x52BVrQlUkhboKBuy5
ZSwINL5JFxGhOysgA7BG3TYzqT93feflT68AK4ubTtVD04Vo4pIbe3aG6uRsM80+EdbeklKLrkKW
Y6hCM+YtMxoo+2ykIbJNc+yrH3YstQq5KVyY4m/Gg8LPMYGPaFQiSSOigBbRDGAngaUXx80ESfaN
EHwNKMgDlvOVBMUOVnaRBW4yNTCJPspDaTwahh3vJ5aRrOqsgt8JhEmMUjPxrG/jT96IiP2uNApN
4zbGW9/Wf7mRnHDne3ZioEpY/trSJzWrzb2Pq+2OeSvx29o9Z0rf1JZx9PhYRax3NJfyGWM0R3QK
M+KXOJvcLekFM/7YYR393/fcIdbASOwbuIQhevl4hKAzrcUFlZYyarpg07UMdYPcy6hHRhcNB+ET
octLlaK2R60buQHq4FZmwBBew0Qhex712CJZDuo5cyLcPtc+wCbOKaLOuEHX3j4Kgt++yyhTP8Fo
XlSOpunEU49TFCr+uj4T6TDhWxln7ozKoMo5vCuQkcTKLZjS0Hnbxzgc82rd67y/8h/NU65ZKPFG
+CDj0VlbdKlBzUi3C6koT5hZbsF5lUkhk2zISRhmha613YeGaUdskeW1syVf4CVOSN66URXZyA4T
Mkt3Qt2gnmXDQr7g8ZkYhnDYIMbqP2hkz6NxXriH4bhe8LPfQOr7JEinl92+6OPx27Oz1Zvd/sBH
pTGxo6sf/p/XmZpSocxGcmXv4cb1d1KKZug7/0S7kd8bRSms65i2vKy2TLkqjrBW7AL3idtCJcSa
QXoYr2hyfWfw+gjK/Tm+7uc59fDqHcYNCYFqnV5j+76YFhLqmPpqCSv6Ze0JJ0Pg9Sz0XjpDS8mj
fRODQqKa5AkmPfvLGA/9fMslK6QV7EA4yVI7M0itwRxK2/696NSxdKpci8qBezTXK3Mr1XlfP/va
v1SdtA067/BC2O9u/XVuTCV2xgo9Jfe8kiX8+y5qaJjeQpD3cYxywsVLlzUaMttnANuyTF76nLGW
F0BngER2PRfXa0HOD+OyJFmXJ4Ll6Q9x1fqNYu02/4VCrm2PYGWEXBRl7Q2X3ugiBXojyJ3i9kBH
8SilaXsp0JlwUpEbn9zjVrA5Q53yAR0gZ7LQkrp9IOA3Zp+vQ6sVjgvSYZq61XVm2eDO7bDhMwLu
kM9ogb4VaxuuFkzTZIj4Fi3Jc0SfggcM+6Tu+UqC4w4XTkWMOTDdF7OFrRfWT6pwaNvhLVbhAiqS
TkY2tZN30coLlcEtszdQrkXH4h/Ky8gKHpLj78bN6sx+Cwt6Y1C9NVrqiR71veaQSM8HF6BWISFp
efuKqJSLQcoedEMlEOXvsFJxta3vqMyxMaj5a0lO5oiC+y+M2wP/YcH0u18iI+OlJUQbIEplCEoX
3w3qbaVw+XJ7n8RjqCKcEwJCuWTicU1UzJa0GmubRpZbpDzQ/YkoE6GYDZLRXisGb8siz/UuMXVJ
cYXXj3xFBZuZzJJvrwvT+xdxDYkZmTw1j6iM8E49QnB9SlPB2htP/2+1rS0+Jh+h7aGRdkxztLbG
bT28CxyETgKCvv/X7KIh+BvcaCfvDUXWztCmYwe109b6IJo2uV4MWkJ0Gf4/bLxMuUTzYAgfZGEO
GTZCdm1s+/x4cGef6nV1VkGBrJFB8G8RLRi42jvVp8pwoFgRu4oWKrnulcUi1X8etGm87XUk6ayU
kp5oMMMSayY/dMXGkjgD+KG4sjCAybsruJd7ZwIwHsr/p/IqbDBKZiU9R00OhiIYjAeNnFDL4oSr
4cjPYTEPjzhuQJmN1JDa2fVXU1fPMA1xrtF+cTcJkABforKBRinFsxKk1nF796v51a9/cqtXiVsz
8mJpkxOvzZriGx40M2NuBP+TA836muUvAQpa6ZTXpa6HPav4ehs+C1PtWqF3hLPWm0JVIAT5H0PC
vcq0M6IYkAaKNgp7N/Mj89qBFtF6Ow26REKxNeN/OLQKdfz5jHy+l/MwDbqQn0ZyYlNVVhh1u6f3
mtpZfwP8WPl+rgTVBakJ+GJqb/4vShYQ0B3TKTyIlso7HVG0jw4xsFVO9QCiU8HDM6ubXNr2xwRK
yzaMfVLeaHvQqvclcglx6UKtJVg45UssR3I4PswFtMRPvRNLCuEbaf5gDMZZZxkqKNvfud7PeZTP
Q8Yz6uJohX8srr8ybaRcaR5QQ8I9wFWPzoaX3mkwiZbfltk/eXSs5Hrep6HmiY+35F3vJShQxYAh
cFFejSd2zhCapbSl9jEkHU8cTrZNcJVlpcRlYsfigN6C0WXXMXMGHiD6XyX8hmT1jssLi0EwPYQb
c0cBsc7TRMk+oJx+MzqCgIQYx7iyWoEfuFmFV+gV/TqVaYfRTEiQeMNqdsvUwsrN7P7J96iMohYN
tHQGhJEicfRE6/kvYg2MkMI5xyOwgZXKBzU3iDno4mq+VAwwqHMTJaUJjA95zEOHjspC0tx9sZKV
q3AwfC5S7DmZ+NbiyQBnpr5kmCPE1vYfGv49GZzcSjgbssHIAC/s0s/v5e5VvyAG1wN20zNgQWQc
xgmlre53YuyzFEZB5wJU60G7xykPwqVPU8xJGmKEvMmr2Ab/63t7GfaO2zFAPODiVZOCKVkVg4DK
gj27I8SE2qRtw3eWn3baj3g2A1NuzuxAEKoY/tKYt48CvAnJr3zVGC5CWe0SughIk1n7HDN3Q2V/
z+z83py+0WNYp7Js2NTdIslyQFPtz5ST6UqFEwyxM8ZzZIaSoFOoFleD528N6JUQc3b2gaS8ID4/
/D2xkC8WtIgmg9H5lOj0eFFWeNF67x7j2AtHYa5FjTaAlY+yh1ciFDl/sBofxezV7n5A2utZS0CJ
iTU87/me9TxFrbYQ0RQr7+mktFrwPq0g4uyFHcw8wKIHYJAgx7K0yFK/neMcN7YYDToYokf/yVkL
gmC537ZzXpV38KWzQFzS7/XEU/yOyiCAwQ0cHGyJ8SDsTQ3+RzlcxXTUBpKodv/pRAdSXCMDoQza
mvNx6zQ6fiLSE8+qAaXlxc8CrgV+MbUjeWwGWD+OpavdZiuqS1jdWGwf8930ju+xZJkJ6cMsaqLr
9tQiPjcYM4xcHxFHpGZATw9NbN8Gdesu68xB4s6ail3rSndm79ORgIjMzIPDjym/h8b51+Jx7E34
1UvV+r8vmjRQwd48qYLK4VINgAG3xF521j9SweqKM9yUY0BwaQGdfcG5xFBG8B3YNyJXN657+VV/
RAccjFb0zFcu1iMcQatHuU5Kf35upjWvgIWII47FmnMaD8HLUguoM4tJ/IlZ4/YcwFFwe9ZmvK1u
czFkHppLr/A0LP9HmzKNUjqv0xcT4gESsApw3oUeGjNR9uNVL0XXovMuUQKO9a3b8Sr6/vNYZVIK
O+8pwFRnyHiRqqxaTZLVzFcMmgch8EQtdj2HMV/xhPMoNnmbFmSlXdJQE2+FvE6Nb4jJyqrLu4Da
jaByScaxaveppaDaZ6vjMdwUW9I8tcOtAsbQ8Ylojqza+ti0UEUnSzPTqBI0JcDKpTR0VsxlzIij
GuADJOYkQ5395ysdBK9eTWmrlQ3Opmy0kKJOcVl+goSQ5N5kSeq2rnAdF08amhm1BSdh8Yg2DROh
irRyCpc5314nl1RIs0CxU4JclQLmK5JPX67v5+ozGJBqiZsFflXwHwBlMOGOc53SsmoF/l4ddkiB
GN0S/HRBouvB/pcg8taILwFQFcwXcPOCv2IZy1t1HpgmY8ZyQebSUP6BkrBeNJGHrPsQIimM/DGi
jiophNwfAI2LhMmqbEi7/Hu1HGZ9AwrFO1EtyoN7S6utNk8cy/t2ZLdSu7pMRuT1Rkx6JDC8GcY8
Sb3LPlec5jITMFRXslaFckRlhDtpsmRZDEXmNHzIQAhsPOuAyVhWeAMd3XecBCmsRTfbC2kcpqqG
Gdv0uDIwO2eFfzmqiVzZpcZEkieOwMfo8YPAXjTLPOXHHk4YRUNPyIvmYhG0ic2Lf1Is1gmz55qc
arWa75rXlx6hphSEozB1mksCaSORY5UV6r03Vk0+rC8fjfw8y1rev0JaIGNsMTxsT65s2kGiFxln
N9kHhybeoccHV5kpZo7F5Dj+Pe2gNMFiuvUzAckockMbXUWaiXuCHSwZ8n1fXtrNXYagy29ox740
yi78cx8oGXRQwzNEYYvPLSEWRLw2Qf5YdOe/ns9GQI4o2XFUhG2i3+15NWf3I4yTTBqp6lG2Pw4b
sA4XZaKfWGAwGWjkizDQ2/Ct/NXOEQgtTK5nzNHUOOwbOoRxxSaqbLscoI0Cim244KuM7xS0Ryb7
+xZZ/Mk4D5rebuY1dfr9w+EUBJKPs17wBrA+mowff4jbyoWhfU42NeO1WILrnVtoH5L4ITpCPWt2
rOyx0mazS6Y3foxOgGwwQwoFosL9lSszxkD7rZcz4h6bJi7x+VvfdeUi9xmbQOi0fJSU3mESAl5f
cxumcqhABoctN4l3S3vdyTCGfUN4PH0B446zi5Tsrai6rFyo2EcsKPRm8MGw1xzo8y4u29gGizpE
4Sah2L07MJ/2DXbwID7dAfzrxIkbA/V9QAaP7kJSwfJiZbfQ0FyLR9Enkr+d96OtTp0SbKiWpwqY
mQ0UNFqY6bF20dyQFBaQdQ4uydAys893OJrk9hh0T+qZllmPlqorCXssy9wJQ56/HhgNjZzTO5ex
osfIOhQ1gv/+xiEnKtg5mxVTL+MqJfZGroL6basIHuOWDtDPagxOGxqpwE0lEcySvZCxj6xGouAB
y3SnucogIByP9SyvO726PP8hOvdCeeKa8UWfPdSXLJUlncFfu1qjcDy81ohLwTHFNBKlOX8DY2Wz
921m8pF4nnj/opZKTU8Co3BNWIChwAouQzpBS653A2EzNq6QfYu8Z393Ko+IZqNjX2uWVlgGmfaW
yOdv8qLeGeGYuycVLR9tD3qUeHagaJuYP+VL5+JTMAlsGOVQo3+6AcUCIuGwFtOW4fsAkeMHoNGL
bXcT4sBSRpEohM68EAv8ASYXRZyWNQ3CgkDp1opD9Py2wazPPg6picNw7gf2Fs+ZpfTK81PNw5xp
2S+WsVpWdUV67ULtu/db39ulrSb/w21tCKxu6L1sGLgmDUsZcUO7U747u8ROlVSmxCvQ4gpfAoL7
jHrrPyrI0YOjPT4jSHecjXt9juH27g+LQ2BSQ9WHbvSwbd5fpunN4ByiPWU1G8swlMJ0SOWP9sg+
LurdaWP+AK9I+CpiySw81eEX0RJV+mGrj5SxSxPnMDp5cE1GCi3jM+f0OXnqq/m4XS0rclUp8p0l
RI4vlxMCPD9OpPpGSNzKQyri9a7kOEWK1JuCZKOCer57DOmiCejAi1zDrdlUccFk9oHabH9vrNrv
EPqB2T9ruipOQCM8mj9e3jIn0uuZ6y7Re4MurI4i6E4Yp3mSYRppWFQLFqgqr3MXn0N98S98b5CE
nWTDRCB3dHhpfDA2WieNKO6xq+aA4JkgLdUS/ukNYbIRSKOJdMN6X2LVG0diQNtJeWRVklpMmipY
ckzRsKLwR+zRC1dEF4EM3c8nGEbCUqz4DFpLN/DTp6soLnzWcAMJlrVNuvKuHXA4NtXtVJ0fWpNf
sRRSyGjhPAAybvd07ghZd7WqAKYJdgTZaCX5yt8yB10k4cyFGL3oFVhZVpmI0Jer3lfjO2ZsVOQx
Ry3WKp8avc668+No7/LETliMe+XFZfQrqZcPMOHB0K2W3zeGDpSe7gW1hbCm8NFpxID1k+W4a1iH
8zy3upPTVJ/cfkIfK1Bn73GbetUBBWEcUATZfR7Tu9p8QKAnW2CryFLiZDoRlGvU79Dt5s/TwgVS
FzQJxz3+eyFdXb4jDlh09YpbdhBMWXvfXSbGDbiZynM+oDEtf3i/U2Rzg8/6TSrwUUxavRmw7xNy
1tCK7DD9bWNsSrQ/sBD/ERUrbuludQWj8fgpq+y1/kpb+jS5qMAeBgx+fPTUcWBagDw1BmbqUpo/
bVOaKNRbNhK27pzAl1O6EjLLaCMHvLGfyk0KEFg53a4tSI/6ijD1UAXLhNBoCGsLbsY2Rt4EwmbF
FU1+6PNov1zSbvuyq/ds18Ma3hvozndZ7VEGdn4mpN72LvcijLScoKH/O0G9HIOdGvxfeKhnCUmJ
603uEZJIHaL37HjGcnKihd2RqWSch7nxd4EPEDmE/VTZKsci/LMb6ABbwLY2RiZrL0jVuyy7+28t
jyeNeZoZAGWlhJxwmN+YnMh22uLmSmx9g7qyRPcGrhJHZFCKJwJ5+k8ilepXoVIOr2+/ZdM4K5AN
CKIKPUHm/Ov7XliZxfKov6K4icLgzasm7SEL8ayvhOIZvl+s1TIrtlFPoUd2J7o2ai6MlVTPa9Ri
pdT37G68Puf8/BCv1mQ3Jux24ia7Dhsg9+ZE9VhFz2RIQhUCb5y9nq3VCEB20ObtAdvzh0K7Fg0V
Pse0maMBHhOJvl5EeV+lbTVCN5XOkv+/ZhmNys/SRgD9fOjfKW5YHl4AJv88D26D6It/JFzr8Xj2
QzivqlfTbvKGwfuEfeMCXJ43QEDS8FTaf4uI0URmi0ot5QN+METTGFOhV/0oGuGzJBnOvJC6gEi6
YzKNDOrf+ENVEVfKXTAWj9wccZbFqx53f9MUXOZbAO7fScgglkwERgp/ljSHJHcFKZTkDIY6reds
a41rcwQBvG8n70PZqcOynCy98NmLLmxWkGXFKfOITU95vUtfcHdzxc18udn+U6XR9opsDA+9DAL2
9rb1z+LEPKl1j1QbyBzzEZ7rI71T7fcr4PgwNZwDPLL7DKNrJDzHx662BOjvMbLFQE9Cgd/9U6L7
9q//itVZPfJWLUTVo1jW1XY+1euPy+8IRg0hgsxSBQ+U9JfnI90WfGQ4fDolbAEoGaIZgsC+3T/l
X50W93pEeD3fOCBLCFXSXcryFFPrLTZ+vZVSwN18I4d0T2syooZQuKIs2g9E9qsOnr1hUSaUy86k
PnytCoAiaDBsDYrib4Hh/snzh8j90FHD/oLs6SNjvfz7CH6RCCyrWxf8QoTulp+jOVLetTbN9tgt
+1UbcxLQbOVja6TcHS+BmHW/FaR8OkBco48vf3FFmZIhclXbNIYpUGN241URLAcwh+uFadPtZ8N3
WXqmga3BG/BACSHGQKzu30v3ipHRrHpynB+Oa0ktfaVOimhZCATzZ8FEeDmd0k4W+JJ/QxQerX6u
R+AFDaEog+GuSm1DmLO/DwiutNCy/nWXc3sivRK0xgeiqImmlq+y/k48LAPnwlPW4mt6XSu+Fgwi
snI5mFjDdQ0u7P+oyi0rE6+3uE82v7EGv0XQuN0NcsTAyqduP8JRaIiHj3+h5lO47oX+kqfzlR9m
at8XraapqI9qYXWPVX5rRHOQGeN6ht4JkJ6370FSk7l0RTWo49B2qaJWTlIBkG0GzGT7LfjZH/ab
SJKKv2aI9igCtxFnUG0e1/px03N6CORyKUwkCnrKSQbLUenhnV8wAGJ9BaxD583srXYd/UYRIKiK
Wbbs3O0d4YD/RVzRWcclVG6s1rBqzfNXi1/7lBovNsXDQKKTELyoTxbNilyFcIi4UaI9SeeZah39
Wa0tOmK+mdQxaIA8rcAz7/foS/htwZgwXoUrytFF31624Ii3wZ4I6+N15r7NHnvQ96FCbVRrRK9S
VqJcLx+OXDuex4Ay+k5XIq7IDB/lCJXcfSLsn79oriDWwx/MXmC/IVHRQkOSNXmIXmBjibk9qDWz
kEUuTnvoug7ZqM9CuLacbihSIsiEm8iSRuPa4lWpmCRj78M7Qww426s3yiLkflARtpqguZsPVvyD
m4sVbk04489trnG+BYMpFdpArU/fmF349hJLomeWg/puuvZ1WmGJHP1yQZuIVAeHJb7xFKzK5Eim
/qEGtlg3Vz5QXh5eJLN005amkyKg5hgYrolGYXiWb5Uq2k1gAlGWrVTW8jn3osmcfMpKTRZ6E23D
MiJmUFtVyXrbG7uD5IsqYWubHa/Goq/bVFiSQZIADqb2o17L4PtmWtwfSRosLV3dV49IojaPC8ko
rDs65HeRJv/Pw7YwuTfQgGCLsYTZzGNQ+ZVTNbiRqSZqRqrwDDl8D+K3N9mz9LU+zciCd6Z9jCw4
fIdnv6e04EhjgULsWBnWrHRbCYfpbRoGLDlTndeymFErSbnWvhr5g9eY0IcAzjb3ihABIh8mc8Ba
WTzzwraVORlVXYeAVYYwkKO/zdCbzXToLMp5UCUrvJGDtLDp2peutwLObHzt+U+soU6py7so4ybS
YJGNFPBmvg5Z2i7NVtStbThZNQIMCCQhHLgCaiF7XyaEh5413xly7oQT2Nthmu2yyhNqnRktytfA
LKjj0n0qus3w9SyRNPpB6pEh2zM/TqbLyz9jrwx430hajSsQmDj+oLsOonCUKgs7WXJe+WFng486
i1xc6OboWE3faYBb8TpmQePVe6OzKlN4LeNfgoCBYjMoigObfgVyvAPTIKBOxYMqtpgNnrTGMEj1
yH7X9a2CMyg8LuE+GiugVnlHmPHIA/ucZ6fu87XZnXL4KeRWYmNnvHlb2+kNw+Nkj1UJasJ5ddcj
soe9w4/jkbEzqgMa+YyTIzFeSYXzwCy7HwbFZsfSUcxLfXhb9WcVZPSGQmrNMCNKkGCV3vpn0Lvz
itxm8HqEbvB1D36miH4ETMvjXsHZk0/plpf78OJgYEItEdgQS01irhnpON6TXz0r8bukru1LvFaE
NmPy4VoT5LoKsqqu+7gP18WzIJ7CUSQfEJtZjDnvArEGx6prAnoSciDjtAub2pBY61sSN2hw9qIV
WKdF8WqF7rqOTRwLorz0vOH4+aK4S4Bta8P+MErVlH+dpiznEx5h99vYTNLDIc07RMWaLeI9I/3w
Pi6Rc34xwhGcGzYQJB7UtE4wUaNV7s9ts8iiJMXp/DCaVt7UxfKk/qZA34ucEQ4HMUDrnLWXimY9
OLXFD9WrhyNY2kZKaN4cslMiqL/yeOkfOop+DKwd0R4KiZ+CDM2/ryWT8Jn38DEkQjiCZk5lKg3C
QSSJR018U5iaDnKOILZhnmGETHgGHG1eLVNps3P8sluQjuqp/n7Q7EezkFwCSAjssJCJYTQquO+G
2S8JRlNSiq6b/GdUhDKCsqBbUCFNm50LvHn/3T1yv0J3FNiGROH+QwtmCM2rcootC2CpZf5wN2NH
c/RgMmvOc7UP8KPdlulA0d/VtSwcM+e/h5mmCLLzNyFvL0C0bZCAYrDD9VAIbmxvAhh0HXCRR1KY
frhFIY4dO0RRlQ4fVeMKHLEBZTWBddX+euWDB2fN6vnbolImIRKlu5HF52LrBMT9vLHWlSfi+23F
8j1/eC//bHXw2iqlrFTKH/oiqxwiITmjlVq/xGveSz6XdotM/Qu3/TBwLXcrBfPlOhYfXf4kidkn
E7cpfUmTb4PjsXiMgpttOIuCW6M46gdE8BTZy54CDjiImDU4hczth4eqIylIy7WTughCy6T1tJdS
wQHxUcSjYFQivAN2Uljmftg/DfECHbWBF0tIfX89gaYEpRGFAz9i9ITZ9G23IYpjyrabO0RSZ3a4
wayEv6dwiTHUE/gVpUy/MtXpzqoP/xuqrHeP4r7n1ERSZIQwFWYpoJEqn8dtCVrcK5Xh33lZcGIA
AT/F3uXI7PP9wYXTKkoZsrJhQaUYSnilDcg83jHsWwj0arKLXvHVGL8Qlabsf9ehiq/j3yYx61zb
WPdnaOJvwfnMLLrVa6FqESUzehusJAdL9zwnYId3BBi4l71mcnlLhaNpQX51Tg7ueeQ0qbseRGkq
yWBdVFAFXClRVwLLf1PlqbsEZllLKsJdNX4SeAOxcVHCd3lq/xrbDsbtC6w+R8dAgI4pHbAHQZ4V
QnGyxt5HIfGqgIBWw8G7TlJaVYUFh1fI6Ff/GN7nsUd0vVWFB6qBihIJ4Vm5oPy7xTOJbVXJ/gnu
RnFdBV9ay4Lx0XMJwE0IRfq2VnrQvLkMSSMTXvKjkszcUATbaRe1+EQBb5tVLVqH7YJex8lWmkJ4
NcZrEHaps7H3yLztfsHRiCzeLDsoly0P7gGpSOfyp2ReqfHhsL88TRTeoHfxAo8DSi38FgjP0BIT
zlEX3MmQgwG36bAi51raIYAGKafgmmn90/QAGIqAXY3uRI//NFnobR8Jbn4QOgN5oQdfjEA+VqqZ
PjPhWuNvMBhXGgA4cJUk/mbX8zCeVs2xZTkCKcUUI82MtpaPn+IK32SGhCHMwJUSyL6O5RzgrIo2
7FmmOi1RdRxzSfOmGvDtKOa/xMctQ0zvaBbZdca4Li0OzYxt4EVotHYRKLrPdi1uFzOAMiwrxKGU
OoF40s7TcIZ8Oj2I72RGQ0mIFbJB6HS2zEIutOs8tbeC4vf0RwxOPAtLVgdoirax3zUCLxolmQNf
dBcdOurACNUcGvS9Tw08ukFTRr6HEU+oj2Y2GSOGoh2qNInfHZQtxJ3UDplnGf1Vv56cPHjl6k7j
zPqUj4jlzXdhFCSlEWD/FmwokEClj/VOy2jxu3rv66B5jX4iMHdMnbYSXu0r/9+1dUILhnr6FAqj
hATCeuADI/2evQdGQiGi8PRa3XCWyA/xwEZ33XWjNK/+osiHaf6YClOOztYk0VXPHA7HrpPoEA4L
+L9LNwNbzFMUfI3+Ti2KRDPa7kuFHazcPWIt/saMVSrJAYKym/GnMaS64hb1tJn2Go5uYC/iwban
GQ0peew/dKXD1c1XxGjVfOOv/G/xLYVbQ6EcEv7Trw+nj0n2+b2f1edrZ4Qdc/oSEp9dKhTbrm+X
ShsemcrmZpvbNC0Z//0nfRkOAKWJML1t6ylLMDr77a0g6AERAlk0Cf5A0rUUP8ong8nOk8BvRtH4
4aqu415G66nwVlX1Tv6xRaIhkZG0GpUwQeDBqtJxi/shwRIPC1aPHp7MohKTWSXT12ez+gjFY0Cy
cIXJg6YhLRJvZE+MKELQD/OpE1a95ETeekEIqmegwz+y+Ck11buooHuxToCHqANmLbaF3O3NLt5H
HHwgEIjiOuUudNa4GfaVZEalxvSEZGxL0s+OF2r8UjK/l91UL42mBY4kry/L2156qAkoqbE9rhGI
lV5e+R9b5rrJJr9tc6M0teeixaNqG64iP/u1j6bPLwo4RIsoCpPDIgV4o62/CIZNSHJOKC5xQhW0
DIBQTOdpGxjjjMMCO7PN9wUgVD3nR/x0dkfYkHpLz+nDIYkDFkWLmvrO97s0dBvGES7FEGLg8zsV
fcj762qpjS1hy0U4/eHnQvrJULi2mku8kFEQvPzFUJv2qmu/bkZOpEewam5YlQB4spWZRc4aSWSK
64ADlqula9GxxBOpXdyjRyZUnMirWVzm0J1nrIk1qWV9W3gH7L8bgMqARypQwLocx5Np61n7Voj0
Y4dw4GqGghuxJ+7LpGdOa0o3Fe7IWqwINEZ9Akm23348RqaGALgqvTzcK4MCOYl7c68giexdN23F
zhY8USc05X4vyGoWQZplT4ChMEUG6bW+eOR6voowVjPVl2xPT6xq50WYYAlIcXj5UJP6ZSwHQNyR
m3YK5UbV7W9rxZt3cYcfqBnQJETo5fax4IEV0u9qSfzez7k9HLxLCf+xxfrpbVAm3It1a3o9fxV7
RNwbBl0JvbUwl08xyGKchq1eByXH0wMnXaYxyEL+QZfJfAkW7L/ygjFufBN1DQuxgiJ0GItsud2b
5NxgOlAF7SIHY2Zq92ejU9d3YyKeaF/4lROvUHIzfUOuM+pisgCzIv4TSd7rzjE7RzULb/Iv8rl3
F4yeX0pGJZ0UUZ1T6kFG5BuXk4FTKSdMEM3m55obAk7IVMQCIJKAspr4RW6vHAnN6oiYPMA5+vOw
JZjIiZS69gu+I67k1v0zFXArFBYPWk+3ytaiBj9tjRsb89yXwANZbSSLfX8kuJG197GmpH+LntRv
bLyaMJuyB9ZkVPLGOfqc3Mtaxr6PGyTd4rjLZQmn6IiskDu8Z/zfFSWkeng2oYFb1LCviPWKMsdw
GOljda192RIfyYrVfZLAZbliKlt6pZboH+1NRHpkRz+N6NOvYpDtBo31w1SD9shE6CyFENawwCur
dfznr6COvg54egILyDXfG92BWvM3DU9zlQXuttvOXw52Yq6fOhw4jY3PZ8WCPqC4XY4Qa1uPjdKC
T1u6QIgweBC2ojY0iee3P6crYPhClv2pFKo6ZD7nMhE2SYtK429pnYj0XpNXdcZtcue6JwoMm+kG
KkX90ICHEBClMCK7pT2UgqaaBwQTC6pQ7X6Q1+RZJYihJiZgDNdRgHWWEwwOJBcrdAOXI72F1PB+
bqTV/braHkIezSbF9tlG7+9gYkpCTBL3Nr2tYKH5upyLGA416XFxbhikBRbopzhwyH680j/Ak66T
i5prBe1uX6VIxwocaq8DvQW9h8HJw+4t+kUsICdDpmnFFByql0v4ymtbJcSqy6c5nKTHv1TZON/w
DVBee3GgNoE4lnzuJMc5RQoGl+IGypPlU31V1fC84BDascMOTszOswBcgvthWen3t0HqZpf9D+Xv
x/kLwReR44Fj0H3Mmg34KJ5ySQr1Deus15xyu+d2UW1FMtvq4RnEUNFTGL2zUR3xuiyRBNEzLuDG
kiOnZOajl2EGq5oX9U7cA89inqxN4/QZ8An6uXupz4jrG5osM6o4se21OxWafukuubqV6yQDhu6M
jBnBiAq9fS5viERePxeeC2umFqUC2/K0n8eyWiltJE4K2wApxPDdhTCIG5XveQjFUXqzmz3QiR7o
kwTcYgrA92Z0IJ9RNvp9REI3+WbfFi+vp8hrO9zE24kd8l/JRDw8EisLyL/2sXirHML3mU90X0Kr
EjRt9Gvm3sCKaTG6AQhY4V79KDWLzVDcwMKkHNWJwc8eZxZdxRBBTHJEIKzcpI6MTglFRQwcCtDt
oJAUxUvFtN+ojJc5w3HgOuulcUH8xj1qpGlo/AzCkYpKfCEEtGtXpTH01ju4nZfudJk2AMQ5gy2G
BpA5laHXCQalpt2xws85LjLTB5NsrnZ+Lk2+x5JQvkBJVYCp4RlB9uYPJ4lqnl4SpJOgYzOseoiv
ICc+6G9k1+Mm7dDgqdRD7alE4poj9dR4+B9ikU2rUnvEKf9jb2OWP8ReYWa/GF4yxFqM7GLaNQBN
oESRBdB8D0TnH18jnFbxGCQbLc+D7B/tZ8ZxWQMqkXAgcU+XNQYIYXqHFZYcMIQ1yz5IP6KaWLfF
zewFC28D+OZnKsQ2wHW7ElggX5VKmxcz3j3viaJprehIh/+/UYnFR6JYAEhA2UrKo7Oz1ot1gVzo
BO4GwagZ0TaCf1Y29rJd5r9LbtgnPPpv0ZceOkfAXma9rMf7QoIWKDL8QNX5kvdJGvwKo3Ah/TxR
MjmiHlFqJmU9v7UeUOpgZCjo+JK9JgoirsR+Uajwh1PrJTTprxJh4Clpb0ev1bWoghw19XmMNt7J
6cHqD1KzVfy1U4mPnV79SOEmsskL6x5ZvMMWNAC1dvo6qAwkhSiz4SyJ2CivgFwy6RLlJUXLsi2W
LpNV2GaHWrRDy1fAoB8kvBzcTkqbXCLjMuos5KZ3DKM2mBVV5JMdGFjDzhE3ymq3sANdxrJEMiC8
BCcFgwyEfP5MdSMX4fh93C0tzEkC5ueEgW5qohjngcDFGGPNqJWk9LMXtb5/eNncDqim85tDmqzv
kCXPsHN3NnONRlaXvroIyJP0FzK26gMSumZAbCPLgfoZA5QwaYD8ewBDSGKhTl3avkdOEyacIUHF
e61qphgNwAjwbO1JxR8gYVp2XmTNhATWH1ZVFr0yQ0VH9GNvk+kfTk2JcIJWmTV36CaojUqxYIOg
xc0yA+KFNvuo4kS8AmO+iXyZgoCS6J4u24gNAU0cduF9lYE+SmEp9gkWMWo14GL7Iwe9vVRBMyIb
dZPpIdo8OaTrEea8+8/ULLkR5niBj/mJP5rcy/T2mgEGVpHddP4ALX4F/9oSX6bqTFpBsIdejkz2
ljORXlkqT033eZIS04zL1qYAIXG7ux3J+9LBmIi6E3nFUC4wzwjjNV+zkQf3/FYaLX7aEsxpbsXL
10pjqx1LP1tgQ0ZLMWOZmYo+TKCweLIjyR4op5Nurk4fEPlfhLaB6Wseau8aHFjY1SUPVWlOTouN
mzayITqmVgbqQAF8v5OUnwmRYFXrIvvpSCSgkjhHmkvPwbRhpEqnRBUYaynsOQRvYPZ9IYxqsFsB
qigJsxcvs2tjLJZngkfMEbT58x/2OyfNOPIVsxPX04c2zOXslsyM83iZ37K/C6xQzlnlXrU/qNMj
E6BEpB5V4LeiVlsUJJoMr9ZwkCGDMxZeEbK3C0wXKcIT0dRK/zrIq/v3BpxPGGuThmam/n+NsdZJ
PQFnZGSVCusk9g00OUMRJcACy87sc9cdEhOjQIMi47IUk/GuFjGMEUztMzllFOKSCdCHipo2agvd
+KAse8PHZv8FZbDVxebVoiwHaUku6YR0UzVDcanpAJrPb2QP+q0IaQWsNa1C4ypbWugajguaJSuJ
l0KVzbrQShIXiiKTav2Da8fjKK/6tNaoF+eBy8UtRaoV/KfI3GiEVyA6e1o8klxPoXILiVuj3LCI
4z/BiV4XOH53AUntS0oUdElzduKeXVfIh03MaYVORTYihtWVM+vzkaK/viUMOUBz7zOUcmWiZ/jg
XpmqXeR7o79M65ZE8T9qDlNWHLQS4tlvPEN+b5g9rs6FkC1yBczj4+lGhwv5k4MHWjqP/8z6LByp
7ISCWhuZoqBm32/oW5KDOcLEx6qE8oY5AhFRqCV68pFoLldajIv7EM4zolfzBA+wvavqs2i54YUM
NHl8Oyc49MOf1CB6ZT2xZa9c2hdflkI6xTS7OJeLbn01TP3HYX9ZIu+2ZDboj/S0IzIdD4CdOhVU
qlzHi27SRMDl6tVJSV92uYyV9PdzvXh6Cfd+OPmD7MdQVHmS57BQvShwRcRHtd4d+V2lLpSJUWeF
xNzsSmCfzvkwxhTM2wPdZAGOhfL9b/+YHVB/iGo/J4OxEr1Wx4pdK8AUF4SVP4Ie2O1GWLaSITKI
hWnPVhn5bfmojJ/ARkfYWmKhT2bm0kN9nJ/oSfNV7MjZhwJ67Gp3F3w4sgDOflYogexmsWkmkwzF
E1S45kxqIksYSzwJI6D7kGu0czgrPpiZAzaO0A7A2TL9gyQIaTTut+D9EPdaPlsIg0ZCoVThEVRH
KLueQsXKGiRI8piz0HNoCqFKktooxDNmkqgtytpzZ4Lx90MOAp73nmoLNUz/kisHu2lZIpqyspdi
1o1OAX9zrNpcC3Ll/nWjGpbBW0GyqDT9pwoaHvGkBCvLSiWooQQP8ttAHEDaDBhyZioquCSF8jvy
aJk1ItfFziWYewCKpLPan5fAgfHQtkjIBRcF+M2yaTvkuuhBcVJ+OArE9McIFYlb/SPx050I8LYy
lE2hThD/0D7KqVAOdZ4CtxSGnLvRdDSCBxr5WfoTrevdJNiRPvc8idg0yWuCLPVL6vjTfw/aQUMe
gmu5l8rXMNqiPedQoQIMTngRMoHyIYWFn++bT6sTF1s6P8s9rgxmmFcEprCWw4uwJ+AMb+Qtjm1E
wlJRsyDYLuvDk9XK4sltseILnos1u4r2G2u5saDOCIOIVF5okWAYObJ3+Sjhnd0cppcdOLaQgvak
2T7Ge/X0kBEvlMxTD01yc9AjpF38Ji06TKfkwgZGSqde4byFFzoim3m879MksD1S537TZURKBycA
efVVoFPL5hBLxDqVHikhzp+ySFJoMLpt9kuS61R+CLdRdAyGP66TXqZjWs3y/XkCdCLFrvInoWGE
SFn0DcnDybJLAZ7GRdhDzOj4dB6wOacPSxTYZACi4qTrD/S0l+zZgE9lO2z9baJpp8aR/5DhIFLC
AjrDrO1GcOtUF2NlInd2wA7XIMsR4+j7BstHSRNe+yxy+KsuSsZ0SmJWEU1aOkKxSJN+oum1xztq
EYTH2iDJKjjwbwGJ2TevxRhOWdYAQZjH9cn/mzE/7Gj26QNgoiYVRqmsDntTMQDkeTux4ISdCiPd
a7XydPQ73S6V1AS3D+ja2P/PrfKAStkLUyzhLGLfRggBK58QQe0dOrwJvwcTt8/F2uxdrPUglHB0
1DDLXShobDMoyEXNIiegBK3hxEbph5+h+uKqOVkbGXn/c0Q7KPEZKEi1AiecGWHZy3QHtpuk2MlQ
V1iEVXpM/NFaliICw/sJ7QFla3p/YIDHKySlm3zIfgHRR+zkW3WMuIXd6ifXv6QBZc9NE3P5HIZa
lQcE8TiuuHQSQXO8CnBcHjoUCRRZJnVjdcxK7atzH8qVuOVVnPfoq6VUWrGXeFbgPHHgZuNP54uT
gzJI5jgnbClpF7KOXjCfqpnqSwc5aR6VIUEzmofdRSZz2oQi2WcyMtIu52b6kaAr2oJDbBiVITrB
VApcS/NrlFIzkplQhz/XbCSdoJK7hMq3JXPSHd9p3jibhNIx9x9/WR2f5IqrhCbFlweu1ba+A76L
B2qXq4arvncGA7zrvZs9p6R2y6O0oJ8CJNP9KaYKHlmZGng6K4z639o9DWO52fKPu+xALxoPgkuF
ScURN6/ukC3mw64/GhXG0MskxSH2L4d9qVPr3k2BsZZYfW6AiihYYopYtQMprHMesDsWajPGoptA
8maX6q4fu91uWyFAJ4usl33flYcrLgtynzT51BFQdJ6vojotX9yAUNGc3WzZQltUUAEQMEMyQzeM
jLKXgkIRqf001nzEhlOXwOPqg9ocPwsJ5ICbh0Qt2Siv7VK53OY5YA/cqfexo8G4FtvB1cfOo0Ts
dqaTwZvnPc4pLtlRS2fcqRIUvXunMm/LKWTbgaihlJ4eJeta/dxuRnXPVbI1wh5qr6TD3dDajvH1
JDaZc+UFHS1ZU5X0MjF8goxUCHMb1UBfXp7Zo+StV9wczM1IdtBm+l4o8JYAhExEWnL5GJveVupF
va5udoFsWaYcX+A9RRP/PpFIC+nczfD6DDku5t//19nGiLNDO5R/WXlbU0K2Q7c5+VuK4Dwo1rT6
FU8tcyE44zzeOnnYy1Q3rMbwsRKzm4oI4UEWDV/N+ooL7rgWzJwhdZG1tjgcDbapmARaD3fHP8TD
X+Q9TUDqU5eh4S3fAbNl1xW/Deu/n3F/nDFeDDMiS+DTjwkFkSC3wpXw3qca0eRus9rRgwxp8IWH
zBPLH+jKL2qK/kNWZq9RqVEtFt/d8Tf76rGsi0tYBtfeerb62psgVfl7R8tF0HGjJW9mxx9RC6F/
cp3XRNNgzs12lFZSKAO8sNO2RtTy+s+VlMHirAr9ZqA8bfR+HqYXXvhdyEh2il8IEY5ASRD8Y+FU
1z3gpYMvLEr+ssVbClbpf1kBxmwyOHFFLlKNhxhWkqMkFqTdx7r+FkqPYKQy8gQOL5a+aA43+WQd
MElcWyXSm7Sl5mwntVy7Lt7Igjcpodskjg8gOPZ+WoeZthAE8EzYThCY+5EvEdCAKTWdZgyuYOIp
0rGjHZVTMX/5+oCb6s1xCwxA8KRC0yRrv0rhSafZusoZGZGe20wcbbPc4bbgumjjuzyHzqiwk2bo
hVWrZvE5NRwYDeIgH1WuwEt9vRUHhXQO/rpAndxvpTCQRL2l6eMXzXY8uiEokfV8amu0gepigHnF
e88NL02LeXPUP+RQqkE1e/o0mnHPWSniUrT50sNvXPEq7zSWx0DmybKnEauBcVhW3rh0fXv/9V+p
XNQSOdnxAxAZe1PZhwcEZZZT7HFmqAn012dz+I6DfaKw/Swm72lQE3Yp3hJFFL1oP09tRrmyQWP6
hV/MeFs0OuI1hIbgAv+JX0FIj6z3VfnNVYwsAaTa8KThpCefbFCLFa3akkbPUT20YZRnB76F5c4h
9lvOD4EQcmmVuqV5U6++MbF+yWIbzWX2GIPVYoTGBt6RSNsIh3jMEoYOANx3mwftnA4uuwwYtIdR
g0UGotmyQeYiQhHcdXVugk99oqDTAAro0FUI29odGuzc69hnnvoe8rVFKHHS5TD6YHcSKPbymTM8
MFoKtGyLVf8qfRVk4jrDSPaNqVMJpQYAJEdyiNo07BWCAUv4VH7z57H3hpYtu0t2Awu0MMYWoNqc
XFj2D0gb5VmoOQhSnddk2QkhMKkPOhStTvplLchf07NrV3LsrA9ZLnNPgpeSkLXIC8VrcHQdypM5
JpUBCl6aCcln2LBz78Esa/hW3Hllkq/FLLkBmYM0dVwPGaGE4dy3Mdju6yODYnJk2O0vll0q1//l
8vsF6k9k8J2FGrFruXa9kbHUS8TZ3SX8gWngb55sI04duTsJ0BnJzTJh6Bi5MdtS+cVIJG06bd1w
ztY34z36lgxC0VVgtDOtTvgSUYAmC9huS/uyGOY6sEQsSAu66Y2xLglWp+hIZ8KRmE8LSTLL+av+
o88eloK/R6KzcRAeCzOL5H0RQ0PWyA5QOECb+eFVJ/gvAQa5j7/aj+U0gwjTFe4p3g3Gcrz4VJEx
oVgrg0+QSz+lz9udqb85JOUKv4/5SQfmLU2EdvyaAQAFXuzWXdoWnUWlGNKLv0pZAhbLuHJUROB3
ljWmlZdjGBBiYWm0paHkp1+A/S5wBjoUuZRll3SVd7wKtJMylXTzky+M9Hrqq49L37++3h9f9Ppe
Rl27Pz+CjCKDlWs0SI1043uZQbY6bHB4LxB7FYTC5BIcNBprlWQD1S37XOmZh9bpD1lkCmHitB7O
CjxH7yaNyQIJqiXjxI7txc1Tt2Nj5zIa6KHLXmZfqyxmMosq2BYaGExWgshic8DPtpgwLIhP2Luj
tp3HGPvH+qlLmbRopEEiX8PLFeJYn45mulEbrx0taVB+a0Q6B/YW6EfD3GBNpDGrQKW6xztALfQq
gqGlm8qgCns+2as73pF8at/qp5RVn9gi1jNh+c5ZQ9xwduJM0ZjqbBQCeQfrHfzkJ0+RzI+HM7rG
09jSPX03G/7lexfqIZjuIZNb8Dygn21qrV3ACLGgMpo+/ZPfkQl4rQ66yj4rOyxEymROnd+mCABj
HlBUcSqNCgx7ITeyev0FHxCBFaiRvoxtwWoukj1kV+E5mdyFbtDV/fNH4mrNqdVCC5MSXttGFG47
DUCJWb3XuUwI07h24+AukP/8WoB01KPISVN1MKvQuqo+Few9IEEcQzgZEQiZgQ91HOa7OdOGwK0+
e+fhYCgsFUW/jOGZamatXNqk1qHKLftrdgt7mkqkdlrjoj0Fu9TZD/OzHLE0VgYa4gWL449j2nf/
mjp7dmsYs9D/qul1xwsJtgKMaqHWqrNp12Tly0w+X13EXSerDVa+Pf2miYFt6OaNI+Mm4QyKhk0c
/iNcutpRn3t2HPgbY0f7GTgbHlPRwhfXRMhMZEF+9oWukPkveXm7/NV3toKdq5oC6P3YCAef2n32
j9NBRblo7JVuw2YBqcma0MpQoT0z3B7isVP2iCtbiZbAD8Qj01k2f4J8vJXoEcTmSpfALl/WYnuj
6l/+DjY+fQ7C1dC0wv2r/Elt7nW06INgETeMESmn5aujtVUU05/Vz15iMQZbxjgvXUlHbkgtDCCN
JUMVVMG/lFCHrBkbZwWoLrItd6dwsqUXvrPwd8z7zl0noUbb7rgrxCO1D4dd9b2uD0l0w1JJpy6S
kX9qv9RtnOcbWgp9bL4IbbGUxZAz8qmO44hJzRz0V+q4OyCqvp3E3HFwjdeEgXRnni7EioBQNKvp
bb8qMTW+IchCQ+km8CFUfZx1kcd6+HD3Fst5MhD1z/RTZsPm/w3hSh2Sxc5GaGKCoW+mVUajaY+I
iIm6mbZnvz997gxfn6Mx0RwA5ItT+U+Zs3hafr8fHEy7r3ZZrls3qX+2R/Whv8UO908BZ0dKVT5G
H3IGWHXUudTxTY/9DMkvFdts351gYDbeL5KVXYZCFA0Cd0jRQ1nQP3qz7b/sgywnglXXFtsf/5K0
ojiAOHTQpen4IqUHvplb4pb7wX04Jkm0YpQ+lKr6nWjex1EBUvqWU1Sqa2nUQfONVlgdOsCgA5ZY
VDME+ECt8os8eUlQ6YwgvQjmOVkpoxpnxKBCzB+61WETaWi7EAq5KSArdsbE7fgr/bVzDkgqOAC5
uD2LTCtM4rPIFsusf69ot4VOP8I25minwWv72qGKb01I7VHttAOb8Fuvwaa4BKZv2xO/lbeGZFNM
5zfs4suGr/c1omU2wwUeGl/tNTsbLUyrHfvRRCZ2hqm52iWR8M5wsZuvvce7YFEMG6282s6je6Ij
4B/p2ZIb6tgSay2RoH9sMdHJ5Ok6vQopSdMhsu/ihLN6yQqXOA52IbaIjyMrqskEsa0gDZjxr9qZ
xaJESp3eOtWEc5fysyRgt1DSw/NwWXI31xydLTKVEJ9gR+p4WdDkFTXc9pIb7VUAF0VGPEJetiX2
AamZzL4qy7thHAlxISKfALowHmV4qzXToFh/dBd4vYInMx8/jivLHExcf7dB4NAgcPX9XMksMpGT
+lbXuX8XK3jSdYz0Af2SdzMV9Uf/1RVvogMbSUIQYIc/dfV8jNs4YLx0ZpX85jPA+JkA8m2mmCp9
7hmdCrhQeBictS/OfroAUsnQe9r8TYX4766LHZxQtsFji2rx/4qqecd7ehCUHAivezeWpEJIdv0K
xPIn1JaGB3STlcNUNHvDotsMtGEO15DIXTZMiageS5gt41q68qdE7e4r2K1VUcQJEW1oSs6tsO8y
zEWxkXd/CKNa0RwfCyhmm4dnixxDF5ZVT0PKkowNKVIPnd14EDkR5151eOQ548QOBkOP7/+oeB5L
cUjj6rll3aHuWyz6Fy4g5mTnE6T7K6Jt6dlslHQopB0dX6oEagxhU7W9+ZiNs+sf2YYQMWBisDZ+
X5qERNVUmesPMrAsdcgcn/XdgH1A3VbV7z5ZiIsa3W1Na7LU/ITH8zKC8tj4+awgn1LIyCNKYheX
3umTBw02+kvSdf3gnp7+R0d2aUA+jZRNPIpsDdfFcYhx62Mc9dQjngAbakAFkoMzscTqOsqNF3W5
GDqGmAUyVlt4hOknQyiJjivCHKfe8bwMOBKyIW9HXa2zdiCbgu9uE2F8S+CsvGm9fKjq68Z2Ik37
zXU0J/lhxC+osgVI9aTwvpsLWd8OlpeMRNNvu9u0vgmBsDuZqVu0EFSCnmlHGgnRke+iiFh9Xd3c
0sFVOtJEA4BlpOs5GL58uiFd5we5QFo19n2/GFK5SuzdVnPI42lYSqPB4zrzSjDu5UeqfcksblN/
U21B2PMYZvdZGmHpK+hj/+L7Bzfty50caKfSfqjtHCWX+Lf+ao9m7KcS8HimLMIj6w4Q2/D+HYFx
DTKHDjZoQZxULqJosRMgximlAJMAs+o9Z9As8LApnS+j0TyA0R9xIujk0wMmkmotYSaVgmPWK+MR
692B4oyHtMrW3isKZD6E3TEVcRkLrnVny7O8fBPv/xSgL3gvOj/3AUwrR2w6QAyVymd/BJfHjuZA
+pF2QKPHr18QvrxWoBoCSoSCGu5hOm4Hshiis12W2kMgEr0H2YrWAxXHwM/Y3CN36Ux1ZHCd9LXc
DZGXF3kP4Q6TCzWJuC3kK9WLeVW/1zJ/ZaEKEGr+7pllLsLZ9ooDypMnn8e22iTdckuCK9U45oem
fvLWXq8OsG+EiyoQjZ3MRTc6QafTJ8eMnrfpboO3Gv5+0eRymluCIOXqPt3I5DOlobyVCxDdFeqq
ywqSdaYQFTTc8O7QSLqH7vpvXlv2/O7KsxwbnGYy+ayeP6KRGyEITDj5ySw1dV0PlanVWhFI6BNX
F67SD1mdiQqt6WiYECoipP6Z76bbRW56sBBV+gO7YS7fIa3RBDgw1ZI4267I4Nc/huWiWCmyCb2r
55sghV4144xx3hu0AmMwCAYzefg6hpZLwj4oFKyfcgDfMl/RPcUaxgSfLt4srjy6v87h21Gu9gAF
MEuIFY37dKffdU/+jLaqBOdXURmYT3YT/YDxmjFY3Tr1nejHRJBkAl0Bze1aUedllIn8y6znK+ZQ
EDuRD3Rxb7UdHYX0rYabOb51UwWo2oeMGZF4M0Mik2dazcuDJDK7QiY5iEhn27G2Z9izZ2iPmbSr
zdJFwFyE+5tycvVxJNlWf80fZII72MLVlW8dcDhMOzruo2giBQ3bx0TXRphufS9jrNfZgWpgZE3i
xPXOwJ3yVtIqYKhrma5X4gxlibGWbI+mU+lB5tJvsVWla5VP2gy5mx5V9FcMmUdgEtdpI54pUF9g
XsRWSum90U1U6AJpTP0T4xAZqEnPM+aRKM4VyvtVEsn5+Lbih9b/SkK3cWLFbphyEh7XEH3L6jfI
q8FtdxLOiB96F+Fpwri7w+Sx4L0KvTptXaf/OOl7wC9JoYSjwWsjvYqPmh0wYnBiIx8R6xTqkDu6
hNSMcdyGFco5Kkr12Hpu2t9WdtdFt0hgEE+dVWStgoxmduASp79PflklvSyEE7MUXvGySMUlNEVX
NbU0eSdkbOg7Xcv6lhcSIFt/pWnrN+29bQKFWs+qunyA1A7tNaPxZZFdlqN0HreguVTjvDgetMr4
1AGd1aHJ28Rw6iyUNzJ8EVXWiSYyS+04TUkeRwjuOKhtEJvv9m58u4ffV+rPbY0/nB0DLtACAO5U
ydWWeM0Xq5lL//P0QXn7cv7Yc7RNS9anJ35sm/LoM2yFSztpjhDzg7dSu50EYKRwNQOLk2PfzQPe
a73IYGz6CJskSuZuvoIO4x7iZQ9tsR5h9/iv0hdHbUY7kq4FP12iiqtBeg6XtVwfIeHhSQN78Dpt
IDFLC+EOntVVyMoD+yYDXsr5zXYPbeMJh49J8se5tNgqSQAe3P7IcskPLPNoNbwPhIrO/zTyxwU7
KvPDplxWYgl/8XQsfn5zl7NxV8L+Lzbp5e3qxYemf3Srb24QFQCTZChlN1UoWLUzrC3TGGUIzFDI
/LImL8jy4R1dogQRwSo2aI0uS7/I35XVucdY2SOq5dFlGlNI+CbJP5ZtdZuPyoUxg6OhuzELDcWi
zrb4NfZlqvK/9w8rPJ+00pUmCxetoqNI7tv92dEMs+xv+ARIugsKcj2l81Y2Xuh377RfRGq4zkPv
AcDfmE6appBA7pIMjS+qQfcNv77GG64zXFTIixzcSPoNq0vZCY27zOzE/nVZfbRNeNtLyYwey58L
KRgcy/XdD0r1UyPxTzgy2Ad+uW/n9ueCVspK906IQnOGYubI6r7biLRa8Vy6zAaB2tlG0lvKPFhm
oBoTcCh12lgPyy2drE2WspIVD914bHNqeIldPb7TCBJbIxFUHctyphAcABQgfB9GB0xygmvUrNRJ
qkZjPNPqHFo5Jh11slXbU0WxLhhyKCKHeKMgdQoHGtzyoWQYvpdEH97mjlaFKj9CHwyGjZRKfAxm
gz7mAzz/bCS4ch6CsnVBHseHvqomxM0q7a+8CKGfQHfw/c1LCFSC7M+DPGnnnQiKWHSdccvUyZo+
MH8jJQPD85LQ4HiwoHjgWL0frk2RWDkWNBJtgYyEAOuHGc+7iqXVAy2nhoS/WeKy0VGb1lU4KscS
MJ49IEBjmdss4YODfOgq3ZHL2hUTP+3oTw/BF/ToyLfU93com6KaBE0d54lAPLrq9N5gP1yb5g+4
o8vcW9ThC3C9wvyDY/m9kQ4d3buN6BGgc0biLoXZmPwm9ky9mIKppOD223UbjCbtDH/pVIWsoW9r
Hc/Ph3VOb2xVbqxqhzZn4Aa01DoSMePwQSqQX46oKGzQ8u7O2ksv6XjMfBKGWaJ1rSNWH8TeCObn
IEX4BM+nELfYA8djXyT6E3pdEzxQkUDzRdI6N3O56d8FjU2dnTDw6KUONR1Weaog2ayURmB6lRWO
ZEM9V7wkxy8wSmsr6DdrxADX9+oul8pze6zq+9rab2gMbJjBUWjA92bg/+mm4sZAcnb2G1VWiKMs
2u3RGBq1kE1R93iH0OgZwfJuBbE7IxhJGY20WMHlOzhs3uuEjxiraGTPfyZf+uy0cfvGuNnenrvF
0C0ADxzXehaOwoHnt4soC5cEB9nsy1S22E9w69ueZ42oW/dYCwfgFCemhMPCTEJiUD2DUp0tSXB9
SYtGKoLnCKitvXzr2hEZjluBuYUq3kYpTkQcP1DOyM5g0DqKfXGxqKQhPxYnlBM7xS3CdfW7dLPG
m2eA1ZU0ytFtaaYggpB33V8MUG89Yd0Gz9qzErpukDoEeawPwtRWR/FOlMtCtaoHjzYj6WddM5bA
4O9KbZRnVQfTvnRWF3X9SFqQ96UkTK3a5W2JdbrGTmcNGZYjHbnDKjZGF+CxUKKluGFBdZNmLFyl
WXUkzqz+68euGT6fqBPNoSTozXYwkvvruju3ubyIgZee133HqZWyYcvl6GbIJP/wSgPIBJVSfkQ8
zXhdx/HfU7tyVQBlH3WscN06SvSjk5spFQb5IVP2gBKeEsXsZhLHnG0dvmRKdU4y7chp4zibukp+
9l5F83ecL2b/RY7TJloE5DbtPIvPMngWNONdrYB4jXv5ayfKHKrOCbVT2kBcLtltVUVCCTUon9/6
5Jmofaf9IUXMMTL5YOQP3Xbjop6c7Whv+S3cm2qLX/PIuWiHQHG9y7ZFziBQIoeUW6HkmUKSH3rf
GZhAW3UVEZObsNLjxrim/8oa4zVsa7qrwDQajZupEsj7a9q+rnP+gvzOxUa3fGY/OOLCqxB9TQyN
qO0MSzi7bSygJHpiCOtzPnSRnkL/8BmCEe/JD89JoICkzBnskMKHurW8luwo6fE2KerW2yaAGW8L
B9ls2yaqh+rMR3sd+sQPB4Wr1SrOmYc1dCOYBgrAQOpF18gpQtXLBhD8cnlWOfr1sWhZasIDmN8K
CHD3eImQXPBJPZbDn3i9HlRBeXLomREAsLlJilEg0bKV33ljWzLBA4sdNQ7DX2i8UYyxaJ/QiBPB
N2utXhfOtqMe+D1LuN9PTPptX0XFVnx+s4karewQKtrD0mdmmOVoAD8vWW4oEsAYtDHxXIuq1Jti
8eo+/MnuMoZMN2M7vsW3+c5sa7t+s9F2wwu6x+vbNQ0A75fyQ67iQEByhWulNkDG+ocqp2wQbWwj
Oquq3AAV7NSuvEk2D5gpvVMpPLIkN29BAlCKsibr3HlB8XUs/TYaaDpoCpD6LPTO87kxv/C7IhHD
N55OBOi6cHveD63GZGNEKgtG2rJCoYxaqJRdkiUiPhs5W5krQXZgzI5kfNbbUh/odoR8BxJ6EfYd
1Di1gFXgmQm7lSc4PLOZftJw62rxYkUCvtIuhNzWF5auy0+/4iXYR+5CG1GlH4bHbZlY+T6NUvVB
Q3qSipaAVaUPMgH5nUjRJP1YZcNW6rXGCeJ7YBJ/NiP8JLk1/sXdd/OlZRPysHkhiubX4jtGF55f
TK/fkNdG25iEkqjxGRV8xGO5jOluWook4cew8Q4ZdGqJKwBN8Cc2UPm3sPjnyfOlFoojjmW7Wf1g
HQh5FWFxf7k9F5QKEIFDMX8S/4+qcWLkYr8WLBYde4ZWeLJ4774bsazK6nivAWeK9aJTTqypK9Ps
cyv15ICs1oaZSM5oc6KX6Zh35eXcTwxo+8F9uHiV3RdbBphNM2a2v6cqf7yCGGHtISuJUZ5YT/uJ
UHp0ILZ8gE+YQBlRcyox4fg+VitZsRwOH631y2Wd0j7hZePI/IkyStTjnfcfOf/8ujsN/IqOqTqE
qCbqlOY6OXxXm/U2OCQXyey3az5TEFOl1l7oScIDjbQRIidVcfJg6C6FiJmjK94O2YIu7ij9hNB1
AkpYE0HLMeeM4PHuQjJ9Sohv+kNVEHKDd49MPHHKyhGk+Chv2HMEdWky2DoIttJVCauk3a7KPlFi
twT3M0cO2y7y2vv9tF4GDx1eDIpi7nEzFLVZS29F21CyV6dVz9pWf88INyu6tnh4yTUBsVtlDk5v
BNu15F0oJdDt0wnAcmalpKiUKjqc5eSjMmJivM7yyD6bXI1olAY4HSd3DOcpjxO3oVtp8ikNIjBG
yFb11VAbNQoGu61W0YHQNk77A+4Y54X6bUleIJK5QQtgBv2x5bzX1XBoxoMWv4flvu4QZXooz2b2
WTxDrFTO86Af0vwPPG7hBE4wgLhaoUxoHNEbgOgYxKWXoN08bE8rFIUGcF/y2YEVzDm4ptzP6XQ8
qW9LxgW0vrw1cAsDWnigDFtanw8AbdbOPfQYIyZfNeCNKZ7cbOis41mZAB8J8xNoo39AhPtyk9XQ
jaF6UC9QbQiQT1NetTTqONdWUrlrdMHT+iAFTCNGYGn+xEKMDkAnMm9gtnZpSICF3/ePzsOFAF75
lDoBgW8z8xfNqYG7J4ubO8nEeIgNGFAC8hsjUmn6wIblFF80Xl8dF4fEAOKXysPS+o1MWKE8mvzV
LOSKvkF2g5K3jXUAFImo4STUS/+dgolO3X/lc6yG25IcfJWvvEgE0qbi1FATbKCM/gxYDVomcxuk
UvvPlsQFcxpz59k/tHQFLvdNKqoVmoEqc8toLXivn0lSi3tHUOOjmR/2MJFH2SLOPviz/OHet9CT
T1qEUzGGuchITYvk7hAEY+pkd28A2TshuyFD3VjhqqyadSgzixnFBVhtW71RKW9BNp3bB5ku7gE9
NsEr3uRKRX7XsCrSr1L4BPib6qb6NApe5QwMsPJSp2s0ofMwFJjqiobNNtdc6y1gMZ8uMmfT0i2u
6yqMGmbGIRxw6RCQOreMQ/sACvnMS+Ls0c+btA5m7zQE7UpIb8iDsqx/g1JpMpW7P9czt6kT7Xnu
mo+Ebm3jzPGiGqHowlifGjxHxcFVNZfJvPFvJYTVWWZokWV6m7dVBkOoXGVGIwR8oAXec4Tcm0wq
NPdzKqNflv+bySyOGGUDZhE8Z1IY7IJUw2X/tLRras+jzRQHBT1scJAQwmLLZGQlTpJzLuGQTJ4l
jPfG71EmlOgiI3F+sHqjwxMjQJUwsYEMWfNZKC+xhkDngylmaUGD68pcx97Ee0Fg7CofmlbMuXak
s3cY0g7+Qc0m7oCnW1idtIDTumaaf/MXb6yMe1V6AVr17RbMU4ThygDfoe9tzhqPjhOjLVuSdTnY
pg0qjeD0/1ZOWjy56dCdaJn8Rpi4bzN3EL2PPBjmCBRPAWhl/Wpa9wSJw53Zl5AQITAQiCKlioBQ
EU+67sJuyyevoGJFN0gnillpZZFUXTkMb4jJd6kl13hSwh+9sQIHOxd9rYUuPl16YCDfdJa8tasa
9C4j46kAbJBtQcPt1cPjT2mSAWysdhAw/HUQ8WIRlnKliOi5EVUYKg5vnOuTE4ctrdG8GKZGgzhf
Ejdaua/k1n76HQoZUY1wE8mL3HB8LwTEn2NDZc4L5n1fBaQhZnz5YxIHM35e+I5uxsaAKcSRse0y
58ZpH9PWOPLWDgRpk8t9ugG5ycJ7Nub3Zdj93tmjYXYZ5QDElaO+bvbKZqrhMLBElml9rt4IPf5v
e+EZlUnCJtCUuY4wZmzijfOrWsxayoi8/4zNSaxVRkmm2gkJ3kjl34XZdttw7X20tw2iOBZjm6Pp
NqreB/XS7ih0wVFIh4BRjnN8c52blGXqGuwJiZNJdi8fihL7Z53oR34JpTPUAVCjmQ1tKwk7pIds
K0f6TY24yBeFsnnMd9VfWdHabv0C4pKxS6dMytvcnbnlRSdFUWog0GVVVZx6+1m01yvvP3MUbshA
Se/srVG3+evSf1/hSx6yB0OGq2A1iMMeT2OmgGpKKZ6hpf8lSb/0iwh83EVWhnXgiUofVS8UWWSq
QkwAX9ubSMzB5DLlVgmspNNhfzY6IDiLtaYmC48ZFiKDsL21C2ykpNM9Xts3tMVdZcZ00k2wAn6I
47qHLjWaXdERAK0oMUgW6DI3r8L/o+p5sDQpJ9FqKcSgFO7F9tGU+Xq91vMp9DvMRnce7Zp7mzYQ
tv04f5y5543rcuFvj/apVFly+aICORVDRMGTm7ocguGwQVr/qpQNHgokl4xFeUxS1c1ITyqeDtfo
aRT41y6ckDnHZev0f39Q58xMI+P6Hisqo02BUykrEFivryR0+ooha7NLR+6cyMsLX1tafjksTei5
UqkbbYPnNvYNba/OeTA46/9ThWNBZFc2CwIEartmnCEYXjM9ZvlbfmoHgUdTE/BtxR3eR7vjmJUq
I9K/X/HjwdaIjFfYfCAaQjBIg+xVeecumx4jeJ0FKh04EtukM63PQS9XsBsxWUoLV3y8z6CJ0z09
Y5/NpWkKkWN0c9euTWfVXHrlbCB9iZeeL5ktNuKmOYT2mto2aNTE56tWUdf75FBwTaLVJQPAbNO2
Fl8uTSNRd515/mX5201dYl0iNDaVJN9vS7Q9Uwc8YsdZK1g8UIh0O+hZaPNnlCZCirK9QGUnbGjY
p5aSHS5zRrseZBCd7SRjtFa6fdQ5BPKY5ye8Fk7C3TF5J/+yxpgTujyZlc6rSQcg1cppa/ZmP6xj
4ZuuWc0AqFSSUdBvDoSCXHA6nmdebE/V4Ym2P4rson8rwpc3VF0ZKLPc+QFjcHUONtYTF4TXpz/C
67p1FZEKN770CdGpypHX+VZ1lpWeRowJCJWuyXi/hrbceRJCtrF0sTSWBRfLPSupG7QATv1O5tkW
ga9IRJyrzY59nXh6TAVFUgCxGcCW+ym1hMPdR4zPJcdT1a7nZlsErDXk00vvSazcHMK6XOZRgFoc
5vbDwSXMwSkiTp6YC4hCKIEDipTxUeSsDOoO7fhYSLPH73q1W0W9fJT0+HaDY/wR3zWR7jh733un
nvLg6LkuwZz3vFUAMO9D8TFrvOz77bevmiwCX+W9WvlZ9Gzkil2BdBJkSQFtxgbu+TluuVJ/7puF
0GTfPXO5aN3Bz5Yslq4WQLpzt+Lbt/pA7PIpw/Ji8wzbIp5UW2N/1baBH1wSYdl3fISx7sQsgtVv
Wdmu7gjfm0XhnFjxrapG1Qa4oZWZbrxSyyz4neE/gT/am8bz83bU57ZOP70hYRX+JP/cVTy4R3JA
lAu5YiysJYBTsgzcmsw1PlANo8hC6UA/9ZkNogfJIMj/wsWo0tRtBXt4SKNNhHg4KBtf8pc6ipv+
joI2/NVY2fQMLlFXKcgXC3coq7ERDsmbtxVM9D4y+D19HGqptfaE5sU0wKGiP5svlX61CM5ktVaw
PAbtir/XxNEKRXMcvWtgOVmYnqW9yKDrh8q2rpXnstDi6PfEiJa6GZcNZ/K+ejDcadHdsyeDha2z
b0kdAx83Omtw/pQ985X1ylViuwep/vNLfJd98Cj4+xTzqveLqMkV764KaFqpeA6w7YUydzMdm40v
f9RckJqjShKp9BEcq9BtVFlEuWS3ozJ9b/3evI8VJYgZt9XKCl8DvRGfK49RHnimfz3oLPBTiDml
/S0EcNb9CIXpAoibyHxkLP2SLNgmxPGXF36wXkmrfqzTzTgpAbbNOObGAC9akG1KANnFPVOABbWg
aRqh6f9zXGiIlEncfMIwu65lg23ea3bBintJYXZZjIqD+CjK4DL43d/9nks4oslmPX6YOv7Z5HxI
mQ9aLjALJ6qCr+ptIsJcwJnYKRD2elDfObpnuPMdJ9Lh59WpOv6UmOjNyEKJNKVgWxfs4MQcoqti
+roYhU2A/7L7FaIVUMpwrVztYBi165mZbg7chPa1DTUkRx/H+SWlQCIOnudA6dgZhywnjArZqi1u
CRCI0/RvlkcJZXqDsSnWm+/cIxqxNXyxn7//zp0Wnd8ZFG66JhKes2lHgRN4GYcmeuJiKIAcWG+/
osF/+Dk/RAQ6ktwMnzCM3b554g3R9ydKTXsFKOUAXCroAiCRps1WqRygd6NCtTNeiPFvPzYkHFbl
F6G2jtH4Bza6tueFN3SMxQbhNYnkTCETwA7h5T67x6UdzBmoSo9TZNZoKvcj5mg3/f29P4F/WPkn
J1SnH3jXFV4nt9Qv6+08tQpr1ZKVoOLAWP7fU/pz1xPw3ubFUj+lCjPE/9LW3gQdA01QZ/CpyEpa
ctWWRH1F9ZLrz85uvLKEbFXAtRvnUB1tCJzWh/kP8//4WnAmx9eGj+ujN84yuGN98z8SkrcDIBvM
2qzyxUmFaUkgcA6BY6BaoCnzsfn9CVY07z0MuZf5lidB5t50iCz5gLt3ID8L5zN58fzJCBgz15Gn
zzaGMAEow6vm3WkClC6s6OxskOJJHBag8AqKnBNmAF2XeWeU8yfd3RM+I36OTrx4ce/9X3o+6iIK
y+NiXWBmbVhsMfT6BrYZg+D/2x9Un8vYzTNJWQlBjvXbGvwOPDUR6vj/ApedUARXCX9ZS8cCoWln
izledtVePtexHHEuN6YoDE7y7vO5DCbPam2k2NfQQOgPipYcS2D4QW8GjLnNIi0tk2jFI1vLcCW9
rO1NYZiFlGwpBBdO7V/LepjKRqyTOErv3T8IhZqH5eTRVaqbdQAltsXTD0SLTGZZw0YEzTBMbU2/
kBmPF/PSu0BaXvOKtUHiPO1RGAvY9S1xBY7QL/vQJzLrA7d261/so0hcZO6AW231gOVhllr+jHRW
E0GYyB0GW/H8eTm3movVytCra2lBKAA4ufwP8gD+BbDqWLeegKyPnGe9w2TBtXlpju5riQG0mqGw
3+6mZoMyuuzHD3PmYe2G7/llBwcMS0N/8gRFdtTeBIHJ12SHSwMJrOG4qsdaihin2Mz5Qia2KxJx
KP0KlkNjrrdmH4yCIRJ7/2tFKMXv7lPjPD/NoyYfvzQahl0XS5YpvK2R+TX17mO1zwnpigEEWq2c
rQeRrfseuhQVfpyoeRe8yLRNO3RQrgRFPyHM567f1km0BMFZ0yFIK2XGyARLJYazfe0uwW3t9XfQ
MeDbk9VEubxP1gt6/GhmPltreWac50abEqf3BZDNl0fOrgsA5bhB2S5GMCLmld5pt4tn1YFbqYbV
qQGTGWzSUlNa97hQIAgnM5+0NtZaqynGg40xDLPShxgSUdo00RcFGVgaCTBUAx2HJdgRXpB6489x
zD4hVtvx8J16DCos3Xnp8U6TUvtL1IizfdKkQMJuAxccnE+a50lq4aDLzy5Jg5lvRxSE1lx8BMu/
BKUjzV61QDykvuY9Ouf89XABzb1oekdcbfFRjrKPqPJ1w6K+BDRYmyChg1+dq2Ax3DpBohwgvXG6
LxPTYd4Daon1OS6zGG5ptZDiNi56w+eT++S451QdL/KryOlLWMyRRQNONz39EldaUCH3MUfv+7qM
NYv9W4OrOegcmuADoIeG2O9BgiQRV4J77Cbwe9OC7qNcO9xQuMXUtcWFo7IxUoy34Il2pDS0KOcO
koTo15wdu8ChfsEmjVBWKsE35fIADhZDQMSTZ63kOQqLWld3i+tWp094YSCCLEcpKZTqh2iMhJwQ
JTvaagZaPygqzDyVaEh1kq8ZPtkwkPvMHRKqAiSxb8SVEpNB8rZuWDyXKyMgljS4y81kNXS43Ako
N1h5T8c2Bpe1J0jLv4eJAqBT7SPf7qY/K2EVX0t4bixY6vn5UQXH/ITT/x40w8qjSdBgkGi4IYxC
X8JI0UxIrt98eKH63jtgJOyKBwV9hpA+i7da7KKVgeCPNUuBZIfQpTf/qaEXelupgdgsE+4gBBHY
4cMp2pW6VbJoC7fR+meQVCurKUCLB0pPtQ4LoImvf9nVrilAtvrPW6iGdFYLIWGD/bYcLWCK1D7H
jj3ydr3r/7V11WUx1/FXyNOIpE651RFm4/0Ni0tDxsM7jHGIWYDZ5n5p1SETJ6fRNA2j6T7u6lI1
6wddiNKbgakGaBzURowxfXEvoBTfz7QT9FeK/vlF+48EU76tJUbPHyvlfKDO0fxeKh9Y353Ga87E
WA4ZgLT0Bd+vrg5YUtH5XD2tNtMOeZl7g/n+phOrSQpxPcIVtgUhzJyfXq28u4U0lCTFeGk/tbUY
gsXKWQ9aOd3DoFRgmQuaoJ7CS3RncY5e9iccYYbfs1xFoESDukTdBaJBipIbLro3rtWxpopK+NFV
2bvwczOf/lh/wbhIcCF0dkj5jC/OBscq7ai8B0amHQ2ZbSxd1uPgQG/ffIj6Y/hHuVRdbxxdhTBE
FX6wd9uiRVSk8PrUNqg5BENugUZhr15KAHoobCD5Q7tS9dP4mJXZCw7iuYwfSlTxVuGI/HmAiXWy
Cs/WLFzbkuWLDxbNbvJ2VHCpa/nQ7GH9VtbgO4sTHkCYh+wZ2YQq9BebCUrr+zPsil8QA/VLuzI+
Ui5nsnUmAsObPUdHSMwbGfbrCMH2+fyY9zrXg9z3cVrCF70Alctr4t780DPj2LCCkbDNHsR93wsp
5+4zeTk/Y1J/xokXdCOmONxnIIrszozQNylRapYBAmc95KkHrhlCRC9jIkEs1Ll/060cqn2puJfl
m1gSpcevCDBhiYJb+9G8eR2mFRRN/O7XQuIDWE7+BQhDlkW6kTJej/Wcfq2JIua2RaAmrsd0DcXh
eVKvwIuTgaVk894HZldsNg7iY9ee/VVet+CVZiTKj/6NW7qDz7Fzl33TMKf/NnclDAENv2THfEn1
02RXUNeslaZYV4wcp3GxRpVTQEQ4Q6smO3BnJ+zWs55qKdiTkKBU7qxAeFmqcCb4aJOdgENf25oX
eNae9ZsUMo3QEtw0yH6JGoRQerS3k6oEwhZYSxBIPgH5XLt3BxIsaUOw5vnYnUlavUGXrFP83t0z
1Bid4YDZ98dPdXCsuql6fpI1WUNs/M4T+d9kyR3/Xu7KAwj9OvRuQeNMJDHDxFkly2j76Z3XLu+z
JjOOqKl6/bs2sO/gVJcWzj0+gjSSmb+UtxHJbzSe/bVnTbscg4sVNnwbezFu4oszWn8GKqxhvhCx
5BSwqbZwwZnX9Fo64N09j+9dXdwK+DC2ofIt7fxTJLtm4XQgG4uE71GMxcA8RVJh7inuJm67/H5R
7U/8oiOoEwBJe2/rN7jpVvyhIBvxX5yr73w5CFX7DlnrBf/g/sBIMN7F1IJafyH0RHH2c8MQM5lS
8OUTwyVCXXVXx0d3/F9AFnSsbMsUs/hKNT9C83GBtvo/MYTESqg/PTb+cz6Ieox+ue5URznJI/b0
Vp2I805bQzXBJYi/b9gXWj8fkwtAiuJr9o7N8CCuL8YzxjfgG5CoW+Dkn/WXayUGhPAJdVCk03Su
2HUvteddQAmm5z+OiiG01HhiuENFrL9t/z8v1t7EUaRB5S+vM+RpgriozrwYpUD71meBQ8Gzc9aJ
aMkh8UrpnYBgOpbcFXxuwRHxgmj4jrx1qXzx84qnE7t42A8ZkaeMJgbV3T2jJSjFme9o7/C/Pxm0
8m0rPwN6QaLo59iDB8SLhSBI8PeYOQseurMX+EmHZChHe86DXE2Dwrw/D3CE+3ifvAT5Je78uwMX
xVJ+u/4am2nnpFEvZGe0ggiNpGEGPUblxW1TaWLdvodR1gIc1J6MH0rXcR8p/Vg2oQhqaLWGHJkN
gVVWBtcQxu51iEjzpppdrUNJevLKD/Ktiz9IvdFq3kPptJTGTamOJdMmvdqyZQ0tO8GCdH6Rfzmx
VkNud/ulUYOaLYXiWI60EJ+iNiQk/MOGWuZ5g7v+ToDayEO63Q6dlhN+rQHrppji8GlDTd5FUkyW
kXkxHHoFIutNWISZOISDAa3kjqlrucbkDBs+kiG+OEvV+4YxX/SjI4guuXf2DTQ6CqGm6bhj+Dc8
8bHvx97xwi2wGo4BZhvb0I8irNd9lLVc4qiaIUi/59D6yT0dXFHVt/NlSKv8Y3woOhAWIZwrc+wE
7gDodhA+H+A+Yvr8S4hxYKBHJokzsJNDz5aihDOMpypkiM6n6O81UzEUQQA75zBV+26Ljk84qpyD
s+D3j+JOSDWsMoG1QMhB/RrL6wxC0qqb+N5hRQbBZvNZz3RlXRi2LIV12VbQszaItvOBg5G/1ec5
sP8tsXckQDY1IGQ9332GMni4NihyV6E0vhraY4eGdELFWz2aU8UJLwalvkuvQyPJEjNzmkWsd3pw
aGjek4/+XmLSIY86l06T7jrgQv8WgMv9B9cmn2/0CTgShKp8nWo+fFbgiXbpwv0zxBLxBVQaaQ2M
4DP0LXnt+vICfiCx7U76XOZ1ZzZozgq+2RUPf79AyrEguzTC/0FQoFjSKd/Xv929w7Sq9SsISNgA
Ioh5sfEGwMrMOJkw1M3KpNha2gLArX5yBpB/r0IvuA1Dkm/o5YDEjqYElLpnyY+oW4FhITyIWBl7
1SfctVdf1N6V5Lohqu3HibQVfLtkda/mGBek4LC69iQUe9lkRE15/ZUDN6Ojg5iPdOSKfmjKEWKg
OByuBa5GcytYypJbBYglwRuRiGcdvj4nnql80diPCiaqlJilYnJT1F32EBjLQArUfC3axxx/NsSN
VlE58TO1emAA8C+H6HykK3rzV+6jR/q2mPPTyeEnmRd/xhhYb/8MI27d1sdOe9EpyFdkEPQLwx1F
d+E7WWgmg8fw6JsWRPQQlsi4nspEvKs6HpzH3oliA7+KYhDlGF8bK5rMZGottlYWsGC9ya25Cjl7
3oRPh1Vl1hMRHLoQeLPIXDNDyXuHyMnK65XwYeKXYkl7Ji6BYm9KmKhydMSVnDzISqUc//E2irWQ
cpv3IrFNHHD7ORg28FLo/esSOubcpWNIlGPZ5qavfyKvQF4i2PhLbZcXz6fVPCFqSz0L248A27J2
3YJLPJk5iwjs63Fynn4+CAZBLKv8l/7cz9vw9sLV7dgsKxCZelJEVQ22Sq1zyRebkfHdlfZMaqtD
Cq1IolheHQ7BP3ev3HKPZk9RF6ZHuZc8LHTXDdw5u7fqMcYgoDhu2Oq1K5Q+fg3qzeRNWt8/BxHA
67TCAnmmMREjwlgUe13ov3mlh4A23BP6qJEevHWuLvl3nlTWmJiOlXazEUlBypfp/hRJ4cVWrn0M
VVRaZkm3i5efnt86hPnzPyjKf1LfYcpoF/APSQFMHkjDIT5ZVn86rxdreEHNlnPvUn8gheHTQwEu
U7gYYfk1ZR0L8FeGpOEwL8Ble/MVJGdDkbc/au2Fo5XSENy7OSR3+AsKDJ1uftOiQcMtIG/2ekkU
VgiqjPkxZoiHZUxzhmAq1Bim/8xKDe80wethCJXot8v+YtYNMfa3HxwfRuB1BGeSN8kGZO0ZavDd
GGeDe3G2YIx2RlzxZQX62s84xUKfTpP3rSJ432wDsa4APH+EocKLmxoQFAv3o9r8INZEP6RjVa1s
0Ww4XTSu5ZFsxXC3BlquNs7zlGbFCMF+PTy7TUAJBebpSPPvDo9s6WWxam0Xl4wCZvdivd9teQDF
G5jq9szlHl6B48iuUNOwj7N+OIXPcZ801wtkvoQymjW8qj53wZwoEJYhk05Z0+AVEDgyFWiSB9Lr
MCECaErURQ25bpJiPwyW39NZQ8xqsLlVF+1sEhxxht8NoIBEZ29d6FcZsH+WjswqbU9wYLEYMe92
pe93TF2fOHdSp5ffPxfnNSifTTXIwePUHi+vJkmFQwdnf+ZkdAD8o9h4pNi2RkyYVsBhnlr/8Kb2
ZggHlwvopAwXlRyrXoGrAXL/CZnaPTvs9nbx9gfpBKasBdTryZU39Ri0oox2cpLBnQ7q3+vb1vM0
SCjXIFIuJN2u4Tt49GhINRm7WKJqTh6aHaaIA4eo62fafOLAvHezupR4Qkq9NLe9KULSjR8SRkNn
Vd/ThX+D8A6yziukBOTcUZLlaj0syYnoqVakQv87ZSMiiZ6NaGAHySDOtcLuYUl1kXFZ5ZyciGBQ
jICBllEc9VjBtS5Oa4C4yClHaRlsYzlWArX8C+nxFyJwOUsBPVzjI0IexLGkScZhj/L7GjbrBFiD
gxyrbzi90X37yuOgV8d4mz0ih0NdCt3j+hYSPuXs+lKq1lAyNUTdAO2/XxsLftotXKWOM9IMkXzB
gO8EIQN+CdAf+TfTBrRFXy4lSOpnh2bd8Z4s4tlQFmGmthrEGDNNVMAl2JwmAW2tWqXj98aaJvJ9
bUkjTA4SjNZAWSPpIPRVqSOo3qy78phcX5/NTXR2KqIRIlYUrVK7KJKKBa8ctgVQAh/ZNzJYdIfh
/GcQpsLpzPZIosP4yGFpHpGwkQBEkFZiF+b33W0a/iqrM1EFEkyl7HpCZWW96pzVozukAVlQQv2S
/LSW1kvp2DHzpm94qnmI0LWBNs973EQ95gUqSuXrdo07h9KhaQZvNfMJCSRvOJtCn/OdZl6rg7zw
j39YpY5vFseI/pkQ/8NAXSnBXEIewsqnA8IDVXUw4hrsgVngJWw5Si3eibCR2u5cPbR8vJQtBEIZ
QS48Y1S09Nv9PvOFhgnAiz+kV28oz9MuD1jAOYlKO3/WsKXe1c5qVRdfGGAoA9901h4TiFz94vPT
cwMX1CeqQCjma5roCRzN0DR0d+gZtAi376aPuUQ083NfxFFj7VYPKwBYoCiCv6J+ZzlBdtHHIonz
O0/h3BV/OjCuV/qbQeGom2Udm3cjiJdw6qTaDi33Qso8NZqDgKcZ1XFW1naeW8/k8vG5bUoURvTG
/OhaDVVCcNfY+DjkPHb6nAF1InQ1x11fi89WtJW+3Q2APOKdzw2KIdV2EEw01nI9vBbbox1HjH7n
ZvpLav7uXZyU20ZjroqQnULWrxp2Ze3pFfSFlTq2E23PBwTrEpX86OF5dDctYLDx2AS8Y9v221eV
Cv3F3Jmh9ae1qx7TaU6kbHTs5ND4Z+xGRRNXjl3b0wFeUqFatEhNtKGUhD90cKGI6pfem/JnJK+t
V0M1biAq9Fkog+qp7IxZ6CbNA3ctxj/wRBLcpzf6p/SGbFAakKl2uv3zhlTkaWvxBgbHpKiwEGwu
6Dj6J0RkBP1ul4j7FER3fWZTsyL82/752tbmKSdgu3IQYAmhXEi/II70bwbOPuabBknasgLX8GO9
c0BhyLdvLaVbqTjQvWKmdY9SCH0xk4Uqp7ryDzQm8Iy2/w6LQDfuj2FMzISMW/ArVyDjminO+bYN
VuIFakWC52FEPyX5ahC3h7DxtY5mVnJYFLcwSDvin/paCKZMFzZ39JfY4yBmiPusmruMY5wWOgI4
2gJ+LVzFwNpZQZhh/4g7iTpeoB7I+AQX8tvXQd5K4T4/tFkNVEn58O5DB5v5p5JrAdVjPNHJYf73
+6V/YXK9t4z581x42EoPt1lDKW6KZUIqTA3pK7Rx0RSgTYLdlDeunrVGrK6ruQghbOB1fsubiHEm
TFebfE9T8mWprDgskM8CQ8f+/aHl4o0KbpGrLiCR53jXT3t7/t/uEawLMxwaBuWVUrHGB1Bvc/gR
nBTafcYGzC6LO+Pb+PskTi7T8ugqjCZJBMA57tlHU5TVk15YBA64teY8ju7Q3nXmkg3xm3uDxf+U
6HM1ONctxlo0k+56P/yrSlpnh2jvF27s0uDAinzoMwkBhKnccdMQteYI2uBc8Ivjr7czV7Evs6L9
rsJWfJOLJuKjcLgyRxEq6U2/4/Wtf4Q7PJ33YAjcXP1+naIs18jGOSNf3BRjveYnlmNviKZfbeOy
YSQ5AzmQssSNQ2IT5+OsT5XKvNHudog3VxLCGWZJA6bXt0wAAEobMgsWen3W1Z9PudZBlf6trqK5
vp18R6gfl5D6uZ3UmNpN6U8CFgkGcTw/XFPbdXbDYvXjJYWrFuWdA93Lv22Q4rFaCzf/mHN23jSP
Q2o0oUIeFHefua315vtu+RXkdNge+KBtjt/NA3QThYVLT2jIbxd7C4KS2N2bA5mmaJBuwwlyOoTx
J0xNAdtuWw1sqM9jp3TU4fNyTaaR+Wt8mPWNy/DA2td23HS4Rz7BJwgq30YUL4Wz0nUsUd3TYFrS
sTYY2J95kArGhPzOFpBWRZCW5ItDNEgFoKZ/FAj3Nvn12/v//aHX23OlDbCZqqI5xOJOtIs31BdX
ANHFN2cWMKlij4NMk1WSTE6ejfAmP3zG7Z7OZVTNj9jJyPnurL29yKQCx0OkLpSQLZuzCGt5qnrC
eMe5KBWTsW+DtmUzn5jbREgD63vXcYk/1yhIoNGIEZCxFgiBJiqpu1YbJik4em+Xk6VjKTCRl/Uy
IZ8g5NE7kubZI2gUv8/2r0V9MI900zAnzgGYbGyhAgk6JWAlSvPm5sYdeeNMt1bSXA4tJyuuwRi0
B55gdHxXb4Cwp4PuEXqQdIllDVW9hGeqpU9YEk4aaxhR2aU8H8N7qsSz3tkQV2qBfGiiex1NFxnL
5mA9cUVWOIJ+HGzrf2fnPeBPJmEmPofk7OtV/UfLGFUd3k8ktIzbTAiOzaBeRkRqEEXLQEX+KvJb
FjBosSNi7UEQuO5ChvBrz5zswBaTnW5UlK+i8KR/2zvNB4PTD66V2HczFASqIAREcekTfc6ru4xO
hd8iv8qFe5xXvk2Ld7VFMLCnzpcjflCm+y3GDGA4NWcDp1oXypj0Aditrrh3kuJ9/eC7yEeGJgQx
r1hWZ+krxiCSW7Pp31ZCFdgo23FjNxR7xgqWHFJbtiC/xC0V3Hai3VHY5ac5+Y9giXmlMlRjyVWD
pUa8B6W6J9BQGmClARJsdv5+UifeZYgGeWKtbm+lDsjMmX4+9dpr/k98Mvp08jC6nQO1eFnIyO35
/L4+E5Hwtcc6mrlEhVi/fMDZgBNDmjWHSr6p2kNn7E4x3wlQZpH5+rAhaAFfCpWtMUN9LBO7iK/u
R3Ge/3994pEZMuM0ImFqu6+7GK//kfgp4olbtLQZ8REpAjqkrbQXeI9FsHsFCZfo/xp3JSNCbk8j
rShHn+t4UyZGnHtnlGaYJi74FUF/1WDvv3lirXj0ACCuSQaT6bczazvNeHMIHKTu3KgCilQD6aMh
Zhk4MKx+PJv7zmFuX8Z3lhmzn0Vz84sEpAEf3OzDotaS8c/u1I4ZxtT5jmEvUeVanpU3GBjxOFt+
p2fvEoLTZ6oIqK0QILOdISqGf4LBFN17KG71yRs85XSpwU4P3BF9PizfVISxdAQLLM5r5QUJe55E
zxE1C86NjVsuqPVC3QXafzs5uKzZvNPX5/yaVY98zPNjM/O45r0aySDp1kAxi9QEYKQaHnD85hnZ
8aL+ykURCr8zmwi7OSnQ37e2h7kuvtCRqp0Mx+A/t5/VicrCqUTc3YPoS2SJ+ILMsvSUKy1qt2iJ
fnqDBTZiR4wYMS9GT2QsqEG+EfzwmylldwLzZTqqfPoOmSZlvEmSKVTOxTButpXVoqnwmTx+E+tg
IQ/jpGKlqGizeGql6fNGKiZdq9zfHTQEoexgwJWhiHFzOAnxifbzbfYAIZAHIHJhByjLNACl7C5S
dzo4WqAs1S7Cu5pECci3Cx/OdhdNQJmkF333JCs1AtQ2vypsWjpUA/50nHpyHkBZmCE4RyOzgecg
FcaFnYmxZm4VfRNiKG0vDxphwohBCJsNepph+1Aml9R6FiChudW6kaMVS1nZiYdY+YQNXgr02O5O
t2pthxT3BTSKJhb2Td8Hsr6hLuwpQGxCu5YAxdjy+avTtkmjAwa8HcVmYdGwG0LGVMqmxTqpssOF
z54Y7tXVKKIYNOZ+Hz8QA3yQLrFej/bUwXNJXfT1nnpb46R7lYXHAmJkzfKRW4ZnFae9nqsbeqY/
BdVeoUF1pRP1s7XPgSNt+f4gkeymEiO3KB2CjtY4mfedqyZ9OaJ35nrXx7ZwoUKO3//VVJOnUyiw
rKTdz0PotobiG5wGim3VI7E0TPcSamCPEJkO+v5YP6xH5LryoLc1/fRdNC11XKh8g9ksFqQ0q3CJ
cZWgfdFp36fuWl1eIdSrixMaWN4mWB1j0WJC+3ZhZvG1PosDAe9RL4FKIvedc8/OrZ837vTZhWnF
8KaDYOKFTuGXAfhNIiBoiEtRbZwdFmnUgFUZdufoZ3ytI577i7Ulk1YR9RXrTUwb50nhum0NQn+m
ihYjovwMquX/Fjm5CsYglukBmeY4mwTWH7Bw2ooIorFJAQmymm66HeWHLspYGjSES4DIyxuBLEF4
FId3AM2+svHetG6G5QACkBLYesdvhy0G8MUlhAavEcz0Fsf/ghM7RaXyw0IAdEoj1y/IZILcEW6b
n8jrCAWM/x8NTS0n7NLnRz58fNK64Y48dcIkuONFhvaUUaAfifaNyKipAEpciwkINtha7HkkTg0d
p3km3HeMAWrPzAgJZ7213NRQA8TbEkDAmeJkR5YzQ+AtqMVQ6EG3mp/UE6wpyd57efpRWU62Jdc1
VyivqLJ6GcPyVAp0jCf7cKoln9U6vhuFIGBSgNx5vU5Iswf524B5xYO4UsufG5wx6N2xt+0NMqDl
W2Epme7uUJ6rtt1ck0QLFfEk/WR8REvXExJPpEccYBtmN1T868e6ZmObe6WlDkLacEbQ/yvLu6Gx
Jjza4jziYia5bjt+g0Nu6pFecJ7fL1mDHpx+vIl2mryPRFc99Uu/VM1Uz7gA4m+kGMBCnglXcdp6
+FfHABhCP77qV2OJJLluzKCFUSkQQ1s0A8GI46H3TNL6K1vOjdWORLmnPUxxrQtbTVeCBByP9xTx
0KWifTczGo3fw0IzsthIQhR3py+HpH+k7CgGRMlYf5s75eHn3+wInMd+H6qBwc3MQVDw0Ew8QjHt
AV1j4i+QGwGA9GdYOIPJFMOcNmrzq78igHGtQsC9o/Ps7NNGZMfiVHrGn5J9Gui6GRx04Y/hhZuR
ZQC9D8Nv0cKeDApXDXh+H/rtftfGjJLvSlOBuGnQ36bus8FwxXcDbeO8A/+Z6SQrhTCDmF+wFaWh
04LVLoKOcqA+u8nXR49iPu02CNIOil4RbXnQFcCFGo9JQzdnbx6vmxYjez0y+XmPapxwBd8VGRe3
Rls26NYg9ThFeumON+x6as3/Sb5jzr51EesUDbMnZR19AJLQyO4cVU0MXFU0XZMP3ApwQJ+iYGfu
8H8tfyDkckm00CHtP7/E35JQMDevIDLwp0kAmGhP3MiF2eL2xcNKbJDzw3bSxyaCRVDYYIjH9Mw2
cxNwPZQCbpyUDxAUG95b9BYsrSFsYlI+Iy34e9VZFwwzIODxilecf63wkCJgGT+Gh3WY0mpvNxMI
hSIQkM1i4p7qKqS+GXzRLQ8Zu3TgBykE4ev08NB2ky0AfLg5vEJrCrKtXOE1+VnjFhJr83q7oVJr
2FGUHAFnMcKKPufX+UxL/3x+xTW5L4a7ZNDJeCxBo4CVE1hnNcveOa7w3PkNHXBYS97sHuhj0g5b
JJhioyjlZWqyyrhXigesOHXlzuYTPzD5y2lvsshqr/vOl9VBD3+rVP8aHt5A7D/pu8qg411b5jlr
VcGqhYWnpjwjNB0xAmFmzWp7cJhyvrNN3QFeLTT2uuyK0bht9bmhoTXp5mwmC3rlzuP7nlYBX1zy
arAZ0kbvda0uuQMk2kxmD+CIw4gCzTXhGaYF/E/CP5MkhHTTkK8+ZWzPXeMWAuAb//HAI2s6bFs4
P2wrYPnvPWoHtIsB8v8ld+UHDhWIvfl6ty5XoZBq15nlSGsqCCZ7ytAbOIiFjuGIdsWFdP1SSf+2
AnlPjeGSFwUywwOwvkXb1snNN8L1pa6+mHKpZI6bh7WmAHL1x4c0CzeTwagGoIyFhRy7xh0mkfPT
StYEo7G0cAnJryARVUP9SdwpVJ9QAUY5OepXaRBW2F0B/erTXbSoJBtDqNXuunnSTKm0p05nH97R
LNWBAloqM1tMnNuMTgvFEUBihFjzVd9MoyXBcvpDEwB9yQpCpm6dkiU8Ms7ADIruDIq+HmOe5+ig
/WdDwCLpUXT5DUMhbGecy6f54DnUKsfuVWPzH93BF5luKaI3D45MRrOMb208IHheiA7583GZPEg9
CzRDdad6Yob0ONyqMECofcqNdtEAR/7UR0XWZLO+2avUW7uTkYMsp9QgZP6d6n7hBhQ7uZrqurXx
cA2fzJRDmIUH6xX3yhjAR/UL7x9Ruh0/rTFR0zKWGhpJikD3BTCo+oRl3nNWuQn02ieaB1Ka/DbL
ayIc/ZSCCDYyTftdmJbE7gn60Qykfu4KRZjwVwwBDbi9HachAvoFdF3GwOUQJSc5QJXlATjagP4G
HMuytBnPfGU5kLESHd8HKe7DrCEk+no4GjBhfqNU7qNVqtRFc3i5ig+IyMhaYsefXzm28Mp+F8ge
ySX3PGa+ZyYd4PZcbyJb7pNR47oGWpoiFeUP6khIYrpt3nkk38Qg3+WRe4haNbTE1BsMkIbVllYl
LVRktXxEGyRd3vBLaw4xHi+xZ43o29f77swbiqPV7TOi3cje/SnxPvtKdqN06IU80sLTe4f0BiQo
f0O6cwnY8I8Q1jw7RE91x/yXZJKHjJx3M8bTagzMbcHPP4s3y5SfCi1hbr8PCIhghBty/+H1lqa0
2AHvL7smGgwq0H4BfwlfU7kfYciNv70bVr91FVBYUzfGER9Ct8gAPK4YulGiIw88XEtG3c1sPWZe
FBQAgx7Vj+Qq7GuOxdx2j7TymyBx3fdbanzQ18uKfaJEz+3QefxrKj00+KS6nw53nGqWqZzsImc+
B8ha5tXceHrTtpCjofijundgOdaliMW8W4VYyK40ZB7wiMsu52HauZnxmVKoXqaRWdbHQFZdl2bE
yK12iVtm1v/PDARHVManOTZ4vHtYJQqocSJhQa2vunwPqkAemJ8o8WoLMnnNC0Ny1MDL/CwuEiUu
4bjRML9RXJws3yRAgvmRlF/0zxde85a4XgkcEPZGpmPKhhlswgZN1KBewle3jSIxVTIBY1yT4niX
9H7sgytLGJDzgmE1qgQtnbwuzeq/miQcSqEmGVfpxVyEv9UorLAQWR9cHwg3Qgh4EN7rvTiwrKbk
Y0N3MYx9Av9xUeynEzROyvrz/xQjrmxN5t39BbyGoDgE/BuJqmwIR72d0ObjfP4g6/plfQ9H/gx8
OyoIByd0E0RfO45BUys/e7FH/SPhBBwmSszWf3yaZbJOUT8I5CLTb+Qrbezl0THiMYLjsfu73+AF
dpINqMzuKWlcr8jpxh4sxHejBeDWWo93jMFRkICeJD6vnAhgIkx75TfQ8KLh+BJw1uEhvguIPP7L
qDYTBhng/6l3p/1vI30bl44Y2M7zRWU0x1Y5X9LJS932K0GUuuNEr4FcsSyBwXM9gRTOkqJW1cH4
FIl9ZGOU2Zr9PuLSzpx/v9G/YRfEB3H9K/3IwUp8+9TOcUzYMVrllokNtJXngzy3UgOVOqGWVO0g
rX4licoVQj7WiXpAv7E6J3RJGLxqTcQD1TVWABe9Wu9/Xx4zi2LktPEwn5jJiu/XnjdvI56N9qPP
bRCY/awp/yKVM6AWD+BIsmrOHSAVrZg8qp8KsCSLEx6HslyGAtvvMHAGlYS0FhATYAFUH392lP14
40EY1AXS6OGAbI9CguhyXyezMyTlEmpQXaQxJlsCskuoMQo8n5h9QuhLzvPuYhkQFNLj6ylESgVH
d66H9cdDiOi2SQnf1vapNeRRiksZCVOq4Y/8Ml4Jh6tJEZmmOCvBkF+OOcsOTYvoJXh6m9g68UAK
yKIHnnXtkxfHBHGoAqHVP0wVRHxjkq0ORiLtvrCZoTR5MER0/dknf8xhLVJmD9RBluEU8p/KkKVR
WrTE6mBeKne/dTvaUn5aoStL1c42v8F0HWMabd/fLLzGzw9V1umq4FI9OOaBl7g8q2vbYP917gII
th1E07LYVY5CNXRwX4OxbPKXtP5xpVAx/duI1fBPZssZ9siCCO2WBjXrki8pcuEU49uve9Cv2fo7
TUqIGvjHwlVcd2dYRCFn/yr9u4+yIqhuqx4O59N1Bz5XXeCz2uylCva1KOiqre3llAnDvfnCU4H1
4Xxh3RlzDm3bn7uJT07mfWHV24+CNJwY/Fu7ShLlbOArlT1CGKIN9IF8PFNLzPgxGluETUttr59S
b5A8J4qZLUTZ8EGaUjS+BC7uRwhx/Y9ZHWCcwv0hfI/tTfTWoSoFauMoz7hToRjPBNGMN9Ea42mm
l50PyZG4oMYIl198UlMvJgCq07comj4N7gD2UMvsX5uN6N0ACB59UEUTA11kN7lOc8qd6yIWoQv7
w2sRoz0fizcEzQieA+hJ6GDQcvsmQ17ThybgVevivPPNovHA0EItIFvxmuiIH4Gc2+z72EANdHi/
CUMD4VokHkx38WS3YBK+yTLD2vIdyvnGTe6B+ItWESEXhUUwofPRRP/AkQBa1g7KxtXiavG3KLe/
YbpNb51ronw2kwHO9+zM9nGk8BxODFYyCMs6+VqYckDWLVmGHP2dzkJndQ8IoJc+pYGKXgKzi3b4
JGDutN145D32rgR5LTmAzahTNkux5Sp12HPBwIsGpxbVrbaIJ34RivcxzhYLbVB2SEBY1w2fxvgw
m4wLbMWkJ21qVyhq717KNU9AZjxYFfimMHK3QnsoL8CTfA04hso3i6vf3EuIN5YrzSPv/UfptaYt
5ZT4R1mJoeay/vdinp2rk6YSwCYBZ+OswysZBBizStjBDwvLX3b3TqYp+zdVFwtAlf7iYGtpjwwu
lNHAYibu37/2jPCjGIDIQet61PPc4KnTD+Xv9DVxWI8nK+/8jJbY/58ffq6ZYcHYUtyO2a6IaTSO
HdcUxQDQt3M+VbBgmcOc2Ve05ScnzWf6BA9IaMwN8i7qFwYWUMtNyakUkhNWsf57yvQpv5wekEvb
gV5S9IK8sKd0LaqAOaitNMYbkTuIsAKhQydPOzC7k/qlImn7ttOOcM35gf6ZBkXYCJuoC4n2OkOT
DCYkL9TVlGu1LwgBUbvgIrFwDtdvN50L1EHXJJpqHZFdX79g/Jrmgi585B6WDI+Y3WlhH5faAcR0
wKladOKxGLkhU1q5borpcmdgibx/K+80JqwS9/wFckYf6zlPWsayPMYCTloZPS16PtWayRDcWM8q
EztumfpmI6poZa1E1KJTigZZ+aj1MBQ3x2zmz9SOLCEvZTEarXOvgaQFqV4OjZ9e6gc4kPwI51l7
PsKaULofa0GCodTBKvyszsk8eSVE/clTH66yU9vX8cQKP/OLWciXAKvfQDzmW3cQzbLMdxuBNx3R
ckMeNV9bgE3aJH3c7zeFjxAgz+koj72ym6z/RA5vDFkc+VjTByIQx67VNEk9ELwJ+cq+ixKcSWxb
5TSI6jR8MObWYtx4hv/5tZt4PiT5gaVjh84UwKmCzNAsGeIIjG1srQahvg5TuPggYBpOW89e8Cud
QtQd5vEJ4ssQPrKurUnA/RqnrpGhnkobXGcqdAVHdfvEo0YbWSAGZ3MXVSi+IkAYH6cQtPrJnZ08
O7Bei+DG6X5yGOAH+BRpMqzg/7pPh+9pbRPuRPWCQhsFJgUucplquwaL7fGDIgDvXD9MnByry9ML
14atRQm4alqlIJV33wl5XwZWqqDT1bTY/Bu/Cot5/fFMxHSsufDQFwpbc3diFwn6ppoxT5nEWfHh
51mf8WbdhOgVOmZq2EXee6mxZf6L+AY5XdedSNlXfQ8K/vCJ+zoKCh5bYWyRr0dtYljeZMBMPJE5
OboKJLo0ZXSEzGJ0geC7h9YVsY62DqbeXAHGWHEsI9nGxb0LIhl594V0t9UXaTAFtOFR4jDY2xrV
PE1aODuYmvA26IEhHT46w47PTAUwlnfSB3JJb6lnaNoW9yc6IAeU3QKH2oGjLHKbPtkTm1xtGD/i
dCH0MfglTMIfhbhskfF5ICPEuL0ntwdXk3MjTPAeB8TE8dsoOSnM4WhErJ4EcgCnC8PeGNS8wwZs
Ny2q8S6DmfModHH2TDdaNTAImZaElGoyODGUpq1bHSpjA2Jj/JhKzKwBDDkVloEh9dyCzHo82BAp
UbEX8vzuaQF/9sFUOJcukpWdAnGlhgz1B26NbBLO5Op9C6KjUaNg8dvBirfMdwEUjZq8xumKP+su
hUXmb+5+qAUt1MpOCQ71cFqP5Pfb/6hAcpv1pXGyFSBCa2TWTY9DsD45aDbJKHUXME7PM+eddgPF
qDHrnlUp003IHifg7E6JW25ZDANmJ+aXznzASmUNoRiDT6qIknaxzywoIO2yIh0yo5fD6uDLY+mb
/i5IK28rAnAo3LInuiFyfW2qgidTSZKNnDAqqqQdg5FJmL9sDOnSjdFscF2NOgqYifjrWxF4EOcl
O7zSybcZ79FtK/LDCKgA5Jq906Ku/KCf8QIW3gkfunvxGOpuhw3dl4rpkYqWm7CuHR9C3DCEmX6Q
g+gwZQ1RrDA55pNuFfHelPyXJTzUbik6BTCY8xHGyV8SO6KEEUJZriHnBshsyy+He/AXU2uL1YdI
EJUNckcySordT9XLRQniDe/WgT83+99aByQkCKRn/IT6l0D/yKkGLJ9+s3x/QP1fGy+As2kS1o4+
csvXQy2YXD+t14fmOCXx5an//l9T57uFx5CgFYtzzq0PBXvEWwGncda2ZZHEZylYnVfF0Rq29rCM
G56OjQFsp1aV2seuNZaCL9rneYxdV7T6YF6M785o4JvKeU7jvMwL487UFZ3B/8s0O44Obg/dVlYs
FwqD3oxn6ofPnw9RVk5WdJikHXl4271LL5cPhtl+WwaTdNLOwNTu2u04o0/C3KXj6Uvw5sGRAYuk
muJDj5dB7Qgg5kjzqwGBwDt7yCx3CoLj+LBVEo8Acee3IHsZosvIPeWkTZpM0zZ/a5GVoidPTTEG
NJ1WQGpf8PZTeNNs3PkvVHBkS/n8fqQeQMGhyBP4BWRQ0+WCUCL2HFV1+WOoYzgow7PmBxWnhgJZ
EQi2D6tOw/b9oRA88oHUwR4G4mV44ACsr4UKkbnd/j8HBQHUJhVmUalH7b0/e6IUcbqG/UeAfQwS
bCQWundhFSWcEjr2JbvInIzdj8JRN2gPI7eKyuYtxwrBAp6TEnOzaFRZOPcElya7RnBhyioIqgwv
UoCBnTq+Sb1Zbsfhu14YBxlvUdvf5DmQRxYO7jGhvwEFkXbuN7JnZLljrjUUuWcbns1x7I3nhkZ8
pJl7soXFEzDhQ12Ps6M7KqUcJ8QrYUoo2k4U9+RKbfL9BTRjlwN3D7/MFLSpKoMzjs5myPdnY2L0
5O8lbN/TPCjTjyAinCE93AkNDkMA9iIof/r+J83MV0RJFO+ACW0pwOyScCX2BZxPBPVzuZ+RFECq
GEN1dBXplX921b1FzU0//aTuu/NWJLixfZ1bh81fXy/Mk1Bj5C42zKx/cRGEkc/13jxofstZVSff
tXnV3iDD/XkDROkPpDBaYWA64IfTrGmXL8ldWnP8HSF8XIlKUpX4ihprj1/qMcoUVc9ZZb8I9SwK
LVd7p9f8+FnSDDk+Vu0Rkeld5z/My/u9uJojtxz73fRauB/9QCdO33Lvwt1E7i67vKH8ueMQ8tFR
TD+i6d331DK7KTcorZmlnu0LhWz3uvvHWKtagkCj7DHWT/zeyMF816UDSAYfrBF8LmvnRixmspny
68x8ts0j/qAHklIEImWHiaOII8i8M7qh6lEXFz9x3JjhetX29G7BO+EyQ1B3ZvoGK5iRgejSLzy6
0I/n4sIUSBaK+llFQLXE7i/rxQg2yacS8jOr4xvq3MWlqnzffF6rJ6CCYy/cAS13/Z9kXJZmFMU0
gGGmfQgxYtdzosPesAQrwtmHxOOy2UwJ4x5yxHoJhpMfzfZcYec03we+jjIp2Hbq9P3A+bEiSOBa
EChmYRKLflJ5QWmhDe+KSKL56d2amiD64CJI8LDDm8eiAk20u4fmfxFUDowwWHbqaoj9hLXDGKCh
8YVZUVg3l9elbcMWfxpW4JjF5hB7HIbRAZ9o5Ur9DfsepG5OzG9jRaYN/MosTI58ToIZgy8hfL0N
l+3b0lKXlvoCF8loMCAqa+GrnaZKmxDhmBzSFVYgFROo+iaOXxfrhSQkpNVqeTPMN/4LUPC0Nyq4
v3FdV7kvtNXm0iYZxGS6YafPqA4wRAqc25St0xpVahpzmcEoKMxBk5FHQfZ3kRa1ee801fcHnD6e
SdjWgn49LLjWa4Bd9te50kO5Guoa2h07alvo/TLAptGbfOpJXisOpM0uUz0sbzhmlT608ka3hbiK
2JoBOS/Avb+UdZDTyN2zwqV4T8Xr/xH6jPz9L1zcYFKS+PHL5Gurt2Hd67LrQTYtl+PL74opoyL+
lE0Q7gffcUEj/IsmyIz1MZRKG5fl5JMcGb/EqzbKKmYoFD2GzdGOvjJgMK7ljGax7sKprOfUzRoP
FZ0LNQbh1Ock5TTM3Ts7MDU4NIMF6Yb1Aj7/NvUm7nfp5to+I4XvyEbu/913ypB1SoCVZgOZ9MDb
3rYR53XhfGd2w7iKFOk2HtyfsZ4YEeUPMY8mSCa2PklqoHOT+0/LroYYzAXIKCM/ukpXxjmgCKQ1
j3CdRpKdCeVQZHRPtaV54Km07PVMDcWO9YY5sjGFbCFix9fjo1l6FQeaEfanT4/zC/2SjUfO3kK3
BO2svgcLzYntZklGv0OcWgka0R2594lgo1sjqkFQNhwIrCnMs8PJH9IJFoTiNy1/cQhKyuUqGC6a
6bqNzPAKIcuHnBKrPVt1I3tKGVsaZbxaDZBoQW8VaT+IGIlEogARB+gsFBsujdsaeNc0MGoKnZ43
D7GaaB+AWB0GzrhKzmVwuGvKokdz00l8gyfEQfW3KgMhejndLjys8NmnZOtfts78mfqaDeGkar8a
sDZXx8zT3+ryT5XODCSiRz4dRGw0rOTyc3GKcveryJ1ri4CXvIBISKR+8Yh9fDvdDLkatMqa8Jd/
shaU5DH1YMl9NYHkE+HDKfHnGI7wwUR7M4iGo9JPC/5XAGQ4Jg/kVETREzXqaBQXgKGi2F4MPD3z
GhZaFmekZZKPDrdbM/Rzfggr5JjhBNsaJ/dR3ZZYQ0VTuK15HBwsWKWmNJG2iPo+0iDYa7CdYTI9
ysP+vCdZUellQkRtx3SHkjekOpoJPRwXoZ9A0qFc6TV9fS+jZ9HzEfjWyuO16F1AfYBPMepO2Pa5
YuByHJdLSxSovZ69zia4i2CpeggXX4623/4YnigyVIkUpOrgiFCtDZXwVPbckIkggKjlIv25XnKw
HBrqxLDtYKrC2p8F08Td0obKb/g+iGXR+JmLwnB8DV9a47yXQGHZIHmBIgPcTD3fiuLU8A1juyiT
gmBDHp2BgGwMR+oaq+TZIGjv38C9fPe2G79TP1+3OB5X3NOlo/YK0AQhpQFfzzusjh/vQuIibFH9
9ZINEfSS0mCxGQvV2JqRvMASDyxqbHrTGX253aaTJPsWQ7XTgB43QExZFmliTphkYwudq4kqvC53
WJ2nnigFF5hpE3TTuMZN/8Xjbg0n4otr9l2v8omfuvl1tLP0LNRBkC4uAqrx/AonUgxw3lJL6yui
uhep8zovTA9jmh79mShuXHqHvEcoeuy1uMVrXdOzmyEH5qc6abfd4M/tMW1a9oAQV+CKp7WaVuXQ
YvKbmeUZWNYWPkqRyyLtOA8Be8x5KXq+BI2LHmPDxYnHuPsRnvbBXu9kxlT6TbDGjgTm3aFdHfKQ
eItee8oUURv1OYRZchI7XMXhzUWJfYHMq8tPYPTzs9L6U0ZBBSs0aju5YWptxIyDx2uwUdvPt314
4yGQ5yB5bfwABJrgs4JyMQKI+H5hItbWDUudwyOSkerx59+EufiKkL14OlAnWJ4U3t80ruD9Nike
YmouQZTBYC0oqAAetiq5wks2DsDD4VDpzRScSId2CRNH6+ax/Qhs3PBiVfjTTz/62+2ea31SbgFy
kwrx3f3mZCxUEoS668RJGVlkgixsbImVDpli11TbRs8ZtX2ZmIlGjAusmAhyIKgAZ1mqgnfw2rNl
OXYGC+tRN5ff/uwxuuylCnav5D6ccQf15S8LNflQgH9y97FfslQ6uh0SPf/A817++9bJjxqe9GTw
qlpq2mJcN3P0Qi8OC2YHxEBTVMYUDFVZS9tjeO41/+b13uHrZLMGuam3bGCon9B9qjmY4ijUyE+v
C68y7U6SUa4J9z/OpNJ+U6LvkUjvAWVNvuSZ+KJP3E/Ge0lpfXikgNbVFwlmbeou+3WYCQOvrAYN
pP9dEAhGVyARCdjWKMUakwayCtJq3QdqbEt1vEICbqBj0j6W9IxQbQsX5G+EnoauAse5244e7Agl
IBXJ4rd3gW+pQiGuBgaq89OZkshNeTbUpt2zzWwNYXUGRcF+tmJxxNqclpfXaoJyTpRJGJbJqyb3
2JLyTN2ewzlQMPtG1OmeOhFIpL28LhjttZNsjyzpplWP06/r+QRdDKRrGqALDucrVHYIZDGr3vgs
5sRgeiCtqBVH8/FIx4GelddmBkyA/BHuvxWPdFRz0hGfyYhwO0RVHhA9R1R52ZeYm9aR0Q3TfZle
YZyehcdtrIk/9Dl//LH90U6ZDVS42Tu+ZBvIDE4uM7xCwoqc9ob1JCERE2Z9LTMQgwmKNywb2Pjl
z+0OYcCptLKW4x0ZVEfvBGZsbEW2bs8FWr61V+03QjClD9KSzVgShG0W/EdfmRy5Gj1mkMAWDk/F
2LjRn3sf2MMnidoaT+PWkdKffrolFdiM++QQTqqyungXlq/v5E6o+x2Fj9yLujhtvkuERRdnmQwy
kcRjqYDF1Ns6blxprbW7iWeQ1iI0/2rFh//C5RG+YtEcrTLbdplbP89xtSg9oQRrKnuHGChE1Y6b
KIHBHCeC0SI7LA6F/8qY/pqZdP7l0uh+oGZQNRoqeq3kVF0W4DBq3E4bFD30f4heFRJ89VOXm9Qm
66ljKw7oqgqP5A9r4R0nHeIELm4ADSYMwO+oq/EHp64luo/PHyJP2axTAUJJzTBc7GygpZ1ZYeRs
XOJV6Wz4azjc1jfbbeZlqI0ijLz9kUgDhFPA0YaLVlKqPv8icdNCXsWuYKbSVKcwD1M5nxhYTioh
uPkI1FKgqZDrrMC6QPa8Ac+KZEQp+iorLiH+GVTWLg4tMlwAWywnIbmlW0vXxYyvmSFlSo+snPP3
bE9x5o0U2RJdTuZd31bZXyorw0fKpMC2sgNKhp2aIOLuiGjcTPxpgIJtu4YDrecSyb/8KhEDUQeX
gen9gouHSd3ugorvEfGMVVzgnivvKfbo6ioMLXzPkZIbrP3vkSZpP6Ll+r/ADjA4H/ArSw8ndtXO
8V8PNOz+YARmcE7Nr38jciOndcbJ1HPC//JJW2FqUue2r4IhcGnjhNxU1IOk1TthUmQ7kFOhw2pj
7XCNSAAK2hYuSeOK9cB2/VAw/vM/qJ+pAVeD6QPoCGfb/nzGkCceEXFtfFtf42tHtfUCOicmMVuw
03560Gj85U/lDnwJy4m9TQn0w4XC/uiFsjmXbsbGNuol0zS60w1HXIxaI0wZptHZd/DnwfZhMe8U
PxhxBAOi4a9Z/mdcCOvz56mi6NOB0nROnKxjOdZA6PrU77vJFy+tW5wOg+RY3G7dwr3rk84xmyG0
JGE2ExAMVPuikTKGTighzX84Kzue9V8HMEYvW9i+quVyZPg9mcSNQVbHSjZwQxD3U92j/qh879n2
KVmTDQEUphR7W31gy0cJIzT5VFYWbkzyOs7PQzAKhqaC31l/Xkl2SUcwdj6ufqV6wzKwdCK8sa8i
6WcnnG40NxH3iXNxVUNE9Z3cAv0z1ln2UDHTamDWetuHzfxlYDwhCqJxF2fTSix7NTrRrZ+45yuZ
zCwcmX8Wn1U5gId5s5prbjm6Gf5ymD7h1rkm2bjS8fbK2Ig2ATGob9ku6GkcOgngpJJoPfxWy4AY
XKe57ZjkzjuxxjyuTpzmHhZh1/Lp1M5tSypJX9j50bhmhPCaYbXMv1Dwt+eYUOMdjUEBaAxg/G4q
f5m05k0pOouaBa1FGSEyYxcfvp3xVMFPwOBHSabIyT1rVbkrng0kuI3mhMXnMkVu6c4IepQ3qdTM
3UhAfUuacPQOUaILkNVW98VJ9CGla7/0VgRwk9E5ozndn8SosWFknw3AazoWrYPq//Q6ExU+1j2C
gwHC6wlg8ZlBYYOpgnxBGyILxI16MyI891J4d0F/VofO2ZFhPVHJhJKiIVJtnYLAevUWcdkKxXZG
vttEU+L46iWvXPnECqJGA/r3wSj3rycsbRHldNJmRJ/Hc+gQU48Q5PJAvexY1yQO8DGoPhjCcw2/
8TlSIAm+7igyV4tfIPhvyXG3rByHcov/98P/XsDfjUpmAbR10KDaRUxP1d7PmfoJGjCstwfVEoda
gVSVvvDl1D+COpWZGojgqSoqXGxTDkooHH4KeLPMQuUVAeaAkGmc0muy//21cA2cF2aZ1xAiMj3w
tvykSQT7tIK/hg6hVOv7a/5VcfbzKEXJIccnQssfcSQF+TGthuH9ETbpTRhDzZXTp/QkUhXJZz4q
303d3y+zfB0l01pPEBPCD7HBbWwhHqwu/oeoJg7SCT3SdeSVBoGCXkODoIxOrfUJIRvSgVDXBkoT
Zrb1HuRSZmOMQOjo5LfWU+TM9NAdU1wBoKwzlj+8ai3xddd+yG7RslAjVtz1IRwmpBIWJSXtCSRH
azNjyiRgDogtWOp+87YZtDkQhUEudXxkOEfzKOxrhCPlKtfB9V/JG5NePhK12nJG1UqJA1LsvlcH
kk4MWquLlEtTRlL0/41zO5R7YvU/BLQ5slameXjfaTo6oHehd1i8kkA76lz5xcislbGcunCFdGWH
tLQ2qjMIVA5mcAWgCXR+TOpg3SZX8nk7MifBhUmi8URkTjhvZlxvRWFzz5FDFsZy/52exQgCSfZ5
y8s55/b2rTRi+hp8eVU5sKfmkUXXKkRHzMkzkRpjsbu/hVKumQ0zDSqsSpiID843m74aLE/sE0xE
scQhx5bquoARd7K9ZSfq9HGzn4DTBXi+5qm1utdaEteMhRZt+LgJ6MXvCHDxdTF1tUBKn4NGHUxU
0onOAlOff5roHJHA3X3EOypbfTlZmbW0egQfW1lsPX/HPsDOSbP+uBGkDfUyfC6kpmiQBy5MQ8Dm
mtAiFm7LINnQ90aX//lF9A2bQEPmC5eEkQP5oa9XoxQO6cUiSUZNMab6OoBXXYd4OLSQebkEO3Qq
Aro5umuBTkpMZTPmNwcL+XIk5T4OmiDOwN5elSNzJvS243H7BEVAnnVwztGte3NxM6tYClzEvqbo
eFUbtv0NS9sBS0+r2qPz4DcshNsxsJFZL0nSJ6fMb6jMPUkTpiu2TmyKC/XlpyPfIo9+h9BxtKqp
ULNjRYwbuhkrisFKl0tnAlDYLq6PZ9caJ1RA2CBMdpMav7LgLW/oIeo4pwa9WSCkMwv3+bOmlZ3W
opfXYdSnyrgfbtVSXT6mxi5srD6+pd6E869vfh6sHnRt7w9QFA7iodcXD4Tg/MTeSxl7cJ89aq9P
UVHt30rWNCMWxCm0Zpwlw3/vWp+N4gE78ZoDhKhAJofOvDSX8Jxl1uEFz8miUuJM2jMawbqeVi49
6Y+AjTTOqNE96cz/5c4SCvDvmsKrbtFojZujRwPRzyKTmrbQNRlg8Skp6KJAPBqKgvO30FFyKEXw
MNcusbIFpdcpPtr9MvClMyatqNlZDP3q1aeZ3gJtdrwhDJZxDuPxu6Q7UQE2chjwcAS/aVyulRaH
91sJQx06bv9SGH8a6HI3dguPTKVLLc6G+6yRpjuvCX58RwK8A/LebAeY4/xerqj7BLL26UM+vNxl
IeDxgaQVub7H9fNsJsUDRw47KjYiH1Wp9+GdtYLTJL/0Rrz7GKSoFbc7e8UJS3KqPurW3X/3S6Ii
k2B5EcUKJfYqfKjW1TLDQAdhRWPe1WBEcO3/gxYPR0gFFFNmb6Jo5QbkWwKWmpdfkS5tA6VtTmD/
IeC2ioTTP96m5T4nqkhVLaeWofo8teP94zot7HF9xbPyaEwi7kYu7pCvo/EcWnxHHDAp9mxq6LeD
2T39nTAN4LdwpFWUC31YKHosVUi84nycMuRAKv+bpWQb8pNXRQqh3RstxfCi2/jMDVn/Zom0ZE8Q
QEAqAv70GIOPscRjf2Doio7vf6VFbXFRZGNcdthBHX0wP8U2YWcklpHwvfU1a1ola6HqmX6xuI8z
wSZJ7ZnLBqBYL8bxH1n+CJwD+2rmPxQTCGcNfEzsVxNpXwc5UVATZKnsEmoWwtl9A05Wi227tBH4
l2Jh4FvF8AvWFGjOFBBItbNow78asKynrKE8VsDNznZtW3R/kJ4u1PxwOA+aie6ePypgF4c8l+33
lyJ2ijaAiaGzf+MuuM5GOfxPQgkODJvEDzjvPQfT7red5g0Cx8oDWKrHVbNTnGwUqT/N81QLbwDc
eyjANn3ZZZqtNLrNs7L3wJFatMgZweJoqrQXm0IAZZvPDx0NoyJspDnVToG+lsT/5iOOD96f8JuI
bmkg4oCsuhuDett4FXoePj41og9MYvMW5Qx+8oc3sYS46Ur1g3vMKIybDe+NJmmk5oRg+ruVAAG/
/npRZZk/QDJ3JtLPVS9jA5TYVofdgGwEzXgBWzekcs18IfCw0QdJADnjPcPmQtG+oe93XgJKrZx/
oJSAIZcLfY9GrZqBAOCC2O+48acnAzUKXeQDMZNaLCnqj4e/HrmJVpHGZZOuom/omqXb9QDaI8Mn
kzSAmF4GYL/H4rM4VpA/6oKSylwDkwLCEyGdXKcpDgtvf6dG2M0VTvJQFbSirv8hF7v+LmSkuNuV
iMBQo3OFc4DCvnbV6HbaK2CAIFUYSxEerjr9rWvfrrcZNNLvPUF3vlG6JW23718Z5WsU8lrG5GFa
hGiRJ9KVvhAD8I/egZAoNfbrswkNqzk4zlrtctVmbKVz2zuAtXCxuZ1lfz4ngBwoeHEaiWJfcWC1
hM7WPkX0f519b2NoWugo0qSieFHiSqzLVlRZDmddY9685J+QwSvffBxPivakj3l8xEekxQ0EE4Ky
RCQFzaGP6eHofiIo282PX8+4dpuTAZdSbwVr4GCYdzB5WalZ9r6v7UPfT+K2E7Bc03nLWyXZYElo
ha6h2AomW8tmGn062pKg0XEyV2Mal4ofgSMYpijZpt5Mp0VS3bTX8xuyKHHaeh0v5PPxG5/DrBBp
q5B4PN+SjugGYU5GVl1ZWMWMrMLr11au5YYM78Cv5BDZp/kZPyqtz3iSNPZ/erOjdXW/B5cBO7JE
DTfkqanPKUvfApq60+omRHLbYgJecJAM8n8ybX+FwvcMOu1PLC5n84Tk9n+2q4Acvc+y3AmJ4bNj
XWB3mbYa8E3/mA7gOoyAEDVNfXmmyFgiGX82fkwYVwzBASXtiXatTUDex8wNNogixGvAz3bCd/i7
zV8w28tBzu1T6mC535eMve4/qqd0FMNrx9wZsOlCPctna9F2IZQv3sTeI9RMmRbRBEqWXRmifSxB
9SoQWmDbO5t15vrCUWfPSOHqqzTdG6Cbm/PDg2XWFbdOwLRRIyJHrc6jeVkfAbwnpxASuOtyLP4f
xuAPAqjdCHXZCwOnaG6HYRRlE3VqfhdQUZVqatNQa29yB3zNDVY6LXrn6YK1WEKuyBBS1rorOIdX
afgbc3gPe9O8HzPfvQZEraC8ACCdLUWq3+WfRdiT4m4m6ksoroG6+EwWhMSaBkH6xSMza1f9mXDY
24m8M5tmFhrwja74L3dCotQcFqPJ4fnpLsG/53/poPezoWxfXLzPMS2rG5EVZIT/FUMEK3yu8se4
2ZHYzD42kQlcVUwLTUw4MOOBoEP9Q3ICW3qLXnKJvStS0BGnaCfbXzmH9FlAYugvRfkwda8FmapN
jZdHypwkQlgiS07f6DNOGFRzn+VP5ognh63Pb133oVUpijTcrpSK19L8MNOCS8obNpAlAvB9E2nR
6SnaFnGv7zTXaIQfHLCfZK+mAFI6o38w4cmDxJfxImtxT3WFKqNy7KvWmugFK5ZAVownXief1/TN
ymzB03fkr32qRl0iSm2UfK3t1RZaAQGGqinapmxYx2H/GFZRrq57fyxWQwVXiUSqGMzIcy+uCDta
OaewqU/qVDIXiW38YXqzsyvIimWRWPpowMdCoc4GQiggScOuf3+7s7xBotBQLfyseWQqXg0mjmX0
uRmha2ugO4buBRgAgcf2Tk0jhrbNHQk+A9fqLooI1pogadvyM67XqVI07jcMYs19Mc19sipxeFRm
CerZUs+XX7kXiIk6MJLBRjYDu/+UmYBVRnRG8rK2Vec8UNrtf8KYs1qzlLuWrhCDei/RsN3IcAxt
l7KQeBIPV/yQytOu+k1BnBrWhzar4y8P1qoG3o7xrN5BuBZO7oClVJbXUyIfdJ4bAF/FBh1OT8xS
r3XpPlM3Hl0i3Uo0UmhKJttHBpw8rPGHESIxpZKTpNExfOSbtkwk7Hs3xjdW/j2FVh8e7fI8Fk76
68HM4x19TDDppIAeeCMXiuX9qYsOLk+YCAImoga7C6nHfrjUmeH498xOeSKxW2b3onAnkdk1NTgz
JvD3N2snOoJtTp4bvVVdYNZkM1g7nqUan/l9QWWysvQwiPJC1Pg/MVlsdTH79QvLlnk0+BFdNXci
75dsBKildBfXQU1ZFyYVmRduESMiZ/KmhHtmo++alkbnaOln/yi2uRLbtatlHpmDgpmRTw2GKkh+
3FqEvblLqjI9rlstxE5zClNH+hvjRbMkNyVPo5tg3Aa5BgbcGBIGPK6It6ciKFYOfxy89i1DZ2z6
zr8AZdLnDsbbGbu1+icltntYJGFYlvzQ0Wb0Vjqe3j2Kqi75WvWs0oaM9pHIAwp8vvRpPl1rLwZo
MSORCALGaj8m844tLNMA4Nny80pg9nI9VrZhXCwyKQOaYEMJE3ix1Qx7EM2bzBQxC8VdcvZfNCDr
WU99pGsExSvuGJ9e3xlxm1amxy0kwjW4jeYmMSzg+r+J6djOJqOK/aq9cUORU7kIz6A6y3DSJ0fU
wG9b8IkAyip3gKZgZ1pJ9YMtdkprbDd5SP7zK1PFPDEY5drsAQ4NF1tmxSuwZCkca0uQSlJP0A1a
pufor3XwBRQxAmxVWgvTuKBjHNT1ii5kuiWm9iZN2tM32x//l2bh6pkUZEFgDGUsO7I2uKSF2wd8
MzpyvsoABd1K3ovwGmnEho7UXmwz+kUyCWRHkNYegyGN7BNEY08+1XleegcDpZsQg2cvVgj/hzX/
L2CpFzC5Alw/HPmfj9dM1HTLWrdXf+TZBIESKq39+s86yM9STxyJ6i+/xYHqjAkL+isNYIXuIUH0
jKjd7WKQIOsYTprHUtrE3GKkZoq3XYsZZAloiRes6YII74ZKLMl3m6k0XcPQOAn82ruE8jjglOX0
dGdc7uUUPP5Gr2/ZqaqkH4bOa0PFQ8FNR2MV2d92XFHevSC/zJZHfkMGjHFJGl+yM/3uoX6H0Tm8
OpoZw91itTyr61eGSSpSHCQlERuNn7lmqf1A563V6EzrDq90ZSQgF2Kp+6k8ZSL+jTkS9Ovq1RI2
+iSfB96aWhy/1mot7LOf2qtTFpPle+SMWMzxcyZFIxlVwDuCPJHHCQgBRJplm6H5Ma+ju/IiUAw2
mXXb6SLRzc26aqhlWayZiSbK2AtV1nsy6P36oSEw3+FYaar9/amA4A913OCG/K2483rAOPFP5NTN
NcVbA4+wWnaptRwBpgMYb1fg68zFcBJe882+ZmDiYSVV48DOHuhF5Ex+OjY35MQfKTzfHZtathAj
/MvwE+qWP5MLBOD7nbttCxjWgyDXuj/TviE0b6EL7qZQrneBxErpdu/QNRpBz54Jv0ifgleCIByM
TQ5bqEcatFOP/rgi/Ln+xuQ9bm6WwqLtJ0pYs5O1Mf9T5wYJVFRyNlO1wBp44caS3Miz62e0jVa3
+wPBSiIWz8X7B7P2vJcWdUsyXVCt44zBngoYcrwEnxKhXXtusqMlIRK2+1k8tlY0jUhTj9JgB9tb
CrVV/Kv03InvXfg7pqImAKgsVv+u6GoHFQLRfRLeuQ8doPl42HrWDfItCFO2ZCgPn1mIh0skr+AP
Nxqmw/S3ULF/GLw24kWionYUOHpgA5OUT9pyrjzTyptk+2A5z4Tri2KIl22WPkU7Mb5dh9b09dGY
NcEqxKlIVhpYJDzOX1+aKW5pVRA5fTEaZ9fye3HITIu0M3LaYe89gj1vorm5tHW/hvRoEbnIQLxG
lYS4f4dwv2WkPkGRQvK6r6QX9XnvxKC2D9nwLVzZrAVDDMT8+1qzRvnd0C3EFNoQIGEsE+ySPWSC
eY8ptYO78XXzfk70IyG06Ka3cTkVr8UhGP6mxuIuupMtsGGSzPJRNt3qDyMXJ2u5G4Erbj7pNZEK
HEiny11qqG8cD8do5GTJmsGaY6/ti4G6HSDh7Dn17X2Shy1D5QzCR4aAKaUHrUFOr4MPePlfp87J
2C20VoG3TgNDEv/GftTRgOUpnaZuC3C7pHCMHVKKvDpEwI7338/rILGQ7UlfwSgvW2dK+EP0JNv5
aUwpD07gZ0Rc1+2U+7tW9DH7ZoJeykIdh7Tnk38Jqw58L4zavegYllmLjOtf5t5SVCQSw+ENSgOa
FwBdrsjCIIUOopz2g/R1HdpOoYL5YnxEnNasgw6oxfcQNX3JvqH58EocgXQdKO8ElBajaGPcfzn3
vxc58ZY/KvjsFElafcr7tfhXa1xDyXjKlXjxZ41zE2YQNgWMnwcUKrFoLMNdWyLJIx6Urq5jAbS0
URmXfD38kvTN+fRgA4aOq2WLx1OZmNUDvGua7Dq4DfFsxCNr+fk+AjttLHOAuNt61hfbWGyGNabn
sCfwszjecUd3Hm8URsj2OHx4zQr1CijPBh+xyc6o3OqwVW5L7X43SIUwiEkHjdVQq3Ivy30QAP+8
bb6mvrmvTJipC8aR3rsMckX21rvfzdJmSonK9aiPJKmFwaSMl5TrjY4FVtSHNpRjyr4NG9f0GMuE
iCHi8lFt/nHidMLbhcWv5tCUxXvrFLg8K7YvVjR4pfHfnyM7qT27+snZq8halHr5P9yk7h8y4h0E
RprZXHa8YZn9e57pqKbAyPW9u97dF1JWn7XhStnt7TDQ/zNhG//uBTCdSdK8sQTMClJEuCinPtLV
uKeSnejJWi6P/95EpEeUouLY9wRaw/SOmhqRXBAG/wRT3AjsM99CPP7f9lK1lNRphHkRhDnu7q9e
ap9BhRno3IAQWfURNQiX7uzPyg4mRnwNbGvY/7nHbt5V2GAz1JnTd54//rMCNIl4M3kFy/ObU98Q
qn/xm4L824+qoEgkSD+CoGiYpDn2oa9pDwWiuTNh7aBEdGeCRDmdxhbQefxhoQZxCjbR1UJoBTuC
uEOHMWy9HGTrCorcOvSloXZ/+cYhl4+hA8qCQsxKWEq/3DOQfIRUB8R6KHFNtwFHeTK50xawsuKD
3PW9sJsllr7a2iihoMhsbZ8XkWEe+75r9blUW9jT170QFZ2QkWLEJKJuftXk3GzYS+0bBQAkpL1c
DiN+Q+Ul43J3daEXjMz0I9RMOdtpXuVCaZAK4YDPZgDZzwBFjt4vBFgHwd9PEtDQc2/0j0itKD62
Izv2hlkndXi3DPhvRN0SMco9ris9K92PhieDTQAw0MAmxxx8C7XrJeLfB/oFYqzEQUHhp/Y7THtS
flhxliTT4aIKsdGLLeO3/rTXQpsWhr8F8dwgPgfvHUUnqjjhK2IULKRCQ0VJXXGXQ61q5WfQVbSh
z0djttwSL3juSXyogQeLJhzalAIYllThPZUR3L/HkTk8CfYDKVxh8O97EfRxmVzharSq6PXMTQXk
qCjeWPiOjky+6oKAka0yFtRVezux4Vkfe6dQqP5oL7yO1nHsj78IZ9SXt6nrnokwDuv96tbvf3/K
6yURrNEzyuEXp7oCFsCyHbZ6LI9oQA/Nzn32SdUMXnATCwDwTEqC3lNd6dmECbHpF6kwO2revhNs
ezcXYWOUZPG0O1r7wA6ZMI52QvnkqHvP8soqcFB7ygaXygM1zb/wJemvqSS60mWc8NshAxeKzzwk
Hn8BVC+eZx7jgxNWKDxDe8tF8CgCJS9LwDsA4iaW3zmhD1axcu0iyBBm5xWdVsTageYYcNToGHz9
dMLJx5eu1AnruknrFELnr01NZt5AuF4neeTxPBJ9ISmrCskZ1pjP+P3f5sq8JU9eJuIJKGkYVc45
Y6OtabQoc1dE3O8HI9vPFQ0YK6r+YbaCCzwGE3nn79fMhvQO0xWhe57mhhXtCTXZXEG7hdaeu1oZ
wiaWLkHu8BLKmJhmlO6nmOf43soWk/JG3yybFh/xu/lqzZm3H6C6dTPFLqTdD5AwjCPADpuizPRu
yZdB6wcJYmTOENGBXZGDitaXMNIj6cRT72SviwOiSYADjia+QqNd3UsJ4LbAURFkP7/e8xF7sN+x
E8TPpkBXyYv43sJv9fw2O+8NfEbDCFPhUqoa27pcvr+OfCVlS/mfPhJk8uv+xCLsnrhAn0ctxgWQ
TRC1kdj5eOq1RUkeWXI2a2QbaoHdiULEnuj4ikWGNV0dqSC8VwQQPCIdQUhm+cuL2GMFfYCod+gN
FRvK+Q3w4r6a9VpgojTDH+FB4jSRIf1jyNZ6ewA/Lc19znBb9n4iyXJRu8XfL89Jg7PvUHUmMdyT
JBmjIhoLIGTP3z/oe72fV0kNuAZ/J1/aml9TtbF8PL+BvQsj4sGPuAPyvQeIbT75pymo2q8YpVuL
2QIW9GTWPyuCtNfIghnBH1sjiDeQiWAT04sbvi6OcrvYsFA558miv3Twmplw13gtK8xjDsFgxIXF
2egxD4Pj6EndtxvVUHj1aPN5b9KonRPKV9vma/Ar3wP3Dykk+fE1C+yf5HyTNsj/oUrC5v3U/dQa
zeOIQUOfc+SFN9DpLbtMX9JrikD8SuqGGHhvgGwD8ougXHS+iKNWsWRRZuqKxdd9HySCfKHX+3LL
4cQWDCbPn50IWWsb/Qz1eLx1m/rfF6zKRRHareEy/tBYQKkeeWooT3VHoLidyJhlQJRQGvnV0/JC
wwOV1+0NOV9g0YhnmgmfemBNUSxLxgu9PD1qSVHt3Ss2ZCTLDyn+Jc5OY0UJzqWfP3WQIy2azZuM
SDlMFIdTX5oXhQ/Fht6hzRAoSqD2Bdn90rpDgFSNJVN6t/YpZzcnyxhDjMngg7KL0P8Msd3Tq2Pe
M4sGJKmkE6AZ5x6W7vKi16357CXt8Njh7/wlGp4dm8wGdlIHc+cf9jw6lgdyB1abnSOU8l2t1749
aJefdfMxHvsj2GmSnxnRmcQ/ciVKuirpV9HGREvy+ch7IHzE6DyCpxu8c4pAnab6kMeEgQhbzWbF
L+I6leNP2f6c1IETyQYPA6hElzUPScsHO3ZkRJv7khGx3R40+ID7KvQSqNxtoDYpYwHe7/EMIHfr
Ep3EwspmhLvmi2Mi6qYiFjNnbuLbLiZGRkoCdAcw64RHubEMSRQCIkWGukYi/QCXaOtjTPFenOwq
E/Lw6uknSwMshLV889GSChf+AsLfJ9TX8BYKLSna5A8nOLiTC3EUsTQdeEqqm/aMOX1bMjWWEiah
VswI25FHeGptRDtR0cB6ml/heMnyokC8CuUck/YP3vQxddlpHZzMwowx/HlSMlxnZkaN50YEgt9T
rhgCaOWgv/ufQ8Hdovnk8BasX5C7hnfvBFH6acm1bVsEGvj5n3vZGH738BGbWsYpSsy+jG/FANck
M6q/QWhPW6bo97H502/4a6t2YNwiqiDwoJJ6lBld++caRSOIHvLam1fwzM3CzjggW8aMtt9DdcW3
Py6bL/CCZxC8X0YJHRNhfqPp11Pc/d2x3lg4ylUH5QDMjAIrtxVyJJB3zzA/LrnOPx45sAaq80wB
w5JVr0FiEHk4W0MjhUrOICTVegCqHHjVOpDUWn4zozk7shR30WGxIOlvI3TDmD2Mow9zhBLl4b0p
4fDaAN7+c+LIngP4hfjmOTOu9j0wcm4jgSTiE0IE7JpumMIaVlRIgJjgd2ux9o58UYZNHtq8heCc
QleyL46jw3r8cP1XgeGB2bNWM2XVsF9d6rUB+dleMro6m/xEjPfCOlsd5UHfzf7q9HMf32hXj7LS
vvTo7++T+H8Fe3OPcxSZ3ZNiszAU8rgOLZ3ghoauj2mBqujFd2T+r27Qo1IDvxZLQGo4cJ/ItKON
eZuDHuxXcn8St+w/cgUczByR1nkJy2H9WzCw+rsmSLpdW5U/TwJvGxYuOMhKG+cF74tm9eBxT3Y8
4EXyzQ5CgDWT5OnCEZ0KytfTjIbivCM7udg58OGtRm0SGFVR8ot8lqPuLFuWlKzzFhl+rid88WJL
0qkBk8GBRneC+viOj9NvNSfdAblSBxzrQz2hWorEgEePPbaB8jRXEsi5vgEGX570erhrz+e3NjYO
nUgrApNJnlBl+xrmAqzC6TS0aUafGa1YenIuTYlUQ85lhzV7xPYb/toAxmywzuLuHviGGQLq+9O8
n70GZh+ah7YNGUE9cx99zCUyYKhUDlsgDmq+F7Kpep9EdFNjrm5BZoakrb8I/rhSpTSQe5LRTYq2
GESn3875rV8K8iydsUR24fEYrwJH7KbVRDv8254HSnvBwd8QCRAJukv0aSjnhO2YzRHiqO5pHBg+
B0qlrn5/x4jF/4+54bV0yVxeCAo1L/gWpYP1o1Hf3SMsuN1QjnQ59MxKZM00SgzgZ9clDoEK5Vq+
eBcii/ElafL1SFxraxVI8TF/oW8pQryJboF3Pcj8d9Uurf+AT/K/46C+Lys3buKAnSIYdB/FDwAg
FC6H+w8Z24Chc91568GU2aqIkGeH+92LikYd3G/K1nwop4dO76CGGw2BcdaIdYBwhOiaJrIXPPda
qQIlhx22V9hfyJhH+YYoVct6Ic03JCeQJkgGnMIr+J49IocuS49FjrNJDM02I0qsLyaw2Poatlvq
8zRBRgBSQVNgE/3OSTcHVkrh3Y51iLg3cCMuf7Ypr454uqg0POaXfoh1M2DSdrAjWpEZcmcI6blC
nVZdvmjeyVXu/AGAY/AKb0y/vrNnWnoVZaiOc0Ttr/YvkMKykxBPmk/QO0H4rdrkuRd3r7uvqLGx
eOK6l2VU6V7R6RPvFHavMvQWgoKrLwmKTRQzjeB7zHjdHoC5nvtw1KkzuN6x8iFw5mp3SC1zsTRE
PX3imDJMqEJJ1xUk9prIg4m7G0NNw6ZfttGSjNMETm16EeebzDCrxKuwbuyBAzkzsis21r9mngND
SaJUOwIGFy5alTQPF/Cori8BQjzendtDIefdUW8uPtjHxM8GlpOo4ejclL7eT8tsGlMLdMz2TYp4
WLHZEZX4PT+34WzjXmLoKAOe4EcklDJFLOUeAoQ6WTc7aoV/++sD366QvHdvJw+Xjz6U7Tw7j0Ru
dp5nqVSLoc+1+o2sK6YN5wwUetNKK5Miyj+Mw9ko0/TEBjT3l3H18XUcho5h4iWK93n0S1r+mBNI
VGuDqMcYzxwqqSKx825VvNxuzl8yF2qmPFHbdqsrNAN9oNY+KMD2hdZKfAZvfO5ijoq/vTrgJHJi
vHIhebZ7glCw0DLWfE8bTge4muDqRVdWqATrnqp2GqlXI9RxhPoDnH/9x6Q1PtoGyhyXsdQESngx
jKD0pzRxVlG72lVoUVXsLeXKI3fNZ95v9MgZXPzD44iGpekorgTW6EnAhtyhDU95nI45O3+wvGTZ
UJz3NRtiGy1C2ryqSAC+eWD6Ho/zvbsBeD9auI+RIo3MOeOvRvAyQSxFKqjQ+xGahMCfc0PFwvq7
By2+pIscy5ofIhRv1x4og4G315w7EpjfCxDBPw/F5CEys6utjBvEXwADkvh7F+JaEBUk3FlxLmjo
4jlxntFE9csYBJDILnLG+2L4yjn+BHcxIaKCvKqZG/BfgZ+uy0JFxW+j8NKhWFrCF9jFmAWzouoM
sAFZoP5ykPh0Mr+sJz4rENJxQGlMfHKfp5OFH0HgrUsfm8l6uuGCiZ6+C8CNB1cogc7r6HWujXZG
I1teS4ihpkD4lp+iZzLw9D+Cf5NiKUpbxEdKGGBpLVf5DNg1DpWBPRi25rk2+eP6fp89ovz4rgyl
dyWb55E7w8jH4c7AtsvQ2/aAr90CN0SwbqA+eWbkIqak+MB+8VN7bep/93QBjUpAPAFpb3RrLImy
4dl8T6+TszdtW71jtPKVqscPvqUek3IBNltsardB+v+Sjo1zPn72lh1182CCeQcc6xoMLt0rn6bd
TVmxJKjg3A5uSiXUPeK5WEVR0G/vlPus4qnV/N1ddr8ww4f9wTMULfXjLHauCCDWwCMxM9uKb/by
XOU/AJsDZqzx1XraByUjtO9/YiUI59Q/Qwo/8PSI9QVRov6xhS9b03z/aJR56wbhlpKkYZGOx+tk
NHeuP+dPZbrJswrJxBN5zUhkbiG5Bv00Wxic0Gk/PsWQF9kmPNoFm8/Crpj3oQW81nzP5e0i5DHZ
Z1ogbzKTGEzVsbX9T3VXUGqdz4CQjquAnPPE+MFHbOjTABY+FiHHE9bfEXuNifW14Z6unlS3jQa0
4o5LAJh1zD3tZ2FYn8VMtS6qOsJ0WqheByeUJPY1/UWURfqh56qo4yraUELCK5NC3tYJDn1YNDKr
TlQDZXQS9JTcY+74+wqQh1tLrwPoMVsqDUz9AVwlNaONA5WxKpC9bk3XKemilvMwdkx92f3D00Qd
n5CzHZ5bYM+p2cchnquS7v+Dxs0bznQEnQu4nei4ZU9Ido7bbNRO+ub9gwnokQtQ4weA2/4HDjX7
QAZlioqh87FeGZT4mLuBNoNyyf393l5H/b2ogKYBf3boO7it/Q0srXKMMjN6luLZMYxzwZMmFysn
6+w67arOHw8pCkc8htm4hhXQ/ciVnBg81t75fXLDhjkaekaWBfZUYC9khZvrfPwuoWwdh0RrQqou
qkrBP8Cu8cGPG+rOqmxSt+9wwuFlNufpBq9RkDse71EulndC4gCyiV6qxmuP3gtTE/1yHexx6AIk
qR1uFizHJaVzv/TWM5RqZ/3jO/dG1D3PHHQfByXWnbRnKxqaG16nOjj8ZBJVIEH6tVexRIkT+XF9
OMth9+//hSpGGPnrMyCpYn9SPXiViP5CMw484Q4oGJJ7AFodTGXjfClvMNZDM2vCtrUAG5gPctNn
FiShfETYRyTNCuxTsneNprI6O2V8nuefnliSifoyJsXHppl56cMLpUpA5MUlvNqCnNWf/Wr3nowo
Dv+zQduRhsldedF32vthuGffXEBZ84QxryM7adZBGo+DQv3sV0mzhhcU4zqK8XD9m5j0mElEkHhv
HljA8rDXejKC0voxbQiZVgNlEezKMrXSTtuSNLA+MnICprH4+Vm1CbjHLb5V7Dy/SmfE3A37p/Y/
ppEDO8sV1KudHnHYzWNpaLi2MiVOSn+zqTs06RwhgDGwWz9AACbjRnfnwcP4uP9qLhwGBVTeLYFe
zKn0OVeAZO4QrZcathhSvsm+NntWbNOk6ZJ7QArObWDRSoJnRo9pnqp761Q5C1wPrSS4y13PwOXd
5RM12wqTCLEiu8zxnhk1jJsBFJqU5wbJfndyVa6CL1t5fgU+/6td56wrE1VTLEuSf/Ei9Q7lZkl+
Cxc5lZRlABThT1cs//WhVLuCCu2vahAGOZB27MQ4EM3en78Eu6rrLYqc0SuJrXuczTlqVEZ56eq6
CUMuNgQbu/ItADNMqsS5qbVgm5RL24uxnSQrAhSPS2t8BOF1iLGOiy0kn2P0+90xbft8hs5859Tj
2YfUizKGdWSmoyVAFm4riy2ij6JsO09FeWTsEA7GnpEr1J99sRJi9KgNya60npK10gM3mYfSkONb
VSZ1owH+nN6FBwQh2ftaWCNPXTlh/J+Ac0e9O5E9Qqs+6h5q4p0njUH7x2ROXi9k26b02MR4aoSf
A0W+QogvsIYMK3qCj8CIzLh0Rr1MJ4d3LbEAYs07GAXNFUtC8SQt6QF7lXcXrU1rYxgPo6LlYvvU
ITg9iwfRRY8wTuqIrunIer9U5hbyZpdEzpk4HlDC/jm4J9ldbEixwe5wru9+a80qgZTMt2tQC0du
JWRimCruS+7BFJPVu7s7EnjRLmFCGK8f76aPh7OOvKn4I0ViTjdhGDjRk+wI3xukIRCSoYhNiNNs
OchApEB1sGrwXcF0dVSmerS+G6OZuczB/EWhU/sk2AzIzmHGjwgBby7S1+2Zo/SZjJP6Pzk9lLpU
a+actu8vxwCRBW8Z7uQue40xeRogPpNofsBedop+fbsomanX3d6HTAX79zasBPlMg5h2I1uqFNqN
cCvXIzQRrIqFOGbdJ8c1sdhcVzwWloEk1XhMTBv3nLjgk8P04VooGbZlwH6oLNZlCBlTSarKW2h2
K4CoVHUHgbFdaTVCuvMSzg3/8rYVAUAogT+XuSWfOTV3IwoUUjVDoc5y8fTDYpW3/LkoX3QgKRoD
Vby/0GDijptc4CfevHnDitEY5+2citvruy1ZGDtqtUJu/tx7CJdr3tLtXeRhdzYuuAvdfu1dExZJ
yjwFa2PgwqZvO2VT1GHSmXPq0J+aOObeaQ2cupV1+o1tvELqwjqnBvI/odQRmE85iBqvYwaTMCzD
yq4uAJ5OEDjvevLkljhWxw3v0TArQMK9wk4soOvGhAUxiGHpe19Tis4V+mBtZyiHU9VtCONk1mlL
5uJcbjcO0LcgTiIb4/BPBLX7u7m6SH3aaWY5SNAwh1LnKLtTa80PswC3URV+NnvDO6FIVcZcsgyE
bEc7z45cf600rW06+jKxbsEHKhj56x4sVqgeS1/kDugm46l9Y0LlWvXyGLyswvqrPW6uC/VL7+VN
BHZaklir+9Sofkc0iYccUPSD6xoyS7r2ukYjxL5q1c6FPciFLQypOMifaSb9qs2soVcQN2d2tpv6
4oqJiX/4pppTPNVrvHg9PWDn9DnXdDE/d9J9qLiDweQwpTF6L791gU03ht9ONTVHN1tquQ76plWN
L+YAubOsNhbvLRGUnK5379SHi2oP8UaIJA+Kqh3TkeUcm8EdKRtrcpRyRoy7fBTqE88PBn5sd2dC
tPWCgJz4u5rFUI5Hipmy4gjbanH2ayKWmAE+BrUcwApr3Z0CKLGo8ZC9QPA1ardUVeEUmaqc2wYN
pA35rpp7vV7pUcMyOYy5ysw5Oftyi+jkvXGoewinW/dMq3RWrKgyAfxJuwswWkMY25uD3M01+N13
Yz6n5v1Xy4/L3MiT1P0FnSHNrjl1Qo7971/kd28BzrSR/iDawHlJARHSPo3ZkylwEBCVEBy38r6x
N8y+Gp/oVtNpHxb8cHleqVrVISBan5NBbZdM9D8pGfjRuw1EXmr7p86NfEv8DUFDGdF0roFn3pD3
CtH4cHyye06klDEAOzgS3u/UpKj90Jqv6EB3hV9mUxMGxxGmnZGDWoMNFttaZaiNOQ0kUpdGXMMa
txOmSslFBWAqGU80YeewOnXIBQZ6ISofBnw8IhhQrdIWp5Ipopo5EW3vTcUFL96zB1LhllRabqQd
Hl7bPach92BTTM7qj2n6heKpBQSnLeJa4y4AMzBDdzhFOr3jNQlr4I6fGVCc1FNigds2GGGnmrSG
X5w9RmNQfsncOMOyCiRNN++NDChIP2XD4JQlmVbmqqD/kDXdFhh2WtGN20LlJcpv9oDB7iMiuES0
EhNtLnGKJSkjZC4JukoqA4IpezP/WZPee/FlejRldDC8GZRbrN5tz9zLZ6TCvPB41dgEIXvkfT1X
ePmyNX8DgUYuOD1I6c3O6oPd07oRYPu0UJ2xMAeUldcagBNIFyMzddU05ggEO4s4RSa+UR/oTHHH
5XTR5oqgM8Q98XeIi/h1BBhHDrUm+tUbO5nJUIb3OXd0erAUQ0HicKBGPP1uVa8u4QeBNMhWQ8EO
zJeBr0Td07p6XGE+u+6e4tfBNRj5+R8yimKNVBWBDl8DImC81yYtY9wiKpBx1HielwjEDTWpT2ZG
94WJid7ndHe0kk+yRDuWHI0xgo8ghNSnonw+YxOqAAElv33eMJtOFhUe8/TLmHgN6ediuODUT4S7
CQHKYe4Obcp8IGnYQvWpJEQo1lsxe5HiCfYkAkhOTapgs6nkbnSmlYwd2at3hQFUcpJn1vO1moF6
OrV70UstZ9YPOYTpf16c1ZfnkKoSApkHhm00D2NBD5OQJrPH5Hq9CDlOxVn931EfOjzTtmXKtksc
eOnRd6cump19Pd4h0pWluVjK2zBa9hP9vV2HkhoEH/OTn3kHPHEe+ZXGB0TqQYUZPfxvFQqAL4de
0vtDwiy6z9bbsJaB+t+Yj2k6rryiTTIA4s9O8rDO9GlAtgkegiNtzwf4wtMksbYeyJmkwniXYRxr
xDdIFyjeswCRrUdRJ7O17u3AE7g8O1qysbKxtQpVApkTcc1m53qT+iWp8ZnrwpprO44Str5Q9Qzv
ggUwyY4Qm1Hk3SVlOMK8gn4UfqaAr7+EDe4sJgYFNhBVir5unk023owFy5d3OMK44PSYT2g2jn6o
WCyrQpOsOBk/zqQKhD+7XGWHGvwCtCIi3mnyz3iRNse9uS6xXPRlDvbVZo/I3DdKNBnNydE4gIjH
BMgAKzL2D3bhfzaZBL7yVCD/+UUNIRNPc80koN3fF5u8TFHuinJJYIEAF5a1nO+8zxYH5sGOdx6y
eBtmQHQ0uY97JrM3DedJLJ8GZjqHgmw2paVaL2Wsr+730g/6b9EFgfHfGLmZHtq/yBQi1XvYnm4I
h0C2QjZAHdTocpvitXBoWOEp53RBToYsz/HzBKveTs0uhg516bKaGmpMwXMwVpvh/CCWg8cVAHXB
91iz6lRmY/DR3X7R4IOiobNJ6g6j5ucKeBBjESaot43OBz+8ei3xW5c9TgMDz33je/142khzjFN0
/ykh578aHYGlcDFaoSjEGsnI3k8ZM+gJhMK1noqywqoe5MIpbKQkzbfyKlIMk8EgeHlUUayBYj9p
hCfvQ1HmAJniOMplNjgLSAm+VKnYBlL32jT80R9/o3oCUsQXG06XPwl/sl3zJEf5uMvz8qLiesxT
N70rXFVy1ebFWrEKXZTdGL0Tht3C9oVly+w4VlQnzTLI/8VD8u0Zr1r1kDQNE4F5KEztpSvcCiVe
a5Isqvk8gidIkV0AVB+/XYV12EpSghp0JSoKfjWgoc0ZdtE7xTon37iuy4mf595wuQC/E1ziaHto
ERPDO/kP2kZ1J0TkIZHkGQOGouZfkQWPJ+G21sGVFchOKng+oY0DH1A3PQAlR87cuxeO9nd7KGM9
yzWhP+Sr60iwZ6zbT0FWbN0jDAwSrOrE8Et3/rNl7NdfGCTFLNVhSoLlDCdHReE59FioYF0STw2h
NN9Ifl0t68oPVwcfgPrgLKyAwm1fjOHCxNG0oNwZM8Zr1wqiHO8K0tpgNHlZOQgyvIjxv9D9HvCP
SBUCOsww98gcVbya04RDYK+XQOolmjtd9l+ugARR4QxrVpmaydmrPRfP/hz9k4bbtiXHWS2gVum8
73MR/l6gt6GgAJaZhsk0ad8qS3QWsGhrYZ7S4GOmsEoc/nvags/PvpuyqlyusfcA+Ne94Q9vg1RV
RG9sZZk+y6X0+c56nKHlIh8ymoOgNHt80OA6bAQyQiteUwPrmqIpfIzCxgiZrgW1MCMpG6zRB128
OUZwFnXglvyMxCmq3I1T7hUnoZnaD7IC8OXkZuqjaqsTlerngjCXFYGqrAik50CliiAMuQU0IIXH
3MTZwuZydE5hOxWcTf/6NdEn7s6CSgM6/x7w5BjFLVBWtkot/x37k+NsUm13YNpCnmQ/1e+Yp4E0
aoo6QThvEhZzpMgCoOGP/shr1VdEjYLfWoqDb6HJl+73FLquC3EVD8m4OlFMDdWXP04MrkqEv32F
7HxZNxdJR9x2ON5Ev9tZTf4jEqsmLftdSdVkD/2i4ipnQO8L/itOHy65OYiILaDJ8AHLhnnDA1sM
f9cL8Ima42l8yHM2ggkBENCjlaVTrKZEWy/QNBCetg8n86OXMlrliuZkp6BZ764L7MBDIdIbmQWo
bz0iDTc9Jmt0k14HSHWCY6aCaZaQ9JfBZ9bKMpBQvEWe5LNr5y1ai79Neol+8ghbmqBvy9CvWb7S
AwdNAdVO7Ocs6GjRlPMefoP4t6c65hbQXHnZYtRZujzUBx/DfPrJKMoFSP0FxMS29lgbSx/6k9fX
Wxu5vlA1Xo9KXevAinADv4rVOQdQUizGiKQhQd3DotD0g6r35/EWqixFML9kH6gn5rUj0h9+EcGv
hoqriFxEbONqsXXCYQ0FcMwuzUiaCzcUtXTn22czekasuI/7ZSdB0s0UupttN/QeRlWwbcguSImM
j7Tl9NPU901cP8sgI77t9a63CcdtTkbXY3aqT0J9Y8l2j9biwMsFDvK3yG0KvaNEIg+fz0CAulOx
weeGgiHRdh/AYJB1CHcdCe9dBtMduF3+Sh+tYb3FDUhaNHF9P2doxJpuBoYYS4FvQzSODd5LLVSR
26Ufx/+zyrzK4BKHyxJ3gL3zradjCp3xounvtSehBy3iYb0zM9hGAasGnae3rE5uBpmO3ZLbMPom
7kYwEOtl0e1uml0G2Lt3z3y8JihX9IMJPhgr3x4DUtZ9jIfYXz0NIkzD06RSScazSj/AsR/izPF5
lJOPcXPYtI7v7wtxS3jLnU2kJQPnQm9NHve11xcrgbFlfVqYfEuXOkmnZb5zYWShiwDu66N0wVbc
VSgnEzeffGq4X8MwWo/b73A/pa95HgjZjZNitEVVRNc0MRF7cJvhNhAkIhZib6AzZDBLtRS3kCLP
LG+Jzxfeu38YjzSXT3DGakXv5aFQltlhLcu9bteAplyD7zRF/nTC4En19+WVko1wHeM8g3VYrDxq
L8mdZ8vlwXDqs6cnm2lS+JETfWwDez8jKiYHpsUbr05kfTkaMfeKoFdMYoSrmnsYbOB6FYOrYVQd
od219OSO19hyBU68iPxiVJCxhQN6SxyhhR4A8SwNSykNO7LlIWuv9owLTk2ZHlgx/7mqg31Acu1H
GjTphPGu2ecoV9jgvvQQabwyno8HEOgtcH2rdsjqpFbZBzuzraaCTPR3MvRZYQ5l2t896Ul5Hnm8
xIHvAgUCs08HoBB97n5Y4GCAvHzNfknwPig0h6ixOrmfuQ2IHPbzrcVbDa7gmby/Cy9XUzXtVoMr
F7VoPMNrMzEi6xMihKSDix+pgHMEy9ZercYZRtX18AM38WoCTe6SKGYtEZni7t9hLSyMcFqJpwnR
EOu8qvXltr8UYtMRYfs1lLKV/nFScBrFpG1ozF0TptnHdY0v4rWM+7RJoccC8nDBX2ZKEjn+2WVr
3EKiWzueGuckD6k3O05VJIik4fF1IK2G+lmoZJ/6dZbSr3m9ZP9cWZikZUy1tZI+SmsvGlX1HTrd
t0Kd+qqGloYoLnpGUCT5pIuqXgPA5WVQS7ktWDLFTTGvgiJxy7EN/AmsapRkKYvfNoMo8anIExvU
ojgj/O0ntrssJR2+gAgr84QbcDvghFSU0fqmgxmglMhfUywlAlVRWObZTl7MXjL2hqoTLpRjJJeS
BDBsAgbFvinBxEOAWUNsL1DmzGkv3HZD66pkXyOY/0z0LPWaDPJoSjrHiP5d1gyuJViENsT1B1jL
5CYu6bG1lnyS/jmY798y2D7vSSjebYye/5HI3KNHjC7KAFjNVfzz9iobKURwiFvGxnASlT7o6jba
gQ0mH/Mieg0kA4+hUVI1310U/wtRjKNqow5sjQgG04HDeswcE6YX1SgdbKP+RseU5+VgUKh+nlln
OXejNlxa+5dHdlbej8uBxfPt7jaxdbrpjn98ZHR9Z6Ji5hbJtGJhGwe1/klefwtsECbQVl0AWdX/
SfEIEGyRXNEP9sRxayngiVwFqGeUwqllQaY9f6PI0SchD7Is7NokYV72rBjQncUJ0AS0/EJbuY5U
r3EYdRJM+L9F2vqxWY8MDoqlwtfYIVbak+8Zp2oFQP+M+Ki865f1NM2DgubXWSZaKbRlWfP9rZ9V
KzxHRNVg0+1ZLPC64QvjxxfbVc74W/i+E7sU8HwUKqeLZUlU9XMsrcORfSvbcMf6FYDPONAAJ6pa
mPZWoWdxUcDumr9lAMhMAigB13r665DJoLyh2mBNO/XkOynDSIP3rYrsNKF6eX3P7UeWYrjpKE5g
oHHybOqbUKYbKLPIQCQ6489G51mJ542N4R9CHsOK0oRQMxg48MmGHKF9HwoRkL0zb8hPpQtSR3S7
erf1xKKBdruLQF84UmEQTOEexBqhnIDl5qkJQNkEuFsBYduul18qN3Zmk1jmoN/7rVg0wJVovGYd
Fdi+mAE4B1vYSYhQQgGvmxDJWc9nrRD0luVuxNs+MHiTBl1CVqf5Ds88jHuAAl1EiVxOkxN7ZYaz
RJnpOuqR/copurYhJS0kF6sYIvMsR8yLxufUWSCd/ydra5hFuDPykoBHRo90y0+/3Kff/kAcGQ6o
bedweZof7CaHh7CivdYgJZpw4WXC7jTsE2FZQsRD6W5ayPN3d2H6cBXQ3HLNs8Hlh8daMQeLcM1x
RtLqLON0fWz1AmYz1X4e5yrhHxdztbVseCOAKl2T/DM3t7MIRPMimupNk925xxwQIZxdPL8zIw1g
vbZYmiMyu3TECX7Xbt4nqQ+/PFsI2m4Lyqos32fsqboil/QZYo0a7LhYaQS1cJXhBcXNwfqkWngp
NSlnTE4Q4VRa2wFx29IN4QWtmwTYZ/3Zr4vtx6lMMna/d0B+Mu0Pkix7bHAcZIOMhrlOld/cQLFx
0SxzRHDYsbrFk0Sb2MZx3GoWojMP0RPKrAbwOzvsXC5yrdeUwMdyQCFT1WTMngclQJXyYksefYNs
mJIEr7xGRqtg6kUCsBM3wF0vZI6wJMHyGvUp+oGxUpW4eaoREBlpoNVGxfWbdSyQLFRzi5E4HlCJ
nPBHHYiWhylPIAjYC8Y1cbLm/XKGpl3W6QgHmULgL9H9FN5Cv523HBR7xHJmCT85K742HKtGvWb0
CMuumecWUpUQFgzqdbXbYTZeqldk96QLIMNHSKFkh2ZOlaLRlJy15fYDDCzpjxV4x4E2590ddwwz
PgAxBYDJVovMXVNZvp16cwlotU8dLSmBpnYkgn2LrTEJ4rIPpxm0Ju+efVCyWs09e5HSvVpqH0n2
p8Cs88uwqc+WNo1+ACPYGwx68aqecFgE/aWB0eHh1vP3yslvMs0oYuuB1ik11ExNN7B6snSOGO3h
nJKDyS5Lfv2xuL4qstwqAcjd4AvZXsOghc+kH9Nk7zFh+734kzCPVA9vT0aWyDyIn/L1MucNNgDB
rhAowiGXXhshoD1yaioK/EcRVi2J8V7z9jweXprG0sJyLkPmrY1aMbtercoq36tBCWlSETZe9yUz
aAgxL26wE2QZkT5i6KrqhxYmlZRmPoNvbGP414fhavV9+NhKDO9zo+WMcDwL8iKb5Z66iyqCvKYz
PkP67Su3aAU77qIMLA4WoKm8xMjBqpQWsuxwVx0tnVEr5fAGLVRoZlQNV1BzRXyawcZlCbFjHTIo
aR3iTJllmUtQfiFB6JDuwonC8jHvFuifz3xVTnSLBHa8yDPEsyPAExNBsOzkMo2zxKVUhObzu3wj
/2HBvLbQZa3ouU/08qqUbuusW22HV2KfK9wH5llBqylXmje0dTCq24XOWEvchFUgtdzSSkBlUdZM
RoPq7Y0PHz2iuvSTeelYAD6FzLCURopAmH1O4mY3vP+78mfnVH+vx9ywuDGDyxUIItSRD5tjFqBL
6mZjlljpZhnK3VQQxKoB9J15NLaJMwwohR6a3psNrFyeUg18xirrMEVKQ+uLyTR5TFvs+2RKVgVx
L7OtWuG0zQfedSCwxw8605CaojD8T2Cny2QBLi0Wnrxkg+p5Rs011piVwyRpwFRoG+J3ZqQ9/L8w
kIOlHPICwPHwZ5dSjcyrsKTwBuwY9AWElDQiAY6Rr6MjzbJC9niqiUMOqLNKtsz3mIVl73pGHP5G
Xht8MKrhviAG/HZa4viiRzhYBx76pt/2DkfdkH9XV6ZJ0CCYt0p50Pidu+IKRHy8SPNHzy3SDd8G
XwJUClA+lbv7SPWCpiWQpn/H2faoG6uacl7JHb8rrtdk+kMsAp37MqGS2YC2Wpz2bNKqfsf25MOk
v5e0CUlGV0PEDh8OUFUN1OSCJzpWFkjeJwvl3vzyK1YQ117mvRbnHPDwbH9dD430LQjPSwKHeyd4
Yg8LcB5zZz+tcBFewxIVHFg0D5PxMU24Z95Ot2Qcb+N4EQOBXysHTBZpj+9q1C6YstyvYQsKIKrg
yQ+f9wwRKlJnfpbIEISm1t0xFaTQuf786FUpcOSMTVZzfMSEG9DxhdO/eSUr1mi/7Fn3069mHnyD
/UOtodE6Ln2XaBwefDnVanea2WHfWX8HJCt5zuyoxNZscPDy9+lIAc3hPg3d1B5v4PxPS+P+Ei60
cP77UBwUYZucrZ8/EHl5K1LBys1wubszx0rrqBW7Vqq0Sne/d8jSrtKXha7Jc6xK6/W81MxoG0tC
pgAG5z4O+GaBhc2QsdAex4/Qx/b9jG1aHqTmKi6tYgk+KxoWC7UIowEopfv2NxAXxIKDfEISNSyY
UmOeCR6STvxCOLVgSW7a0ewENWy16O47emwa0Y3bycM3C31rRBvgtGgNS3Jb1P7mpzGrQJZCMx6t
+zlGAfVppxW/7qGdSwaI8RibcyhAl1upOA44EvmTN3AAbcAIEBcwU5zwFyX95KdAapcOVOHhebII
l8RjC2O/62oMeusuRD3V04MThvs7Y496vE8mB50F+GAAVQnBYMfWS3Cnk5lHujkdLQUqqCM9Kj+t
O4FfAfThT5Ud1Ly1KDKZf3IpoAeZvJHVf/fkLao5tb6gQ+VwFjoMZjhyKen05mVtTTpOmp+hraJ/
8HdAdSkmvPwsSLM25VHiPKH0Juv9ZsN7qScULT3de1zvI+6qkKm1l3fuVCh/wDbEB9bz1o/n5KKV
elpl9+7Uk4TzJMgvuP7bwHYBXXMsNX/chbVJ2/cFAdvMhJXOsBLCDKi5IfwAMyjJygUIfyennnS9
b0uh3Mbhl6NXPrEe/JPpfEwu5gnUoa1OX96fBbfJTFceMu30vrjl3KEDYrE8WB5G2T0ozYSpeP1+
0/vuG65tLSSLTFY4tHHdTyTnagowPyBr25xvBTOTMMp5EnFO8E3miUFx9A3yXWv1mJkUkmFujOQO
xp5tfBIImN/3nkpJUKBgK1qgBbTXIuqJ7ra3cIaafzPRjY+dBiPad47uxW6VaWlaB6Ad9a3CUgO8
y1qK93zsuBDWh5uFavaus8iFTIwNJqbPoe3amHXbYUBaCRYWYr7wYww1AfEAeIbH3a4YFJHhphew
y3u3U85XzscSzkiWDDnMIc4UywCyHKrSvvHqtqmOfFIYSC/svxJogDTd/+jBScvyxMtIg+Qvs/qE
obAzUYZRxBbf6KEBn41nZkczNI+n8G0CdLMUzdyVSVFlksGq7FaPsHP1CsAPvHpce0cF1/laBzar
Ajr/rGSZJ5J9PW4quvA93SWit54g+KOmWIBa801Of3bW7ku3lYj5m/sCFIV5uEHK9z+WJnnygy98
fxm//1tr4AcPFo/54epAXh5EohFyfJIRbQjlZa9CPdxQnR2p7pR1KW4Cr3nn4Ap5vvoIVwk4EAUf
9EeeaYFcX2Lv0zHs+QQ0FMwio0trA/zeobiQtCRLzXiOSi9Sq+vlb4hzuW/fO8dfWCVh20ryjcYr
MKWH8VPx6CulbXvL0ZxkyJuLbesNWBhl999QpCncYJ7xsXBOzVEKB99KFc/GuZRofNkDcy/yN8u/
XXYIrj5KJ91EmmiOnHCe+KyqA6wLXrCW1RlkPET8HvFInNnuXAV+Qn1UlIaV/NnB+4ZM7WgT98U5
3pQH+irGBsN9rgXBkKS5j1clp0XzX+FJS97Yewf4kLnHa5J4LuKtBG2FjDpcnujaF5AD4uDUFNPP
qUO62cKYR8MoSc/d9YycUku+jkgsJMJLwvhi5IfFrWsWO0jPgVFrkcoPWevJJ5ftfd8W189gKlvN
06NYP0C9z5nG1sKqPA5eyjedqAXGYp5xv31CKy69RDAtgRwgqQP0QrCzlR5f2Et566YfInS22ak6
AzcrakXItF6L4DfNpqxLVq2Mca3uuhyRRGwHpJLGh7Xqy5fNiIpu6WGYh9/bo7iF9GfcblPI/Z1F
PuZ3OquB+yuUpJfpjqA6AwTRcrO76w36QoLPQ8lVNE736rvSOJbrKFHwFIA61IRQknQdsxsKVgR1
hz3TURIvz6Q2W+BZ1h+ehxc+Vj++cuogVjsGTAiSUanwSj8V9yZTdbPbPf2+5K0AdhE4H2uR3vpq
RcfGtIoqdvk1OEqtr2+geahqxhsXmQ7Xs/od6SBbg3/LIcUHwRxJi90k4ozbr8uDX2kw1PkKC8g1
AIEqrdc1rhfTQQegM1re5QuVgDYqv7FesbOSSl5PI7+5Pnlvh30VP5572sqez7hxgT0oRMzUr2VR
0q8ONMqSru2kRb2MA1wCY8g64Wnvp6y+py7SFWPUU8jYZnFQ1FtwzSQfGlIIq7rGKl7gkTP0/oT8
5qfehkWvXh2OSp2JOLOttYj59W4FgaSHjGPvfpIqq4NVgJOcYkOpBSOvpJF7TSQDahonrGbA558/
3U7nRZOT9rwEup7nJl1Xg/UwXqSnTM2sbmyE8+Wt8MPViDQjgJJOOMi39uo4GPqgWZZXWOm416ne
1afbodBrVDItwXVW15MoUPxgPBnWPAw2MWG+KLQ4CpyCrvx0rcXfni/lCw0tvt/uAbIbItWbnIN0
VQm2584DOWuSDw0QRF0EcSDrZ13jGcoJGaTMzl9kaAX8XQjmYu9zKxUEMzutBZOqU6eAVv67XtQZ
Vj1X29okDwCPi4J1hr2P2ZKwezIZeugFN7lyBph8IxCW85T8aPsDr8M2Cdzn4+qENHI45bii5ZTU
JeyTLF373Vu9UdVu9VGq5aFaK6TKSyQmtL6/nTyWe1ODO1B+R+IuPU5b6CZZfMjtSWxsNbKEZVPY
eUURCAir7YpQ8Boa7tkJtIlrB4DA2sQLZ1lwmHIUaLG0ti1/YVsl9UFIwZWCk49UEgvcbZZEnD9t
p4LsgGK1ol04+qmyT0jXNOMqLQC3YGvDpEEYvA+s5+EFaHN8Xxred5/Ig7Oe+1/9WiSAYCTQvEDx
cvRNd9paOz5CONNeceNOifSOAquJHzlSlwLfCUEidYXIuN1AG1+NCTR6nNK0xvSwzp7Jo7ifSvfH
E0Us4+2hRInakOLmNSC+SKSsRGuqLn4oKGJdvCBHbJ/8tdBc7Lw2vNgByS9XLeZF0wJ43xikswdp
S7D+B/4YFihgt04R8K1fBY//02DhVV2VwCxD5req5Pk3tCs2iWx+izz9++TWHUgl4ul+kxS9CIc4
ZT2Qi+Wb1+4vrQqglxX1rXsWU+j5x+lI0J6t4m26oxhIARjInzKKoQYfUA+vjaX0tDyHs90lpVeB
vPehF/XFeQlTS/LOLKMDF1si2CRY3sgziD2yY/HnvFXYLeNtLEjxoSD7M8+3tiiHmY/zXLQHSpqb
y6qPxT7ZeqwLcSr3C+JHgpUl6FADCGyyo+pmmqE7O3OFbZu/fykaHwoXB/DeIEG3v9p4XVc98vz8
J440YB+LmKjhYtXForhcu9E+6Idy6p3wb/I9NYexolN21DJj4+28ekPGl2Fe/au+hR+qZu+erWyF
XK1mI68W3TLIJ2AiA4dfn8AE9HCDzyecL4+c2fSbfRz6vZY3ssu5GEzASUSToSuSCzb0MFJ7Jtu/
fGFvbQMDsx3/OvKACoi47gPAMPmw1enwoFyOCB4W/TqRNNGSLY462i4dT/hDbF4wf0K8nFH5+d0y
ky+CNf25rW2R1JrskQFdUeQN1htkk02Rz6VWgedbotdNx7cryIoaPn41yPlQ2hLG9Vbm7sYHcxnp
qK5MwM8bH3avy45bneLei1ZvOt7NWKx2QzVjifTB2ihI8MivqdNLJvrAc0mYHmpOoTuNGuc/qwmz
vHI5lbLVQkRml/Vq3RgeHd463zVuomdw9DyOfrf9Nyf4BoxhUVy3/wCou7FUm7Papr/6yTChj6W5
VM8fUk35T4mPFIDIpbGlVawhkwmztAnO9Qzse8eqvCvNkKmRx2dZ0p4LWM8a3L7iSF0aW7WRnsuf
86WS58SFuF+SH5xkiUHvkk3N1iznRXdRuNkO/eTi+/sUN4IlTCtWnNeVqScwK/C+ukp37npFOQRL
vsqGyXi9I7pHS94nLYRnsyIEpurznrgEBQChRlL4Xayd5N7N+PZMNf2QPrsKbQes9/Bn8XqjP/4t
7FfhQHCP4IMSUtgmR9X9Gb3Zmr93w5zjHVkl6IUHLCs16vrGyVGRHZV8SSVwAZdjePDmHCJzJChf
Wpa8R8DkLSsp1v320j4ciw0q3+Rnz29tIQaMio2J5T5NK4wS60yLrlifRjN1zIiYBi4NPIDEyXEy
3Afz9rzzqLp06/8KbsBdh/yKNOKyVaTYDjPpv4hHXxUtPGo6ERv3Ee0b69R9Zv+PDWDp8eXJBZpe
bP+y3bqs3NpwuMp4QAJ6+kQJVGvnb/beogbf1AlR7oxMdDcWt+dws6pJEO+Rxmw5x98z/2oFm2EN
ZFVFrupasMeyeEC9hTPV72fv5kWhVqaAfsM213oyqm0pdSbqvSgQaJkigvEAG5m0Sx7PKkVabP9V
LFqdxtwEawYJiUdYqJSfS7rcTM2yO7ONUfZM87PRBCekA/TcDJqo/osJvPJftkwxca2401Xp+wiJ
qzsUbixjQtGOtSWHImqs/WylBqzLjW0MFnUQEM5+AZUianw/Q92vZJoS7E/dzct7SPmHpiYZ9lZe
9+mojSJHUfWfPnKX+yIOkmiezmTT3GFND3CXlfjHsds4AHpHvp8Hi5GnYbhnq5bFp0uSfbxvsSuR
PMKEMfrRLkPL973SJRoaVsjziEFkMCyq2Jad5HJFD52GgRsVj+A8QNBV8XHHRUXBDyB6/1TV5ggo
Xs47bvWvMgeMI2UDW6iEpLO1DyKjUIHGNfYXVcWIHbg/61jSKUXJyA5K/xsW3CTZNip9R7mpoJVS
y7GchKZInjfWE+bEmni7M1M/BeAlY+8/0ryfejZ8Kyd2XeMAyUkW6upqEFg85HeAb2RQCKbOzYiS
2IwGWPkde+uA+yObnkhvKDpo7Onn2U28PcQEohLiqUnMCUT0VOqkMSskcKYPWwIcuMPOUo66wYma
mrJdayexXdC3j2/AQEbFESnzdiZHcSuBMZJ9Qx6HvxYoZJgW8pqGw7c1A14AbzGP+Y5UBvUc26W0
J31HjmQYIdUsoS/aLeOScm+HEM7VmHbr5vuKeXRImWjdo1N25RnDfJb5Fe0UnG0QzfA2NxFrf2yv
ychICyk2TOwQYsKP0L8aGnAxlRP/riACY5JHh+mfI8O29OXtjy/jfbNbYvuNSMYhE4Yvu2hiNsDG
p3z87imeWgaXpKEekQbLAoJXPAMSqXlWQ8fhaGwRmcGUOAFCs4fs13nAqee6n/usoA+61fUPjZE7
YcU30SY700VMON+PUgwcdBiGTHM2fTraeo8+D4sAA2451TiZ+pIaQ9Q7ii6WCizct9ISEzJey29M
iGiRPRKzz+mZL/CTrRydTlaWzy/EjskyK+oENcsuBud7h3VhCBQL3fvq/17HC75xhuIpG5prr45J
zt24YbXGceNZU1smuevzCw3XJzq6+oBQNB0aYx/ZOURpmaZG4FpidalGRrC6OoGfkGJyWp4K3EzO
cyoEZD1/oDM3zD08+ZQD/2NoxsTmV7oP9qbtf2ZhmYm3FUzjU6JjVTxKvvPFfnKBoHR/c459WrRb
Efk+Bdbnyk9lW5Fhw+DNRfqrU6Uvh0E0M4BdD83FQlmKYZaN+YwjIYxXHqeHLkO/UJZeEXRG7K2g
oUUoXepPhgMkQPMrqdz5Rug6eRRHcz5Eyh0151SulQeRFtOOEUAuht3eSrNUXUEzr8VsY9p/Ktug
H1hUdlMNqVrhszlhX76YqSqg5JqD0QmsvliMnd2aVuFR53BrGkRmUepNNauBfgaaFen0a+9kSSdO
7ESDdg4db8pFW9WPaoe2DLyMy9Ko7ndHIPQnTs+A4Soi2AsGs4E0OZXdIPcEVHslWnjC2CJ38QTe
FdYTYf74L5nU+3nVzPUgBnug4JRd0B6g3GDSmQLIMG0koFhFfINhFGl5BnMrApAajEAqyy9bTS77
jMr6POxOpcDyFiXguVO4gG0IWNQzmHsvdhA4Q746zp5wMt6DOdZCyH/iPunZkC2KVNSEdwW48knG
0Uxs/EvN2lt0ObnmL49CJEUmcfvPhgaxfwi0RV2OOwZHFTW58poOMTM8ttyBvQdsXWlD5s9c0dwJ
CXFo6xXqje555h3rnZ5wdfEKnOKdItpEGdm5r0AX0oZk1r8UPlIsBjaPjro7yTynyOx3ze66XE6m
x6Wae0SE8v+bq6o71pBjoSskfHKDuD4tsD3DYzZRqlUrxfEeSwGbUFNBPEqBya+wPzjh0Rf4HYTV
4wcdi4N/QKkHwV6oK8Lzr1Onb2oeFUHeT9EyBuph/jPu1GrPJCR59LDlV+omFpvZzop7sqB7dx1V
5DtVOMQd1sIkZVVjRN4QiLkCSiCHBGtI4Unzff2X1lfZZW3Je7Wh6g3TbqxHBnjf0XqFx+WJHjDF
d303quNXi9wmf3rs8z/OUrl9U2HVSNjHQow7kMsTwIOzVL2isndRf5uF28mZh6zrmEL6M5Phjx35
IJCv0zYNOIuNWWmx+rCe9W89CLWNcc2wwAZeoY6ZPkpKcKAA56FbSq5zj4PRFx8G7n/JsGxWNWiu
CNzqoPasnp477LBcxio0araON2u4AE3elgCOAMjnnaWoJ7KkGeyj7BiwMGM6BAt0uZKObBTQ+3Wn
9dJdcrbe63qySYDX9nC/JB8xUrGE/aDBDFW3RljxzRgtA61Yd+nVn7Kodb9jsqW4Zru3I/OQJhL1
XDTn8htRGABKrt2EqFo788wqeQM9sHFMtCmJSnpuRAT+K0FNj6QWXAsxB42OhiwXywhzYgSV/Mby
TuImEensgis+s/pljBGnpJvjaulNnEbBp9km7J5kdqKazUqCbzSYy/RIv1qa2KAvHFdCsK36WLQX
Vy2IrPPWpSbadSKkhHBkqmmw8zvKYiE4ASzYC+OTBuYLK3t6koqAafXd2kHTrr/mv4rdLjcaitX2
AAHN0HEEw37/Rq7lwPjejC2rayDJo5yUyGFJGvq+IOvzp3RrWqLfXbZ1bnv7J4Zr6VPhX386DyGG
RP63b9zPgByY1COikhPbIVcsVAzb+Gxs7Ap5XUuIsEirnzq7YYqVLiSMTQGSCRpC1VSzthx+AspK
bH5gBh5EIa9ZtUn7D3qqLZ72OLWhSRrQxXn/86qCw1yns7LZRYV9S/OWDR3ABkdF9lYoYfyAcKYE
IGZTDBCyMPbAFyBPHeEbsHEVvMNc2xmbWNSorJAHd7aXJz3kGo5AEiPCnvTTwy5xEbUBn/ADootS
z/4CF3kCGt04Y4pCab+39WVC6waF8eRo+0QzkZS3Qg8wJIsniG6GK6g5DPBLa33m7ZotBWEZPQjS
0olKtzLEYLXNP1OC602nwHt350d/npDiTaYLgu3p4iBerWxSjOBXzc81l3RG3OQCk/ZvH9Ph3dRB
+kKBp8I5Jb71X6SESD2N2gmt5gyR3xeP3v0wHBIFJdfgJRmPy46TGlab9cDWrzFu53+7uhlMXTJ0
HWusD2uvglh2Hnj+Iimb5dS7gTaSWRro9uK74/DbxGzJuRFv2X+Yowr1Yb6AUmRIj0hLGxeWgqH+
ECXManTgWppIAZyXjgVesIntPyOac76pmpMwwK42Ep+3+EYBWa1jDHWKmJxc3QF9R0DJGaeJwIJ3
WeH47oAV+t8hUQK+XKoKLipGaOFxYePesRvslhc0B0izWgPi1rVI3U0Q9ED/OrUGg7dhypxMBUlc
xQOUkfIUp3YeUensztIRyYTwtQg8UiuHK/zLkc+wvpPLYIEVNohlmJNhIC/EhQ68rQWf7DbKTZxA
sY91PNI/SG8lw71zum0kJzwxZncADFz43p55+sXMf/bjiS3EpSl0JavDuoOnGlnq3+DKzkMuOX7N
39Yw/WuaYIbrt0xcC1Q4lsQ9BmZpXQLddLU9pHrjrlZLl2KLb/WwzQNAIlqduwf7cmZ2kntEXsjx
7gyZTplM85NQMKZve8ISMPTkoDVutt2tUUMhpWo0TJPgxCYUWuAB+9q8hfKQa1ZeOZa7D3hciaHM
/Tt3BREKU3OIi1Nuwlx4IUYOkYn2d0Gxtlu8AN5WJxJeiYMqeJ73ZbEiIYsL/fANFJx/+Dxa/Ql0
vhIQJOBjy8DLaYR3JXfIUatUJxxg100AEFy/TKZbTOev9S0LzM4dvc6PBbq17UP7BGmT8LAiq+bG
Fh1UoxnKT8AeisOPLkht0+hw8byQ35ldpCSzi986iyjCXvSOJnOpytQ9ztEO9Ak6elENFrJ1mCiX
QdXDgxkOjWtrFnPmoYscdvAWaIZV8gjsE4fLqacEaHun8MTrpv2gEy24kUq7nmLHzHRS1gslofIC
3N+eYfMV6gBcKvClRFtztuswO/zFcP4uV02fHKjY7wrRWHRi4bR224cHltfub/djsyVKptNIr6h9
4IbCoS9J37QMBTKuzjmGSU7n/9JpwPIMfFX+arFsH4H+Y78cmTOzBa232WLV+FjIOvEh9+ise80O
S+NlFpNyZ5lrdHpabugJiJX5guOKLIt++Qq7yBJI9wm8l+dxPDIV7X/47RwzmBHfzu8ejTwAOa3Z
EWlS8n8RCBGx9vQtiAgPBZ9UoNyuWz6mZKkzZnvpcyUqC0m3g8BN27+Ii/cETgPru447crSjG6lE
m39jE+XdGsdfeqzQ11SIriDfiVSngO7kgQxnAcSvjN3S3x9XB1r4o4d6lulEcrUnNsSiPlcCyZfs
IE0D3ktOuJ/Ag1uOTjVWzt5tnkT8MgFneY9BCQ4jRQdfDup9mi1ox6KurhxpYG0ak/Q3QYmSDnfI
7q86L7L5m7hn/IfBEcEX4oDDTB9v33HwgAvedl7TkuNGD63OaP/KKvw3hU96tJmyC12W3dTkPPdM
SZM1OgaW1eA/cQlOT/WqKym0YIVP+u9ESk+HRTkkXKj9xXBdZ7hifV5HjfRuwLvzMaDcB1pV+7JH
qbbUQ2ZqPRyGo25Ii2hBAkEGj9L09vgHcHrJj0kf4m9NEFmLK4OhhVXlgdMXgpDiBpo5b33fIYaG
sYWkUHQmsNmcSpJLg1besHCYp1NyabyN07q0nM+sIIfo7BI9HqrQp50/5dP+rfnOxfxfRF/xrmL0
R55Oogq1OalBPuqqkXzWg92h7z1j7ssSHMSqgh4gwrak4mxvy2i67blw1GacVmprcuu8BjV6GZq1
PLCl7sGZsecgoEvt4Dd5DlHXc3Kq1/KLZGO8TeOhqZzeP4wARJOZM1kCSLxBUT39cXF+X+uyy91u
dtFGs8wXQHzJ73iWdg6gb5aOid2bZt1Kxz5b7mBr3cKasbsZm2QbLxxZkdVgdnz6a+SQED4Nfe1r
6sbsOFK2NI5XBtN6Ef2FZGjkvOLtDbBpPtyIUhricWW9FcgpO/LlUHbO9QR0ux9pN2YcJXEKehpx
C3WLKs9r8tDvt4ElrYcalxM1xkMWAPJOCg/jS2LEsJ3PrDUhRl/KMT47eumzOATEMZn3m88OiVpJ
MSFEr/nmweALNgXy+bauxAgwB4+xnmiP/xxjNQrleUNHi3VDHpO1f4MuIsOHCiBrr0+x9+F/PshP
3chDIyTosENlwJidEALmnVJVkbsSKoYPaa//fjc2XDlzvOpSBw8mNHo0iIHJYjgu5UrM9euqE7lm
nw/CriPeqOQiuBFvW0D3G5qNbGbxCuBRMBhKLFmYur78QK/pHuvTzMEX2gdJKaYqJcTJ5aVSaWmR
H0Jm9t1ZUA0kJg6JRRcmu2pw6s2UEs4i4QIuC2li9b7xHqB0+EVeX46YfGH4vYWYHScLJASjjYtV
dNQQwotH84va5CApul/DkhkkP5uoqz6RHRUM4qLhtZGlrMMvaNGapylB3fbUWHqjKS5b2QjxwWkS
IhKqNqPIZq6mM/9ejAuKdLzACEak4F8w4c/VV0uhjwDY7W01ToHsrjbjZTWgGyhpkS4mb/7yR4Qb
VrnwUZ1U0MBtBk1U2Ku3NmFwrFXXsGcdB2EMHVO6AdQRZCNW2h5UrKSulQGSRNn7aBGgpzE+2y40
+n/ASRzWkfBRbjHX/753eL3uZ3O/fOi1i1JNbV0f1YmgCRDreqvbLrwLa6agzdAQct6mrJJTl5Cy
3ab17n0lGMm0TI5ThQEke7sKQKKIyCS79qd+S/l0CFQms4l6BNpL62LGNYDJ739A7KCCkVXLNtwM
H4Hx0/8p5Je+dYrP7tHKfpHDIt+NgafEej+yqQo6/RnJvgefshLF480gkOEW551BcXA3lfMgcMlI
mJYUaI/FrmKJygmUt4Vg7/9wGC/apDHPAuMYUNrPbkajfNPoJHG4nRLdhFr9pPutLCkWMQylBxPZ
NZ3/ZGyxIJooWNnZLKASXT9jI9qVUCd/mEBw0wVMwbq+vHZiUbkR5LqqdJemO0oRQsZOZednDDDf
AIVwb/w6ph7rnaJ/jedrcQ/D28z4GSaq3edv8m6v6xLtYGCTrZh8BmJ9VL5A6GMGmjamQlOL7j8S
PyKSRjYb9LY5pNxLSXJTGPWGXAiV0Nun8ZkSYsLIRlb9FosHelkruRQVxLt7o3M876+SUKEDdTMt
karCSb0VxURpcWgHnyqP4xbhn75VNmfpiLPt81etlSNxHnbRJL55v9EncnrPfrIZ7oPQaaT7WyCf
z+7pktP7ZY3GCyJFg/N7AkcLCOXZ8RsG61zFikFq/XOQ+MPy3iGRrrirepuvFpvg0aOklahtTOYC
sj0pezF1a+IqsXMBbTHmmqeIDbNVjjjWN990PB7gD3knewSMI6XyY1fDhe50RtF/kcLg2I9JvUw4
cgSFrG4zJ931nyZOfl5CZy/W+EQDVd1K/pNQ2O8uMaJFRA8aInsP26TbIY9+ZCKbnWNR6rwNWVl2
YbqbG0CMmQvghjcgNj9+tknIhAVTEk9hLGOfLgzKldzP0xiS5Bf0ORZ9QQzPlqZdgTHwed3hpk6C
LHe9BALSIHOiwF0aEge+PHBWKtxTYlMiAHFIzp2AmiLOK5bYJn12qtSgd15Limi/So8U8TOzzPIY
XaZTbccNslYH2eWTH+5t9eiCmKT1itulPFJ5nhDQEUmDUGsggLaZqp6MPb9EpFnmmwyMY77UQDnc
zhTIifo4bjGsJfA1TpaitEeiJohMDPTHPDXE3V/tfGb90bofDFn/zZ8+Ror/CLV2mM7H3v4KXsQb
OkCmbbLk6YjcYhuAcpvtcXGf4+ul/+qzr06fMuS+khEwnl5dhL30s3PY85MrH7mT8WG2bgkLD0HO
XRxHCxNEdstCIjS+bzqfkTiCcaLvyuUBe9R2MFzh3XT4g56CpFImt/SN9A2z2qsjaUASlSr3rhUo
OymPIkQyC6QaIEHmidYAjiwX4/98+B0K0aAEMBFqcGABuUaowIbLdiBkzcygF7AGPTxtUwfhV8Sd
4u+7VDiys284cCFCVpp2c978LS1gfoPXXbzU4HGvFO77tGnqEGLvk4sJEFIwYbADvUj0onvyKSuc
+/pcWAfvxDV5LZI6ygcrXPuvMhpZNnPKkAvQdkVSOVN2bHHMXQo3XDS6yDrP3FB7Ax044cULb8we
GthAzQcPzhtuiIgdAFiuhVurMwqi0U6nuIfWzFe3L+VhH6i1nCa8yqFqHvuMRW75KIFbTReHU2cZ
4oxJ2bAJnVkQm2pTwLGi4Rqujg2eGwxLawgW7txOBU/mj54MNBMjJRPtzUcgEZVXLP5SEJhT3YsO
9Aqy2UhxURsQw41o9CrRsqB9qDQeLuyRt8xB6K0IfbYd4kCJGRA5S2XSgNA3givcBK6IeaGs6bHV
Sk2xz85ILyr58ooG9k7u7ARzhCgEmz8jm1/xhUFmPGKNSG4mIYteLanGcmjU4KTG1su1Vt+qPQCz
olDrEQr3xlGu20uGiLL1TE9zRoaTweybZbnKiNLNaGSjBqlos48/sdViAtSlWSMzbe39LtPSdwyV
JKLGtKIaRb8cS4sDXMdGiqFaFG+E2CZADH1GThapg93EirDctoW7Xi/cSg7s0D+/5WaCB98IMy++
5JjdIVJaN38IimgzgFvgabCwjHHh0rEh8lgr95vL119VIZI+ZYfoHoKpaDR9lxSg89zVhDKbLHwE
+vHroLpJ1S0g2qUgZytFoEmVuNbj5zqfM+7Xm0JrrbsKvzMU0wPSVmEZO3qt+E7ZLchWJ/boxnIp
aCrUS5SVjVYdiaQvb/yngfwnAbxPAwmenukXajFU3o0qt2pJ1KUk9XwQgj3AY5Y5DtlgkkFAPrU/
9ajccojAzaWe3s//ERuhrWnGIAngnRADqgViFXwHt+J5+d555JNtHh4HizHmrzjyNytvKhfNkc4H
hzAUB5Ci+95xJfnfbLHfUNQ+RDKGywV6DQ0loeC6SmpC4XEj2Og292TTcIRZzntmRbw6hVMuRm9l
ecEye+LeKTbTUUhwl4TXgJ2k+hlK5Cl6g8rW7QuyNKzpfeRrPp9yYXU/lxqdij3n5zKVUZ0pH0YP
DaHFbNMiqXNnirbXL5OleWtpj3AM/E3sge4dwqM9lopqM10xUphZig4iuHunTv2kmsZ+rEnnmPhb
Xul+Be9oD3a4A9VvFH3QKk+5W5eazd7ToBe+fukcVM67HZVsnyXpNRCo0WqJyu+tqqzL77XBD4Wr
cEpP0DhTAk9bfkaGLTSdUn4PA2/B6moFJELT4KuV738IFnIifmHRLGpWLJN8y4lCvmT/uUlsgCgs
UFQa9eQr5hP0QWZtrJvwZSuJfG37FCsdK4l6vIFoYThY88YCn2KjBSmQEQ+1SXYmge6gjL+9SR1x
S8jeyE7yvWs91mAZBhG5lHntKB9yKr3IhN/sfVsDASfUpBlaiE8ILVYebXKolMZzCrVjElsY82v7
EJjqc2FP/qbq2gawoPbvohU2ZmO7j3d+AIFPkpx4ZQAUW87aFQzmvY/kufg4ynE2fYZzo95t4JUX
8UJquMDzoVZSNM2IoJtwZujtJRh+lmn01g3oM0uxDwDf1mlM/29F95CEk6M7WcCNgNUYz/wbVrBa
CGpdoVE26Zy0hXc0EqZE8ggeiGREWsC4gACiJA/JLWK0Olo+gVbcCx07W1K8vqAxe6W0Vkw10iYA
5TAPJKKiH2SkGAEJidl8U4dnoy4roFYUpLjZ8vbzIwDAn2x8SUpmVlncWh5PdiCREh+/5dFJZQ/1
zm1dYblBRMF/U7RHPvA2mjs0AWwOtU4Bng7q23+tK75IWQlSRx/yGyx2PdXBbni6KT4GMaHFmjgU
J147ZzGepItVpy9TCowRASzGBeQNVlY8t8hObSNxNeZool/4sL/CrozAkPKzVZ+Q0RJwVoweR563
hwaik8mXxob+YY8Yd0BJRt1oEGB7PJzG6D9bQFdEE/EAdi5MnZWyfIDfRLQAlmWSYdz2Imd7IlqV
TUoQuWXNii0KHDC/CKLeOsbxbkxK2YXqJetMozZOwbbWn+2LxQQGLskUjuXQ956orcH9s1D//lY3
poWP7Mcn4EUxA0TV42B/g4HSm+z0VeO3TG2liRfKLYqjTFXl8wk4rxEIc/Q+ErsHa9lFJb+NhAEH
2kLWYGQxa32FNBEkzz0GothOoRL2LTAxMurd2glfHN1jSpEVmyEbgG4OZd9ebysE/QaBmakYM2Di
8k2HtDYZfYxzpA57KpjUG5xz8GZ3Ea2eke+LmfpWZhWpB/0RczdP3gAw4RvsRpTPOqZGavIvhf4o
5ZFmxB9fbWl37FN5pPhRtqaFKbCUAePQ3LtV7AI5xW7cqGOIlyfOkE7+VGJTxXSSPXmGwErHt0Ir
oRjIBqzoMyVrbWJzlFTDWqWmT80xIeBFi3zPkauQmnJJlJSDTv8teUd3f9y5LQ9+VdlfnnbAwckQ
0xDgHao6ARU0R1aN9ev6OrZAd2w6O3X88g5e232AuRZj8A83L/XX4bEB6HoYXIHlmqbm6b+eUdsn
0efjBMu5tzfcEc3vLdHlvncXHewjKUzA8wkzpFInTIDfSwCzYfnvRCcxewJ6+/TW0d7PdwV69yAg
uRIOjnWJLwHOoMnHJnQjL/sadlrQb+lw586iYJ+hKBj5IeCv7uwVUx5H/s/JPy8A80GewtVlt67w
Xvifcks4Ci1mbJvHLa9Ewkajg0bnyuwIhnajDirzXuoKdWBmqTnIWGFmoGU7I67klQBFO/pApUqy
xInuxiGUujbictMIK4QNj4iuZE+oh5podDbBtX+FrcLXtqQiqGk53UsYCIvbatRvdlCrkXs8wLxd
J6F4eiUk2nkupf+LXnKrGGJjoemogbywFEytf5U7NscfJUaRLZS4V9KOZtCG98qqSr/kVVQqmgPs
vDsnsjyzOz2vnyCGStgYpB/4qd2lKWBOoXRpv5XxEm1pvX0gO+cDAcyP9Zp57XWGS9ipOhyCjgnP
9Cb94G6McP1l4RTkKNNH724HXdn1qyXPzuE8WeqREI/rPKdNICOjlVNiYHmfmxZJbXbOdow2TgWb
xFO1f49xtr1q4IjwpkeuAVZVWbnKl695VEbBIXGWeHXqAALzrWgcbE9dyA6YuXVfA1J6B9n8gg0Y
ZRLuwxT2Sdhzc4xqBlKn+YHYvPq54+u9jlcK7c3oH1D2SpNnKWJoctLVLu5eiJMTb/cvZVWMuWwM
vCf9UyUE1n/ytrQbLNbKR7hX+HQn+3USd2yPKt+MIMUlx3qg8Qjlf6UqDiDB0lZLXMxW9/UCqE1d
wQO0Sc8+zUXR7MTUYegc8QiBo3+w/RLVqPP3ojoeOg57K8pnRx1Rn/gZQVviDMhvIkrxogKEFxhj
kwWTISv1NQpy8/yGtuXRkreS7g3C2Yh4H3i4Muz9NTxNlxCAjPkD56erz61jzqtJGkLttlkC1J5u
a7mvdqDgoSYWUivgXfo/5IDQ9C7HeRUFUFD02mB9XeScAuIbnQpOczGJi+G6c0GAsTf56uI4epkb
vqcDysiz0UjcHMMGtWYQ7Tn7Cq8/opKbligB9+m+DWOl20AErJBKmrUJwlwFW3SGBzqpcYLBdqsK
jFGFwdQtGwliVcGa+6sf11iNZ8gMmrAirDyG16UQaESFZppqqWojzJqN+oVYrdD/ug2464srZZhF
ajoTMinwTCNj+ZhSVL1a+jnZtxO4adrvgxoT8hEexO4oiQsLz8JIGP9BEtoEbgqFr4m8MNYm+dHE
678SZX3KoG/TbliDOni/wcvkd8FUpfPS/FYxDIgBkztPDdGtvMwJNn5OYxevZW4XXZ6s26QYcfWL
XKBBSv9PaZd9hVq233GTx/sb4X8zX8aP/6nHha8wCjVVWOiwnqi175xHV0maXIzUEs1uqf1cPU1g
eYURm04/yqyyh5T64PXp5N2CJbLYbhKU6stUQX7M/Hl9cK5Q/OC8VLrH9D8xLrrf7uU5hNVmx2kp
o+uw5uNvIH4y+QfMS7mLYSWvV4aeyLaKzVpIXcHfYvDsn7vx3cij/dzUWbfVQkivg8qIlzqE+LqT
X4bbcrt9vUVSN9ac7EpeKs4dI3M7zEhtguxnoP8jYPFQ07nthHVDh7ze/W8kZN9dIQYywPy4X3IK
QUwH2VCu8XJ/geOPv5I1KkbzmHP9JQdvvXCiq11JNEleP4t8zkcy/n8JG9h3XAIfdnVM5yuw1C9P
DDO68CMtZp9/mpGRQg6+DIgLkBsCv1HCcrn3BjBLRa8pPIhtZtV3ned+0BsAhRAxs14HRSDC1oKG
sd03aImAM14jyv4LkvDeFky84qH8jQm5OSUlI0WWjR6vs1SyXr0kFE3KDM9oaJAn2YHGwuK0RDuo
xfabJHibcPQinSj/II3soQKqPNjOI38nr5X+Sz3TB9B+ZYFICi69YE4d6R0MVrTh+gP2RDPnP7XH
RuCLnvNJWFpmdUVpi7/vv+ScWb4g8bHXIZOOyL0hoHk5+CEti5ybO0rNACS7mD7NfdKcFfOA/n+A
3/fzE2VPHKqk+Xg8U7IzY1HyexaJBFRZPdgNlZHsxWqeA8VVixxUKDAJLg6ueqNsAHKI6LulA8cC
fEpJx2Ywn2BexjGd+w+E+ksL6l32U5iC4a75+n1j75TrMP/HOCyJ7AqOXY/1kAGM/8q388pKyBsb
2ks2sVsUWoCC2m/dFbgnh1ovXaQ2XIqobtc0i0gDGE4IYnZw2aKk2kKQECQdkuJ2A8QF8KnT8wJM
2urQ5o7VZXMs1yBZ1sX/QfJOur2GG4tdw7FNElTBN2kojuhFoPNEafWsZFtkJv3acv6gbVbNoYB/
AlN51wg8n/Xc5/Q+Ue0ELElYx5tugyMsTJUGOc70GR+Pj9l9h2U7nU4Ho4zZVA4Gtvkxp+cTlC0p
W5UiZHBjwB4mBkNiUfta1qpUpoCUaI6XBHtWJ+SrjkRrGg/FEgDROUq/L7Q6jNYsXrGV7twW8Jti
3RkibtuB7gHyIG7iS9TWhWG8K6fFd1uq3EtFOBxiScrKH7/yeuRvxiWiEFSIZzkx0B77yk1i2GYE
v+PJyXfyf40AJ6FxW9Ou7JRFroT0wcHPuPEGoTLgU11u4m5MfAuTU8nXMAl1GYCxMoX1LDzlFGcp
kp7h0xK/F9uThsJIj31JvVTt4sCLj2moYQglqAlqTDpdIFn2w5siDyBc5/6n/dtrJs+puGqRFV+O
YOp8LVxpfV7JFOZ/kYgfA8otzEA4bluYQCSXtMR+SeBaUfNvlufzBz6Z7czRMfn4re5suerKWuuw
Tg86fVP1WrqZzT118GuqLTwvIONd3ObhKYQFRHKOMhTw/PRyIugIbxDzDdQTg38ObisVNDXZCbAp
Vkyi71sO5RbfHvUXm2RmCL5GZXxmcUFfeeRUuKjmZ3yoMBtHctvqtr5ryn+3TSq9syYUZ23K/4hD
Y7QD8PLqa5xkNMY1T8WVGBoHvQDmPQJUKUxdgxeWIMR5C1PAIsfqJ9z9jZbAQ12zDQIUdljPUQsh
wEJE9GxohKgPTEr/6L9tLojTjalAnpjQGvLrfXVRHwxFO06dXV2mj5uO2iFDAJ6IwoUJPRkCMpZJ
2jSne/PhAccOgM1zqziO1TrpTVDbay0Z+AMCtxQFxoiUXG5II6JMA7fHLJtUBpA2dWnYYGtko5cP
BKgennFe6NjIY10tTqU+t3jVgacwVERCak8Z6WEMYbmWQmvnsL/smv574Yb1mcLPx/xKzbLqjidp
07gd8Yg8Wsv60cuG6+nc7nB+uove3U+wGW2r4GMcOgsWtAGfvJYCGtb/kiZ/ZmMzvBSYU08xa53D
g3J+gHZ0GDH93yFh8aayo/DElDEfe6S8gR9bs+G+TxPNEYh8z5CjWUiIZRJj2K+Z/04LAsy7DsQW
1LI5f8sx4p1LI6KRRDfz53M4+jKONAe3CIf4GvUoQ1hmJXh0/KViao9Y5u6e1aJ32nm2Docd1G5v
64QzIUJOZpDUAGuw5HyfJyV/RZS+ZYtEVFBSqdYJ/mmrtWvjxxeQ0XEx7MP5WJM+gjGWIXn0O/DN
fuLmU9+HGAk8R1mlD4+n/oWMekVpOxbUJ2upg4DkuQ9/uW7akcewwob/h7u3uxWngA+8K5gsa1gF
FVZXw7zKMy1zVlAbfwGWy1g6ogyg+pP1TxvjrGT/Hs+UisknfsGVdD2bM8dooJ06XSA1xnW8bLG7
vJiufXTysKR3EUCypdERsSandsK0kEvaDEfqy83Iw9uu75uYquqCGDMSsci8AU2MyCztjRhRDJm0
vw6UmV5w99o6fuZKi8yPb9GLvaG/5TszpUSM0UjHY9ysBGozWsnq3I/Y5Y0xge8p2egRjqU45yZz
BbLjpGXkS0wDcf8/3a0dG9MH+csXQkz5sNpkXAl+g4eS39BdNxpqrdTCtg/mwMKmXcTaHJM8B/gS
kVFG6ZwWKv0njehBdV3c6A7fN5FesurGBQxYDGaBzJdZIDs8NNfeXgYaxqvYWdUSphdF5q3FJoi9
8UMv5r4Jl/hjCiFq9jfHOw4Jskq+x9QmL949CMgdpJHN9EhOTYqmjs86SjNHdMUuBS7C2uOggouW
70yBYnjpMQVfCJho0NbYmduzlTjU1VJZnPs2/7qM5JOqzZLz2/l/RMgGcCLMZle0lbNI0w7fo2br
z7uiKe133D4/tqBabVfRzxfCZx0mXTIScrAPQfhz9+Qy8ZNT4yX4UgT/89n7cQjRaZgKktqWLVJT
48+XKB08fOVexxBXiX3W1zsdGQiq9BPaDj1mkwbP5lD8RIPdjLa/Dt78Uct2UKK84NaTlj9bZuOc
bGkHMK7QL3FwEa3DU+ZyveBlVoOs47jFFjUh+vIxFunVPq3407Rjw0TaX2Te6HArr0W4y8G3sTqC
c/rrBtsqUdg4mWnsIueN8TU6YF3Drt1CokdrQahja6TP4yRA/W/2lrkB0T182WR/SrZHWsUR0g/3
vkS2QAN1G67v4BnJTttYtBtkmu6+hJE8eMzGP3yAcO9LDBS9S8Etw4qhCX6bQbeTLAr/+JiLxZrf
J00btgoE9/4jWd2fmjnUgM50zdMhpsHnHak9MCUGBOt7kCUBFPbm8Adt7y32m7weyK+yMDRB8h83
Acqlw0zivwSuxM33p1m2Nf1jvVWgBF7197VpKneCMAvxA7kZG0WM9TgGDRIecfx5kRMqGbjvaSxj
5voMwHI7Qz2BeVSBxhqVadX34IORQSSnjCQbuIV2bfbERfqS62neaY8+eNyVgKX+OnQhy4+MkNyq
oX6TgPw+RkmCX/QLe96pa0P9sfPvdtKpm1NbkONs3PG6C8D5yT3m7UNTO37rn3NH/BLWSCtyDAuj
kHvqbpnXnQWhM/WBo14pzI9QklcjcZrZeadeFV/OaFX0fC4O+gAFZl/CzthlVvB4578bNDAn3Dbf
m7fVS/x1ATQksWltftz91yRn73RBHG6dCbCT6g7Q3m/2XuZgzi+x1v2WIj17Vnjy+7sKTQbubf8t
76i9s8YdC/zsvF3+g6z7iLKMh8/DHNdb077rA4H5tziDIV3ZZPh7cKd2c0bXzS5GFXdWbEVEEPoo
2gACnVPRWP6Y2iDYzOsl020oVuX/q4pMATKkdXqkZFctwGCdr+B0EkoW3+ns1uzkKe+8/ahSHjdn
acqql0sM6pg/nnYXgi8vAoA9kdZyU0LylfAsZwsomyzGv0I9YjbII9PLexhyihnF/NNP/XJ6zoEV
pi+qXJ3EmDvbz/FAAp+g9++iLA/0C4zGe/2Y8aZHua9Ty6+8pIaD+/FLI03E1Utvc+uZyBAF9Byh
UE2MBhDkC9gCmprPJgyn2K32oBMio+1HG7PvptjIaTccPyhXTBBRlOjmrLwH/KFoA9Y7WtHREXiH
aD2q5zp/yW1rNELCATJ4sLQWXlbKy2rLvFdkXN9waQQ+QiS8kLSATDkjiMXOeU0MldnKljF3sXIq
rVyex/5FU8WIEDiJyBXyS4jvOBYcDiLMECBWsvH4hBopqzNaFuWdoj1jhhUgW0YP8HS+xgadQMjs
SigLwr1rNPX4VPLYWS8bdOlZjgQGfR/f4A56JjnZFV6Tdjts/L+25Wxr4ZGrDFijlBXU2fTs50uz
bF/cqvhEerA3cBQiX881/LQxuNqat7C4kB3/awu8WFnQyyMKwjyCNzKlbBwS4zmEVXXsYWWzdnla
4wvdznrJuTXk4in6Q+kuqHFxJpqfwgrnDAY52QZ+4sfddY8sTnPHP/ixVWBysUoBIfFGeBLoEtgo
Yvev0yBHnyGSF4VQ5tt31UoUkJoTesqMiAIcgLP3NwROTo2ficwvAk2FzzhqlJKIh/N2aeIZlGtY
ZLKa53njrHZA66eI4X1IqvCKLkI60nh+/7aYlWALKjZEJ6i7B3V4XZ544IlMxercMY7T9UFPjxgz
IUL10qD/u7yxZaokAyit3qpvukDaUf+qviKciGLxVI13i7Jbm0miN9F0vPOdQuqwxIoR2gyu7dTX
LG3D1syDyA1ZL6JV4KgWbc504Bnt9aBN70hrQth6fiF1R031OM65Q2tjgt4VVwWy8iXMbk7eDCfr
iziwOO1088b93Hg+x+OqS/FEtLt0tPdeBAsw8luwoP7gdygzIpFdqPJWC4cMuUauQnHkpgFvTSoS
Q2d4lb0gGbSQ/RU7/4qvqmnzmrUjIxi3z+o4Hgexg5OWOCLUqLNDa5Ne2pxVKbxzWGYTyIqGxm8s
uYHD7QExdvVcExaqXYMNTXz/2dGvXsH1FAnFN42oH/3SQN/MD4YOT8X73CCL1z1A44j91KXwSqis
0mCWhBiSWLhRQX24G9sTcExKhsfY/xLcSYSmztP0NIKd3x6chrAU+vaPdHU+Xw38qhEsyBK+0kQJ
buwoulCXhO0pbocPSnZ0QQ6OidT+nddNNpd4idbENYLb+LuHpeasbHABn2s57LAQblUDUT1A980w
4PkIiVVzTPQtrLd6k4M0QU8XZfRiFinO8cc0w/8BQgyBjrZ3CLpccRGi++dipKYAYuaMRwTIn9lA
G69rGjeYdKVnkeolikLGq8WaqDsIB1I/6AJPg4U4KGYvksODOyi2w2R02PB9ThVOg8PMAk0KpYl6
Ni1CDMAFxvC1dxEIxvqpZR76joA+aK0Qc0es7mZh12Xu2rw9iI26E1hblzuVXr1rzHCDHZgczuSr
4+s6zOEz7nfm8jRTUu0lpdo6fW6ghZ0neUCXxAnJrUizTzU9jBzaShxKPe8ioOjSf6/5t+Fuva1m
nTZtUWXWew81BH+sB8/nsScO2+1EEsvRRt0GNxeduyDhfgkHmNKMHkHJDEMKE5Aa6BO//C3cnhTj
Lbhyh/ew+S+yHkXNRGnS06D15I9e6DQbbTU44CeQz/bhPKdNBCLeJE0HK4HdQUL6lFeaz9ZsQMwW
es3IYa0xyihQ5GrbxR3MctW2VNd0nAqY1kPcY2+dLSX7sX3hQSWRGd/XZ7XdRPJnHLsuUNW5vL//
1Drg17uDLngTGnHG5Y8QDkm/tRgncAY4bJnmtXjk0U8Nkf3LBWNQzN2V/GVZpdALiEk/WZ+noLvn
C1OFiczrrW7FDQSX6ClBF+BSxoWrbCHgADsLqdecjDGxSmsD5EBzyOLDEKUB4zXR/L8gYnoUC5+5
Uccu8gMRXHaR3nrYwGFOMeQ2Oag4NImoucYVzcXf42orPV12Q1u1iqGn//3lV6rBZFvfL+l04qAz
xDb1vIP6ic/m4ZQ71C3i1jNPBgVR9vEn8KSWzO95WzwuPubOXp9Cf46OwBnrOeaJ+I+USmJk8kgd
PRDAlk/SqBozhGZSP7qx4ciseyQBpRTJ6MtKkr5gt8By17dkEL7EaKPtJPGH1Q2PF0SLer9cgp/C
ZFn3VNyQEHeeog8VMAGUqqSUn/HawQhpePEI53zycGm3Si6QDDDsLFbQfS21sp7sWbdbTX2QWBOP
7AV/N0ntOQX0cA5RmI0U1EY5L4S7iY+zPaeqHd8WQ3ygoTVB3FHbIKpWtcFN6nXqCpJ9d53+a+Ex
GHSc3Dsa0sin0BsjXfc1f3Aw1xSr4sjsT1f3MvlX4xlMVGCTFDH+4jSYHBXp11teKW9dhE1ug/pE
nn4l/r/ZnhPjiIowmPv77rjMtu1uZPMYJyrrV75vM+QJ1vddAaTaIqUz+dIDd+3aoTi4VaysbxeV
bpayWW3oq68zjjgGkxQGNKTrOVVB/SnhZ5RgGvYhpQbpAMz3eo2B0mQw0Z7GjIWrHl+0MVt5QwAf
owdv8i25MQZKQmAgkQ4+K6TVHUclOJsHFvUiO4d9hRjqA1LK16NnRFHSjSMyO5k8WEk4+JJeeq/5
JcsIMns3HurQ+ela8/GqK43z25xQuG1ECbG5JduRN+YycuDXmZq/h31YTqFQx7IdG4yDuG6Hi+w7
XYuVr73iHqCkGdCeaNVGpHkcUoLE6j+PWEtpCc34yK0/oZRL5pX9RQ3dnXKO6fh0Jjk+7UTg9YmE
PF9/2cW98+YZ/NwuvlblS6Ys7/1E1O10LsVcarh0ShBD65mhxqwHZJrT9yYtm497flmHZuXC5D+O
CAcRJ20UMpJZDQeVq/dsAvlePOl8vteIrsT89lXWx4LVteUsfgkX18W7aU+/HHtXureaSQ99NOa4
DuVgmNcuwAnXypgaXiYMJR9hTfLFpAEj0bciJlDqyvYQhxSW7sqNN3BdsAn0MgBhpks2b5inOdzn
k0P49uKV6sXG6oNmttVOAQrXkU4RJVkm7Hd47V3k2FKPz0hgeaOQNagMnetAfGbuAaYhfeI0Euvx
TUlJ50YE5yNH6Vcz0VipTkQnWMOUKsM7rJyyvjjBme89iaSqiNzqElivkEa7KuFKPwfJnW0vlI4H
UpGKfTQBEByWCL2BsDENM928iApjER9N8Txlx+XvAnenh1y6q+CH7js7rd+z0WTWnv3Y2llImiRe
3KPJWm7wT7Zft4oqewu4ndY03cXcarKa3MIxJvyIWWIZXcJW1hRsx+MtVUNKu1y4D5Dw4vuovQVe
QPnR6GpJxAszDmz1ZGB9eJSEE8MMxXhmexwV6uhX0lKR59AIOqJwlLMmWORcuodW45TfyQsVDjo3
0vg0SjynrH5/Lhc9XFEPkKt0CYu/7enupl1/na7dn7b1IFmuGTeWuE69qCPHRA+NOwT8pATUSJ60
nqodUOx4JUdQ5mk7ZIrnXXsCF1w+jnNQiNyzoWl0RaLtEKXPpV0LShM738sIDW6qeS7nCj3jo/ib
bW0zcJtx7rtpFhUHq02grUl17s7HF/iYXUGIwKfqYgOLpNHE/frJ8OWPGFiNqv9KKr/HItEeeF14
m3nq8K1f3J5XIblsRc9Pa/TLk2CtT0NMtpMH2rpGdOO4nQsmTU+fzX6V1jM5Dj0DSditamINfecX
ObYKaJAIfblcmIUj9ViTwkSucBq5fAhj+3lvVfuIxGdnBqOfF+5KIyMHIxB/g8mthmkmNOm5i0Tb
dxcvFpcDGsLxLDFExFvFTet5RRbbq58ZpId/RDm2Rw+rYoDCuO/ccPyGCKbEZEWyhd8Z3voy8amU
vTviG1fqO5z62IKL/Uaps3Az71AAFQUkPvup3ypkPkQVEPhlI9GkAIpBxkXEKQSkr5Ts/On6QJHB
u/bq/ETCA5bB/2D/4EkAZ28cYd5/w/v9ls6474zx3sG+uDo8x/h4CPbmqtF/teIR5qKHBiKgcOv7
EJXyPHoo03vl7JfhQPMrkLrc9luLm1rruOzKVTjpnTStRma+ZhP+XALuc4K807zj1BQ8zSzBwJRJ
wMK6NXmOgQzro4DDjC8THQE9ZoNbAZP7eghIuAD+WdIww1MKXgvXF4akn2nrT5mALQwzL38YxOEh
Qn62wRgCyKVXdmNW3S9k36STuGyogft/p5UIPWivonTMXGgGSwt1+BfFkh9blGgMcpHs53JXz+Iw
s3yZPSGy5COvUWixqRe/5q10uLy2WblCLTX15fZPm1u0e1GiIsgkqKAuUMn9mrOl2enxQJQyCxcx
qNcDqy8iCMN1W9mLsme6JWwFEnwTpdCBhMXER+ytKaNUuoyx34hYBaS7BkoS4mhxHbhO5w7sbUbW
E/Bd+Yk5h4xniKcVpEZHFaHfc7gs4q/JM0EptGyO9TDjluS++ySpxv1ED+zvbxon5pTqI825Uz0d
e9Ux6olqoP8JntlufYkNnFzZKgnvgQaWgWqsy7vteIL3yqZxOiP9eVgS9jcsFZAp/1O/BCGXCWwT
uCctnVck5hM0WmtI5IVtcxbdMhDb01lJFw6SoymHLHuN1aczo0qAry0daHmuKFAmn36/SJ8MoVLO
eAi/zWwRYU7gSUP9ICPtdXuKCNhBPKuX3pftN5e6hg2DPw2LUKBoDhlib+ana8gfVox+LT3lf18z
VhiqLGKS7DMjWO/U4TFxJHuUa3010l4BqYd3jwrjEzalbGbvAK02VM4pfbHJVPem2aG6azqss+PH
HHgQbSHmqjWgQkCsXTN3PRNrs+Zy2kmNoZFh36gwugaLwWigc4McSyGDGkCKKV1BKLdEqNNYBL4Q
jYuqOYiY34StngeJ2J6b2qo/dVtPeyF0OC2qtjJENpy9aYeyr2eP6cqpMQFs2/a1Y9bMLCimS6tc
XH4923Dp5painI5Wu9n/lFxq2R1YMVrHRtlQ56CIAee2kaT+T5800VGobVTqgwQ5bQPKIAOcnv88
v4+sqCxKY6zq9q7/t9kysDCQSxlR1emVAxXPB+knKRpwDUsS+ktuxLF9vAL5SNRiZ4z15XS1LUNF
0QLNoqRCjC1Fv7bgNAI98idWz1qHFfqvw70sNu9DFGzDwnEDim1DEITroylyeX57JqzR6ZeNtDHw
PQuXhnH2JT7sNJxOF8PrL7YvDqy9RsXGV503JWuaW7tjIye4nCpvHdHfQb28tr2d+yYq6bkY5hKf
f1KVg8i4LoktGA2Oupkx7rxavsuvtqa+0SZIV0iio62E/7LUNGohyzlNldpRhCc3a1YJ1o5kd0nB
GsxW1xcS6hOJrNHZ6jon/VKH+Q30XAeHU24a2ffg5Qem74dZ61WnJMk+Il1rkHh5oZU4999ZsUSz
qmErMxXrS9g7894zjf4X8lH0OIfAWFPO24dXxoUicMm8X2OTcOkv8Vf2BO6+RUOrjhwI6izpoY3M
MlA87ptFUMPRsdQG4J7IkfY5WJsE6lppOArIvhQcV5/bTZj2Dh++/22biwWZXtrjiaVqmV9AFKYK
RLFZG2gwJNoTJnvGTENTSWEbelQOgO8bkU5DPqY7KL4kVZgtNPn2+adIthzdZgT2J6yH2XSGTHOW
90+A1jVcsoCQ8UlnJ1AYFwmH8mb18kZBRSkrAVb8Y7VHhd1rEdI3kehbgJXVQ1hTnaH3tq6N5/Sa
t1NAEhx/yr7SX01Vgh9m5CEUB0vsJJE3eUwrHAg6t41FLdDhJdB8lgkrbmJcAPidFgSb4/3QOwTr
ja8lzqUM/GXm3ZYJe5DHuTsxn24u3SXrN3UsQtir3xO00UKZ65P1o1EJRhFFxXBR72znjsXV27ZJ
+U9n3MQ1sd5xzl+cMs9kYAmRyQVnWsUPI7mmQF0nCg9yvbHqrTMDbUly/tC6983XiKh4TXZ+Jprf
VPXBAQ7TA5hCcI9OtM2/OYUDpCBbw6KN1KG53gJX4+Ozoo2OpBLwYXdy4zNcVXoJDygTkWlzi5a0
iZGGQhBIw/PrnmG684XCuIHqEtFoi9thUCXJV6INh0WjjSbDJ+Qg50yR8Ef33aUj6icsRBy1QyuH
FPKbVvN1qr0DPqs2RgWF6WG0dNyPQ7W1Keq7LOzY8VbfW2kKqJ+k+wOVtVM9P1ZSgEUYZ+6wBo6E
mh0M9uSVp4nvl3G25ho8BCGJBjuwMhk6wiUElTfH9AqZOpSIuE161qKm16sCvnKKKZ+qJJKHACHr
GXo/JCmtgozNkz06SuOpNbbsTlvDCe5DJ9TbarsnKlPHhT0swPTn8wl1LjlHTRqj21QXeeeMrst6
rz8TWwS8Z9/kbTa+DkdtSWx3pwOf6UJfHo2nWx0s5XYc1vRPeKxjolACQxxQmblZVVRDYnbzq9DS
HSsf3X1tMvq60nl88ZGBe4Vd69M3MbGta2me43Nv0OdUy7VXM+ab7HBrOxAWv4GHmgd2DT+aBadO
nsgbCXT2Xfttcmn3wP/5hx9qVCe6PqvqNtq31iLGogteT4exDk0B/vOM6Sqy6xVhP/OjW7M8eGg8
My6+NZOoT4D+wgRnI2c/Z1Xyr0W2Nh0rILMSv7j8ydTTjGrV1Ibb+J5rHdpk0Mrjway8YLiVptfF
h/SlB+kAosVg76m5Dx3Z5LH1ht+pVKKOECj9sYhG25yf5A9FNiPzw4hz6jKdiYQcR9ikw+T8YN2e
zaRwlrOAXFyd4NV6RCC/Bx/34++KIsEqmFXOPQ9Y8xT63iclar2wE4mCYxVf0Ib3dVZvZhDKK6B0
RgOD4fZyTkiyfa0c4JpXlXi343NiiXB52bEhCz1dHYmlHn5oP3W1Lfk/a921vyvL1j9cxt/6sydz
5WIZdH3xZ6yiX5D7Ju/hKb7hF4mtVcof+qBmXUW74SRLlqUJ0L/liyN6KYTe55Zaws67gvE+deK0
AB8zHJ18DEr1JjJwZxMdkMJJbUQQMK22qYV4rS+7PJL4INk/mgo+QCu6eX9/oRykeIMK9bezUyMh
8Bx/fUZg5d2pLQbH6dBJg0uvb3t/apSEa/NHJhTZ56GDgoTRs64DdYmvCHhRUN7ZN5gMHnblcy4q
a6YglUC1J3krOeA/swxCXHu2kLXSaITnGvdp3OWBfz2jw2pFzEty1GLy0J4H2EnhIlh8ao2fF3lN
TzEarr99cC0y2PaU5rjT61vpWc2oMLCZBmexpPQBP3V8Cy8VojO/tSJgRhQSdbavmXCikyeVDy4i
RE9cf9nurqDyGnNFtEk/e450iszMwtKWKzHjCTa3gNTFq0zJti6n7LwwCgNtT7esn321NIbJcAgv
vNWXsM665Azgeisl/rpnPHDUI5oY6E9iFTWLim2A0KsCUVfRLee0W1rRfJKTeF+w2sgx+pmbgyOG
4fsh44nFhug8rH6xl4d6Z0H8chjDB2ov6EqFuwlDXbaf2D//uuQpuhVbyk169VEuBlSfPwhtQnF5
pI0hIZeOvZfyHKJZ8qnYW5jc7sbuylP/aKIfcjhd8EeXlquMuLPAAMcpnOawu4iTu2mRsvZTXse2
EBZoyzN2UmZGZmGb8q81XqRrfx1byRfAoA1PL9EK7kz3pAdymC7HlhPDmBCMnOw7MrpS77xlyxLW
zIEqzg1syYIx1g3seCbMLVapHx6CEqJpQLtWJF48UbtW3HVZgPdmRnqkkLj3wFeX/Hf051k2oTsA
rj7nG4KYHxs63E3ffDpMoDCzsCFl95lYuc6TdXSmztByO7WpxoSCCIiMfZ1/kk5cDQ/D/RgEYn+3
GWDYrpvwBTY9U740CEyOZF2hzqRH9AJnE2mIN+UYv615mhdRmYIo3DrSwW38LGHmcDsY6LvfFXo+
r5DAbecEowt/BK9jlaQn8bpk339QKiTeD8rxNORYXhAIPds/QbLOCJBFcT2KdLfqXpb5lJH33/Sc
M7xLNElmNLMmYlBxWSSeNnAMPMAebdLeOveKKiRiMb3cr5cNpUzTx1dsIi912OWbEsGVOunEtTux
GzzgPw82fJwbwPJSWhTU4WhMnGkCEuQ9+fWa5r+Qj+6fU8qblBU6jyTbTCcYu/aNS/4z9oPWotCm
bXoGnEgYS4B4/vdmU3gnahQoFAFF8yPG1Nfwvtt7WuL7660aclF4FW8SJlHG6mKAEjIX/dcZhMVb
FXn1/Ut/d9zEGmLcbVIuG1P7VCZz4r3R41zsraoKmNj+3B/EeYBUhPmcHzzX1b01PfoQQ0YfPATL
3/A9IQ8qfZ1WuEL0bioujwiXRGIxsOujITaB/hijpF6GB4MLjQgPDrd5l9ZN69Hkj8C9KEtlTfaT
G6Ip/c5tF8elXoIgZPmD/OpIEhvT/SFDIRbHsqeCUoy+8xbN7eIGGWuoAm93VPqpWVix9BGTTxA1
CliGgQO7jK2P+OucbBEpEnCY4c3208xc+YnFrB3Q2+r0GzewU5V6Q0o2+kmLTQ4Mh3FxDvhMisjp
/PGI9/HCp39nhR5ic3sL7BcuRrJBIgwOrp7h45AIoN6uFeyf02CrKi4IojgjsuHQ+gAZDUuMhKdH
zTDA7LxsKM9DiARfp/ur9LZzWUjeimrhfNM5bm2DPDUPugMGUz2rRnyIACwp1LDjXVkhRQrN9foj
7QcUn4825XL0qAWN5Py67urOduZGq4XS4lR4ylHeG/9/tFaWg1Wasfj0aK1IVpSvELJgxM+nXl/p
SbQj0//ssszrOkRZ46yoIl/yFTKcI7pPRQGaaFXefLRgyEDcTkZlbtsh97Ev4mvjOkZ5bvFFtNot
B0yTvNF7DPA4HOmBPhafC6cUaWP4Ae5bDWkarOQoPxco8fTUjTzQqYYl/kRbAyBdo6GpDOwyOupN
V+RwAg3ObTxe0hhDbaJBqhuo3w5NTylFez6RDMEhed04HQ1y2ThOc2FuFFcMDGhdsJCWv8Lol1Ym
Z+18a9aD777kPQADqltfldzrl1bR0Th8sYVsm4b1+6hNGFvB1u4iUutFrBP+/9pa9l5wWE3d13O4
UvNqw9LbMV2ussZZGEgV9GccT6A/eL4fr0RmRwM6KT7aLjLAXrHSqH41Xz0Ro8u3kmsYIeSMWkb+
ywGT8AXokjpm6M0eOPbzsiNaMrrHleuSMknSPspN3fAG68gsKu4ODj00xdKcvEqrjGxVEpqTSTRb
y59ldev3dzswya6d0zKvG6WhcNBgihJRDxtJ0g5oWRtL3tzP2jHkZtBfQh3Dxyor2QVMmbM5c0fp
0IYlzXoV4ohsL5K/QH1Br3UeAvcBPpYcC10vSvHF8VKqsglEmsMydDnpijMNPcTmsHUfm4WcQhb6
498gjVg0kNMKkgltJHwM1X5lEVa3/E/cCB4Yk/ovg7NDVs4pl30wvJdpAHByN0R59KE+r8DVoR6t
thMfigHvbcE7D9YQv/ZIH64WEPCDJ098eJJ1VLDFCKfSRb2GOCCHrp+G1uhkTG1wKWFE8E/uLBeS
mPO4yvriQATK0dAjf5lczkE0bzuPBnYPQcP1WPNt3uqsh+/ko5r1sTjQC+9lt2WJlGRTntseCs6h
tNQKImdiWXudraQ96540kG7PJpTyqB6gPH1SEBa9TQqmO+SpQ4/5x51KB42Vc1Je6hzetvQXJwcY
4CGDkN8oAAE0lRHFipAZtDTn/1FS4uKZyN6WM2kXybr/mpE3lF+CrhCf2oCHVh4c13KRsf0Z8IIf
tYpculobWkR5sR8rnHmTwyQEngxkbEVbN79TJzw858NsvZMr7bBkr9KgsmLDFCd7SosMv3LEfhAE
26DOu4mAs2HmnNzS1BVzTExerUS0r1J2b5nlVfJ4xUDrCvm71SYmJYmlNdkTKk1ES0NMgSiEQoz6
Q4SEDZchkcRz2myYhyzz4L62ULlDNAEsqwKPV2wzj6ULbNwhW4ZRAGMaYZfMPSOz7z0VNEZSw684
Q8mx9Gs7E6XhTQcMjXoNsAjDDcuoGeqnUuqjFJ7vc9NSI2B/7EKCcP90xigs2qMEvri53gP+YWTM
byD0u6RDXMan264MT26Ag+RNvotfq5mIjVNEhh1+5Qds41UlsxUfa+Sc1mEWw2q7z/LFTgW3JV3W
MOPqF5JfBVPXZUPOuH2TWh4QFRuefichQPYq7AX0ldBWP5rBSsB+iWXfxT5ZDqSuRJgQNWvPtNGT
Rhi0wl23WOgK7LcLMcukp8/bjhncf55i2E3Xb0XY+p4U3yCVXzJn9Jhq6vv3iCChhypuz+TeSJXi
1Vm564v8cbnamBWEPX2oXapFrs7GohNRJkHjfA5YCfhHcM5mChEzQ5uG1Upikq7UANN4WhhOYlGO
Sj7Xgbkj3yypjKgCrf83BsotiES/gXq4H2CJnfXvY/TwfPaL/fKL2euANfAjkchmjNhoxJFvMdiq
8XGPtBwIYNojBYym/g3KKRe8u8N0asyZGxETyUcAff5uQQfxV1EOT4lgQdY3b8Ylisoj/Dlc1zpF
cH+KHHufZ/JBrbwkurrYFb7dRCJ0jGpb4/2jHJYdqtLMeHuqojwmtwXTXS0Oo1403LGWAbWdn/sg
Rw2T0lkbR7OKZds27P08EmjJcr3nkmSaSeYr96yxj1PZfLjLogVThuEFQ1+9Li35qoapCoCbxvvL
J8Yg9nt+HUyUqUCfIFdkMaynnoU+dje/NwkPwUjkw0/GYp55EAy1G2raAp64b0lujQDXJBNJr3yV
mlzXTOfYUh3cCO8/f9RgpynUGH4cscMBTK0/bjgYEVe6xYSA/mohv7ToJUmFNOIy/IXidd72tGkp
MT+tBgwWQl1mfLU1Kc5QT4qjriU7BqpRHScYzCFLIEnG6yb7UXpZ+4QOnNCQ+srvRLOePlj/NzPF
yRGWqmEpyXLmFD5Z14UUDHIBRfisDx3K7gF45L/bf6MJU0OwLrzXK6TGvtO1uN4ZdR95j5BeA/WW
IFtVFaSZ/CuI15J+6u4Fq2KHxDB6eS9+QqpxAm8iABmRzuIqAhKRDmQqHbHghd1fHLgYDcGvd/c1
9317K6ycYng6kLrcQQN41Ni3S8NUzb/JeLqQL5f27bQpaA+ryFlct+0xquGOAWh2clyckMIYt7gV
h+g8WVRmm1CuULDPg8CwKp9rLVSuQJRkwQTUTkseyvRI7n+ONfx5/4u28n2ZFAjRMDitUdw/Kwz/
L2EtTjO/5YbTO4/iBNGH3KxZKvZ/UPJECFZSsFiyquebwhNa4tfdSh5pa23m18fmdacMLDsMeOh4
kznp5YfnluNimzfKqYKMDo0EC+WI6C1eSFfgbi6eakUh/bx5UhoMcgoVkdXCRyUNP6BGgT1ilPXv
f+nyhIjQLEDRhWIBJ0gjnqbWARAFJEU+igjoBDuSsQigdydDUXp1veI4UKgJGilA6OOoY/FZCj4W
hkMEQuFBREselBwWJE87WarGdWpEtoxtAtzitdQQch2GLsIilROgUtpd35wAUIocD0pW0nkyoFIR
7uiL8ld1u0KmgyA9Vz5Ks3bkL8CVaXmkxWjPcayAXqkhdlA4i3dGYX6CgcqSI3qUBk3JKHS6MpAn
TiJkqFP8NArmIoX3WPemp//Al++FOPSyooi6q6a7QvMAkDP/AUS4MYUfX/F0tyTGrLfn+tUUagoy
TU1ui9T3vovmaywP3II6DZqkoln2+9O3o74tYmZNUG72g6euPnb8QA1eYkg29n4d+XTPWuG7Ws0j
fEIqSi4ow12sTytKXL7OXLKi+L7BgZNe8ywaBVZrmeFaY8C/g1sRL1cABaiEKIgLz7C3kvA3zQT7
7wQU9Wne0GVUJrxaujhGzDh93/xltGXOhP6Mh16DX9lxyjp8eZvd6FGTSj+v3yTBolC7hwBLAKGh
aNz6/EsIipJJdIEPxDG/pPpBknRk+E6CUsqsmqbDazzy5Fz8EtV++DrfFX/Wjvnc95vIUEXoMSxi
XNGQszQ8VbWUBZjQfBsh+SdNAFOlSXqnr6tzL3KopSB9IKK+dv17ecRQ4hWtF2s+v70bflTUBrjx
Q7VlUCCfhN/1AD4RMODfu5f94xOlWgW+tSSLnhYNqCI7xngBudn2Px8NwQL9PvuD/YHKoNq+PKt1
F/kCqI2eg7DLmeC7WrodoyPp9zHO1LGCrBc2jVUqkajUxZQXK4Y3OESEdHYPSatsIO8OudX3EKeG
2MuFNNYEeoCbP89HdDHn1YAaHGpnaWFojZn1BCYGnzQIct6TSEQUEXAvW4nekG3RPv1vuRW78C0N
IAPh6huCB8JHLy34s+Rh0ZlFcRWFjX8TQwtHMuwa8MOFyiNWBL3P2sM1SQjL8dUsELT4xfmwvRPU
vJx0kn7gNHw76PExlpEafegfBc5gHGPdgi4PR8sCuGGl+jF1xbtTnttpG5Yn1DiirxwsQ83Kku7m
g0MmHY8dwkgmGyjdE3sqnVXGVlX2nptLG6OGXUtuFWqQ2ky+n2mbmPpwmD9kMU6e8oHO6BDFcU+S
YtmiC+0OjXBec1P8RhF8ubXm/gDmUk80prfKid5IfxNfdLgyST+Mpk4A4oPNbe2htmR2zjodnl5z
6AHW0Feym4AJB31lfyVxX/XuRhgQLusV8OGiPmMWz2GUirXt3Qn0nCXnA0T5zu35eM9xKAFPYL6W
TaZyJ3xNxdS7qfukW0E5OmuulkJCHkx+rtp74h5OkAk+Likh8P5YB/+MVVw/PGOkhNk/b/zGMgHb
B+LoVaxWP2zJe57SZ750f7a47LzH5+MYAgeVfcV4MG3BxVVPZIeCis+zsPhPQy+Z3ytERQ7jUejz
rrFxSe7KUiOCWKR3VbK0JxU8jzAJ6wy9RsRrGradGUB49Rk7d48wh2YY+BbYzbTPvbuMgcONCYqx
rj9N/oxUhf1DTdrbnxQQivjnBq0kdgT3ukxjXWrg/LV98dcQ2SsrYCKw2p1q2bwd7jpsIipWygp3
Zo4Pwu5EjrHRpQ8CXPiBaPJ/AiWIuS+bkAAMpfacz8EgAdu61lL8gxOdBW2DI72pyoiFjTsmb0B7
S3r2/qaJE/8bnetIaaxQxx07kuC7SVW59tFI/BDvbZps2FkeiwMRpHZUWVIewzFr3sqWHx8xHM1L
x5yUSUz5A+ubbNCcuyfrLh0NkNjcvCQ+tuLj7Ws8rIfrDrBs2N81rRoM/Fn8JLBobeJIB7nhLVj9
wHAA88RjCs3o3ZJCgZ84dVLScIg+kuqSeY03IaTy7O2pJyk6bBsEKj2XIwsvL5mTPboB6K41qbVj
WIN4XZJnvdU5llJnr/Rz0vqi2za1byvUPpbYPaNxnvNIBW3+JBbj0LJqbnXckZkTkVz2btp0RXlD
C0bxfKnSUsN3/wyX7LwA4sbVBjUE9FWPh/XEI/JnVLzdXjx6pp2U+7n24VNRsEAVuqOmWSV49Faq
iLPJjikDwPeV3RDqCEZFNq/oHlEBBdaCIk3spyaFWEpfZRX7Dlv+rWvRdNBGGPunwNlPeZBiLArI
Miy+s0OP9p0nltw15N/EDiQRnpDdUu4xyw8NqpYZmdUhsIJY9X6ODVHIW5sm6BIsnDxV0CXN9vKv
jbt4haLHRZdpeeBGiKKyx/h7yHwwA3PuaCfCrVas8/s7c7BhaRIg8dA7EuDNFqZJ42q/OwNtpzbL
Ux78L6Xlp2qIuYJOIlOJs3wRKjPykIQ2mhdMAO/cn4AvTlXyd/Z/Agyu2hQ0T5cwXgLj1pyExZT1
Giebcs1V9Hm1wuOrNhhwRurkR7ZkaNoiGAss7VeXVqFHi+w2M+gFlPXz9ALkyc4xJYxvH0RTNfrO
xV9giQEPCt5aejBMXdFO+J8a0m/2Gf40yiemHR8EGSmlGAv/yb1OAS18NgJEPS5jn92yU25TrF5G
jgoaVjalZW1BGXnKRlR7FCmi7YiyfY+wgZl21Gv0SoRXUiNgMtFp4bSZzTNrcpG6duFHaqhEw++L
Sv/wabVfK9CtoQaYyZE+LLuE2ojzHTKqc3fADpR6CpjcU/wsceT/eeDS4P/m4yC9VcY9tVn7WeEW
uHKe16cwoarQP/Vs5LgqFw1cNf522duucS9ChfnvZzab8MfxzYNzAOvsYNNjh1R8UHgUhZQjNLMS
ZrsCJeOw6rNGkfQk2syIhSVgEmrHc2kvmhEPCPKhp/1b/IFAac1zKpdJz0aWvORIfbu/O7tDzZ1o
7Hlk3Zag/HfoqxtoUH7Ium6jAO6aGgLt5lzS12mdPAxWeeSOLGdx42Vh8Iitb78dl6+7dYi420bP
asufXdv720BKzSBIEuMjm/tWbbYl4IXCBA9iAzFbue4w6hhME0MhTTSE2KkgfSReBo7Tc0YTriSo
WZ+w3rKZy+ngcSA4MY0W+j8W0T8vH0R2XwJdFpjmQth3TyqUDSGZp0bE0CrN0go4qPt18N6m9t/2
bE5OUuQnKymyUDghPIr52nU/b+o25lr2KFb3TQ7NyHz1y5wZOzcXziAnzY+/0zEnCKoUWHbo97AN
2FDamtEJ4G36rrzWAXq/6se+nN8AGhcxG84bvuhJjfaLfUQL580uQfAa+3tjbIs2N50ZDwnwNiw4
TNcaayin3FE+uHru6dJt3ScjNmodlWLUeu1rRV+HclwiPXYV0X3yKLUA1RpOmH4R6XkuhSNlEwLk
W2gpQiG0F+AfNh7LPesbX1oEGbT0fDOCEAsOgPOS+K7Dp5I0NDk1M6VrKJJH0lx+k2cKYtUEYC5z
gPL1+oFho8fqcU1IJzFANtHEp2/rnlRtPDgFwYKagEsSWkBZBZxsH25gl7owfPva2/ZfXSLJ6h4e
qyoo9TVIcdHFs6LXd17lW8SGI2zGN8JugssUxZcS5+WyACJbC/mLLbDR8doEYjU2mlkuTD4BH8xJ
eTiCc6P5NuxiJN7gejzypU0wigL10G+Erp/+h6vQv1mZ3BTBVO8H19+52QogpHm6V7rr45HlMf5D
2hI+dIM9AH7Wccd3QHmAZD+m1oeMzwo32TU/nJ85ldBAUBVlq9VsQpCDv44+eBxoib9Ax+HaDU/g
kGnWlI09tRWmfmyXSuVXtOqaOnZnfXZ52jLIg3NHn6+TFVx22xMaarwvKF2LlswZfqYVivL4ECtd
9pTQ1+2UsqJNkBS1vjYvdIiBf8cBcvhrg7KnCS4J/muojooj85fDs9Si0bGOyKQPsEPE01XAcEWO
HJNOhW+svTxUPNZ4kSAc0rFRsNDz0imZDbQdOHXdkdD9aeSOA+RqRm3e9kN21g1XoK3gJbD+cy48
n6W0VRX7A1JBfbLLIWIZfW1cw8o1H0UIaCKhHybMcFZWa6hzUS/YcoJrZqI0cSt8zHDXZ0lI5PVR
6mtZODZs9I3J9E6TCE9tVrZIITpedQ2vOJtYAF4dleDKMJt823EmCekbXNoaYll02rL29hxlZSWa
DE0QDD5nDNevPvLeX1G+zM1QoK4u+M8OKjz9LRR2uYrgr+kptpjX8OT28HMABsCyUhu46PjI8h3g
j5dQzacJRo8HXgPPhxXv9ixLWdENOkMRH2Wux9huPd1ttU7HubMXj9kWg7BaDP8megfLBeZ6i5Ym
n3TERtIfZgreiDY1Vm2VetTl2CGCrsD1QqNiHNlZVS+vJSvvRGlXRIF2cxIjDYEKckqQytxZHKMv
5ZdYl7XnTBOSvdp9jo6RZTyq0rFBGD6dxO4b8bBKcjuL8epBU/whVRwzfe9Rbrint4A2hBD3CPCx
/8hDIT1LZszJiAix9f4Z0DqwbxCvpUk2pScXugdF0JtLn4v8u+x1UChxQprIu4TYwdCntwlDF2m7
1McTEDvm9s611y5SxIjoBh6qCbDa2/fmn0meTIBHeO4aomlHY/ZnGZECW1d2vpcPH6eRT2vYpkXa
RnXLiNi6Lp+0A0Qr+oKOK4UGwlXH1A4QzeyD+gbTBsEKlpAdNOt92CE/ELhJXLCaVRe+3+pDydcK
P4OsnoO4IZjueOSlagFQBmxURK69aJR8MSzNt+UwbZQHVloXQAXZi7fPU2OZ7sspMB2AyOFlNZzu
iJ0T9mqPqgQ9NPQbu1WKhBKSSv4CBOo9gWR85pZzkmX/tIERtPNK6AEd1fZCR3VLxhfH6b5Ak1Rh
0qQX1yMqspnw1VoXISezwh9vgCPhtx5o02wXJFTaupZ054KBKsaK29b4ps/xICWaohCeCGd7PBkW
smC6IDhLER6tCcbwBT703H2Ng9rD4IVotOOe92Nj+Nf8zNGfy7nFLxDuou1mXTmOcAUAU0ppZIOc
lxxOCX+4OEmogcPoh743p97tT18MM4Zy8H1DF/ri1tkV5VvonzTuCPzTDoefMtEP5MNzGwSdQ/ed
fSTbzoaJp6LyR5pPoCoY/ArxinxqT7oWNA4JFm/n7z3yg5Wiy/h71GXvApFm2ZiF5vZ64KJeBt1+
LpQhChaiDguKmR87dqgDIYVudJRw69WGc+/X118s/VJlQ0PjoVe//WBPExk+Pwqe+pRS9HuUNpQb
yPY3rEDz+LiUzayHgZMNjwCZDepTL4naSV/0w0cQM1HJVEtkwTaf41tzZy6xwz3bdEwIzRyUDhlz
8fBzpKo0Z3H8MOx2yEowXuh2pHDOvbg2EGHddvlXXk4X694QoNakNul+vvPw0M7A6daxJmrIOVnW
3ANTds4erLY2t4nFRtsisYeYN/G8qumuBAYLMD6UemB7pCfZQ+Ia2YEys7/Z7iNVHy9L4v5sZRjg
z9yeI8Pq+Rt4SADj+ujj/KTJ+sNLwVBpMWfxq3nCddk7cJ7QYGP9hsUPqehJmShxPV32rx0dIjUy
T6He0O63LoQCJf2qvQVZfePMMAbxCWNUTSfx9pb1qMwpwYblYaaC4iuKHjISY0fdnjrWuK4bm+SH
D81woGW/SwteFXy+1A+8/3ye4BRdvXLhX5inodevCpLgDgFPGEjfsrZdwzGgu/e8OAJg9fFCJwb3
4CfeRg8KCfLAkHKDdv8zlKPKJuqokTOSn1SF4jCnnzMJm/WysqBay33ALpD3WBHLGn6oJ24KO405
NGJAclRDgUOyykXlnuqXEPW/m8l2rUhbhmXlE/mGUkX+QdL4+OlDX0sLhdVfSt1Nu19WIvqhkV3t
4qGkkjaiPdLEhiyX0+FWHsgyNr69SBW+Cs8+oYIlDkAHyeV7B4EX4NnXJsTF0/1uRTBIspwdVOv1
GxoVFXL9PTXWmGmqJLaKXET0x+HKoe3D6CjIaFQKB2HOU2NCRfIfu1fMUrM704RJYpOmQtpHxF/G
CKryyxfMPSNKXyLbwIFVHJ6idjCRFSn4XS4YumIWAQWGT8/wPIiJLeP3qe2WstKyI6cf2/dn5t2d
K8qlStBpMEdBRoNHgGUSFbUz8/ftBck2T/vXW+mlK3sGKHAzBkn/Ecbrr5g/4mINLvtro7LVUmAx
mp4zBjeDAsyM6+BsZB0MwcZNePhtoYaJ83qGNp7aQfW8+GP59xe4QNaLU2PsicgjkJL1lZiLQMXB
dNBdzUntdqg8UNPbPI75TN8lnBsNjX3e+v8MR3fDcPg6SX3ehWP6oXARXsNJwDi+sDa7WC/0cCuc
tMRO2R48C9k3uGUyjikuExSE4tq+wpDv4hBI+L9ejHrkSwx4sbyYir/P8TpXDJbSoPUjcPrfzXzu
jt0afS0hwRppb7T5p2w3uK9R+uyVdvOgQyCrPZNDWKj2DQJPdYYPvnz0oADGirm3iFWpvZit5YJK
KRFrrvLhwOO1FNvOexp1tQC1zPHZoOK2UH8zQ2mU4HnPbL48j704D5LzH5RgGfs7KA8eb+ZldQ7G
hmjWFGf2tpULsKQn2gIofOw6j73DHdf7vcpqUTFtxtOwC/dUU2LrcNvMWqNyHVaUS56LfXIjL34+
xFODsviX7iA0ueolzREINC7ZtpRObvo20maRFWAXq1tl7WJs8vhHXvW9E8/A95pda46dRrRXWdKe
NFLks3Rs15ypcJWc+ic/LIKL2VHm1UOSOpPmJsxi38jfB0XX+TNycCX8Za7wcXbYmSC2sLUbuhAY
DgwM5zHnBjqjLC801dfhHiVVOtOHcBq+Gk4rZNcJWj8u+HsBeQfQJ3JBFl7hqrCdE30/TybglULx
meIGx9LcEzKYAg52vCcIpt93fUIpuuDzYJF7ps8RYV+UGLROyqGMlUyKae9aW/gaHHQaBZIL4nwd
lb1wPcBNf/w2mc8olsR8awTbvn2vuynM7XaDi0DWSBxfLtwY2112WzvBURZBO3ODPplU5f5YY2OT
QopV9slSwzh16y+fqPICJe5cIJm3MATn2GjlzKpkGyJ4zP9mOIhjPoLc3O2U56Ycx7Vj9GwdTHiS
kbKeKeOuK2J0q0aCkPRnnc8/FsjRg7npG4ZSMhjmVmpx27EaxEnQKzS0jSP+KFINjmkY53+4ZzT1
VvRsplfsB0eK2qQaoeX6ZAdAS1idUccbNkhQJYNl12Q6qyOpE8QrKh54x77RhvZLFy/9fsgZ4AoX
vt2CD7o1nvKPXXuY5xmuHMltglpARYxtZq3tQVtHYQyJhxYrYmKq0hDtYDbZI4qvxiz9aMwvFEIv
R5SXI1W3GMv5L1uLSAnw8+6cDoY3s0rPMyylpMiqIATKFu706t+nmORG0r7uom1HVDey6EFcBeS4
y+Qt04yyxxZc7FfNEF1bLN1lxbXO9p/rERmkcOUJNS7jNwSY9/NL6LEU4krTBnla4npNrHvrSX3s
NUVtKxE4ExsxHOabzayyqogYpicJzdo6k3w969JCcR4QsuuF+VTmnVZ+iokkifMZEP4McZdu+OIH
tMNb+ziHk35Mle0CfmcUCxghdlf4eTLJCh4+xk1BaN5Zi4+Kob7dLNBuaO4UXNaXbU+Vul9lfmD+
B2voB9nQEJ+/vMIM2fuNl22nQzxP/1PZHYRLItuhdy66t6NJKApwNGq/gIE3nyi47XdYYkxMZj5r
LIoMr7YTb2VOUbSl4FEeqawXUoQidKHg8/aW8/w4KFZNbRTSoeTgT3/V+7f3b30Bg0mUnNx4r+HM
zISr1ho0NKDXQr7cTwcAh7KWV2URLWwyfuoN7A0RD/3oSV2afBGMAVKFp3CN+PQjaBF0EZGofmf+
FasqnRuMeYuWnz6QvrJhT09kXdEIkYENIdYAQxAkOXx7x206MmdKQ7rXqQfYfhxfvl3lRX/wvDz+
5vhvQCXUOrulvqgsd10Eu5ITiwdyV7AI9Tv0OUWG/ZtBay6/aD5YpVtGpCkBVjDgaScvUYK6klqD
sToHpJ66obtnhJE9IWwzyU1HBrN/TWRWDDQ7kbgvrzC8VY/1qkdJI3xqQhI2wiFpT6d2BEY4u78k
bq+4+B14RaSLsmtb4KKGBxeQeL6nZ1MBARwmQUsE7LCj1P2hIAAkxwvBsUAUzQ1kQV+F6WY9hDOn
ayRK8BknHxGyQkp6DVPOh8lvkdPcplqKcGYlsEpbc7lVxw5IHB4icgnrZipIDsIIKIYIQC3rEt5r
gV9j/5UfKwPVgGe4J9DRs5ScUj7Jc+gQmjyNws+ghsQmSO3SVYiycbRDadulERPY2u73mP3c5Z83
WzfmbNqE4EVwpAgHb/Zx9kyMqCcHMSP7BEN3CBNemB3JOLjPG5xY21HezraL29UToc5tyxenmbr+
S6Rq5WfLY3d09cVcWCLGCLAuyp/TbRxWXSxh3/KuneIkVhMgyvbcltXFoiyUC3WKEu/GlCKfUoNH
wHN1VSOtNUjosO2iPlbV0QQfqdikV6QKzpEEQS6xHGOZSM+xJ63FviZL4Z0lDRNSj3zjSC4K76YH
uwFM5sf8JJFGLq9nRl+tC0Zpgy7iJXcGDqpSh/02aoXW6CMi6ky6VsHbuonVkepp5XT4BMk3Az8F
Wxw5jc0ZgudHXZ04LphlvvCpa2kzsKEZnujFBf1f3f0GGU+5uVIHzxRW+unrZPQsJ/0ZDxjAW63X
3W1KhojZBdr7rZnqmaJB8Pc/b7gd4QIuSAtpN31orL7TRm+xJJenT7PNq6+pu0tquYul0ux6HnqQ
jXmVyPHndeVlCWqKOEsCqtcNDXUNTvPU+g1RMW+xMB1mwk4K25vC4NBlirS9/Nl/rfLbLu774uYt
zJqqs5bwSxKX4nSBGDlic+X6wdO9w+MGU/CNLQo7WJV9bECBwA3XTOXqii8Obos7N/uycm/aGobS
cp2/tUUHNdtAsKWoaHZen+uB50/rOK6rsgvIANDvFIsbvcw1YKM5SBCwWfJH+xlMO7RFZfkE52UF
vhmT5LiDPHGhuLpjC7AITUGXeHPVkFrLBcvr/WM1nVYBBy+FLnFGQfq8qHAaHWjoA9AdzhEw+NBr
5MHnCdwX3HrgK43bCZxsMjdxbxMR6uV++i3X+td3ACWKT+rji0KtDOytdDSOsLwnEWJ6qvoamowN
61RRv8wh12Vj1zUbDid6stoksYnWLpsn5kkonvzcDik5R/7Bsatx7Jko3+ZD7kdBiRSbBSSNJ7os
Ja9g0oOrqI6b6ZKqlsc3w9anCEsvLzVNRlLrs9W0KCHSVOT20MbJmQOP1YeqClLqAnwBGJyl3n4O
6hL51/gPm0Y8uSRrnmwBZhxev55aPaoxuop9Uig2sqxdnd1uUGl8yJrJr61Gy3JV7sGclR/tM4uX
6toyu4SaThGNpUjc1D6hIh1SaAKAJ4xRz2ZpAQ1ddxLW+MFmbjZ5FkyrswPYcXgy3CmflsB+N2sB
wClbFd4FnU3cjtZdKw0X5t+jqVLxrpZm9Hm19RIdt7lggnSXb4x7mvWZzNxtYisrJTESn53v85Tx
jBDt8IxWi3XM9w7zS2byVupKzZ8Khfk9zNj8/J4Coyo03oBnJg7uFLOVxEsozMB7VMutCzSOu7Q2
+EdbYXIT8yhZb6/2zNrScKCFMYkB5R3D/lwYcxJRKpiOD9mZI/2mUnX0s6qpSVbCSqGlEsjS/VGi
Bkq8FbhptoChoj2A7XvuUCtkceWN7ZmLEbIFDAbs6INBmPHyJPg7u2B+WdtvAfhqzrhEhSD7q2um
/84RG1odIDCpcb4VFCrUVCNjTlk3Y1AhB1P3dEa/YlGDLz5xa5vsqw4RooZ6oltDSeMe9mrELFTB
JmEo3ZnWI1zV8POXDf6U0vjJgAYhTLQbtSjuGST7ZcADEMCPj4BB1LQD7pKLlFwsEMZpXPWcWCbZ
i2q0YxlCLzwsBnIKxPumGh5NmopHtSS3QSSyLH3fieRvPsmUHLUYj6SclealrbBqKmZ1+FWnC/y6
ZXd7bJ7LYtkstP+Cglv5N2hcQ/IZ1b73BM1TX8YLoXH00Xq1zRQsXIyyzefT/WP4DN23mG0GEN7O
MZqov/uIvmdU5JxsGfzyrcFlALSFn2rQiqKxg9NVn8K0d4BnrtgZSUBnUg8ZZAqs1E7WkCZdXZGU
0pALaMl/EM02XNiG879gBtfwK9QE77pPY1BJ9P2w4ZO/9fgncHZ5EUqLF95W+UTGXZnOpR20sIUb
f4XBxMhOny/6Ojyt6/JQQmXsUc/T9ul9cXtFO+tyQEi6uvkdQ45YtrynH+ZIfmyBCAUg6X+XZLvH
kRbSi+KCmTDfHYHV4plOS1YCK3pFJJ7WGA7jIDqPOAlsZCneBJcHNnMi7eFSHIiuEprkJAQQKFGn
iQuwgiaxZZSm7g3AOSpCyl+GTvYivIgxOZU5vczmCr8Y12yfzJRYzorqkHC/9DXvDyLLtwjhlJPf
PI1DXqhq/JGT1JK7RXJk1Phtc4NWQdgWqKIB11z1zf3C7QQRH7Dh6MeMdH4GOPjfj2Hdp8MijEbR
+I3I/bW9PRGmVvsky6MjDfgiRz9U6C6PuMYJzKaMSCR4kj2d1hV8Ooorieor8vgFGYar5fMEsndE
oj87Wik3K4MEiF64wIC4VOhiRewy22tDPKOhZvf7kJn+oYLuwe9YR+IRd1z4cyr9sWeAcu+C5IPZ
jhCihiWsInxIHJjir4Md36DGhUGk/ct53YpicmukkojyQ6NsE5K3VgaCIw1XutMzzJrz+sdh4G3D
LMh/K3bO+fZEu8QOlvoT53Vcavgpx3ONmvwUFEmAW4sJL4HUNzmizxf4vclqfD9k8XZEkDyvOUec
wL8daI1EJ213jr6+cYVonMF/UxAYjXjfoXNHEOlfoOrP2zc0crdtv2oI1BxWUFch+Emz15QPlZ4f
jB2iWMZ+kISRC2cpyO2OXc5L8JatL7XYQQCsh52TukPQWHYShF/UjVwNwZpVios+N52EOJSe0+Gu
Mju6GMh0XV6WtU0MnzGmsLb5xQJSc5iCaccIkNa3zbp2MsdY2eCrM6rkmHNyP9RazYGUVS/Z9TvE
+wp0pIphcfynlhy3ik/nv8SEDywKaOmCPeI/JSKb0mt69Y/peQTofU7CLdRFPZsXu6TtZKqkNM2S
39yNV0NFwgS5UQ/BwZq9sDKh90A48hvX7/7PlWxbpU9RM6sllUIHPz7fG5+oTv3s28IVi04Qgrx1
8zNNULnG+C2yNQfQ1X2P4llcBu/1byBcrGkBcWA5YQbeTNfMrfxHJQZYLgKEgvEtUSgXnXqWSbEV
holeaCvoqCN99xynL0QyEpn2okErn0V/F5ImlW+28QxlMBG1JFtOnadjSseLsnEK8ien1KOPMaFo
37/0y61pqscbGw+yrzh2QVz6sLxuLs0Ia1V8ITiAlZmvahLj0oYuqtsdTBG8X7jz/v/Iff/r7OpU
fpGM0iz9YPaE+mw+6Zt06lxRC8GutKzLjio+ePCyUieLBz8a026Aveyl4Ir95vHqhpeJxOmE/YyI
NJqmdXT1jyGr4vfaiwL8kh4Cj6bJC1nQVktSkUSoRCLIbbjje96hCRXI3lFX6PUJViOV9FXF1k9l
rHQDydHTJGLxNB9ul+YW2xeqRLRcw+10oaUu7WGRn9AlDVqlJtAHxU0zdPs6tcVNsH+0d1b7TolU
xbaxmIHvn8WRYuQI50BBc34334ulHfteB3GeHFieUXsBKuvJ0Psze5TIMmVZdto/kCKuUGDbWQnw
AILhQdrOdfWnFvUuHYREEfoZ2Rk+/hKeJO2g3DYapXKIZLhC19A7xO/NZ89sDG0wSJzm2ga3SyTO
DeOh5NZNMU9RILyl68CI0iKGFudmhDY/y0o8OkP3LhIj9NF9OCovz4iEshIXlrTIA3l2SYEEbNtb
t0WufTHPzu+fmFt0h5oFKpz5SSMKSIgDfP3f2YfvVGMm2mPJa6e+AjdkyfnADS/gD35PpKHompdS
BfLOA7A+US/SP5DrSR1NTDo8RYT82gRa1+YASsrohmi33fuKg/1cPrI/36pIhICwvNM98WPXF2/Y
F0eyr/girwg8SvjjRY1j+9HbPwajkbixSK9PBq/fghwQuYZEp0icpHFnU+dLWB5VebDwcc/eLDXV
uP4+wrpGOcHy46F0akWlR6UqhZm03LfYUFnSTBGAqjmCkIwybHA5AWmN9AMpYjjzbqDTjSXpP3zv
cmjvzNOwvTYaOxOoQ+f63evSu2IKnnL9UBks0z+2OLiRe9TYlNc3xfcI8y2zJLvMkv5OOtMIbPH2
MZnBEXFRVJdbBXm9nAKSY2pERNf4eepOJ3ifYEboAj4RtquJDMQ+0cxFyTjXHmT+19h5WmB6Cmhs
X0wERrK405nH9Neas119eBj4zqY2lOOWsv8nqgEbary2TYAQ0F5RzqzkoOacWr5ELPClnIOjugZ2
Zw4d5USUW+4DyF6khC1Fz0G3DmEKhTtIUOuDDBYdD1GbqQp3RnlJMzkerR6pU2SRVQgbUdQlte9v
aIdSNp0/tutsuSDrtYLwC5S+PzRoChelAgIurwFfmP9pUAtngMAmrBhk/HYRB2JOEQcgr93cwBfE
F11eziTnMbjdnLJJGQ6u/fDD2l9NbBJPDLWkM/kxRNkQm5VCm955nYafyMwafXIQOoNskBmCPYK8
yoAGHOP6xJcUtOoXfhoddVqvlfGcKvUh9yc8PI6c626B+RThK29MrHCR7t2GZk0O2Tv7ZWpdH6hU
35AyAS73daicvNcK6E4e6IUeE0xAr+I7uz7D+EM87y2BsKdCbtSr3M3q2UTT+sk6nMR72hqurAf6
pGoxk4ZRcdc/5HGx624eyVtpTCoANfJ6NLGctrPvByI/E2wxgOnvrbabmMpwG/Q5FryaN909gANO
kvk3DGHndKiV3Gblw8IErqG0Lm6J9U+F6U1WmkU7I4UpZ5me8K6CG6wDv3yOzn/gQBqr4WwU/8b6
gAfcXQ7jGg+HSovZ81Ynb4Qzozd0H2lZWS5pftByUe/PDm9wSDXRPEgezkNChNfL2j4LkZxVRzsz
nPuVyz45X/Awg7mXF9XKLGZCHn8hb3mJap/84Ut72eImcch7NbP+oDGOanY0j2l/Mau3AocJ1Hfw
GC1yJux9HrHPc3Ua9M1psfiKUFIEsjJN7eLAgxLtp+8xZSVARVO5qVo+0DjLK1XF/PJaQIm2tV4H
uys0Ezz5yA7LUhP1YYy+FXoNKrxBS6e+U/gXkZ5o+wXyx/qB8hwJ9JoERbOcl21cktP8ONHP/lmh
0/tks6JMk4HDn9I+TT8RrLBdXQH9cHzrr4Ks+2NXZNH3TcuHdaD5wsl5zo2ksDrtHKScVrJ6mnK4
S6XGsH/HuvqSoQhNh/fbk6YXBLWQZ/miS1+E0GXxUbI9ts/Ox9ib1jbMKl8ZugNVZSkzDbMCJtFf
sgQO+uIp21IFEYwoPrcH3O8TvXPLhvIzUCQkJJ3NdU/3ou0Y++fTPSAJvaLDWTr5ftxWto2jMTFw
waDgriuPbegBbr9OKSXu57q2nAzmMIIsxQPzLgUIgM9qJw5lqG0ykbVjfwVPIwwtPNA4x8lxQ2T0
Wgo2OGpl83xBW5DpcoZAe3m9N/pYRiQbayQ256SgpVImDcdTz1crGDaIphKMFxtl5RB+1+DJRClo
byFX+wpxvKJ/0YNsWppmLZbHoylNH0PlfoTnZ4kt5TNHfCy2CDD/Gema2wf/O1n96A+cgNDVKMkN
W/TvKwREOmbu61YABv7FPZGHriedySscRof79TMlK+3+WpDLTGQFEEF3TBlIzt9RDFJprF0NfdxP
UjPSCR3LBdrrQkdE9xT9ERpZd+ORQbHrYVnxrI1zMXqktuZLtz2DGlv+imzN20fo4z02lCjgj1rF
uNjj4dtOuZ/bPhMTtW7sc6suwKGT2MkCPy3r4FVThtOyWOViPwC00E/3nRRCD8FGrvq/MgOV4jH8
+ks0e7chfFHsJ1J6RMa1TecmjE6CJcLEKwSXAZG1y9utIf1Ba7D+HYc+t+NolLjpWE8cgl3k9pGS
7QNwbVbWSqzCPmiM0+YmhJ5s31UGEDvrZhddUlsWzx3Dkm4F2/yKeZMdgORpbVqtY/miYoZyE/ll
Rar4l5qTmVOCrqQE70G9D9NVzgkEoj75YnCLlBdRaomN51Te+SB7jzUQlYDSen0XgfuZ8dtjSllu
c7CJc+Z3jvMnQGaqWcHWYKvfjI3o8ROCj/hT+Qehz0k2FFGLFOefayhxQdZ5gdAuLwvWqz5UwhW5
SEEQszOck3ovQ2XJwsE1GgLJNQqvZiVpFON177kt07lH05Yx0/6WjGxU/JsRTkGAo3jTKm8NSEQa
BzNWXS81h7u9i4AuOmSklnghFKF1mDDp37NTZ2L24hCpsbtA4B9v8s1D180lgD74J0i4t4N+pkHq
D9Ipwx6PHWyejXqAkg6iTJ7xQgSQxxPmWONUmVwiNbjU8CsO+w18kPbm1m1hrZ1kF5vktfNG+nJV
cwxqP0ILeNn35+DgXcgtmPNOVdO3xn8UUTPqwYCV2P2JBqu5igySSDk+tmeasYAMW5xEFNjS5JEf
8R/yFaHOCON7i/WEY1G4QIk0GGL3+3Xsyi9pxoB7Da/OO5xv+A02hdproU11oVZL0HNbwf8Wuc6V
MFalUQlVI7qXX8FQeCAu3JBNK/EEz5NiPbg5ewCdqwn0VxxKTOyxvpOuLqOVQqdI05eTS15CH2GR
rXwh3K2tj/fP3LnsOxgrwWiFrqJ8rCTp/kHO7OSgyWXtI4oU7JFMUwiPRvmCGbOFqqe00UpGfCel
qB/PuhsfIZZTeKHM4WGjnAAh1dIrik7UpCxYjUMN9kJqJI8baI68+BIntQa8zGI1U3yV1cF/3ufe
GoiSzXVzJgs5drLAFB/GFZswY6OFrmRCLnkCJIW1fDi5tGbd2ktsJC3S1rJdrYKPEYF3ZfhAGYEp
JLDquXoYIhDcvqS29sizRwic5vPH6BHNxRt7zMY6Bzi5QW3cdxtyKITmFlX5Q1vNLSDV/W66sV5t
syZ8fqbYVqqAq0p6XW1ovE00xeliL0fkvALh7Hrnz7JAS7j9ASxuwAJJuC/r7a4ynQY1fsQlrUgj
viiQlJFzwhCX9KEzU0Ubb94BM0UjbzY9SPQP8s/ZRMiW6XcLrWV8mHoZkxZjiCZEyJxmhrRt+8ty
yqBzL3JStzDGdFO0qDhkyhsqMM1naWj73NHQS+Ts9DJXYF1vhtW5khAjVPPyQNRn8P0IelVTGmD0
uA6Cli3pjcgFB8Uhg69NyrxaBgzMdFdwYMhcWtCWdSxlDjljyXhrMlc4P9B60uTIi244lxbIiBul
EF7Lr9UOeIWhrr0x5L3YPmh/QJtVBZLHBdyVSourhYpJKUmWz3tWsFGc5imBTyANz8zSNpe/gcPc
Uo/qu67tH/JVnT5OotYD9ylL6dOULgjY1P3TYXbAoGMiLRwP+qNbZtHLWQ9qM6XoBVlEnR95DHO8
4YyVAGhZz7Qjy+zMb4XcRk6uhKVv+S36UCHY0GxBhiWMGVB8BlBEiM07skK113QHXtr3s4LOEK7z
GIbusMkLKi/v1nVnXzQt9Ws03LZPDDAp67yVPOEh/YFJ9F7iPo/Voe/8pcgbEOgV5537/FT/nxi6
MNz8UmIIOHXl8vDbRY1UrZULfD5encCp2NaXgpjfBaDQN6PsSENWr8JkKBm9Lp+IfECyUEobptwi
to3m/QKt6nZReivFZLn05h8fEdXc1ZUQ4qVd8Ct1ZcE7dZCpgqeuJK9YLzKkQaulxQPRCaGF4/Xk
48NJKL1+A/iIVJyQjf3JVj2CKUdimOC2kurOo1CCuYUaZCPgA37h8D+ZhDC9xbqAQnyEVTGAbQ86
dqZ8MBUuKqVOLYjvzOG/QS6V0OjcIsBIS5A8GmL4OgDvST/NZoMr2hF78Zr+KGaf1eG/2yWD7MU6
qcbu2l1ws7UUQBIsHeo7ntFg+WzSq3WFnYeYgixs1/2JMIfb0NKL4Jkyj2nua/jZMdL8tUzgL43n
Mm+y8G0FN4F8ehw6OOGHabzym+7hvjxN8fJVixICG5xkoGp/gwGya9uIDBnCiXniIgQ/GkPF3WmA
VxipbFeQ4EqM7UcnVzQNwpeMCxrSxeKy6uVXkvBAH82wB2Q62hf39dzAHPNruBUNZLvU3+ZeOmcl
auE6tXkq3ka0qv5h83qpDBRtYmVJwUJR9av6YtUyXYyle6jfhSP4aqDChbAlY64b7I4nxqOUaGZ5
WIc/D1SFFnGu2Ve2O7xeGqIOU5crfjKrGfVvthIWXq5ZHkSPzBdWVbuAhBURypd2zG+FREhrYEFq
qeAPnE8jlr+2ZoKJbn7FFl+KPAuOi3lOJzGgkPZtSd4sh8JG4BJGNJJJJZSK3DksydItlcYqsha8
hcAj7Ol55r123xl+15HUFiH+/Tjk4c2ch+QNehgDnjtSVH+fM5e7U4lmhHifZhX7+jlEYA6Pk4OR
IT3YWYU9JNHCBwpkmSJkymiUQabdSSWlLIlJlHzV50Ap63fAfPcusPSLMxbQBn49dBgamIxWnb6b
+tnXAbc8iKEYGlaXt0SFIi4g4tblKmcE4/+SuWV5Dm8QLXuabvAxQXtKPVLA42fEjNw1euTC/cQ1
Qbs4Ve9iGfETvKOoL7BR2/R+uQt+4Fmo7quU+NXrMGG62uSQxMXIIagdOxFwFkm0ivQENQeYPFGy
jbX5JzlHEDTHyoWgxRApp98rZouGN18O5fblgOXJ+TbnTSti4BdRwFt6tKsWCtWSn6kDhuzol03W
UGZv1Ev/El3IkHoN76ReaMy+Y/ybCZtWG4oNHlu7rtBXlIk1hsixoxM7xCKIOzGEsfx3aEPdqhZ+
7QUEP5HAh44eJiQt2yOiHOXyj+URe6e72GdDev15n4AWeAMclcTX7J+77fAiOp88NApOjBJKrXhI
zDNPdfUcZLITILiO79pib8XRqLbYyXRmyg/iuBQPUPTLUnw+NZ8G2zLaUPYNU5v5saGlhzAbrZxU
hyykS6AEuUdCsCjySTtb0nCkEiOHEsaukYw1qV7ZPB2LFvb9ouP1ytCavYvEszvjrgFf+t2sAkRx
Mu7aXhlo/bLyzm04I9pYpS3vPcShP2E9OuTklQmALMogJfUjU4TZJ4LqWeaRa3JBEXq2SFUHgy0R
BvUAaszffVgYWxY9cmw7IndQVi3So2+8Eq1fEMGNPxcMqPEJNi2Q/vp9xm9M9yA++wdZfAHO9LS1
WXYKhHseiJWgiN5GzE7TgnsVz/vqoJ1PhbBXLdYZdx0vEqmWNElqTfFuvPpuJg8VctpayaVLqAjp
CGHaw0RzwLhLyuQ/gYyXg+1wGxWfOW4a1jUju4TYfv7fSHjW1t0R+nKjTcBGd2PEtNoj9W9Vsoos
zbPcgDFqTdzcl+wsCPNZaOYxUCbkDq16vnhEBAenUSfFW8efUpyah1Wgi5aAwO3s3yxy/DQDoBIC
nsYvmhJolZuLmT1MioGeMnAtxOhxoyu+ujWNGNOuppEKdMJbJvERG5pwsTnT5hYiLZGXZzHbz5pr
/4ObKUBHSI7wB4xMswfCZMI8SZQ7hyv4BiUXEJrhe0M+DeSxmIM02g7NnZ3hf91ZiNM4xE6N/HoY
1XD58DldBex0CCDu2FaDBEJ3pic4asqwBvJcKfOAzi+WNkgAESD1YCSU3EG40PesAFMqqqlN3wWs
Fay52roH61eHdJZJ6MJjmU1Xl5XZKGiq4xDqXrEUjrBd6aQSLllZuvC6XWUyvw50Ap+nj1tUEuIl
XM9ZvvUKFWg1xJ3/TvBkdJcAL8+49cyfPbUb5wZ2Xm2xyP1IR9jDH7LVYhN7ZFWjb0QF2BYdMr0e
CsZfqX9qxRPnkCdc1xkrZsHZEx1edTI0g301nRGyaXvV+uOtAWUd0R54K799fPkBwof7sOc5Jsdg
pUneq9Jch/7i1hGeEsP3xVrNAtHua3tmYJO7eieoAMCtxLLuL8aEjbgpQFVYw9IhHm+Vpkl3gTEH
HNbfYdt9b4MGu4v2jtfYxTerY6iurCdipQbx68OzLyOOVKyym7OInJIECweBfIZ+5mJzrDPGRyGb
7IQI+cNhMAvFvflLvu8jBOFY2cE+eAeYPq53BccAt1f5Tj2qAIi47r2UtNJZI1mlfwytuT62569/
b1xHFD0L1ipl+K4FcM5bsW/+aERkXZLQpmLWCOBgp8TBq0xv33SCRjZOBrBl8+HEe/n2I7c676xn
Y7TTyobq03DjD4ETnFbspqZHxnPG1evEmuPi6yE29STx9boR4noGKX5rdF31ifPlV+s7I8bmw5YO
F4hJz4s4/aCcQbvlMGPyZu4Vm9+6ahqTwppm4SBp98Q/vqv5djBMtrmoQs708/xFEEuMwY/Y35Qu
TsZA7AwaKuNSe8V7ghLKIL/iXxYALifo4j0oI0zZ1NgNjBN1i68xC6Vc/J2bnDK0rizvWqTJqxIM
VIXjPya10bMzWA8+VBFjE5fOu4rnfKj0rkzvr5igdX/TYmIkZNAnFi33D2qVLAnVQSuj7v/x1q7x
9MQxs1ezBgaTxP0yiXZTdKg9obNJcrT6beQD5kv9raYY76cxzK13cJ2TU6nWR4xA7L1R6EJ245gC
KOa9IhWrTlPu98pSi9hjLjwFO9N12kSfvanMUuTP80cx+UVLa7Xb8Lh5wGu307LLQDw/Bjw25W4G
GfY5BqgrxbuHoa5/LL3g/bcfGmRvbNyEoe9VxhE+r65hg5ghqEneyBnw20DREgQ5a6IPpBb8Z8pC
tmQJMIgENc7oErvsZbJpNrJk0bmpjTQpey54Dz4AeoKDbUu1ys2dNKiYtN+SRtGTa6oNhrK8K437
+Kzd0yCUFmQlOVKLwnRd2s3GBQM5jKI3Fk5SQCOI0LjAfRv1oofE8H51AwptDJBYNOzZt+aEYn4I
K2WB5xdsoNqyFFRRZEZ1UwJvKdBG1GHOLVKnjUNw4cgPnVNIPZHaOTR3la7BP9PjlGTcF/4sxZNX
lhXHdzO2fs4KaaIxGS0os1cWAg7scdEW9egWshocsxcME7RCHAtMoejJyCam3MtBTZY2hy51QflI
dQGwDDR7N2CzJWtkcD3i5QysEKFUsiCIJS0FgdP6Sd1YaCfB+QwPem5yp6aFbWJ3Gp6H+bQS5ODM
huTbwRaEFKOknP9KDevnWhqC49adFq98BPvaO7bcVsWChoiF1naLhSbx4xbGHYQmHzbZNEchRhci
nA7jzMdcRNEgkZDBlQZReWaSnetxNnJj16KlzWOSBa6VmmYkvEICqMpkbuIbOO+cmwMmGRNi1LSh
KCKX5E2InfVuvNHaTvkDR+0YjEbVlqd5pV/yuDfoNlhuvH8YAYQTiO0kJbLDR9c9lhxDrYL3hcJR
jit285hYI6fuA+ee3K/NLqZrPaaTpENc/Rie15zvvgs+E0iKnlSg1bOFHfLip6MhngfewurviQek
Axb/WFeN4baHMEv4s+fPJylDza8IC7y69Jh11fFQQi5kT4EdA927X3g1l4Uv1ykB8XG7SkIKbthw
3hOA0XecTrzicMs2QFPIS7wPleynChgN/7RGqDSG0pg0lcfqz9r4X6xac1znCvbvdS7j9zcBOesp
l3q8dJ34SXqCbUd3rhf7/rmXUA/pbKfr3zGYQYRxnqE5HGx52q2saZ4BDK0fsUMUiz2wyCIONNoL
ZYT1jO6zhJFsw5MgEdKEXSFIwka2U8Im5rCI6g/z6R6HDswEZ/Q3P6bYtsixwy7SikE2/TNhmIWF
7qz21G7JvfDY7mfyPLeVEFLh4CgEVSAipyypp7mTHU31wX5U9ip5XudJmCycsRz1aaXlegW0FQzJ
Dv1KxSUNwRrxA1wN6Rzjfq13W3fjXsfygczujmGIywHW7146ze26B4aybKoD3NSuwvTHlHmU46AX
EP2ZHkedKsZ5vHjPBFPZGIRdOo9GAkXLFRlD/DvEVCrtED1Liu7FOQ5ylxo2LGI+ZME+6AI+gQCD
Mk8C84IwXaKWenJDowP5/munUjjAvyVdlWESgcEyTP8abKOE8SxK4NgvJdvxJWC1YVL67cpuFx8e
pV8dbxLRUBtKKhKzY9b9WqNDLWt0V1aFwi2/HhTOM5Zbe2e/XVqV9v/eRWhmjD4+zYvz11woqlv3
SxNWVamP42lyS4sSMDXJLlo2w/MIimiV4Hj/fIMI4glChqpw6DlUt2dy4IWZ50KOQ1K3VWFNaJM7
CpX3EdfsD3ninJjQ/fRRfcCUsiKoM2/366Qo1VN36bzjgbd/wD4YhSNV97YHBdZj/fuW1TR4tob4
cuYBREvBNhMhWAGDzz4/r4H+fARZX5nUS11W+dLevA8TtJdQ9Mhru6+qwfMF7FK4uy3/PBVNltlf
u3r9wMd4uNNuPLoShNTtMF9697vRHYc40jzOKeEx69VW8cZ1XvGFoH7HsQOeFfGVT571/mrgLvoN
KL94SD356kt8ybm/4t7LtnVSsS3H530Sd6XIIVgzP9FnSCJwmMbIFqt27wuVLQ31zAhxbf+9KruJ
0ggDaWm+DOmkLoYipS7aCBikby1Q+86xmbtEkYU+5VqsqGHR0pFGnLN5BTK8pMaX0qqCcaONvDau
gjy6/5w7kbTi0mlNLF4hnucJKQIRA+mg4rfiRktAIR02sVjQkpdnHFzNtXSocvOBUlhLR9vD8LWN
c8+hX8nD3DLQ2xLFNk7690JXdptcIbaSPmL0hoRnneMU/yZIiSgQup6GDwoovclzFYsiCmxa88L8
9GrXmAVBGr3+IbBapovpDduPTvzp88zCh3GYkjmHOin6LCKhg4ivVqKCOALKRpgShhaD2TtpZ3o9
JqtNGtrbUFIiobCNnaBjpPnvwc9oruNG71EKuT+bee9K9r/MQHEa0O5q6oHq5dxy0rQAo3EslGPl
kjO3+W6VXzvs66MlBVRUQF/bx8yVECSZbDqcgsnzdHIh+wNZRr/KggaVV5WkyM4GhpBb5OYeYVgA
/TV0NV3B68wh4QgbGSb+khc5kEi1X97TjRZx0o5snQMkstkLMrcGOIvVNLQ/hASG8wVuoJOS7MQ0
8T42cz2e/S2Qelpqpd0iBFXesCu1RRMnwLEo4itKL5q1h3C72FcLJYgImiyU5S3Xp29ODYPBdWLq
SO5mfZLfYkQzOOvmocdEEfHA/a8TlqwWWqf+QeU1NzKu9J41MymY0R1SbfKE1dH43zpeUQu2L3/G
guGxlcHx+0/7XM7UWqOYw3ktV2aH0HS18L409Dlbn6KDLwOk4y/veNgt6VbTvpSlPSTm9fw7Tz2L
5XJTbwgw8dwty3pC04W0WvUKd4tU5NNZL8gr8WDq3/SgS12xyHl9r5l3wpFIpk35AppFotL4aaoR
8cxq8AkKwAAVGQohuc1lqtsxEGn5WcGaCyecKx/J6dxLfbneXoLp7XaEYEtolXmDO88NHaOid7lC
h85tY1YEkQC1/r1lypiAnwI7ZcXwy++jE2q/pAsnzTLf5GNk+JqOk0dj6GrR47opFR9IhCXhGkta
WJFBrp4PsDiOAXUuKOt7lNggjhmYe4mJxocflDDa5h9n8FDooYDMOjxy6TcuHuP8I9SllsHi56Ce
z/aPmw1u6eLZeXlBZ86LlVhp0Who7sKPyX+zEhtdVJsbncLljCMfWQs6uRxspBJo5bOJXa+DhJTB
xQHOSvZbliAdUgAbWGplkTWOf8jMiyD0osCibdcfFovjuROzB3ssEUtvNPJaiQn3vaxUz5Vob5fm
7o7C3fgxn7MkT6bY2n2hV81+ffx512e2p16y+60iNlJ/EZOphDqwqr0RBhcByDoi/720CvHtoRBN
tPp6Rj28macEfdHMPpDHKW7/57oq/R/HA/pcDoMHJOHwTjB+kcdqkvXF7PKV4Qj4gCL08hzaV4pe
juxxJ9zt2jpz7ugmWa0xZC7P7E5Dc97gV71pXfU5T6BCIgGNGB0+ZA3PnFP2NwvDhUyonH2ZNaUp
Gm0V3uHeRvdRt1y7aiio1+4xDcezpP9H4Uh5oTdZASIUWjfXMHUSHzvT3E/hV9F0Uy7kPkMxJnFT
ApTimr4ZJSNZysByLv0GYvmeta7dGNFdE3/DJIEn5FrLI+N1cWK1C+muKRjZtnEJFC0HX7bD2c8C
dTHvxn6dRKhQMAV/RUV5vneZbti9a4xvib02r30W+KK1JgbvaMSd5nXDVKl9z7j5L96xP01Tqtj+
lyhVZqvfMaYhsPwagbUJVCoQ8h/0f22eOsfzH0QQYry8D6dzkXIjHQReQw7ydqOlfutxK0afuRji
Amg3PVH1JloU7VZx3kW1hDdBVPPXV7hGkehDmXYLMn/gxIP8WNJuov15Ajlio/aZ4KVnfcYGVKo7
tsWtgFYtM6aX9TGmvUKe3kVQ1ISJnxll11fN8W+TID4S+nLLqZpe2jQ1QOSHXcay8ktIv+DXcFrP
vgqQIdFgS3QEZRYXlXTiZf7uCWWwuEaj90DDXsnTE7YEQFXt/lNO46Qta/CvWadyVMcl+hBP/Qn4
yz9aSEV/AtR/sYTnUD0rVnxGKNbpGwdy8A1MUq1oHHIGd650fAuh+z/aGFK2mJd7G4L/VVnn/QhE
PESIRlM+FD4r3pNkOahRDGB1JPwpgpryLEJ4ufGaFi/DLdcdCNbfCwXLrBjqGSlngAL51y4DBYrP
7QhifpwSb2oUfj8p4a56leAS0vcbYWXYkBB8yYiRbx41pi1qVXXLHycyFlY0RNLvNfhDxKJEAxmn
WL8sfIB4hV2McgbQIvmzLNakb4urupd7lXcJEhadpErXCdk2vQtxrK/zxNo35actT19iKgRFOMFG
YS4CPVmyelP5oR9Mom/dJWUt0FFmengmN5Mf2a6t5el91BVKdlVAS9CYrySWnALF5hFvDFMWtvgd
dTRJRrnqrOx+70rL5odbbSL61viHqpMMNJ1lpi01bzKjIe7lZj9/aa8sVEr4TTt7yDMGqbUYrB63
077+I9kqJUf5q2nOVHMYBtfVMNy2DUInEQdTIhxINEuXwzzsOVp5So30ouLg5q32MnGB0OD/LtdY
47c9h2Oj8jjK80+RWyYe4nX1gz+M6mrMeSvSTArIw9qR7I6V+3xcHqQ1TPwXLbTHcEPk6SP6ZkxW
tBHlGCVy/SFrcDHP8QjOKRYKTqHIUaE1tHiYuLqvs55TypVX7fqQfX62LkP/gwTiQXTdKw3eBA4e
8fMDuwq/upxQpOWH4qJRKMeJHdI5T52bKbXnvAy39riFwS2pDb2WjqkHMjMVm6cs1yiXXypdBjyo
EMcK8jXBR7lwZlGBUiQONaETY9ZoQcm1TUoCVu0qyMY/11Zy7EtPzmKdg9Z7vFZOKD7ogZ5L5rXv
c4pwaexSoRtvKAtASTLCXg3mAaCYD4TCwBZ8zGcbAp3u/MANyVBKD4jdLpooVSUvkfngroOSJiAN
q09elX/ibnHRQ/lHsvZHME/UvUkGeMRLoVhKtoJgkJYIHt4GsFw6bRErke3NY4FefHY2BsntCpGO
MeykNKbffc7JyqxLOqmT17B6i1y+gjcsSN9g6Xq8RZyBVdfaZFUMhByLNw0sejFXCyzDPdplY3ay
GldUa+P/Oe6eqn73ROY1vzCyZGeI0D8nYhQHDfrrf6894I/HmcIlDUKa57BFxXGAPKyMnAaSQANm
jaz1PSfEWmw/nU38gxw3Nn51qXTk9ne4N3Hok66n+FMa9KZ5FdaJMC/4AMs4dq7Xu/tN/8LRcktM
ve1e4hZ02D2OHtenaRl2U7oSo8H9PZmqFFsM2tIa/QN29XdI+zYdi3C1HY5rz44aj2PInhPGtlsU
LJEkaWxxboW8VUZMbZvXOTpPWKMwvrswv6HXUWc/+XnW/T4okKIqAPimRyJkFm0TUBjYM23lb6OV
Yx+pmHymEkDBxhIUB6qerRBbGQN5L511ce4dRiL92aV86c04Gi5FblTjCaI2VMmanObuR7014KMx
WIpghx+26YzUXqT6eKlAxz2qLkO4+ihOYxdWi7cHXJLVsfgK3LyVpMVPf7drh8fODXq9zHE/kaeS
DaBTN33Y2mlpgn6zNefyifhDHo6lJWZMiU7s7B+Md0q5wPeXGD9GkgsWbiWXsdQ7u7pKIuauO2xY
HUltxoVxPLcqmezCvs7LxrB+CNCaMhRtDJuTJS2c3IYDiFOw3nsEGw3+g3H4oqPAp082draZPOOJ
PXOggGwpzjeI419wwKdUZieVItRLqSrl9pKSBsvqd1HWgznIMZ80wIp2BPYQ6+ogoHWrAafitRM2
b6Y8dzQoUxTmRa/MXt12fMFy+XvBwfvhJ8uw8FQ3r+C/q8MsrcCbZYBUQdB0Wj89pCeggv18D4d2
lTLU5kroo6ptO0d9GnawjirRDS7tcxpBQDz3s1eEu1tE/4mGKJ+gpvQjqpwTxVcb0xCb6VYQhBVY
IncEpxe62xkk42B59w2ckZ+kCmEbz7nMNIrTNZ4Z+TO5f9KCKkmWuzF9VRtpjKUd92rk7kouYKib
NH0nH6NrIQy1dd9mNm7vEaWq/P8KOqBUtYjyV6AStkNK55rnkOWO/piCpBQogmedSXeoBpEvil/A
L9t9Z9+tgTUzscuv0pcltV1MvrIlT35GsQXoHDqq4Ky4XG/tbPmWL9iu+tbT9asRQg13qjurNghr
YhE3GsO/4WoUE23bNWjsQOuJoUsvYnJkH97lcaeDhswr8MvhftfpWZ1k31j12Jx7XzRX9BcnZpyq
LIsysK7uzhtg0JQdmeQ5ROrWrjBTyj/6QTG+3uSCwCM2AV0rIto1k0hNJ4CA8xmA01811jodRnMR
23Yw7irNVVJq5tPk+aKA9coJyhVXOqNgNkw8qm6IciLrGo9EYqHFm7v0xWvl8RSI0l0T8TM+HbVB
hsXARCJgMcloLL/IEwgsQjwW3egPiZQCghKIPMRBw1qO2+sxri+Lub6ssiirbLTLrPC6c73fYgB6
p6uZQVR0cVYIiC7mEwvWHXVCeapYZAkc+SgF6WGhoDJ7WxCDykssNHVKdDu+VJFijB0CtAHXon3Z
vERjdciAHLcR0aIT+OAJrQ5h0y1R7rtSRw1BeP2nyR8G8VrUUFC2auXaZgCu8ZEVQR2qZZ1KgmJI
f0fewP9VKyDh0IFoAf/QwLm/m2S/q5WNxaAwcnBQR/akTIydwFX+5rTmNKTz+BpVE9Ns0rhJJtqk
6xV1uuF5pOPf3I/MKqbl/xcmijUkNZRofAABDKXfrp49bDrm0xHzH0TI6dtBtoaM0+VXU3X1aqF/
lfr1ekxAvQcgOJxZTUBDYaSV0Bafd0VifBL3+fbSxlFmop9PYEZT8SRTmIn6LYE1nbESPBuPrvD5
YfeFpX+gDhQhHp6t/WaxCgYo1ihKNnubRTymKNCd84X+iKEILbwPoFPMbnkqrI8kWwMduteyazXN
ZWBynmBu0lr3Xh6G+R8dgdxHJvGhq57YoRawVnuMxuveknQv24BG6NCx3EajiytLIgYO1v8LrZwJ
yVyF+IgvCn18Se8dSq5jeTlK03qfKPIjvZd5MnBe153zLzOADRKhAHk8JwjInPWbO5bvhP3TGgEO
lQ3yP7A/KZnmyGAiQr3vqOjgC+Q2p+eD/O4Cr6o00TcEQooBhbyCi0IMCCt4JwrFa5aTus2owCgf
bGq9mJ2PMQfJC7L+2LQfuCLvc648c7cX4bsMPmXtbn34t3devKrlyFZwV8N7LBT1ms26w8A1e+2y
J3EMZBR2TGacmn6k8htKhdtUSJsnEByg9DdRm1by8PrhGu1IHw0qmwsUffExlUvltJOgXqNtSRhG
2wdU2SQFDmjqgl71WGkPmobxni0SPc6sk0QD/gV8l/ekzUBWsGF4iQfQ5SITYaSdBFgiP22FF+Qx
VVkR/3VV2gAThBYG7PkTk+Znd/QfW7pCtYx5fD5sJjzXMVJx0KehdUl9yC5Tnzb3r3UfSB33/9So
DWd3BsyxfseOh5h2UvDkIia+ipd7rj0xEFN0KTlewtMiSZ+aJVgphoEejPTNsRtvwnEergbA7HWZ
c+/0ESCuptw/utHQMWea+ny5/YPBghhe6mIEknzdnT6v8G86QGY2bvuqsGDu3Klu0Z3QfOTuq3Bb
cBwBxDd1YyGrEnMOhGqffzP7CJpPd4xiWjIFGevG9tXu+ocAj1FutpngE+EvS5tz8CymT197KXVN
rl/pOnlOs6/T2/UaiA2JAgf0MPklqygMGCFs8KIocqQhcrT50zT4jl2q5DV2fDfksFqoQUGu31tj
bzPyRlORo76YqIPXUN/WFGU0Jq0BnwtwwIt4eTlNx60mfNLQzoe4valS++7lERZtEI0GeKUEoxW/
+3akU2cyMxKKBf72wmyX/3oPh/efL/9JyDoTHbx1vYgbTrpXZrQIuC4sHdpHO6GLcvEtU+OEwF1I
rfkyuxfatLczpdp0Kp59FdMbG9J3hWdaDFXQS1998/j1enpjdQNcdGkCr5JZDZ0KHxM6ecxOy8S8
yAEY0O5aRdsZuywzEeOQSIuPgx7jkXj7F9mOO3qMnsgAjbT6O/C7P3yrkFK0bpog/k5n+46aSxq8
jqQADwVcBFf/WsZRNEp8aKEwJ9w5TGnicQh8BwHs7iFgMFfk2eNTFc0ruaO6rzJaWr7wftjkqhnV
LenqflszwvXEh6gP18MU4ye6PleX1kGUGxefJTdxSpyd1a6t428FguMEuFNioNjK7ejPq3ccZono
s8hpko/i45QW1pS+UHM7Ddvz6jCoOcMl5TK8ab3Z8o2FZwvaqog/hR4aI7DwqDG5vONgapkEKJf1
1gZb7IQtC37RUtHbaBGDv2JbtmpwZZ8/90qOKOUksjiLscw4vR7L+/07sIMEAqwqyn38G0nLWTeZ
6aOENizxFepDqscSxMLaAjY7e8nFmjm58RS/0iOxrbI4q15WEI8wBZFI/WL2EztkU7pHm5jFk8uH
oBIiBQ6ZbnvhmHssDrqF8n3CINEMCR3OnrWL6OT6G+zB3iEeR0P7KoYYr38m8L5K/DCb0qzFZGH5
K57qi4HdQIyVOMyalubyyeXNN4xFYX9nWp+i5K1XyjOEESQuc0udO6kUT5cINTs9s71OKLhPgTkZ
kD8R0lsTuyJX5pNmtVoB7ePQ5C5G4jyza3LnARMNELuMuzVjJXgh4InGRzRi2h6OiPYJn8zd0R+W
Ax2DnIlBbXzNeag/1tl8wYt3UX5qoEpg2Luo7PxihwG5VE5FTVfKrjzbVcseEtq43k69gI31gfSR
ZMbiq/tLqA3T1NzwHK0LJY8SsGA+srNMcFr1RTMUX28MjKBCDDu/2S5Jrq4JpRvcRrjeF96VWpxv
0x2+vhpv2GCp6cCpADQ1PrzPwbdVU5zmUBuvKelES7zbYFW+woV2KOkyn2e5XCxioxlqoiH8/TYz
8qVgqY2ezZg9Jgd1Q2G7rlQu8ABCJlbeEUimtlQ36p/ATHmSx4Z3jk/mf8Z7Z4/D5rGuuMS0X9LN
N+0jHqFyKyYDE09cVYtN8FRHXHyJOENHInx2ETHxXITkhwcUhEd1xot5FYPwBXsBqown5VWgCrzm
8ggpk9CgeBIquOvkcFd0Q2vTVjnWYS5qdjo2v5YxTsBBZc79nTFkNO6M6YWTYvamBT5cdkg++sVg
G2aAWwypig87HqWZvdRDbA4vHyK5VwuGBlenLlOz/slfE9gKEI3ZMiBz99zeSFoDtn8W/cYdNG25
sT54vbkwDQxTRGiwA9Ezrj+LEiAegC5TnaTVS5vRWmEBBHp42IT2aGla1po4wgL0ZzeyadCPP3A2
S8pYgNwsUZDznauwoZhOCPU+fNgTuMBV2c0S29JiQt2gxU+o+tv9WVUkSRSulMM6WwwOIjWH7uMk
guBomsmzF7MZ6Ng05Km99I41SF4LXK+HsIW1eioRdo/y++2vRULH4OkG1/mFxj8ssFcM9TTyguL9
bwM5OA1xOL5wVQSlGTq9zpkAyy7dxLRxXUsYnosoKCe/NVSdW70eLBv9EGEXkvUvbEYxVYFgVNmi
/58MGmL7aGLR7iAt64vLwnwqijZu86XDDEhfU6YFrYaJld0Uil0SigOore78lKzqQe9tVHY2umQf
U5pJgUba7zwuJ8mdiTtuuGkRmPPQ1R3IUPD0/bHw3Mu0k6EYdHG0EaC3dwzediwMPOJwHXG+Mg49
4Uis8uSpTKSC2lDOJ8rkobND4wZZwfw2oh7x7Nn3M5i+5fjwGvIV9t6P3LzrYaCjcTw+0hQ1TtZC
bCTw01oUSHWwkUGBAT9Jjx677lfjBOeB2jHuqdVBn0Zgzb+At2XvdUYHTRTq/3RmSo7wXJfK2alc
9psbfAiM4IhKN0ftu6PMBUsPym+5KehDxsKz801Aa+q29Fhcll7yOekJKqbJNeyEwhULZfuAMDHm
+MgZka+LiE8HntbqpPadssBjV9VKz7XCMasZamcDkWU1gOUeDZ1OwLYxlki6VT9gtP4w8SsBOeop
xyYXzKhx0q8FlCAo7qQfTG7jUzBuCRrV8vRRZWzFEItzU4NuGZFYrqPb6qo0slm6uAhLEZ+FXfBP
Mm6IrAAQx5b266eAgoKGZeK9hctkRv3ucmNrNlCanTZYw+IA9vgDc9ZCq0FxwDz03MV2kks9OcZt
BqVSHp0Ri67huUbdgr+qPDe5R+oZmQMw7zfeFRNf5++qtO6J4vz+nxSO7s1hPCHSCtwdzF0YQ1Pj
uSRE93SGbOH4AkX93BWYJuatEd4lbWCVCAaKpvMGceLA1vBb7l8WgHLZUTeBusf5wo5gEFSwcGQ/
eVH7qJAruemQzptVauitjzZZwIYMuaxholjNwee6brCpqb/0R1bqguSBKMa8oYovI7UUYVMxxJBM
uI2VVlTSxg9IIComsugqY6KBnSs7ZeFOp86UJnEiixIUHzZdYUmE9MUOFJlcmCn1AOIRnvcedKaW
JDobkaG2Ja1psNlOtfUaigqEcAdHL7NHe27rgra934Z2ktlyjbRvmuf453ooC1NO0oEekQ3Pqhd9
GZ+X+d50Tu8txGX1DwOvRxT1rhcxbDpNwg7XVE+4z1+vEl/XadHjH/H9Fye3dLnKc/VdizrxCkk1
GFilJfAWNdiwbFe8lyRgPZKNRyrrP0HcW2yYRE7x6CyHGHQta5nfZqSarbdDSwhKWyuTZfrxlEhd
2gOfcPJgU8+sL5fMgci1JGYX5vT3T7yH+LrxgkFn6x2KCmScZENv6Xfn3G1nxDS4b6IAlEWeFhkQ
m7MJnBXR6usKNuU8napX/Pyhp4f82yWVDcszigftzMvaDOXwNzA59NCpGCmUl+K7NC+XHemFOOkW
5CzhLrl6bQxMKkUKvnV/VtRB+5PcM506QbYBImwFde25BMJ0gcO2bFq9IP5qZ4zxJH0GYKdsmYLf
6/cp0upn2tFnBoPsDjue94FM6zifOWCoM+08CQLzcP8/q9NFIaAwcAPuDUiIOt1Rz4qA3HY6LbPa
S/thsyXInAv8zskZ/hIrI8w+HlTMuU2IwBdLVnIchflTNkhUVeo7z710fM3vaKhwnyZDGGJ/w1to
oNW/bXwHZozZVVZaadzJsV9N0ZCs6+AkmahAMcTlQH8xT6rtX3QorCeFsMATL6hf0vtOYI5RQfOI
1QfEqckIR6hHR6FQMqYgtaYmlV+n3+SeHnJfbM6KKTTRJzB52Gk7OgXCmEF5vv2Z4dkjmghjFJ4V
9qdhuaY7JMFrmdireh7ClYD1WnWy7NeyeeULx+OM2I+Vrl4AP6AuEx8RwfhwnrzwzuDDfUNwn3Jo
S4JP/HuUcUxUzJC25MSMdFIEqWiLtRfz1Q5qdleuUd/MfbYQH+iAZdazw3aDN8MQsbwIi1gCKGHd
tGJQ/FIAyXC96gnWEURdXoyr+TIMQsjYLy9QenIuVsKXdFRjAwjSu54Fxu1jPQUtFw9bOQsvyTVj
/Nl7a7AP1U7vHJtLiel84pRdIMBx7QoBqwXgpjjJnrVbQbPn30llnDdfcs+HkNBORkg3j4WVOw8N
BKQma5n9StnePZFDPvMG40F0veJv6jPWAnngsc7WOdCq5z6LXmBnFBVq6megcOUix/5EArBWGBvU
bYB9C8Ew1sk3C8DIBMKLwNpc9Ok0BM54Greh5BGtLws5HEiVsNakRRqdTu//MODBNnL8ICSxVtDu
zmZR6mF/kE2XCH40RMEOPvHFvA4JXZjCgsgbjK5GjyMQzMH/omdZkCSXA2UmmtoSwNN4O5gEVqri
6nk2PPuaSXN5oVJUVkoGBah8hbPj7P/mNZCBptTUvn8vLElZ4QcCQkF7SBgWZBQmpyTILmyXZM/f
h7n+OBcWCTnf4FECWAyNXhMxCqs/AV4VOPBcT5YJfdgLFPVyIGDhj6nN2gmnjlVshYhs0PdVEBdt
OmU3FShqkeBFAElBvQoESiiLSFa+cIXvmVCOzC4MSP/2DlCU9QSyZSJdo8sZCSjYOxkO6UkzSjB7
QjBADynxBXmWcimqnlD9MWoSjs4g7CwTlrSkIccDIIysknHDd3doVPVb6mwXHczLx4IQxMyGE4uh
wRBRd2L5jBW8DdFIoKHF1P4a1hU5DkpQvLO/2SF0RFBKIfhSjBJC45zNe1BS5Kx+xpsl6yEjr+PQ
EIOwDiNspO25nbNH7Tb73XJU2ReqJOiPTAb1ygdL1sEAiGXamM0oH34H2S1WX9CZmLYnO6ElxcvO
isAzVrxRqRDl86xo0LGAvDK9H8f+GdViZYY5emrqgx2LHZwn2OwLT3+n+IstKXs0f31dOKlRlHdh
+jfTI7Puc27QGuSrYoB3K0/cbqw33gWY7coQrrqpdiEod+7RLXtCTYLhnCFi3GH+PZnZzkP3ltwu
YOec2t3SuGzbyxnoW2YQoJGWx2yBgnwxhaRT6G7xcw0kAfaCDmeuQe64Up5OU0kg3Pca/qlUuHv9
7ffgMV1d1RTM8lS3wQwSBCt9P4Y2yHPUI22yv/QFGEhSv45ms8fvL7N0Aw7q1HQZC/UTCo1KymNa
pmniVa8K7PmCh0dQoMeCLLfVuAfblfj1Mu8rraPAIZ/YwKbE9fGNOtFhVTeCmD+/Wf9RkOeOUquJ
2hYJ23/jApbDenwHXfOBrgUD/7aBdOuQx1Cm9YRwJiftSDJllrqYf/AI5gsAI7twVhvs7LX0ecOZ
It8rUMycH34h2zhVP5HNZgaSBub5YFT4+ALwbPNx2FdZElKRlRZyGnzonI/QG6cSGuQ+wR0j6X/k
zdmNVKtYGEnmbOdHy3P2XoByv45ReXKfpsbK3t/mOS9nVM/8u9CNCNpvkI0fkFYr4PALwtQ+UcB3
z6SlE1xkAM63foZUGr/WOAumw2OP04HuWtpBT/6zNVcAZNAWrJI7t3uM4dhmPvRw1itIch2basG2
dDaBEEa1Nv94yiKIRBJvKOUTZSUyS1t5LSVjtnIJwpMLoWZCnmGEW4RuKeq7KkRybriwnDPWCPsB
tGULJdavGS+KKRx0UfQ2MIzsMre+Rl+NOrUlx33BI8R1z7uBVLOUGCfNKyafIbSUOzDdrFqQ9Kub
+9T0cu60NZ65ZwcMipxxP8/YhtzdpBKyegr9MZMmdA2v3WrsfzaP7J9Vy90L7wKEK4ESvR/EYeAm
vKY5lKmMxMt7OhIOL6kij9QmPLTP7pksGXDJJRIuLql8cHxsDkLoZTOQMsdD2dmRkUj+ZVOPU8El
toLY6UIuAGa+Zim8hF8dHC+g/bah9PBfVlQ+uX5uZiSH+XNDn1UpAAeJ3ZQKDG3ep64NS/14VZiL
7Vx+Mrzhj94NjE1gFalIhwGPs204clUSsQZO27CtPYytg/HyI5OTT6NK4wb1eDAYYPEwLPFCKDdc
pwXWo/DDyk/bPqNCy5Rt7D/wj7AuZPdqEffwudeaG+ENeT55cSuBSAaDsDrEDe++eey/sUueJdmk
PHmtclqvLWsvT8hw2MmAPpJtXw3efp7dL5I03CV1jZ2VuIE1tWbl/t02PyqQ8RftiCN2VA5nOxWA
41oVIDJnOTv+sLKnlyjGrwziIbVPXvchG1187SvL8+UPsApVlka/kJppXoAvcp6D/C8MmpyYlmlt
0YK6/ukoqyd61J5h2RupPMgAltl71Hf2XoTPVczGHALazQ012TZ+2nfcurHL2szKc562ZsNcq7Gw
KZRw6thzWrBSJfZ3Fh2y7i/6i8GwrB46Z4trWJ3UKwx+O32NjX2gDV8T5o7l2EA8d6S7+obewB8q
feGydeaXvJ56zvM+yEBYfg0mC1DFUeOtP56FH0RzT10n+ktyXr9pBcjN3DVsO6BFva83Y+KoYlXX
cNqIO0f5xh3SIM/VznEBJKysVH7kgtWwcpI/ibWKXn+H5DtpKIMt9DHMpwnt1QG6kfmo4c5YsAsb
gHcYYtpkcf5opIy3bGbwlPHKKXb/JuIQP7tGURpQ4iriTeYos5kkXO0E7qFoGU9vTzHtqMb3CoOp
q7PWDvfTYD76qKQkOZ9wZQTy3hI1NxsnNJ5DvC5GKVcd4UoCW55RSM2+0FnA/Me2XgOsM9BhOy1G
YNXwnA+dGJrD1kvFqJh8GZFbTWsQS5pj4lk/00igFbgB53m79nIaT+qU9AqobXWEJYV4jc2NDJRK
/pArmLAmS9P6aeH/S/xWt+QnODVbWOqEbWVovEsT95mK1D7MC1CFO7cBi6nZyo0ypU0veFuOCL9r
1R/kOrksX9Y3hH1ExW2/jo9sGo+j7j2JOTkOk4eEI4h9a2eBTEZXgv+1Hw523tgEH5m56HFq3Eul
vBGApxjC3QPO5na5hDN2JkoWPZ+1ZHDba5cWihJsImJo0OY/5LrJACzq5lqvFkgaVnMI6KmSTdu0
aZnta/Rjnwt1kDapQyJO/Zy/QFttw2wgCd9obXUaz9xljfxlrlqiyPUUf2oLXCt5inf5vwynUPD3
WlxRPqJvMDlFZjFLOGlOOgQG2fVaUvfqB5RmryNTibEscSD/MLDgMkGzdW9uZLvQ8Hyd9yuNwABL
4G25CKybJIjNbTNTorDcYqlyA0kfu+4RCN+Tkf7W2jwD9AKZEG2viIWwl09lvQKfiONf2bkm+oeM
Ct2f34q2H/u93SltF3yPEbbCIOE1OV0gRaiSpxxD4zw8j+P9SiTvHVOF6NpLGYzSY7fYNWlHBpD4
VdN2fUFi6tfiY+uz5ig3kt3Ly1ahTWseBtgspHw28cnpcoq30q/1fFBGp+4hpi0jCfH0zbYuaOfe
VsTcp58rgY08uF3fHBHgHC8VEFBv+0KtXVUOHId7Y6RmKSo9oTGU9uFB+Utso2Qr5U7SPh/SLwhq
5oqtB/j+uYuYAAN76C4e+Edq1YY4KEhWVJddIuHUoF7/JLqHLiiQ0knsXxPYGJUvhDCIlCCCm6fA
ylcDVta42tTzSXP42mdDWAqtsJyCKlPozc5IRjHm63OlJRsLWerpnScoW5Tipra7YYlB2n9IzOAp
s3rx2WSDjbFIkgEORG45sIYtzI2baGF/29xOPp5VTjltoXuCpUbjiIroLSLN5F3SRedfl/nsRZ1H
UvWeRZs5LyhTPv2HCPNN6k/CGtlHKgvvCoJtu6WWMei32BeC0BDnuKtT1N4v8PtkSve+QcvEEMN8
J/JMGM25/1MQSlj3saddeIKNDf9qYMke2qaDuxaWjn1QeI4XJYKQsX8NNJpMlwvVOnkTT5329XTM
6o7sEEPuJm8vd9VqgNFxsdDtA5EViuTUR0rlIIWJsMshkKzfFQ8GYjVJUhq1Ubzhy0jAMJtINz71
DkpMPUdgDT79gyJTMk9Dfsjh0s9n+kLrVu7JUetrWQgA4uJ2RN42FR9jhLUUeqKE4gsF0C+JJSLg
qEKsJP1kxPhuoGZO/i1kAnWt7d1pdSJV4ZSetyDGS6Dq2H0RNSowgMSyK65wA+Y9P4TaLfrF2omx
ZM9MC3QLQX3/jGUjlLGvxSf4hAVWQaJ6AAqipkSKaRIQG56IXuhfth5NrstDkfr95i6cB151UHvc
BBwHy87QlmpPAm0Ge8AtG4M7hDA2bG83JBg++iz03fWa5cYBomlxhRkjSJkwSODhA2s8PTLl6oY0
kyatvunzBCG+M9j+uaZcYeM03y91Qv2zJWc3aHxy8J0vvMhH1MjIrWAQ1bKlI6zoXNDzGT29nZhi
GSJSx4bZbo6I8/QJJ9oDv1D2OSnHV/xacYCxFLziUKWH4U1Aij6g4uWt0UpCGoePVmVqEyN7AANm
NeiaBdvBwJ+AeMQVi01hzInNjDWLtAhjF3dpjMODSj9pCFikTJrLBJfP15nvzWHq42oxfkLnQOYl
ppzFZpPb5aLj+FaeBiwkMdOD449t3uL5Ao2fRtygWiBIgH+SuEcjXW9Vq+MjJ1+/0N+9llNGIOKB
EQTFetwN2q55gATlYAuRdzAoLuGHG5A/Byxu5+F2JelGZDwm3Qry1qQrqwXGnQAnDZHEgg0zxdMu
DX3xbLd5xNxogGLISOXTO3eKi7zR+721tNcjVjdXd1s8yCOv8khkSIJuB08l9Ouxp7ECHmus0l4G
piV3bCxIUvhJgEh4ZRlb25h/zjstM1xUInsMYP5mTM0DGtp2kSwfKKhU/6moH+WD4x7HOcz0tEmL
vuyNNFe5Qah0J/YI60yEfl++uPO/DMEe2Z7wJeydSHgTPrgJJZv8Ju+G5cA5Yj1oG0fNJdOJv5Cv
2APRIo+IomvP7T2wkK3z1zItBzgfKk3Tmy5coe471M5Jp6aBUlRnDzuo+e2bEPG2zDkCAuG1jRko
IogF7sfkSfxwloh1Xcc/0gAUYgv1EpZkHsH9h5wv5c37AegbVAKLnxVppxwh/OlhtUMoOA1T3kCA
eFcS5MaerM7fFKloyXIv2WF58aoB5Vmbp29XSlikbdvaSqDbTS5nzyLzr5BAW1efzqCuSf+Ac0q0
BsvRDIp7CZ2ZppT0ROBJqLR198B9br9NlrQkf2fWK6g9R/nG4Q6/ONA8MxX01OAmqA/FgDm+DTKF
5fxy4RxKDUyEYNEicCtq9Qzr920WAhqqfjxJcGy7T29PRFF+ArAe2Z/7iQSiMwTS6jE/5CEBzg0c
kNZhRlGAGMlozZk3nyC9/ktaMft2VSTWM/i2yvFoEPnOi14HJWNtHBTybHcDGTO9SgPL33ZPsyYN
CtR43GnSOPxA6zrLM+jCSrt1lEBkWJ8KQZEW98JleLEam2VqYZTsZ6X/njvUpB0Vothj0dlH3x5E
pnyGnYhj9FlWH2DmvhNKiI4zNpqKmDOHxP2emobBr4+wTOStW7WCcox6yOW2I4wV1Tvhvwt4SR/b
oyyPNQpoxP7ekXM3QSnQkx6PIyeQ7uFrjiavwI7p9U5MBWi5gcIMggBZStyiBTqMjNWObM8ntHSD
gIy59KrHlaLvjaaAughc8o8pPiJL3xSeHt1JT8Bnrp9m0eSk1qrolW4rt/9QoZtjNuAaYwQrWayD
SlR0ji4JFz81s2k/NEtsOU0jD7QYO8GopffA7LzHoR9N/XSViKb7p2etP/p8Cc9WveS4DHAPjFdC
SFEHHNT/NPO2CKba5NSZpkIeHJ76PjEEhEkzRHekRj89oDpQ6+w+Y+/Ex4gEW2sHuxSKfE2WTZ4M
4VDrHXMjpezslopPzXgkDUOR5EgNbxP0aFj9aG4HqLOIyQl1YtKUg/oz4xl+MrSbFtqD/KUs1w8i
mzbHdUwN23/Trys1Xin5/sFKtdKxNSw1nRjlRLXN4APsPgdTCv2rhEQFXs0jQZcHgC4TxdhWbsdS
xyGn7cuuz2Crs4hBwlInmkMC77/OEwBTT+cAwuiPNfHnRQf9Krlt4R39vPKrBkdlzeTC6qlaKjkw
t7wCxSjEhH6MhbPAYQfmb/aWf0bHIBxRcZEBiU0JeOJsVgxpe/dRZdC8dSC3sTncbRY3A0hsvaDF
y+MlY2ikzGCV6TPw7KD8UIylv8dAstm5F4EcdmoZpOvf2qC/z/QxhFNlo70S/Hofkp/BmtBl87iV
rOYvbqm8hIJCAmk8vLu5PypIJRuNLFv7LU/qh38ZE1kloZGrHKxQOu98wK1t/lxHfFClsjwVam2x
jWwzG32mkZU/XXw7PU68AKoHgc36EQEe3GR/Q8Tr7JDoq2z06dNUhakw5Vx/yOV71zBRDhEikQDz
NTNjPLSw8N8nxvGXGi/pnWjz1A6PVDCt978B1/1lDNs8o1xKujKgCI1JYm63Kfe5V28C2oSZkSdI
klFCcFogtvKPfBcioEBAFrvKCXQxtbLjI4Yjz6JS7q+RqJiAR28Fvy7JjoIIchlw5bJMlPN34t07
Q+3xHgI9JAAGUrs64+zRLB1IyrkXW5rjaeF/EnZZtCYcg0MoCRFnsTH5IWMw79sxwiQ/0XugfhM7
IlY1/Cy3okLi51w5E0v/ZZ0s4EigMK1SpcQR2SUQwNqw4GBskKpihI22QeGYpauNP09vJYfvkRgZ
BQ6oa9YlXZgQkoU2xE1SJTiRlH3P7er/pVzdBtwvQ6zgfIVeqOMPGniB615dfDERAQTPrtjdtv2/
8mcGTHjIqITdb1SGWsmN7dycAAiuC+O8R1wbYp8moJ/J+NCmyobCWP4LeH1lxMWzyZY6HMqx0/BA
o1DfPRlukblMk8ZxwLWYmvLKodMrYxk62MQftneeqoWRqv2o8JnT/NZl2hrQ8p+okcHFK8hXzGR7
dwHVgTn4YT+Nhx7BZN+9arQVJLcyA1KEmAXatQcOPELl/w3mkAtsXZxH0ggm2ugX3boOCNn0roUx
9uQzDPcsCUryK7u4gcpk7cWShwP/gkPNuPax72cPRGLpmkWRtUupfFJ+KPnY59uHQ3GfoR/MlZPq
KwLc1dcqruDqEcJzkCCbpbV417zhERMikNdQEKQ4KJANcdhj9QSNc/N12xAMzVl5bS4QVjYBLVcW
CuA9w7sgId5nNNiGIyuA0koTrsRNipxSgbstRTyeez13cWKWL/W1v/WzZbPQ3PSAqtCLGOGMgSFc
C3SlPljJCDApaMj+UbF5OMBpIaBbVFO6yG1KrlzbVo+Ha6Ipw5IlQPvWpbTvPHt9PheMdROOV0w9
y6J1SeZaFP0GlZhBNxRGw3tC+Pst75bUK/wh17/HmErZyjvWHetEdbJiK2PB1VJdVtbbVszaHLNF
V8yvhpTez3A41B2zf6hgmZye/YnOEx3ZYuoQD3hznTlavwWFkxnVrGRK8u3cvdiykuRMe2myz+jA
+7yKqze2qrh3YixIowi0umr78hHlXAxTwpHilmI2sS8iFsXcao/Tv/CYGfSNXkMqn9Zw9YSvQiFm
thu8E8CV3GCxzkT23H5EYthCeW6eGSPW4ebQztwE4b1BlhyiTJ/9jkmDK/hTqA2bvjOgL6chI/1j
NrdikZz8NMUJKbx/ixIeWxy7tpCTKxMhL6sXv4Ta6o1iCeACCX2Dn21iwtZq5MXu150WhSx+AbUF
iZe1CAx/w3nidYGAVztCBQ/rWYriMNY8ydx25OtBhSOoohFQ4iuPXszyI4x6vpjKY9TZIQGQ5nse
2xV7YrKSALmzh5JC+Mlzbcd0Njep95dwgDt+N2mh8MGxRmu7No9T/2eiMTxz6j/FVOgJAW7R8ZN5
zulSHXzfLIQ1uWZyEvDmlDVVQhyh16In6Ut5vBAGc8US1JECppmXj2Wr4VbS8Wl5OfrgS94l3ABS
71Qecoj8ieR0LNPuLS/cn/fFSbj8tfNmPOw+F6r8/Bzq08nSvpuntE832Qi2ze69Pp0n8279aoUw
+evkTBpeZDm837VamTmqs5zzdHxGsgAcmK8j8o9VPZuiMBBEVPYzJEmXphYLWHZacx5bIqF4Hp53
kY4dhvn8AvOt2nCQGcDOFE84TmQe4nv1G77lUdhsWS9t+9FuKKcFIjDVGoNSzzLWYjPfrIuczrxm
5nCFn/EgQa5c1lKIpQT45IDk4HWtAwXhlcbI+AWqMAz/84+E7LbWJ9xRVFvsgvIdU7VROj2OD8DB
G2p85l2eqi65b4gPFnXuFkhjXktfmxi0HSzBgUVs6XwrCc1TsMP+sxl6w1+wNfKuwDnib4g2vmAk
mwARlFIYBCgNF9ayba1wB3IofroGM9gs4E8e8bdEe4BwHVItBGtde2pea4TCQRTzAz8mUiLHoBgY
Uzi+1pV6WR2SwowA3NTgqw3O/0UY4USnCuWMRCXObsPJCXodjIZoNVCvZGDhuBA7yZQreITGbTr0
QXi4yzvRrg/nvTJzyMH8MOk+TtOJzZ8J5MykdjCGOa2nbMPgBAmg0T48aTbAL55uWbPZbLkP4Llw
IiFWitTpYQ/EDIaXavy8/8m43VA1qkkPlBpsErBQ/8raXyeG7kpDKD1++p+sF1dLaGtmnv7pN6I1
vo+JAiUKoKwyMnSPgDv3y/JEAoc4E1vg0M4REWLzyiM0hFWYre1Zn2oZR5uIXiDEZlFcudxwPLuQ
rQr6Ih3g1+dn7nzZkyl5qr9mKQlA9agkf5wQo4oYdV0AWuXZHbKv3LGW1jXM9RKgGY+yXTDcKwZm
R66xkhYPlTNKgCzElde7+2QxvRKqJ+StXUpOkDX7EPtzwx8apYwcsb3tVre/STjFIfUaGsPpMtG2
uTnlBjLlLchD04aZTPU242v0Dqp6kSqa1jun2GiEt07g+jxh96qp3dneBy5gCLQ/DwfouCiLqkoN
QzNb0PsQDm1oGwfMm90nY3X1am7kggg0t5nv42iMfB8MfEHtRHXeZOBMS2WJJKpRRfvuUNFHCHUQ
lYwWE8lyGYRCVv40C9/j8pyumaam/0iTfs5evjKL5xXsk2tVBT5uGHl1S2jzDPbRnzxVxB+spAPG
vIsA5hv1iQB+ztbJ+HOd11pTd2Ci/ViEtc96gvh1OCZEKcfcu92J0EbSg/4Jqgg3qxsAH4Cq7Jtl
KwALV17jj+C7AcMnWtOTzw195b9pQIloXL5pLfvS8zONX5xo+Uv//wvpU1kc6HMLH0WNcJGd9q/G
ig9plP/YVxXf62e4FVi9+ANX8h7uYQREZL0noR4eEvciGlfFYHlO5dirQD5VGX/EJPnoxulvJs92
YZHbmaCPkCfD7A2CcKEQcJ9mJ9Pti8VmG8f1K9FZF2BCL6cXjSzm5zenwS+Vbz27zeF6ff64XgeG
f70ej62XnVZF00fOJjrk2qnXJp4RN6uj8B+RiHB8uLcB02d0CKgIbo+K/ge06/Z2qqJD09r/BgAe
ou+XWHZCLtsDyUQxEVXV1rMeiJN6Fxwelp9UpY+Sczd39/i7M/hPgkNZEu4v2jU5G5ufxwh+iUhe
gWUQj8hwzgU4gaMHwBA89fOpGqCYPU1avbpfpJ8mP8nfTrNanxpHX1u/rakpP0/fVbF8cLFTJbIN
eU9mSxVpafytJLO+VFGh5fivD7DEWVuwcHbuQIdlDFbhzFf8cRnR846Lz9Mju4gD+Qo8VO5izjWU
zYg0J1ZZI9rPSCWIT5zyCGHdguG/Vi7fU/ApWIYOonPsmP10N1MBWzyI6GaKUCG0hwtHr+2vSllr
SWTo7d4zjHfi5FlPcQSYhrgs/1hrsXzHLjHo97VbedPwflzaV35dW2kvC5KktkbnMdeO3cyeA5wq
R4IkS1snGDOJrqCwXPxJpLlND9e/Xcnj2v+qhMU6wuSSRn09fMzAKUuo3aX2eqOlRqvj2y9KKHia
ZoZND4ZW+wjIS+v98qNLVqYUaIvD4xcA6raxhQVk14+bP42X+JQ4iPYAuWyW44kzZCU0nMHXJi0k
4fixysweZ2AyzICXiGprnyBLCPxpPGhDmLGY9c59Piiw0+ehddAle25WAguG5q9bZPU1nuibKwMj
zMRftWzHD6Xkc4ARAosIpx7IlvLJNiHIbo0KDy5yMdKTBLJ58reYl270GSxQKHJCBDrrQl5VMLK3
6uccWXgSrqI+QakdgUdA4igMX0fvQb5neXJdE0clVn2KjVsrTEYwcPpOwX7lW8d4/tGiAzuBseTQ
JX0ySLiCK1m8lWPPJ31e1JK2gPp8H8pEKNuO2Tyqn16YPepII5VKUFIasi++rneG+yFB0LnsU6LJ
gY8abuhzxUqQM0j/BV56D0KQo6zG6V6wIbRZ8+jrqtTCae3Wznkqb6uekhZkExLSDjPPdqqE49vE
oCD+5OR4wpq+yDZzza2+LoPb8hzg+NtpkxzQjD/sBhzzjG7Kq6H7ecrmCIQeyfJkH1uBRhIGx2FM
TetcneEb2d9710icj0YNtQJZdh9dfGgDUFP8ZkrXsWhFj1rN6kDvR2bWOjqlCzG4zdpS7/YxxBTp
FeEXKIl1BQ1przR1phegB+5VGm1cTbaWgcqekKbFrEadByBccJ4IHr2PcTqVlmwdg46d5JONzkJd
un82tmhGu6SvzYqEdJw0j8U/XGP24OxNqDuWrZXVwmnVKw52KXhZAjjqZ2qUBZnD5FuXyFWqlVmX
yeUYI2G5B076Fk15c6P0UI+SyQT1VSwSmsqf0w6cTFKslpJBk2f/dJ5HH4nJzyJZfgNCh7WNhynO
D4RNpRV/Npy+yjJ/ADdnVV4wyV24phYyTPaewD3pj4fCAmz7TTwwonwt/OjuObjqybV1Lh9QKOMW
BSyLUd3VuB9hj0GlLwM5mVGG7SytCIDqDOj4dZfEdt6wOAPgRVJ7SdUCU4XcFdtTMFPCMPHg8Icd
GFk+T6NqU8VLx74yoMs2VzPBJQ95MUkk7Erfd70VAiWY6HD/3Qr/rEA9TXJ7OnbGM+K0GW5EIOqV
neX2xpOoAp143Ziobd/aU/06/mOVRDIiXngecCrPRlVm5yPEO0z/Bv06IGTpQUyct8V+ShScQBBU
9mfwhR43f3wIwXHfQYVt58Lvr2aT7m1XtEZiw3ZUuqHQNZjjHnjK9UTOYp1lj+1SkRc4ofoK2n07
4+MzJEfQLI9DoBdqT2f6jCK34LWMd1x9kW7eCwTxA3fAFdRV78z2jAuiZPMsWnpdu007bs7MiQj5
oNCXOZHzclIg7EvJLitWzretD4zhe2WiODgAl9xpDHkVyIeX7Pv+x8OZ2CVLfIeFyTkbvyqicBuI
98oIPf2vYIfyK2maRzQKCaPPlx5hbavZvou2yGQfHesRc7tPtiOiPq44DCgmOOCqtojCyd+ysrXw
1SuiDke8Nu41u6aqET71ccxLTlvSjO4t2jWn2v/oTmBrzcUuKGQ8tQTEPyId0cDWJY9BA2d+5SaV
EhaonDiP7SC+1i0aGta58QYjJFF/Em1loWehawLuCztpAqg/tf6IASEyPEWGMesRVfvIrT8HTpmg
mcb1usQMOqFD+9hLBFv7Bh06FnvUTQ6iAQp9tLLyEwL5bWrF/kWGFmZtsEKwD8DXw2JHNEcfzhDm
xySfbhZf6B/3MGuSWWITDdGjVQJqsi5j4wcDnMqI4JyosE/YH9vImDQUZtS9TUBgLaYi1+v2pvG5
UiatMas8vy46HNWhlLq45lsWBETdDJFCSHDVCcJSwMrxWQk1XJ8uhu79Vo3xAq2cb5gxZUyLabnc
1lJFCjtIoMz1mpKtWYRtgWxDXAhsSEQvjCgnfSJeg4K08kmY0l0KtvMuZFz0LIbSGMxS81lvmw5q
d14A9LdXiuQrRHWd5wCBqOJS5aw45OoGOxxmBAQDKdp/wItJXuLBvdz0c27xl0i6IaU9INatr8YK
Sf07sErMwK7RKVX+dX0yJDj8FU/N/RA/Y/fJ5vhib6kYxtKqKywjQn8CcVWK0hyX1fzujFW7re4k
GvYqIF7i/ukwm7KkWHzbsYQg9T504tDfiR+xDRnoveLeu40WZfEe8r+PklnY4ERBuL3/1k3jaPLl
kkwNq3wWHxNJW0s6TR2sxtLeEx6VykUpZzyYsmLRkywQCTTMYZ7ymzetxEG6hEhrTyFRsZI0FEYJ
uQ1OjawbtEldW/q6FRkMGPaZBPJGiRdIq+otneW46S3aynnD1a+FOa6JcJ+0ldTHv3r8q1uF5h2C
n1LcLA+mKZiO0tjNzw09ZNv5R9cuUfEn4ooFx7buO715O8T8OxIaBGiJm0Z8aRqP0JBtOf8EiCAt
aQwhoK/QuWAHrW4Jkms0BVmoXvnx1pN/4CZrL6Ks178ALTvm+qtN8iJdya/V4zPcr+3MtHqstHrz
UZJCywYele3pSW2CMbDvEyrKWeSbbSeZbJ1eusan0z7S3/xBHOoolnBoYKb1hZzHUkABKFXYxapd
7A5rGf3Zr4ZlnODZPKQ77owkOCdQyMootuZVXTSSaBkHw4Bvul/q86Abm66H2c+qpqWtr0aupluS
IjJCE4/IF4wo0DVqVhUD4zJM2BEk9oUTRlOKgVc7lgzeMAsUy2A54bbovTk2jiollibgwRZ+G0IG
YitPWfmwnyaw291rCo34w3FL03TbsVXFk1KUI3HLKB9k07bopg+uaO9AjfoDQgHbXC3q0Hoij9YJ
civtPbtbMKxRzsi6ha94P7honZM6tHZNKqeciVokNkKnVvkTXdE5T8Uw9dl5fUJeymP6Xqj0jTht
X8B0LE+6RnmjdW1QkxVRQKj0b4Wj1C3YpzasF/dBSQ90HZp0FtfHZTYGwSzw/dIOVLuNEzHT59rf
XkyQlTACRpt72LuMUOECl0vzWd5w8Xw4SsyCVglKsWithqdJ1MsQ1zDHLmzfrWamwgWs5LJTPoMf
TXsuwgdT1a75E8N0JpWSkqzOyq0weZxcATAv3Piq/dbVvX4n6avqY1Oe2sKcJvzFgurGgUe1TCF7
Ax0HlEpvy4+epht/K33o7e+ZyQpOm7H1QMfoDFbaHgb7yIuJOyaJtDzFqHIHZdXbvZuDHhmxMSUg
fWkxyqz1D/NiATgeZTR24U9izHBd8trEbJ5XvhmoYqQUrGS7760gSTgmn0Egf5ydjUM7F9PoEXx8
Drl05yfdyZaf2e4dbW+onMIc1oceHYmYCS0Nn/vRwKDtXclhGNqH2Y8Ar7GyF2JVZM9Jg4aHtSSz
HxRr4kIGDMjBOd8klrd1m6qMUt0J5neaGfD/4cIUU0+chLV6YlNEmmeWby7U641+yIk675/N9KZu
0TqjQ/K0uW2g7i0KLpf0u6jU3L09/YNw4GJYfITMw42/syZ4KmrwyrbnqlkiwDGEd6w35du4YvI6
teMWAA3MMbOG4eZdJ721sZjo4u7SOBbJCX/OqpEPrk+4+JnZto0K2iLrB5QTc2dr+YAGv9oKi7SJ
zldLiQ4w6srBDfbhbL8gZHv7RMFhV5yTyZtG6tU8KkK+Ixp9xfCfSA42YAHR6UIHBK0pNp/U+yza
r/2mWSO3Njpv8EnG4XZEbVEVgsBq24pZTBrcPa0kJLGJR7l1ZXNsl1rtkoVmvqCxO/ttoHagkoBN
R6zP3CtqD/D9E03oAgE64GMTeTvxSAbDn8vgZR0P1dhZcS0aMd3elb6sLR/WmsnpjCZ1wsW2G/ZS
vGj//biZAK8w9yg5fX0tBwYxaRHpQ8/4bKo7tF1PXRdB1zpv9614G+hP2phCYSgTpMZ+i87lLm+G
O44XeoyeIM4XnbidcdF+Sbe55SG0iQft/ddcWFgZ4DD3mwur7VK8LE5ZH7l2DKeWLc2W8HDgCorD
TUJ0/6ykC9dkp+ki/CaF5tmEajA+m8OBofMT5fVZQ2rKp1AiM/GfI2+hSFB2OagWyJyYuCQRDV/X
u8F8/YsjuLjSZWKh8Kgurrfaa4foLMzno1Kti4Zoon1QwwKUTFLZudU3GOnZ4q31UDh1jjwLYXwb
TmFRqdw9GPq7cNo2rAqdb5wM3KnfmqbiyFMeUJBhTUuR9Azdh1RuGyc1wOVEAeBl8uITCQ04FR7K
lqJWmI9ad5KTwC2WNUNms7hy+Z4d7zuhs5ENxgVJuQm0xTxDkUehk1PekWaH89LqAr5s5LT5xf4G
FMwL53XO1kW6CA36GDyMa98S6OCbSZPQBoQ7VSKgrVd6gAXvSrmh9VtrPRc/nB+U5hR6gYtRIx0s
zJ10jyw/LhwbHVClLocWUdmL/ac1CmXnrpAehKJoZQXiGCHxMo8rwsZ2YiUU/CiiCHOmdTHmTVCD
PujjC/KjCWzH/fz9nbIBIxNtsuokNhXjK+VvsV6bR2rrnTVlrsNoWbXh/modjZm+c70WHy2AQMmF
QS7R+hHODekNdQoN/nxP0RHjEGN52tcnpeY2InK4nyTRYKXoDAeIzpNjZTgja8dmZzBuuBp1i5gT
hpy0UHjoBZHjQZj0ubiWl0+TtXXKTz743WQ3jW2i4kN/lCxmYX/n3vrv+UDlIXLe+LLSpzB89pbT
ABvKZiKJcagwXMWiH/4f89JXtmsWxuWco96bgSIIh1+zPwWMDewb7YK1uIv7pG+WamnrGEFR4o9U
+Z6NdXhqESIDLLew6/q4EdD8vpkarSyOT38PKjfYU3HwfNEpQfoVmPxFGTJEs7rzRPQkJe3vAZLF
n5AmBW/mGCw2JbWvXvbyCZ/dU8Scd8p5UPBeOIjXpnDdxfxvgMPQekmX7GFP+uMcpVoA6zCPqfHD
21Pp80nM3YiSZsTnK/x0mo16ZqoUDK1zr2AXHg2TeEDZFdqwER43Nj/h2aqwVEQJp6BRv6Wd4ijz
yM9ucyq3GTWS5N7NJ+X6D65tfbcTXoyDElI/u5GDuSVw1pR6HQYgJCVx0ufbdro+ZAYiBHvq85Lj
YI/fMxSy7ulxb+vaVyD+ZZOV7aH1j143dPNY6ncD3lOyfYWkaQa0Cx/JE05/ZY9b4Hb2/Fk0dzve
0C2vVPPnxZEQXDdsyQb6TIrfqlDbwLuokM8o1g5gUamPYY0Nx1KFbo6pwu/TTHBR8WbI4/bndGxO
EHN0S7Bi7dAL7HEi+AE8X+WDlP3p2r7BQlE68BtCPahiCp5z5myEBOfk710OS3obv/2h2RQaKNH4
6RwRya27xbUBazn9zaVRDHbNS8NnexoW3UkcIyOg9rZ3viteesVeFEr7vIibx7lBb8k0v9wiGsAp
fBBxCuc19HT3Se6FL03ujqsdaNzwSYyo7YvJMUE76hjDXs21CJoQCM0LU6ZM4QDPFsDT7jXXnEhj
pd8Hha5hHkI+J8qrkutJeDF8ziGmN3mRm5DEz3wBj3Jcvvj7PcJUJ1cHIO2lPndNIfVTME0x8l3u
OgT1iMZ4aW3veWvpPPS4LsF+EVj6zHTaUg0D3859Bi/3wSLRsSzJ8A+mNvavZYrMsPdl3bkUbOGO
RTxsRsSmz+A/ZLp2g+KptYmZ9jcT2QR8y67DNqG6xT0p0Fv556vHfbBxickolli76GNedjB5nt55
ZcznjmX58t5sfdfiG4bEBrzVHwKZ/BF9u4I625DKm+YAb9OlUbWD8/SiUxk4/2a4UNhY8oxWUuoT
BjYYCvYzWqvAQhFoCPApUqKZPIGieP0lXBiBXvLnKTBrEQzbyTn0for2oSJ/Ba75qEZ8g55EoRPs
SkBTw16Rqqa21pMDvj0sLRhlSDFIhV7Xpt5lymxtOf8hdWQcT8ZefCnf9XhofbFXUomWeEl9tTgV
lxiN1Mf/OAXmigcF5tOeYeLKSEb7saT1lZdxu8yQJFAf+Qld6l1sop8WU/MoLNrc8PcJTI/vFHKg
jdQVNUAMDrarAFwSj0aR4I5KofgHtqXlAFAtTppHUOICSXTBtqEgT2fVt+1slnwUg6R8F7IyS+Qz
thDccBaKCfNdN0Qv1Zdx1BVoCPxDTR9mx2u9Tr5eXbbnNDOPtc2ebFCAaqREhC26h1X1lOX/OAAu
aryyBm2S1QG9FFoQzx3lFdShHFPQ016gfBfcl6SpfZxojtdozS2moFch0r8q3x9mXUhe5REXmNv6
YAgtKi0AeQE23O3uCVU4NmYdk4CAbMOBsDlJjhXWajMOrPOQwCu1EXDZ++x7aSU22vo8DmM2ts0U
n9CR/WNCkwKS6a2TCKv/HwoHrOXZUlcNR2Vv+2xDTNh0PNBWYsxY9xeS+wfV2TGN84fpvsu8bXKM
EX8GAgf8QnBJnID+oqlL7dmjH3r1IEElam1ksZJpVN6h8RSMgfZRRx12zjElfT1t5RT2ccC6uUC9
C75/Y2UmC7L+G87GHO046pCaPpkOstauzVmJw0vvCWPQQ6BRYPnAT0DVVgYRg2dAbZYOz+wUhrQh
RBbdqNbm2G/yc0U1wQlxFg/RYn+aV80hYpbyXKKzINdAtQjmaNczFUvQAfIGZ01wbS4lQ+RM2+Wc
r1N41aR82LO8FA1OOmbK7PT3IEETA86UnPy81TxrdHqaMtSaIzS3EQSN1XBkAFsClwKiwyHO0XiC
VBuj16uNlKaXot+Cb69Pz5hdxVd8fM0eN4ZcrXdL3IHltQidg0stNXVx0XqNF0y8vpvzXFBk4J/X
PO8VNmtE6WXdZI16Rw+Z3pDHFka79RnJQnvS6k54uIO/vfJ8rRVz5/7FlkbQ/hZr4QiWGr3Mvjug
bvWb6TmMiA/mSLWq/Dw/5Qi/RepV8inq4CcE7YsFtpEnU7a9bnIi9W2rsMXQKVhhEZ3sx+SD93Cd
m/3PqbIwco3D1BJtzqCohZwHgdxmwn0/kQSgFBt2TcEt4GMZRUdJfJSXC7y3SUS7qF6AfLe4YSyh
UJOAeas9terK6FRN3jyl6OomjWnec+/qjPlRRCXqD1ERUjkBcvHMo2GwnfHgX2BuFmqr1XCQpjIo
SdpZllx2Dwjxqi7u5hzFG3ft5vITlE6dK9IPVoIQHlOnC8+W06/Vd3BsCl1eXnjqMIUY10Q8LDN5
2HCyN6I96Nz5rvF2gzKcFuE7CD2pKEcrRbiNQ18Q1D4r9DJeMo5MhnA2No6vOLVnAXHnx1awcODf
OzUh+HeQ1HylMIeQivtukgcFVeUOn6IYqMRH0KeZjHcyKU3NZRYnPQX8K0Tcu60p71Eb2dx2+89j
Otr60tMLeNEpar5jU/aQqgwNrskcXWb5LR1CJKwhNzQlOPx/hptoYCiZSdMjCnoxnAq3+3kLPNbS
cUfnssByl531ltchu4jZlwyg7UJLWOqzD+J4aNyhgdWJ0w/+D/3TmHggQ35WWRiRVTwlQWrbkYKO
VIeH8ZJmVqAVxs5Wym36t+AJwz6rUw3a15l1pUheI+IB3sdDR5pAYqewwjIXHOFp2QFiUjgl0E+X
0K+iEYQtidMYGBLvyecWkmzTGyQWiN1xMqgR541XGgmKl7Pe4Vi3qw+khGC5SM3QiWYlRQjiSO9M
LPUGglbP9mPYz+xB+fMgVPGy5W05Aw3o/Qq9V4kxJOSr6uZmV0nYGT0Ok6pCoPOUmuZDZKsEx3F7
BJ4JcXySVdRgMQ19uLfw7dh3gJlzhU5Y+K3VQ1R+Cz7iJn66wYkGECLA20YxcFlvQQf3Ly04hPj7
ULEIOZ+Ag7R2srUQcKSajGbHFCIF5Reycnb711/nyuNelOThBZgLVd77EfkkLzb6IK0Tz1Cw1Zrn
y6UaRpNHp7FbKhW7N3caLKIxc/OLzD+xy/bbQE9j36pdVRCmIddbO15sjDGSEn5UxEO1pivZw7X9
YWE9yqDSe67gs4OJyQDDmUcxQi3mDCbb9Vn91k5E/0aHzzBVFSxytxx771xKWROKwSJ0LCGFS+dX
+K1F2LzGmbBVL1O4y5sb7nN/1UtoJd43x+TY6W43SZWI/4mlnDtQqQcs+Su2PWFPv2ZcouHF1SuC
0NmgHXnDZOiHEIsBIrp64z9nVXO2SWJGTlG+GtCit6rCYvAsn3vlJN6K9giDFvQ6bnSRFTONOCAb
ln5KF6F4fqESPMV/WiLLP5ZtVDBeIEntgLE6jOF+L7nAEb+NMo5ftZqCgsQqu2HhLoD1dyRw+OB+
i2zyKK7G7lTn7h7sEunIpc8z/SEULff0QoSReDa5no6IotS5xMOF+CMEekpoSBh00rdRMfqqJWQQ
X51ZLJryBalUkzqumSD5juvjmtc4XLHsJ6wF0K1ht74+5wGeCdNyRdZk337LQ+gj2csSjcHZswvu
VeOWjqm5FvnKtNfhntWp6CEnO3dEJ4wprpVscemzoOZk5dMnyhvfqtTq6hBrDvSTDxQztw3w+b5h
xKqH7goAlxexNY1UGA17SCo+ODS0/UGeFfXQFGmpxXN6efrCEusWPdjn03I+p8tFZP8b/oqK9b5m
TDXwQ+6G3oHIAvv6nB0KFEFRNgSdV1DeMNyT5f2uLFXlboJJEBkl9CfDEyelAHo6DYso/Ck64NI6
g2Yt1txJYJHsPhkq/I9Y1Yn+etcq0ntB9Qd9kvVWREfVO9crExJ/nl4mInnDmVpqeB9Ycgp6XHto
nYb/zhP5rimxFnGuYuZwSGFvlxjifjlDS7on9ujdXdty/AHHIh9JkJNpDmjWriGGRRRw6gyKg0B2
9Y2MhnrmIVFF9vM+E9M/73/PfQJm1KxDZR+WifYEgHcHYwGt4LJw0Vm0NSEa9yB4AnzbYDHZOZAa
rL5zuJvia3nYNdkr7QWrjSzKQAp16fSWoAb3gPCh44yQKlAfcjZukMoZ7Xw0/DftejHIdwF2FGwF
o8C9OeAjlila3Vicr8cgO7VY56a0NglLWpry97p38fB6Y2NtFUxC0j6RXJiTPwoP2vyTzEY7fUTu
ZrvllDvQy1g5MsrMDD2/yZmwAQN1qW2q8Hzsp2bWSow/enK7heuEIGymeoGoRT18FFjlnLQp+Bhq
zG75Saf98ynqOJoZEF3fxghm9sitMyhmA8eYazGET8xDla5+gutaIxQgHT9l98Hi6M3i5OjC0RCX
wTM7CvZTSQ2vRUs73IUmpn4EPXCNnHP2X3OjPqjJxePeL82qEnjyAa2Dq2ItnbbKlKGyGTRsE7sQ
4e6l9mZop0cFYz4Nnjd7eH2fzra5fgCcnnD8m4kQvGy/cbWUpQWaL/BFVOcP9+qnIZ4NakI8/Fv9
vLDpp5hIvoq7BY9tugmTD4Js6//h1NJa6Vaq6vf++m8o+nOWxho2dDt5lKYzOCUJ7Nqrd6Zj683v
x5zzwXYfDjJAFGJ+WnrlmqdN0b9+zL598IabbngkogTCDB6f4nr/nwP145WwuGrZLrzkN0DEisIX
5Ovu6P4GRyaKo+ppY4qOnZz3S2L90LhzLWTcnuzwYVO+QG5Xg88Z1+mZcPsbNtN/94C9vRCzCMEM
49uHxN5PWPlTu79YbzFGvSs8CwOcT4rzPpP5/Nl43qRqK3Y/1u3SyhQC3cCBNHF7cLbPxpnR3Vv/
3+pFwh1sZ39m6eb2uqmRNBs5o051+V35RAC7yM6o8ralkJEVpfDR5i9YtT4r3VSCkO+HByNwE/sh
J2Tm+cC/YQcz9JBhySGlZbF6vqQGhyBClfWVxAoKoR4HssRG4cH0mRCYzIzg1veRn+hsefqQMqAf
IYXvaZjQcKCYHejs4y9SL0KISBBTZolPyNZVKBgtjq6cmgHQLwWAgjdBiRHPQEruYmvH/odaOXFh
zuHxmPPqh1kEY4H2I+Uq2CVWc3XgewX39PppAT4IQ2KQfla8QuT9zKajDMF0OkFTlNIsEBIb7jIB
WeednTR+yY7htBS/IOIIIaaSFzxgwvEHdN/ne/UM+lZJTC5NY2/q26o/U4mVfEnbJRty4R1PO4bG
Q/HSTHwz+WPenC5+YKRix624EVEtb3y4Z66Mt5hGSOrZDGWHgZIH7fFSukR+aBdPjfXPVMn2QkGq
BNXuL0QsSBpBrC1Sl7ob54/ucDf3Bt/vEa9ZussqQHsognvGlERaopkxPM5duVkXkrm4+CkrL/Ic
FFgyzjsd25ACHGnHLpUww9CR99lSVJTRwNeq54aopqdP4L7FUdC6gt7ODuk31zx9PS2yE/Mj4If6
Y/TyTcCxn95YJ1yUg7z7jeG6W9FxnTTkf/Q8aLh9v2klQXy7lsAMZ7yXGngXvPfZlP52lx2HjrGL
l/B7RXWE3M9HlxVH4fJT88ht3vZO5JLF5TLrmZitPABrIDyYqvJ0Ebks0QxdKFgQeJvIwalfI557
tOIzX9kG+6yFYcjkPZlXT+bgfju0pzI0XXpsEwDspdaLGuyzVtPnqQs8mtZn3s6C4WbMMvC72g7X
Tj/hh3OBWDrSSNDNRyShdUbrnhWVZdQC3V56L4Jtiv3BLAcJ6/kJy+s8yqfa3WDbjMf1xC8A046P
sIEdr15gYYRLDEK3awefaYwuszogNFvxB8iZcssgcM9/0aLI7/MtzQwgAh7R7JQEiioPr7hxH0VD
htdnWPMSR8A2mDYkndQvgVJv9pVV5gfbyk7MIHPAiqeFG2ctUUMOdH9gr5i3w3AASB5PDA94yUwX
daHULdhGPpChvMdMvCqFn/oQJZpC6mhFHUaUDGXD2xSVViLtTQUr/NdzzbWj6svRAvWKo8MZGcgy
pr8y0Di4JeQ9e5jI9NlmC40VZAvP89Arc/4MIiyQR4fYZkNcX9VXdcRHqHzLcvpQkRS8aKex4Ecx
IUi0OnDlOluQEEaaUzRPDkCTjUqU71jVWGt7wFzMfRYaq1oKqxY+Lb6mHaP/LG3P6UPr7HgURCU/
HZDJGTldkqtnOqAk+d+2+SqBZH+sXz+kfOvbl3IZpfKwul1E/xXR8peVW/r0bXtIZcwym8CV6djf
D1cUoqKttNuW5jXHWpzU93hGRMkEauxKUMVTVWwnK0Z9hcon02+K2atGXuptFElamFciXYXVd89E
gNEYi8uQtaJb694AzMHztWK1gEOIyMCFwOSt+qZEOUMdw1yu2rdor5RM08ugWRtm38U3rJbyH1On
H8AjEecRzonKcMLFrpqlqkEYL044L1G6ej8nYHsTWWb4VCBxkdup6h1MQbHhyLH9dFrTtdWLN4Ue
TcbVwn+HoGoM0j8iqYqBEotXTMn3Su7RVy9bXO/MsmXd7uwBus/dUQv/MP5c+TpZp43hUvscmRik
1mz2tJHjcCbmSWpJ8RX60ieOq6bUx1cPZoFFYk+vl8dBW8Qz+Wnxt1bxCqcqVlcbjOWrzv6hNYrT
1F6tS2H5haU7MlRJJzPt0+ClM3MJiIRuXoYdSMSOko/plyGbGAM3BJOuApB32zr8EStXT6UxSXTd
62ZXyiRIXmQiKJlXAR2sdZr5IoJJE87dbF3gskgJpp+7GBXAhgRwaMGGb3f0K/Nd+wwJCtt3ooFt
MbFxV5vzhjOESkq5zO+hO9/0v7kZk3GtoriCqGbva66BB8Tpv60aYEgZtIlhK3z26NNUNRaOBRfb
huNvsLdX34TJYLYNliMJI86ITj58pFdKA6EorsoTuGGgdsqeoAu4lKv37qtetQayEaGnrjpZGvJZ
JI7x30Y7Fi8jdqlkWXi1xd5JHGlC+Fh1l/3PJitpYM9SqyqpIlG4CgGT5SyJNMR5/1x3pr7xbrhi
XH7ECy0dpf8bKNqcwB34/Tj8F6I3Z+3rZLDwuCYKXzo31iK+L+N3Fu+tN45uH+7G5woCYXF88Pla
Zw0q9i/jQ8TAMnCfYbfgYqvW24b6TQioFBwqY6aBfvSDD4yScrxl4xoGsBqNQMe+J0RmCHG0wb6H
4pwLfOiEMRe9ZaQy+0L5RX0qgHQMTaE/OMzZ7vHAq+Jc0M05TSvrbg9RKSmGrb5nqVP7t2aH2Rkc
fm9n6k+WlXDpRGgYPnVNwJqITRLSFJRyeHxU/gDP6/mdoObx21MrqYvdNPBalOKwmFF8T9CSi3yN
P/i/ISRxyNdi9c+EEkV2+QvVYl8lj0BEumJZiEyPb0Qr8CXt6/XAjo3nzFNV5t0M1ktwDhE8SFkf
5lE3uXvMAFoA9lO1WvauZXTfkulnRiL8LQyKBOh9eUI49hEZs3OIQDl/7ltYVDVUr5XJuveS2vXw
E/Ry3InsIdRl5LA8Of3APl583JJE7U5fk2kr08QITTNOohiMeH9qOeVej1K0M75PONtbiqeQ1LAN
IFwnlVHPTvi7kFrISkP3Zy4GNqchgzadWpUFHkapYcBt9Mwx3l2p+hNmV07+rUnZ34yngPswcHHU
YA0EFWiR6S0f3ragvRWcDEFnCBVOSi1QU0sQcGIciBDSsU7ibeyBh9cHbAMbmrpdyabTYpflEI1u
zSjb8gbzmNB3pnEUzKjJ1R2j+mKic6E5mlORXeXcc+ZYhOlhtOrOv24Qsf1qlcC/Tvzz6Gr0bVKD
8hMyM4Zdgh0mKA59aCg1NUuCiUMz3ssZA1pl77r5VLxX4RBDJ3LI91x4Y99cEDsfwBPK1oSmTDyf
9gtga0Wg2DY7eE6bq1VS6f9nWwdsFklazuK2acFVZr9+WF9oL+ooT7Oxj3CtFwinwh3F7pfwcc8e
Lm2hR65MkRXAjCdFFGg5NdKmL4E+lDiOMnIopy6/L42JKzj9nvHs2XPf65xrUR13wX7B28w9jW7O
g8Fi/L6gvhRQO1gngZQKa0+D11tzo8tplRszNmyn5YCq1kGcRaCaOEvzIgdH7UoCJw+kecUYEgkR
kEOYWxI0luXFB6AoQwbJNDgQGV4C1XNv7tbXI7YpOmGggPMSUsQ9u1Gl4FrylGWIh813RSI4rbTM
kQ2c4bMJ+iTmHlaYTEuMNn80U2ad7dNaaZAK14TJJTl2IFKXJ8JyayllEMySqDDRkcUvUGj81uFY
u6d8Ga9dM7Ci7evcUsQGi2enEeFfNaxTigcyc7ytnAZO3q0LGKy4/VFfJYybfHDjy0zjOOXMxDaK
uAnyLYb5MWluToRcVv/XbYTRmOvGUyQYSAS9Rl7UUJOsISLa344uyc9v0SoVwczYLCfRRbd/5F8b
mFA4tow75LN+O0ObmaWeQ+MkDppVS//YUbEzDXhQpvDbvCgdfY9p3nbG/t3sBwEcmjWWGHaHR0JZ
iXFK6GuEsQ8UrWdU4ajBvGaS2OPYNjyds5sv/7hJYm2a7EE5XTY9M586aaLEnozp9zDy0Bj97QGi
njbtxmVX/mJC2BlypOmNmiQw5WTUAshW7BOljazF6GH0zZxRSNc2yUNldQ+Ltgv0lc87nfLD9OSc
Z3M3RDGCBeGnGM3bGZSGCGs7n+7OYMKi8LncM6lG9DeONET0dIpNis/IgPTRYCLQQAy3gj9X3a4x
//HIYzLApJF3L6dNz+VRTtTQcAVSZtod3/rPxAsyhn5bzKgXQEGFjMPPqBZshh0SVLBw2ud+lYim
rXHNelCrJWggoQn0Zb1NVUCMdsoFC8hWh+TQCbKN3l1VxmvS6tYVAGwmM0QPNat/PWliQN0r1Mij
M4KF1RjUbdjE170aQCTcNZq1cX4pjOSD3Gij5I9DhjLXFacJjpqdC7NlAKAaIo2WIno1mUNb8mhP
ArsmaDM2oElJCZVLtOM+buONR79x64gCeywBWFlbQBm1Q5zf9YyIZPdIp0QeGQxTYEIDynvQQH2S
8ie9Wsl8ZahSS080aRLhsQMLgND56I05M9JHQuxBgdhoxWDtLALw61vX7nz4mlzPlJtuPq9gZO7f
A3T6R8P3qWXhwSD82nLiZofEWVfEXQI00iVBDw1LeUOZPMpGtJaupAXEunrjd2fFvQB6R6WTvqXP
pI02BbdYATn3OKAXYNm/yA0k8bRqpQBrwty8SD2Cu4nNt8DAVyOXjahGPjnWpF0phX3R0Yn9jc2D
wBvsMkxhkaLBPwPSlfJcGzsUSbAglLZ0BUm3FuYC/9Sy6G0bYQ/efEcaeeWa1XAjmgaY4M+Vwxal
66g2HTJg5fBzePbt6JSDFJKdRwM3y19Q5IBa1rx+V5S/t1lVQoLPifFKR5z68nlF8yArQyeSZi2+
xT8EunktZSRVot3lXICEOr2ZxHcUw3/+ZMOHnHUKn0pNhSYuFElY4vinv6MstvZPJE0gafHf+TWS
Vb+sFKjWsYdXKGgx5sx0aw3JErwRbAC2l+fLKLRRvBNxVGRfj0Att0RjidS9/0fqhygagXVp2Gj7
UqRc4Em0DPMj8hqaxLwWgzWWAWBzM+f8nZkpWFOr7WMM4ozaVUwk9DYmbtIuuGCV6+jGrE7rLSxJ
2UFCM8wlZfrnZVzoOsp3isxxgAOIckmXU4HDViLfxYYMa+JUzeuco/Fr8J+kzuW0SmT4cdVjcrgz
5hOfoLJv1x4pCmMZcqMfxGLrw9QTOjeUe24N0JglAQ5v9YsU+U/F6g0rLdo/6u2mUgtyTaVIW2dE
OWX+hxVw/QgRlIpjSS13U5/l2jEZd7FnVa/1o/Hmk7u+tfM0tzz/KD5hpP2x6VAm6zQzad6y6nux
pyS+7KMSAv4iMoXvbge3aXIVyOSmlfUSnawQ3sBwEjEnrjzg0lylnkCuJ6GOTwpDHe3tj0r7D5ed
U1vpk8NZIZBDGOO+wZe4eeaE8TRYzDyjBn0zh3j3ICZ4xkmZxjhwkw1onagXpNk4Q9D1i2bAGQ3+
ocZSNRqVKlixV9RbOdMJjnyYnAkBylYnJ1yBkUbE2u64dqtdGqV7InRGNXjrj8SF3v6ZCiM/oi4n
ack6QEfnE740dQGIfRsShT3X2Cid2PVqmYy9vgl9p2aC76iWB3hNMpG8VjIoWmJjiLMSf0LJQ6yk
shSSw3faclgQGf6yRQ9xJVtS6V61DP5omaHdXt/58tVnBqd/FegxfpqNLR5ZsTEGy3sqB9L1vK/V
pXmwjvoJ1dw6B6sBMOkyc1mLQWxs+x3fYn8LwnF6ltUJyYAUgi/kuCA0pSRQ6Drze7h2/Wmq7kWt
Tt0bxLd+P9CdOxtlsOS0vOdofGCGm28nQ3AfiXkTa9SYXX/vYTm3oEd5JZUv7IMAIVMMFTczPcSz
/uD7jtPLZYR+Pnqk51y7obq5iv+fTjK7+aToaKqxUpDT5fvWTQstKQra9a0ENDaOR9uaocIRvDFk
wfL5Oi1voOXlcxCecmSdz5KwvcxdmKLWfZjKFd6RFgqo7/7405/jhpL/J0OxwG1iBHm7MBdXVF//
nFVs+wotcoSPo8vPhUigxgnV/d9p/gKZ4R2shjR6UJSXwcQYaekhwloHHZC+Vdpg23mo2Yvf1T/p
QPDiCL0i/hT44/pf9Ze3f5HQoY4cWfCgSlQhDIqRhEGBCHK2IQwNYOxvfQ/UvaF6DZ9AA7azCu1g
Lsju2WNb/UM6Xw1+Ua3Sp2Jw9CBg2rQDQMzeXCQD7sQPhLBxpP4nnAfept2bEXasWnx5PtBK1vq2
jt8ep695RBSqpyySzlMcXsnTCwYqsU9oQoPEZYpx/dMsrd9/hp9hyTM49YSNQ4lib+qblrFLp3zC
SxkSxLKAJkUHLopCM+0CpqHxlPN2BBTwF+0M/6rqAY6mj9uDPV1FECgXAnW3ur0GDCpnZgyw/nzA
K9gmaAZRSzl1jFDNQD24MADsYKSjYuJeLrvQFBHidP4rZJwSTaFAyFHlNLuMovGA12r9HcE8qTXY
ygVHKij2szPrTCOfI++AHEB8Ws1rOxzxuoKRsgGDsq5EcKOkgeCew31MmtJAID5QRzVLRsL93MAB
mKaVGL7CNxfn4bnFgzVgvMza6rQFGgOi6dh8BvZzNoc/VXak4IfaPAX/79KIFo3rQahBjTr12rwG
y1h8nhTpUzU50eLvj6eLUFrdhCQTLw+HO3S07lIV+jfbhblX51Lz38F+u8fvreB1jXggPhHfwwtu
QARc6R6ZVn/u9AKd1sJKtVt4jgacEOG1K28uZIqMqT3zZ5zRZ4E1Uwwlz/p8zTpJQc43BSIjD5d/
TZOkTY6fC50W+3yT9JqfaZQ7fQZkYaYQaaYdkxbcdi26hJH4PoMqcPSCIUCAfX3SO9qW2ggnihCQ
QecsqmnqH5QSxuGoMLRQJ+GbYN7DsMMbyalwdn65dn+wl0y/nuSGo9P5al9IFdLnrxLJHPUF2WAD
qY9WmeSlVGlpYy4+rb9MA4QA5d73H96WULrTNK6/UPe5/at0/kiIZWNiDtgq7ANgOPtB9vjzXtVq
QwniySNtO/Pqr0VKTQdSce8ZvVgU8xgMdyd8oYJ7OHoy7s3LPPGFK4kgFVzvtHdbBilXuIeiq/vj
TlfQOq6BDhWeTSYHUD5wN+qL/BI9cA0GLRumDYWHY95d6uGs+atY1jq6r5yK0uPtNvTf/f2ZR0C2
f2+yuhAZt4iFM9wyPO15FTGLnPE6BTRSh1Ht9sQKQ52fANpJGzUhLqE+7mJlsV1N55nECNuqZCm0
v4Sy4wQufAqaBTk++9WJYmz7b094i74wt73AfEpJQflj0gRD9QGmqRLwDB6DwhkNAfwdLqceC1y0
/ULE/lJ459GgEd3uJEL8ZvsppPn2zR0M4akIwCEGz68RquVynHhuJK18oCIak+RB5KJcLEMhfIUu
c+miWD9K47LOhEWuXSSpK7+qgfkyUnA8cvf2ddyT1DvLLvz6ihJRwj/US7ikgWiS3ju7R8xVe2z/
WkWEZt2i8ektmvWo/vlTHiI2OFXWXWaBXShw7juUN65UjTGomps8Jah+k4bnP9bB/ilESMG0rMhu
4fORd7+/rGKThkh71yjGtHzq/SFT7Cx/n7GtyfNLjeHYEmVITXoElOFY1bG9mzt6Gq/2JBaUyco/
qRaifJVoDZWoGOhhcPQq3tsyNZ6lC4vXHr7sBpeDJ4c0vTZlvqsJsmuAsyTE0WMh4KZKEOfKE7Ut
P/oByKY5u51X9RUyqdeI62HdTdW1fTdzam+t8FHZrWVmFdvbZCGlUPDUs3fIA8bRklIYiMSK8COE
FXmAMSDMUh5ckfPwqoqbxR6ddxWrjtLajyaxpZpOQwF6cmnautPqKo0PRy8eapLiQ7IV8QtJrdXT
ckHbbZW/CErmNkn0H5H079JxDikJJerUJVBAhOnXtqfT6gPGO2OlpsuVjtT3XICyt61noOj3x5oL
mEoXXiKEsuEUsSgutTP8s6YLEMjHdxGAzf1dpnEWA/OYlsrWjBPqv0CFttCciaWpxeUkFWnujjpj
Upn04yc0JYp+R+CUmy98ZQr4dszqHn/eH9Mo1Ox/fnxpJh+g336nIx/A8/NHLpxrSTCXET93Z1oa
E52MInCUwTLbfRYSawN4oNoKAys5+4pA3OKFqcvzulCao78LJ7YYmr/Ux1Zs04GxUutY+BHgg7Hk
l8EfibcV6oJIg1WS8Y9Vl7lzeDeuGvpUCxCw94p3CDseqiHl+z6ksq94i4vLNviIenA1HloXdyah
n/cnzCPk05ED5vll+tv7zpDOSHswV21I/oHbPaeqp4/+3K+Z6RptupXHNuA6XFmSwwWv3RUEofcQ
a3m939pbHA4TbeVR7KVBmOqMEq9KQW6L7/qlwNeEgNiKlatWIhvqSMji72iIVkboLkvz1KHXpN3r
34AQyQNGmXn9QIicbHXL0IfiezuAycnUWwmOibb0YY3O5EKwno686ozgjJPcrPm25+RRGeMcZ9qR
V+B3dlwZFdVlP7YeepplDfQXRSXQ1/rR9X13M40JKccuGDVIlDHU5+nHg6iTpSNLWX84VdiRMKnD
uuZicavSD1tqJdtaGVhidAV8PKatPb+0AxKPuPl1wgz4UjZaunAfuFxTq5n5+VHw4Esp1uBLlvzM
HIvIDZFcVV3nmwLU/P5oCLgkWzVtPEjr6Oypjt+jFil3N7iaSDD8o5B0D0oN2/LKGH9JejuRabmm
wyadd0ZlHlmNVCVAh0EZk+e8VdaOYTXlaYMkDhebj3KJJi3NFfXbp8Oy4br1hVdoMudA45nxXB1I
BP2sRg25bDxj1vBaYnZpN+8LDrIOL8ncDRHhjeePUwJc7R99sZY0OUGZC60EvBUyY80+xx6ROp6b
X7ylTpBPalY+KdVEqPPwVLYDdZv3Y8GTwrKzZSJjO3Ze7OxvFJKa5GvAJwwr8G/ntc1ofIPDogw8
W2ybYD+KnCGCJwUT4ZwYh0CMB4TWQ8RAPjyzBPu+MGPqoly8wAJOEtKSQlJBBogvcC5aieogKOo0
37EUeler+ubTwh/hpv0FV4PrLKuC+x5BR5yrNW2upS4e46b7PtG0Qdifk0D9yv/stKUcfZV/EjbP
/20exzvn7IAgb0kpF7b3MsUifb7CKAVr6g6RDy9JdeDPam9zuuwro/y+ZEWy1ls9cE4RYK3M/qwE
NB8cEVA85YJ+If7b0QRxyIcMhWXh0ZPCs1QRucToNU8v3Mf8JyWLrcd9meTQ716QK5EUx6+x9dOk
ugP1jSMSiEGoswuKwBjoZM+u1Lz/p8grkGhOY5rp7YGdjcvl30nTxTtyXo4a3xN8zM2pzXr8hvHf
qCOgSgT8ehir8M2JtGf9dKS1tvP5zKS0OLTS32sIXJz8gE0qs7S1UDaxOE+KoeMZXMsNVSAo44Yc
skmR/s24omR2rrbdqPkIKUNVah0F6tPd2PPz5REpxXwuMHXBQKO1Q0dcUsIHL8W/hKOn1v5b5N85
B4e8PMy/ww9gk7GzVdLPfbAAmK/Oa1Bgobr6w0bBYfcYn7lfq39yXFU6MCc/h+aHB9hIEYsgOg96
H3tj4xqx680AB7kgDRBqZFtMqrDCdLSG92P0AhSzqzx3YYjLYuFJSe/pXm0w17RxQYGn1jrd5fpH
5pgTpIZyjQv7OKkEvaDkg91GG7VK7taX9NvuNRft5R0BmzAFRQ4gzhJuPegJKhxmBprajJebSJ55
d/st8P4HBITfAWkLTBByAXipE+tLSrRo8v33c9u4OzFLi2h+T+x/8QyOfcbxifZ6khwjGDAthdd7
s86fValLtWuOhvm6xn8YojXVIl2DEtZPT+X7kQE8F/R8rplN4h9WNEAWjGvS3K32a9kCLCjhACV7
nUQr+ED5XAa+P825uMmppFBhlVcBknCSCcND5luOTqyZExzqwtA1d04mIVr/h3eSogpzAKPrfzEG
ORk5bUNVhSg2NmlgkLYNkM2u3VhlJan/cqyWvAOzKvLv4rqrhSfLRk7XjHGSI3Ky3QZggQOkxx0e
w9o3CFv8WwSoP/7ZrDmNM597CIZpofJWl8HcV4oRFXKszUzwzLM3SVcIrPIotJ9xPQ9Pwwz7gzPt
rDkrwRCKYSE+ybCqD7yijqe0Ike8m3XrkUk0OJ9IK7dhUIqxRxYOoO4Iq0Yg8Y+dROEhPo+8g9ph
6vuB2lpB4BhlcUcOgnV5MV7H18zg50SWplsNJ/qHszfm9K8dFzkWdajyNQxh2d12b6vNA7hHXTMq
M8SshULEwBTUrabPeZJg5jLuBPSfzK5edqbVQhpKdCLQ42gxrRKneHobKJ4dgrl7EgvhRg/fSI8T
RGkdI7bkKL93MHScbcyYtPSb9Jg+MQ75L1aOlKn8cYBLftUMoNWur0Unhrza6EdDW6m+QuNdEb4k
XStYtaFLz1uq88HFBmKvv2W4M+BjW+9iBUr17pS13oYzViMz4jtOhvoMy9c0yofYwyPn3wS/Z1F3
zW+piLuZdRioC6lNOiBo9+27Qe/UblP25k7V7h6NIunbqubFgfz5WUupjlZbcEnsdCd3gj7RFO3Z
chUkzIxr5PkAvq/WnzeAiXNiL9/Qnj3hW4r/slMycndVa7NgALPDg6OrrMh3rkXW6/XoBdjUvUZg
nA2jZdpgCHvci0CUlj5Lj7lVggM66mULzTPwpzCf0sLB0EtifpiUGlDbDCewKI1SkULJO8/+oc8U
78kxjPeyMmRmjLdIeu4VhDgepyUqeZzdku+8qVpLdwxiewrgNz7WZsPhScMKp1xX3WMIVCrcmVbh
nZVeDQ9cOkMx6reE+TZcgmGMpHGhdA70ngl+2fOP+fjtF4h6wKu4HCCa5Qj6S+sGhp/c2LCCZSCH
kVhic7VDAnCDJTu+auq8yaRzcKnYRiiIslRjl+7+isZs+7Q+B2DLUyxmHkKu3G/53kzVt/lkO3aV
7q1HyRdaVd9L3bFytZnq3s3Q4r/wyXUYHeu67uGujdzf9rhvxtsmB/6z5o3puqaUBafgi4ISd3h3
P1MCBEAbj6b2OJ4ea+4KWBIGeySiMq2C60XFR6O6aEXFd5b4wiy8NKwMT84cF2bR+uI59VG8SGF2
D8IObNwavt8ZTE9KvRbks3R1Zbagh8DPl+iRigYaPlvviTJYpAikMoO5J25xre0HlzOoVcODlVR1
PBrGvbXytBGB2aenr5AAuttqhi9Kgb1yAxWe6ee9e4BRogi5vj1CRJmWM/UD5qEXbEjh9ad7jATr
oLir2YSzyHP3dAT3SVqBBqibG+/BMBVCIrnwJyoOEAqr15VlL9Tb4xBiVsD/oebcLCy8o9jv8+Y2
Xp9hCz/VWyE8AZt/cXWZ6acyQRKRHpUeI4VK0svB2i9FncAPf6eDtxduBXbnKt4iPKIiyM0bztzE
lVtFXtUtwRvr6xogenA+l3t9EwoXvWpOntz97aVnHSY9YRVfPKANwjXtCLX8ezoSa4+qRm3jM75A
9t3ePYBXKqwVI6y4kV1s5IS6UgBMYwO+RlA8u2nBF5uc9N/BpQeINFPkg/l0XRd4Zrv2bI+rUMds
alr/Sz/Xv2+Jegb6aRFIlIZIQdzjy7nUHTYTcMLXZK6Z2Vo5C8hxcDtdWEAwnzAmnbwxV2XzMAeH
lu5+uQG0aqTgWC6PmP7nNg34yip1WCbugB9/m+And+0jlpeLMwGaD29Gla8jnEeUfsuaCx0RQT0x
dbYaHCNwoDCBwTCVJ8je16shJXPE+PcJqxGC6FHE7B0njIcRMrqkLBM80MjSqNuIUP+jSUPLDy28
qsJ0OqIIL+keeXY4IaDmQNU5jr2zFzfITlurZcVtkf/+MUrctHjXk6k8vJZ1y+SeLzFhaeG5uQE/
XwID/no3nj6IzjoT0Oj1S5L6oHd1iBBM6WhmGDzWmCss/1mKewncMcNg5OXdXGu9OWc3TPosroYl
ax2qjbjg+UI+2MOQsfYiJEXd+C7VreQuo1J+3R1Cj9t6hP1iafHxbgzqkzCTrRQfJ/k+GeBOUJ/w
LS7ZzmjvEVkZJmY9eIvu8vvvOx0uZxKE9MdWuCyWfyqT6xU/MhzHjOtqCZK8ZQHxaWP9ToOj8w9V
HgebxQ2JJekE1zJta+jCEXQp8Hrh2so19DXeyvnjV0EmLMvVeoIU4s9P9wpeBKKmUfFJoTnlSu1w
zb3p2Y0+I7Yr8Sy5421EnvswNbh0A43yxcoKK2qklEUHj3JM07yNKmseJ2PFDAiMwmvA8bib1nnC
UV2Dl8sPoJ9HjwMLjcxbwdM3lxCXU4C6xpAi/sdVRAFI8WZO5ouUAgUEm8mjg9N/YmrqO+W4LHpB
v0yT4ueAHJaICUe189zUY+o67Z2PIFprvSYvLm0xWUz6HIjVQoVp+dMRXnICkjmmWqF6sX7A7tgA
BJdON8d2dtmqUOpMfFgFxoch7sI+qImgQLZj//MurjJDBdrx6S3xwOmX3NWVOjsL+zaJLWE1MyJ6
gr9Gg1KsECigyOT5Qi8ab0Gv773dwRi2QRQcvy0at/7de8EnJA8i6RzoSoYEXOnxaZRlCJVuI9aY
SoI/VueXNyZKvPZ+8olaifKCAMMcwiHFClvpGIFQhO6MdS6Zk3mI8QlNgEQzZDNeSUsLKtLD+xF5
CjHRxoGnXMojdqCsF+41uGAyEvpZB4X3DlqK3AuY4l78Cj5LEWF20T4kENW0oW5jKL5C7dJhM/CB
0CGNDbt2oR7emxg40y7yDsVeRghGtZHCmrHFaoPQyjB26VBKsv8bEKDH/SQA2SwrekjAFD3MTyVQ
ye5AGgFRyC9pfo1c7Y/brSW3f6BmTSj5hnXLSaQRCmHDzr0cKD3WI1gmRhDtU75MBatOFRvuJSqh
3w7OrNfWdDABGTyS0TYYB2EQ204XubWhFjCgRUxWJyELrGns6CRFBY/v8ctKtFPyIf9oQn7cgwu8
WOcbrEqDd0lQVkzeWjhx3Lf270aKQqYUtidbzdhKdejMMY/zgubX/Qft3uYlpT3OyrmWgFjU3uuc
Uj7lRi0Vq14N1iziWvU+4SBRUWbVuXik58Jdrisy9cSycCDmIF2REhNCiDwP1rjRyBVRzWQWIjVf
u9HoP7EQnJxPUiUYwfjVdsF8Zo9bh6tAMQ8MoKahDSQcuCqlxjiWHOalgqq9SBKTZmyzWHH/QI6u
3dEBDOFRGMAKpO7d0jJs9UNo6RY4vk/TYvFXajGhhcHGqUyVv6AjxvjwEiqh8LIC+cwope8QJiWs
m0SQN4Re+sIyF0P46ZP6zKIWbfne9eewBbM8AOSHmEu9EHkGY4TdTooTqHNiSqNGLNjc+hAMBngG
oVf1YuW+2lEroah/p8G5y6AeTRVXV9vJqU9WsKCwQ/OVWu6zVEWpmmC94vSTovCopPHHh6N3QRjS
pIdV6xM8ljBCMDQvz6fV+vDrAh8w9qVeE+MpeBTAjZhWtYo0QAROq+JiigUeqjgmJrC/0kV9E4Sl
PDHpIbIxmCZsUxFDEUtNQBEDzsyP9dO1WEX7SnhrpgtGqZW9Z6BjzhTO2T0H4PaULXOvTUem/6qK
+caDQFL5D4cxf3GOdBRiqSj7c8vAE/CvwFxJlW1loqjkBlZeCq4ysuOE09mC54HDnAUjytGqP/NA
iN13D62wQE2bSDTL5ZzCVJku42uJHrArw0fh1yqCM+SOgw0M/0n0k4GoaaN0XRJvT7/OwNe3VBqT
ZEapFj4e0TWZ55BVFiz0Iv07seVIZhdzKRlqybAx+/c2szcWod2+S5IsbiKYp44ZyeaKKO0uWAnC
LMqGnd6WblWHWvvQeGwMQAuX5wnhwllkw1zFufv9ge6DVog5Tj+GD2ccU2D23S4HLZz8P4U3X79c
RwqlpTlCn31l5n+/LyHTr3U96Ho6wd6QOavAPUBj4tLhIAL+UvwFjORT7PMq8DJnQq1DTi2mOlNn
kMatotX0akUZ7QPpr49vbJmsfhKWUjim3gKhMG29xNj7Lv+7FXR3njf1tqXOoqeFq/lHEXqoGlz7
gT2QorpYrBTIQmH7jUCyO/WldCSSkbYVxzQ1XPGYnnt6wghse9DTG7rmqKehiph70Fv2VIhmNGWx
bdHQNF6o2u/Nl8BMNpLZF6Cbg1ULSB2AaakAoC7yKRJcIznZhYeVGg0M51C62XV1mGJTMfm/P4qH
KIyU+uS7I2BGCNLWNYReU7YtWe9i6cFZB8PL2EofhtRQ+Lhk7iJXxuZc6WDlc4T6KRTaRX68+RYB
c6Kb0bfBS0a04vyDPTvSsguNCZlFCjMYrXFdqmFRqC+RU+G9jj/38tFDE/8R5UbVKmtpfal+2dfS
f3ivcEmX4tJHl3yA/pZ16DqHecfUhKJW+WJqh66blikRZV3FP99mHDapNo6WdioE5sm9tL+k4NxR
pQbvjj7L49tmimP3940tWzVGaHlbs37mp2o93fgLHxU7wAITT2n4pVPVJfHpwew4T5cfoj4iS6+5
uqV8ds4OghN5PrXbxMOlUasJMRP500IM5H7TfK1L6t9EHub/EKhbYnL7iWNDtayu6xLGhqTvszQH
YZics96giSpIPLY+oqm/8ICi/Yc+YifMyo2BPtav++cFJghr0hQAa5pG9zHj34/dEKjCGdQV4k+C
LC8He/qvYatn8Gl8WrPHQU4wPLPp6pyYRyMwIhu6Eo2L4+wqudhf/smoCIhhzhoJDt8gHXmX2DbJ
c8J+KFOr0lzH+RNb3iPa4yl4TjA642xvLTF1WT0obohFICLNFCm5/DjefMH2DRouk4hjIy2KW9w5
UcyHlEyfZbYKPo8mBaJFZ+AABN2kOBkA6fUJeOI4ioQWusUWuIaHNsaGx1OggwUxlN3hhMYd0X7q
e3DGKs0LxuhRuib0F6pIgTC3fZYKGjM6IMzU8JuK9LQg9w4y3tRqZMUDggzRHrUMAYjiaCI4vWQo
ULxUMVYgxKsVrDSqLngk2WaD/7qRdA3mx328wRuXo6kJTNbFxCGam7UmA0LMrUaGD07DdrkBRlyE
AjiY8SNs8IaenpVv3r8AmhL7QC+QBxieVBYCR4xpY8GpnsOVairZIUIAYyhBry6rBvGeEr0APMxk
N28OQh69CfaK03Wi1ohR1xCH3+7FQ0P5AuhWMn/eax/0Ofzddc+BECLkFnHX2P3BPE1df745V8L1
SeYgXIMRcc9OZpHnBbZ5l+JlTZtznMmBoDAmlhiGa1bsnXogmrxZ0lhKIwaS53tpSFARq+p7nuPA
SCX9pSIw8Q02U17FdbQMqPZ1eSQDp46zEYa5MfRysjKVdaIGB1/40hq8MiaJ3fGE+4JU3LtTiwjS
pg05cIBUknKj8YEamIVjVvICEMpJBK02OOA2j1YmojP/pRgt+CR/weIeafiY8dPJvu6vorWxFNdq
Xp2zXVwW11Iw0ryzinfsOnAGbMN/6RmPAFSOmtIFheKqZ9bM1RJqEntRlc4FzrLUwkIgYifSd8pz
vmFZMuaPAdgPE6orBbaRegbQdV7Rjd3ewXLp1Tqp7aCmTB3509mf1aBcF9sFDhVfxGMZCLQGM5Rf
Kclg0BCzUwYQO5Kg671cLWuEyJDlmpwgan67qDlOH7QJm85Jj3ZAxUMon8lTNXmwpMXOhlfH0gjH
NKMIRcvLHKsw2LcXwLdzN2N0T6/F7Ywe85epMptYvcwh+dzq5wErx/bwroUrCuqTrohQS0XALYom
FUjpX8oEMZ3lfWyuf3+KxRkbIr44iDT5L/8nkn7gbx0wKIsW2uYlSLLeQELH4YSDxklkSDl3fAxN
fHP0Ozr7DvqEoFWtWSd9iYBlpPfVbxwL41THf/bscTetD3Y7dR2X9ltb/yRr1v3S+/fr+JXQbtDU
PzhAwtaM7jT4XS34KD3cxki8U0UqqbfULtxyKSF+erYnXBAvqrRGMuzd5Q7OxfsYYWBpQKR/wixF
qqqXcSLDkDZfKsPEGSrsvBuEAZKlxdFsHp8/55b2wG9lnIVHOygRyn/726CtJr90ZudC/t3Qv7Iw
Ja3TpQidEgp+mKJuMF/AVrw3JoutOxHG7EuoFj5nmDuMjnTkE8XTWeoE/nQzUOaLfHJBxXYckMn8
SXaWzdyLCdN6QZqeJOnDk9fHwr5Gh37q8RpXoDQpyOBeHchbk1t3vxJtwB2bKloSlyofp5hTuaA2
vJDW4JeeSuMezUfRyOM7p9yfWgLW4jwsdButxleJII70+Xg+XXKf36FMbPG/m/L7ssHeBw/Mdd9s
Om/yYo/wgOCUu+kT8KpdqMUaLfMoqrgFn2zD4cGX/Fh39dWaneOc+du6m+91Il/m1LE0FHQRWapY
s2r9Fg8azwbCvzwduTZFt0j+lWWwj4Y5q4Bk7s7A1TDa8uG9tgndMyq4oltdDOLgYpLM1FBxZbVR
xhlhhyqVbQdOVNASBDA64FV3DtJ577Tj9bGeUc/hUZjGa3sHb8pkvYHKTAzKZ6xK67ZQnCSMf7OQ
Fp/+eb8wErK9P7oGIx4ZKQZAd0rzi9zF8DoplE3k9UcO6favK0sWdH8OwUzC43gJwfPMg27CavCf
HZHGCY8ZXB9M2Bv1Nh0uwziXchpl5ExPY2x7am9z96ORz3n6ioG2oRuc+hvtD9/K2JmK0glRYYf0
uO3C1lbYAbELISp8kQzsaftuJm2YPq3j+ctoX1ikfaaYTVBXVHJsDD4gX0nz9WqSdjtRXBEx2+y2
R2N8pjnNXZu41FXmnIaadelkY7rcykKOclSyY6FhrrwrSI36/U9uITluLgkdRJUkNp5zPVGjDBYL
Ha3ktyOFBVCEjKgVg542/9k1oCzqicEInap8evbOb81BC5Cqqag9aK4qVU+ZFYLZqo7O4rhVH2nr
qFsWjLW3rwtvKnxYbhO7KkesyLoqXYR9gZxHsubgq8aJHU6s9/Qd5yCj1MBPsl9thBWJPzn9iHeY
mHvJmhua6ZB34N2aNwml60yV/keyyJmUlpL3JwcUei2kzz1ZmVm83a/o0xjWkdIXHFCLWbRXzcYr
lFUQHzSOHvNAi5gReOs73AkOYkYT+I19bUt79Cd+5upOvcA1Ya4ZtKv794ycGbd+7wrrdYzuwE/E
P3aszXV8UUPBsiRUWcPvSgRmBAXAjyx6sGc/A8yFKSt6Dw1lF/+W/kXmwLlkfFn43AObff4xhWFE
H8/+82DOWrej7m++iS/EP/29NVWTKfnTumv4A5jZVsi2OXA2eBkDdbXudqIGP5YlHt5ogNiNRMs3
7JCz7RDo9g9K4pam1JI9aRsuPulg0qgCSv5vnkkAtFhp80RmVtiNLV9mHSLD0wKFw6pHUnlIu0iy
s9fEMXDAcZXTR7c8rw8h7A8Tqpu/A+3oZhGOBquNuMoZwpUp8OhQy5cei1B1KnEqwthofQ9d9DPr
65ifQVeyoPLsdQyJw4rE+fsrWfMXoNQeLemED/BkL58XTjEAMmosPMnCcemwlJzJHEbJbzVYZwwm
RUMBlSDX6o9gti76whaD9KbYSOAFuV2wyMos+d4gj1rgtjSogxmwXXXHe3DzLarH006MQL962Gk6
avKir9nPYVWC1lRrkcW8g8ogSr5nTAXWF/GAUSGqc36FFMYM77NOp+mS5tnh363Nvd1ZZWSRLJdY
MypP/LM1RG/UWVhGnCoAS+lGsDA4kwB+eaqxeYcXPP2Es6JZEXCrKwfYHwwiEZwQshZ9ADQXz9WQ
jF/4KE4ACe0P8LCoEuTUPP0IbwAju7S0sQh/bj1Wga/WsE9R1ZzkrfTubgjzCAIIG7Cgga75Bz9Z
pJn2+PcVC+7qzv2LNn2rfnmgoOTmNGae72jL6piedgnnQoArWhSujk3c8dAchFz6ge5zpm9mglCU
Sr1TerPvlKxBweFcqG8riDAOWwejehBKkR6b7yXoOrFLD6YheS2cy7h+Mfi7ZbrMgWqgd3ziUDFY
1ZLIohKboxWJsB6r8rJ41BsZdc4F+NbfHenuvGtcuJa2JrkmoD3nmjRiwSOq4tp4XbUpNYDRzkW/
L6j0V++XJAytMquZ/wPoB2TxWNoDu+IuN8W1XLsR9187SDJ1FC2+3h7W8/soTz8VqCRUxHRD5QWK
G8Ff6AGe/Etqr8/+8/M9o55pbFu9FVdlVsrq9Lg7sWQpL8S7GGqDtOpSuCcUVzVwPEGvOZ3mS1Id
F5RVe14ljZ/Xe7MRB44/5+t2+DtdC16SrbFmGZe0Tn0lpoR0wJv3qtfkKnW9/nx1ckzCP9XxOiiR
jGnNHmWdH0nluA7LUAfHwiI4xZhrHoAFLlufQfYqZYRGZz9ZW/Wp/gwYzXhj7uiB7b8RwQDhoVgf
psHYTf+PK3bLS72R3UGUzP8gn97tFlMvjfoNcI9fbBvAOvSOIPveI5c1CvN2Azxn9GOZfOpJMy8B
B87hBrS1PaLp8H+wMDx1lJshaHJCi0c/pWebehvAz1azyv3uo9Kq/RLkBRGoGceB9UYDjmlBEgi7
msPwlLDAzWf5qQaYn+5jLT2kJevGDa4xt0YFYmp0F17kbKKWy2lDyV9WNon7JxC2/6uAYW3idF2S
UCHbEBjI4CooJUbi+A9QXtzNw90X+6lGPqYU+4PB2kK2+D271AMrD0ubECJAvz+TVZtNFwCpz3PH
D1VMKeXbMExB0uxPfQJ+t2qNHZRjxQTUuozICkgzMU5ZHn0IphyoccnVTNunQWzz08HNIchTMctU
PDrUPeSN/y4h3lWcKSrEA5DY5tWqsk/aKT6RbjxjW/R9fM8LoKuv1dJJ2N87QxFDyXMHOpE8ziyX
gLqCYmfRkI3HFJxHCllv9x78xxm6bCo4aKUUCpcleKA9536QWBBKC3Tot7vWbRDgQhMnML+25z/n
GIBCml+uG49Ulxyo0HGJfd5rh0CUOI8lzeWNYBcT96vMpfO/dHc2mAXEV3NCj0MkJCLgkVdbVfaE
wcEey2O346Y1m2iQgY4M6DAkoqUqrScx65/U86PaYq1FOEsVf1D36HszWH+VlO2bb3OvSv6EEEbc
7UglLO4nNXjonKYcd6SMw3qCuhxV9lgNRT87B10jtM9nx/n0HO08sVs6KGiQDdPGhpQ/Il5VyVZp
9L20FqWXS1SuNAf3zUj1CsDV9VEn8j+xULFc34M84MicPp8VuF3Gvv39AjuXjSAy/qNLHGDJ9aY9
WU8o1ZFjpEJFHUVkcwHc1CRias1PyiSr3K0ZXs5xOYvHs64oE7IHOxd8TJYviGZrUfaVpuC6dq87
BbcCnKQ/aYhl+ymjo0ZniQWS9ENCupR+0r/uu5eyimr/0FMZTqqslxKh81FjsX5N28mCNck8NLwK
9qxz0JECuDmf8vtVRYRBAnugnnB/Xa+hHMVYC6ylqhjqUWWZlsYSRi/dGcHddcrVZa9S+cacdM91
8JLqsvv+4oNck2YXX55eILqdSKll7h/bjHn1hNnNminFcIMA6qzv/raE8QtGaeCQ+TtLIT73QvgH
Ej0aBntnTREByE1SYe/Nl9tdW6GCe8CzSTn1eSfdgitqDfbupu/qU14jNho/Ja+QhtYfvRIvqzMa
CRZYXmBYmre6iXAaNhQdVkHFvUH2vhPK9J32gLwDDxRQliXkeE9a28+/i2SvUotXoZW5N/tiDoAJ
+RYu8YYaHyygNSvzsU7YH2ou+j9WiLk4Ga+I6vXFP9BrPjP9FMtlT0ma7zo2rv+YSI0iOy28jncG
AHtGwLCSo1LCAlvd+fhyHnlCuQolEozK0QtVgdMeKN6SBokdK9oEDXfuBPdzoJINvSrSDYc7dCh2
UOTH2ymgwBy67ETAxaP4ouITh5GtWWBBm9bHV0sfHYQflGV9NO+ebgecnFN2JaZ7OWRtzbFVaLdY
VtqapDS9Qf7f3ArKppnBbRBzAsfdV7b6wHpA64hdMxwVhBk4Nz+drnwVXNtnGkq3eYSognSVwSki
bPrw5CNu0xF6xR5Y2IN8JWyHJD3AvPLdssTiGG8BRlIzl6oowh9Qgsc+hciZoDn3cKKSgq7rs456
qPixF7kLzNkd9Z7Bz+z2dPnl5JxKMDtEX36Y2rQ/4hRPcAbWM+1RsgmHIuqqgFAyw/i/EzJPbvC+
5Q5oCVXNy2CGUaFHjrC1SD0gP8eq7bgk8bTVdhR481KWLvTMSPjHvUhyG/Vf2UO6j9y845Rio22q
JKyp4B3ZiB5dHdfckBbsL1W+y2NpGl4Uk17Q1AJJI/GysggzS0o29SPZjFhqPKYMKeY1i/Qyqgni
ep04nHbKxXlzHfXVspYywkRrb5bWyPTX42chclsbL+xZp3bt5G1XHR/dIq6E4vE9gEqmotH1scJU
aHTJcQYn5wJO+Rrp4JfVrls42pUD7SrsN4/VEfGPYUk69A+ZXpeP4HS3g3K1k2qZ041fOnNlIg8x
j5Peh4ZgVlpwgGw7qx5JLsBPJRsjiGcFyAmmBFwwHxgqYDSnLGGieD/GUGVNNGqJSzRFf/ZWpAKP
QlmoQ8rbMzXM+07Gr4vsPSwZS0OFz4SdEI8AEEWoh9tqlgSEcB2C23516tTP+aksGVW8kWw94dc6
RdJg23HFsKG1BiVkEldXL6H2ziyopG3ZaKLUdc4bQIqI8BlBDeKqdmoZof2O42Q0bxgotIkwkgSt
ZLG9pda41rou9EkoRYXP7DJx35VplI11wsUXqqAR/BaxXTOEYc8VDLI2BavMcBoTE2kFX5mRi1Gg
LoU+6wRZlVXpBT3O6vog6RLZ4VmbG+Wz0f7BS89kpFJqrDyBiT7YUzguwhKuBoOX6UztLlQk2y+K
bR3jZXfuaCXKteg5tq9tfQj6/YKIeZ4u9GWaahH7jGIuRoh7WbmQrNeP2o2JIq9rPWNPTqdu24uI
qQhxb41ooqb6oQ57S90KZy+m2kgdzuD+Xjjt3rkhT5WqJx2xABfq6IYh0yZNi6PYUWy5GXDTEOzG
XnWa6A1bqfjdC1z341J56AwMh23TtLrA21n2169AcEr/xs4ZlixYEK10Sz8pXyz+cd/nVn+rfKKK
xPHPWdxizy43Id63IttnRIMfnkTdWTyBEk29yK6AoVcVoDb8BHtUsK3znpQELEO/6pcTcbkopgiM
edZTDw7HLmHS5Dk7VeprwgNinEd/hEc3JX477V6role9+O0mWVQmvRFOck9F7Zho8R2CCOZCrUD2
YNBEd4E5ekMosBt9+XuCdA2gR/7fy9wAu9xuW0Wd1/Xe+kPxK8NUwydVdinsq3u0PrBTgkcw8/g3
b8l4jgpD2jrH5v8IFRFoTTfkJe1899FOn8KfhSjtlBEn4U6ZJCUpaRIJ61VsUx6DtGWlpN2nkPnq
9iw8MLDSHxUhCsaG+1BbRuJFkarP+8YuXgurX4VVZXMlAl7l1F3qb8PY79R7jMn1yRmtJuyfQfvh
N0cRVC+KIrYlcUnLRClzJMs3rbC33a2YXxBPxoQirbwDTk2tSKEF9xLMHWXbCj6oHlH/BgKboTTu
3V1lPxOfETxUyoGzRc56FXBfS713hJcCg8RN11tJjXtS6z5GUznCMFcy2e+snnxZmJNA+IuYvW5h
VR5zmIgwoEt4xANnY8t/EtHH2+fGvJ+bsjSkNRP9jdu4BicFacWpTQOAiIyoTRlYKxESEgbsCCqZ
3EsG9Bq1I4myEh5m9PaB7IPsXh/GHb6Oh6VN/qvUQkQvNgQ/8U0ldAGsxT0MnhKgsCEvvBX7SZBM
QMpCEIC2IdPjMx/hHniNnJKNIjs1L7VkI+KvWF8pStI4m5f9MW4yU29DGwGzhDzb2t6hpcyXrSPF
xIAayZTHOWZpOcGXMbWL9r6pxdc3Z6xjRLc+tJNWykSvtcuB7EX4bZTtuPbu0eYiEfYC/rOLXJja
K6Ibh1+bkvL7tqNA1Ox0CYo1VKe+68W7TbVwCUspjckmtlo1fs2ayum5MipTgmN8E9cQra8CNeoS
i22feyuXUd23vy6uuMvPULcLOfLa5A4ulN5k5aj36CtjH8LBs1P2T77wYwtcyGxcvJOfjpHyTTAI
kjAYbqgxmCiLXfCiik+xbFBZ0wxk/Vb/RK0s4U6e21WeXYrF5Scy4NBUTbB41A4LZH0GroMqeXgo
t7m0tVoDy4BB87N9uiUCLERn6uTzJPaNvN+AIjazJxxM1n4dADlTAYw9UYA8GAGZA9HVeDQpEex6
aAzvWP+IlgzjaSH4XNhEHMWxX6jwm94N/P2aunjzk7M6XXc2+FR56m4h2+1nl4v8+OoZLJ0TNxPs
1ElVkcIEtOUDjvs72fK1/Zy2dYEyeCSA27Yx2oJkufjoLNO38RepS5Jqa+24CkruUWuYtwxo/XoB
fyEzpAdbhUVgllp/eHkO/2rm4JxweFmS/Su7u/R3g4bopbgU1rgMxFwiJ/zUub6C44IQCVaQ8lJA
bYhP/VU/bVkNAK3KYR0oWNS/NTGqEStE/z5WHnK2ima6RKHtAm4TM0f4Xe03+zGyK5cXB8N1/KpG
mKTVKcUuk0cTbcJwJsLw30HQpezBkmXs6D3siyjufVGWDr8sTVtE74k36kK7EIZDJXfZK4h58BlB
FbE3hmhev7qMBaFXYxtroqVOIcAyuS6wdcX1NC4vtVebQLnPjQkXg9JWG1W/sKCBDStrjQS6FMep
eThffCS4CgdT5ZaN1HhZZxQw86TBWB5I4B1qH/ewdyZnqXgLk5IAotX58LhYHo699El2GJDpmi5A
PsplmdYoBOVydsLonMgj6VlQlUt3WUPe38ulvnM6UUkHCrfyO1pV0q8RnNj4yi/K4oCuquyY3zog
pQKA9IcgfDH/bxzpZZfCIf9y8fUnaOuWBv3AI4ECSAlHf5iJy4xfe4Rkc/9xCjyUcPH3N4gD7iia
c2d6KH2L40xPzR+xRNvx1FrIcAlvriUA3w/UwSXVldMbptBgS3xVUdElq9UHkmrlWxaocc//vdLO
FSa26rsjS+VMpMHGWMiFwpzI/eYkS33v+rzJGrPvvWwc/1Uodk+LwDN79brtdKlKxzhC4yg8XLBj
DUUwKjievj1J2VDQSr02AqivSwU28j0DTNzJZTskMaKWQ5r4j86MkXqiMnGz5ZHOuK61dj/PM4pG
VVDg0wRAcX1nsiy9lpFZVjlaE2nOaoYW70tE2tdCnBJSNd1if1bDImkO9FYy68vxhuSZQMUkCXOS
6LFUOvsffjPzyQ0LW+ORzDDmH2PN3mBTCHlCLEDOVDT0ilE5+ATE4SLa4EvKL0A5iW6iQwA9E6MY
I7kdlyRqI4289Caa7jRPNyUEyxQyJ/LA9VuMB93T3AaH6eAo8HLMBRQpcsdxDVw4uMCgCaQdcoo3
3AqHtdPX+EktZ2J0WeBaGFCFlnaDS5TtJS5oTqszbp9r/BJyLEB9w8+wRZcDJVveeagGhHJB2mhI
+urJ3JtLgAwd0CIXnX6Jo58mwXcgbNb9Xu/REZdvcFLyxH8e4f9WxWB/1UnQM/eWYs/LQQDskXKM
g+WvMvk9Crp6u3n7c4Vvpw1J0G/AyrOk/I0sb7IbEB+S4WivxWJBcrOpKiM7WZzg2Vj2LoFe3B+D
/ph+a814ij/DFhnhOe6YzI8OE99FEdYNH2feywPgrKhHwzd2kavossUKmLcvk7toX5CsyLBFEmR6
H/3GjFEeF2urfBumFJcihh6GJYgzk64CtiySqzSrYRf8GT2zkW+fDvMi6bp2kx3loroo51uPZFW9
/GpKtNqGjz7suZF4hbctudED5qWfNZycQ09EIW5inH0MDU/DhgdqledfRzNeLVCudUMEqJemfmMQ
66+LdYPM1BbdE9F3jx0vYoynkr1p7/qd7XsuY3ZnoYbSQ3btvC3xE1EDUpHLQueLdXE8i1qzjVkM
qg3yiG0rX/DC7wwe/ZZVs4aQovwgUBUBlUF2nOMDB8vQBnG+/9nLfzaNXvcGMbydgSRfMAxoKMAX
X3NOH6ToYnWHaXgGPqLW+batwQs+VYQNp+e4vQXRjNb/LIiQZppI9uDTS0bvOqK0HZ9cIsABCisB
fLSgbpds58J9edG9hEt6F+TQu1VDcSWn+7aiBiwGNgWycVuzJWQesco/BSaLdf77dcBSvn3dVPKH
w67tVQ4jWDsjV4DEtuoe79lXPO1pKW+U0YNjaGfKvuaa5ESNouQXPMNOeoWx6SVTu1T2iIrJBQLV
7ofYDp3O85iF8oVyjqAYSf7nu/YmAajKhsYBGnMocFvnPhCgwbt245mSghbffDRx0cksl0U8UB0y
XHc+jtLFz+MeXPtdSoFW90m/NahD90V93qWmV/AAMIhFPb9i35Typ3zuotxtLEYpbf9nMmCwA5Jz
9ijYVvkv6m0YtOillwC7XaYK5VINhmc/5SpxhB/HP9cx9nGwXFnNVr/5msRVooVagk0TYpVSBS3s
MitWC3R6heJ02xMV/Rnl5owjvrOd7qMR3202vc+h0FXi2gN/fn45Tg/yyiYGm3ZowbPu/1gxUJkb
vqNOnEh1oqBEWXxVL1O6ws0F1X7M+MnLZpDjGX8jdYDv5X+6rwWhyNtAywpu5QTIXnGWv0yZLAzq
zaGcU4SNfexMX9+gtC04c9DttYzPAuzCTaJGpPtRUtxnetmfgW1ggzwXCYVIf3lR/0gzsmtl4VTg
zl2x4QiK3/pnxbUUEgNV/bPT0bUTDwJR16LiOfq3e1xrZmKOtyyiS9QaJW9+3NDfYjEDtnbeFnsv
dTZYwusQmm0BmT65Djb7ODsQGQWdx5cFwpDw0w+FmpGzGo4tbs097o04UbYITCUHps9/J8YQwRUx
ck0OxZbnl1X2fnobz3ADpCkiw3rVM8pWou7KQ4vcE4Vsz5RcqwxyCIOV1JUea9/z8PGDUNPVVRab
bOabydsxb7WhpZ6il6Uiz2jtl+qWIh4CnYuJdjrBzOpOs8oC+G5vgEPM2eDFLW0nITZhkq1x5n8w
Bs0nePKFJ/8RFB9XCro8kAksCnjztbC/9MR8tBHhcHbxaiYvDvYZm/+qknumdE31+xrzwjWABh/n
tdUds7UY2LOqXEseFw6uPNGp80/qaBjLmaRa26UHLy+HiYXlQkxPQs6Uzu/RRI3ya8j1ngTZfz+c
Dz0oeAscU2c/Vwqbjov04vD5RtKUlia2JFvQ9AYyUQy8A+8D5kLJuiDikEtixWotynmqw1sm6ZB3
gDPXV+6iL6t+HbMcPOWfvrXEs8ACcuIVdmElbQZ/s0V1GJss+YJRsktuE0LzcU/lVAaeri5m8oPz
B8blm4aWimi8XaUfq6JaqqRn09CBU4amXP/RHWHH7rvC14bEikHpAazRTrqztuzKjTzfCU/npjdR
CwQ1IRW+c1OLTlZBiFnIXEtTzgfSIu8T/mCXnO0Zz1Lo6YRmh+gviuT/kSBb7N5050TTBd4uTq84
zPPYTRnHUjOTrFJvTUzoW5JpHqo/cc6zaycr1UCNKLsx7ZRQrhZhrpRIIwvGBXM8AtQeEG1QAJqP
Iu1viA/039dT5ADx42VWb5/k4Ov90bBuEN2EEmAlJleBdhPR+YX4MuQtk41OYZAbF1LPjx2E9Oeb
MJbaYsgimDL/P3JAZvHU3V252MLK+BIP86GPKpZuDh1sK5YgfpWbWpEdAZcZLzG02tdxPXzYDLLX
1IARAwKj+BuBHkDwyNEVen6xRjQsyJFF21VDWroabuz63v7nit2NXjgAzu5vd8u69BbwiUjnWOSu
KXHcgYVJcY0M/T2K7NG0WBpvEIiQat9BBBNFZsMqHjnEan7icVJUyQPdzNEOrWkeHVelxLvhq4d8
k8hosF3r2tRVkRByNDMJFv+tYwwGT1kcYjh0yLyV+ztLoke93R6cdLgq4KDbvx8ysVcXxOqyaSxt
7+pMeHhAO6nEd+Jcj/0WIhO2uMKSrXCQMvLOWupqwrHf+VrfAcQWU+nDe8womF+7C+BwIYnqijAZ
dskp7AHBFMyd2irgrg0yH0zNns3EKx0Kc2sPKhnFFN3D822sgpC8HO3jncrtvVF6B+3S27iiVDv5
otYWU4WKc75cdN0OwPJvQP8St5R1GEkEUAtS5Ho4kP1CvZN9mzYdK1YupEFBHW9suGNxdgu77nhe
Pml/YIT7IBVULUVuq60NEKj+GAYnhBPN+ItwIT2s1hkpIx/2yBGgS5K4xLr0WSyRDY6LXgiQR60T
ZEvHZ6J8JbIPozZxKqUo6NfTd6YDZ2uVXBkwe+jw00BDVIhBkQA7yig4iLIQz3W6xz+TeF02azLI
GN4Ve24ekcsIUe/jGHFH3+VQZnzyZYNwJigxuvn1TA8v9eInplj+o7wlmSyS92SQWlL03gWz9O8z
5wJ+ceiJ8QNdo6LFh5B/NWOpqmmp6n4RFSoDWdsiUQwoADcJMG4bYpH+JPj4s+KYiTsQtaZk40uE
T47rheN0IGB/3HDuYu1hUBuK2IMiZ8ys9n9NQ2ZWMy9Mvg7gk9Nce2IztfsrmXRp/HxcesiwbT+9
WiuNVPuds4vswyRL9KM2+PTbVFN7ba7RBLeueaSoKdLF3A6OIu3KKCTLVh10hpPz3PdfaefsNco9
AijV6alHpZYNJ0F/gmniHgFk47p3WyhO9DTiT5T+viTER6jLQ9cTo7F/8uy4eAXe84DXuxUxHAHi
6f0OqJT2GFXXt4yV2OEBRfH9a4TPi9u5SdfmUDIOBXDBAsFB4iL6oGblHwjqPJwLtB7hP0qcVsZZ
Hx3GLnkn9gqBNoTucO0ScvJt9jCj9FRpIlqngVgHOb1T3qsfPXFbtiD4Km5UbS+sBvpyRkV/LmVk
sh2mK0RRbpCtgIgOgYURGpx0zmfcYGcm3cGIqhxvtScBhrnARO8xZkypRYsXybkdTFeAFrsqx33i
jsCDPBy7oYwlIm7bPMne4rn/I0hP8AYmtzLWYsRSOv3wOAGyxazlgZMS+RAIP73hGxknTU54yzDc
yk/tCc3PBcosogBJbzLP7DM2GG62my3HO4DSoSL3reoMf1KTwJ0qS25iiP9aTLJlp5xPMt5xUjXR
P+3PEbexhgTyzZdvk1nKlME+KDjBhhyJPbJ1aUe4gWK88PE1x+2ZWDJrbpv31c+VfiWnIbHugzLd
HwRDZxBoLsSwDTNQVuRv/rvIi5RBYtuYREBNxThWrS1Qqn2kpE/4BzViBOHRzM6Tgx6q0lFmXpOj
msl+wbFdU83J1nJMMQ2HNDTdba5T0yKt0zCtDbj+4XqHLQaZdENxrpDER0g6PL7iyfV3vK7kFJSd
gljcj98H4dpf59JPdfR6blNQWu5dw+PaWuYr+Fs4Yi5gJjN3Hfn5/FKldEQREeRh3noNqaweUZnj
+P7BdWl66MdcftKbJ7KhwQZppA2kd7Ca25vET6BErl+Ze5Rg07A6H8mNQMoEi9oHake9dRkMBZgc
nnB0qwP2dw+MJzXIVttzlfP5LuMXskuGoERP06rylliXguPLT7JxTTl3myu/hMLqa+ns+vUYO6A7
xBc5i5sXcPTdyKvbHQMCFY7AEX0PXnpDUDb49b54m9th9nCwJw7HUsX/OrB/5pgzuCfnOLxOBFlm
8aV55OH4OjGjcTZfaVpQYQ/PUmoaDGaeO/pqrg/R84s1r3DYT4Lm0+9kXn/qT8zHLI+Hr+lukIYM
6voRms9TNG5gW9M8yWxB4DTQx4nQzJv0nKPWcFrpttZOWwxjKBc6d1kNaABZBrkSgd/lHWL9NS4l
E2/bFnRzxkcftA/U+Tz52UxuiToWk4b6POzRxvhyylPoM7sM82dQAbjcrS+sUAj2Gx13/LPnIjks
8mnyAswI5/2c1Sn7mRFrIMoT2JfUHFzfHjMITV1onUawvUKhZVsMx40LNIaPLIYau2Om0OrahCk1
AHFLm4rxJPZ/8TVekXgT49inrlk7trqCNSVvlCMfhHAPwUNp5PbeGe3vkaEflG/HRUMc1AmkfizF
Ch8BnPPZZqlSGRpKY5fz8KBZZeXXreCZcHBPVwc6VqdrJHgqpxDwElRb9M8aa5Ri52mgOe7rTV/V
UiBK/cZTO6LQbuAmiI/37ndWTH3++9C+leTuI6m+LawKnBoUPR6f02f9aJt/6dzItH/cm3XwlYNd
PpyjAmJJSU/B08SdXaYlb1+BB3HsWsaAdGsTnE9HsKiG6mc0O5kdcvHCl5Xseu0/AeGzANsfeCbV
0SGrjTTa1Mz50r9hr6qSrINfT3DsxM/IUgYnRfmukm9kF4lkxL4NUZC9l1lQxozYf6ePBQ0jUPQS
CxuVDEtEIlLynTc0tXetwXt2Qco6DV66ito5Zagpfa7hWMXL1quzhnrLtJ+l8Su5R1s8WzXfsNdj
+eVq6jSBYtc5enA5YDCUJTPWamYm+MdY265eCm8CVdudmE6OKS+gon8z9LmV6lkBD5jW7o15dvbi
DTOtHMPbUSnsbd6A+WJbZMTswjCZgGW9nkKUxPDbOe2hz8AZBKvQQJMqYWOir/O21PprwacpFJUp
j4IJC64hSuNESWhiGVtRIWTVP6rHGHPE1bdjI+lbnZ1iqtNvU/JepEr9i0/BYLjudr+iMcV82HDv
6OURfWNDWK4Pmr7WyhkXZbpv3CiorI18jIanBaUXlI/r2xaZ7yeP/ftSeLQxGUVK0juj6LNUwWFD
Te6MvuoJs+LKbvYAEnHRTxlOV9RY6KJvCcj/TMCvqXJ6aCmanGwoFo67LQIes0kd35PfxhF++lHQ
qudyN27DBZ8g5L2CSEn1UQL6b3GU0N89IJAG/gOxmx+NP4edorvBLAKRs7Aa8im1mbUVbZbTohaL
tSY03nOMkD9nEBqfJe2wdUz8w2XC+IpvxLh3mPYaKJDkh7qObVW5yz6H+wu9yQh6eoImiAdWHafE
xgZsk8jz06xz3zs1Q2AubPEsI/N7Y6vLN3+J/YXNNpv2qGwb4oLNFSkFuRN5cTO1ps0tdI7Rq7HA
8dWfQP1JgPJpK0U796y5l6cpOGX3Egl1DFoonI4iylbAJICbaYvqUI6LDqRPrkYLKxlYeSfbDS5e
b2xhFYrHka44Fk6VKnbZWjKJrCwcJM0AOHjYGNxUM2Grc5FXZ4sKKfYSUQ9nz6ujBLp9h5SfVq3W
bAb6gwxwxc4KfL11VFCD+AKcyWVbh0YZ6HnITmhRWMrYcn8hdEfqsd5P9pr6MIWwel6vqx2RABbc
5+TbqTrh3RoROZQ2eUGO1rcbGPwd/nzYwRa+xKJMKDtsE7cX/r1WwJ/UWDIuIc8YH1aF2y+QwZED
ZkFRng3dj4/CE1snF2E+meLSVHbUAvAUZjjYReGB8Ryr1QjTAhrWsNCgccaCVxwsDG8g8kfSmYO/
MzaDRWhg45k75aWpZJ5Ng2i4AKqD8vBtUPDckkoFxT+Kro3H7RDxMjirUJYpoRExfvT576Afd1Vq
qda8cTgp/+fmwM9pCyOO0mau2KYg5tVqcTqMoHt5Yw90UhLhZn63d0UcrMRyPcL5YPMkaKPPA1OE
0RpNsqNi/PYbuqX7PkjVKUJtlJt271LnjtHCmzpyr1q+C8+oG2jd8j457FdL8yBDmmRIbFcKxwSD
HmUS5Q+i8017EYNXs1zFZzJTXKDZ1QW/Nh+4JQvlHs8z0Ebtp7LvX0pi699CbXFSCuz4cvjMAwMn
qEYo/ATwnpDkfjRINYxaBpvNplI132gOpGT6jC6t6rAuqUG8zsv3BooSMQ4FTCx2trklVtIhz1pL
8Zm8Pxgdk4WbxHOkYTkOUlUlvEUsvZ+idjJG6tMyRLmvr3O0Q6Nqm8cY+LatyxVWIHW9+cF8lRW7
qQQK8+yqheeuJKcdnhVID3aVmCD7ec6y50+wns5Imw2DeHAZz8JFyCAfIrWIYxDh0i4Yeglzxhoe
2OfBTcinVK0A6YQUCGDRxxPX7oJIrplwo/MUO/T7idMAWdYmAwyZePlcy+wIMpp2GLOvF8tox412
3dyfnBAhAiVTkFnUMoZbB/lTczssrzOhtHjcTWZNXie9AZhnbz8qrOA+9i8i108A4UUSytT3NPt1
kCrhBoHkR6O2YZIkhYQJhpTAmQwJxZLI8b6MLqiHhqhclnekSRtjfEN0t2MLFVRNZ6AI7NJfQfOU
wffcKCbuKOZptc8TPtLTt3N0IG4B5G9oXhewB9+eoJZcuh0B5g70ah5vKdG6T5z9sRqye3CLW+99
mpWFqrkB+719mXKKDiv9WDLa0RyAM338HhANIFB3zbhFkMGyQRIDLdwr+iT/URqKGYEigA39Zz0p
EdyYhasBRJamctENOaEd8Euoi8NtA5rb/FtQ96FaWoeVd+myf5eM6grI/atkmaMoCIT2nV0a0Zkf
el6dqSHJ4cetGGs5Uel/l6LGcDfOninJss7sse25ij/HTZtVQq5Tg3X62N5rrfaSgPMEPDgrtKm/
nPOYOXRUCjn+QKwkqVGi18pHjjsQHfI35tjDtsqWKWB3ntU4Fg/dFSERgup9nSwaa610i9UPnZSI
BMvFGFwxLUBevgpwIKK89Crf9wXsde+ilOt0kvBUyi5Twve631ZDMCGHwCJgdf1zKHLJxBEjx3sV
Cw2efTIs6j64p4GO7DmmiEYvMsE7NZXblxsXh/N+5UdvRCINCKsqr1rP2je5YZrUmCTb1VAyM2lk
j/IBjs83b5C2t0YyZFCL0eH9Mp3keA3HDqFoPVSZd5lhGdTkXSaE4fipckASFFoTI5n3v2P3t0aY
tK5k94/mH1lIKkjjhyw3HfEihWwaD7NB4zI+ydqdYAuavsqcrf4rH7y2N21dcuvPomFmOCdksHWa
KixxB/03XpoAsaJNGgNApvgeQ0XWNV4AZZDO7btovc/8o13E2YMVvIHh/HQO/+ICyqlu2A4OgCq5
LaGDoUkQ9Ce8Kt+I9LPs/dSC/hdyn0BXcAqXEEVP3O7CAECPSd7eL9HPkEPNUHHipHF66YY/0ONz
f0wtgcQwsudAHueMm6AFKjnS0ZdbzgXIOZnUsJCP+IiNt4cs5cxBkLGFIXw6CgQFdFX5sPiTOb2X
lUuGhe17zmHWMmxQtxCk80P7cQftV78HA3sJr9M14EaG6Auy2qix5DUL3pGy8OzwiheUbbDnffLa
BWgzMfs07cIZGeIb761kkNFSZznTwhCq9JPI8Fxovn/h/E2T6/PFdWofEJtJAUbOQUBQDDoGQtoa
240oueB6KiFZDe+KTgB+WgZP1rE5MauIyfv5vql5L31Np0zb0Rb1iJTn8DPl+E8bZfnSK6HkxWy6
F8qsLXjKK8ER+Spm/BSEGUbMJd0s50XRsCPCJxxoAjzcg5EP7jSfnjqSRJwQd9/DiQzd0J1+zzlM
NUMAJd2K9/9NNoWeB3dwp3YasioojyuABTCV3PZDmdzHrfafRLYfducoqYbcipmdRKN8OJJRnMvP
CyAkqgRgfqfvmixBlEZJyaGwP1c8OwQtStyxYJYkrooAtByctLY5cdI3zSaMl8ENMvDM3xQWRElR
cWkKo+AOT09yw/V68z6WgNm0j86f917XGOhbuN+T+rPBALnP279RCG1mHgQpFamRfyiNf+XRWaa5
bCPKhGGvzro/QO0RZFw8j6j8p/Zt0vvhGkW7bhgD+ChG+ogX4HkZRi4LbfvnwT1aU6GMCMqFSBbg
v4S/ndGdfM8xu5OO3th77qj0Zi/bLF0NyrXc1x/7RsVKpiqO/KVy2FpaFfsAztctlzjlxvlzocLK
UDEDtLK6B4Ff6KFBLc+1GApHpGAhHuL/nAGF54D0NoP36BIbpiIBP8g7CNRPjDYi983QQrh4vpMm
SBVgPAfOlLNQeDQnzQ2W67MXgxjeHGStE5RrwsqV1ym1xxgoKlvxds/xyAEEwfIRxr8Ss5cC1DA2
we0j26TdYnfvlYSYJzHDuNTHHaX+kOfORGuO5YneMEiq7rsRimxsgUKg/6je0w2eL/wZwqIBKkig
336pBG+dW5jrxWpcLHZjuy8B4WwygtQnZZ5wg6rz7FJcxvzrKJ9u9OWgD8emPhYubiec0FbfBdIe
LnWnpCJIb9S9n8eTP+6W+u2EvlD1fKzoCcjqG5+hO+7PG4WVSZu+m2VlNGbYtzdgduk6Me7wI4p2
bzmq01WBj3YlKVpaieUHoHcBb69tIJVXI8EEVvSz0HKHZ9O1CRKhA6fthuwixGhXCaXdBxo99odC
Th5P9Wf3tnLGnXSSQ6MReFwERV7mxHp5tbsZksOnaoNTaDcLoq3mS7yqtuR+7qSkNhm9NWHE0/ho
nweg1SdTlSfioyDcw4GkDHhRtkiAeq4x14ikyWYdHRyMPvkOzvDxsa+wpUs38LQ6K3+wncXl/i6k
OYrxKbu+MWZpSHnm0kVn2CkMNK62XtDO49Ti74OBtSsapQHJVVQL1QJzbKn9/vzIyJDHa1m89xF0
jQOqiULR0geA8+d8AlvrzpCm7AvyzvvDk+Jv/hmEPF79FpxI2pTonEChP2vB77EHwDeAeg+lS0uF
HDWkZf3xd8WZEUsjCMxKh81ObLaaLMHpAM3C46NlhPmKkQJ8P3qahiY051FRkJx898g042F/qZTA
/hC9OyVL71mcyEHGV0oVMexQzBu7o/QibFYPmYCQhT+UnpH6suwkl0LSqnXPvgtGizttbN4gNusc
OIb8rHJ+Sl5bKOx2pTL/qkd47UcSEGXLpRDwc1dQjsKbcZwgne+q+rmwyVj34t9EHYrvAEsQ5s/s
rded+r8WX1UVoPTdT/XFrNiMjr7WbuGihd35lz/c96Yeo+bjXuRjN7b5gRDl/uYbWgDymtCUcrQ0
xrOiNd6NXlzMvr85ANHZCLwt1rz9eaHwIoETGJzAMXRNZL1BmVBgZwjPL0qvvSClext43b/EEju1
VoJzRduyFtYvnku4ztgFo68IiicGLCJGsRUCQOJNJ9UGLsf00nS2p9TjwPENOECQFXPV4d+Hrfle
8l1LCFtSbsx62YylQFITgCngDnO3rLnfVJpWOnHyuvDKspTsKvy8z1LlqWQvnWFcnU8LM875UJc4
VAFPv/jJCIBKG0sij2oxfPrcxJQOFOLtjJKrEq8Pj7gVgEV1A9yFnEWc4+YjJngLC3pu02kdqWti
Ef5Ctbziv0HA09rKFcAWqGVH6+Y0eeeH+JC+aNaguO3Qkc38ZWR+DOjaoOGCqbXN5QP4oFvEsMns
fPaPRtnrp1OIQRD7MLFWktfh2gSSITJP2ttb82a9qD79v0mS5T+4njqivRDGwqb97sEyAHfQM4k7
soFAAo1r1ExCXnrKppcPrF+qvylIb2wylUclwliWM3nOHi9DjdLTBbYxE+fM8U09pANt+5xfYYJQ
aM3F18YP5q5oMxvm9fpNC+0eju7K52lsVyrIoYntCm6mm9x9/3kTpLSyR6+XNlwri4y1P0iScvci
DJ8EhgvsbXgRmumYrS5LOQc0l6CN2YS8zhUQncaHHzD5h+a0a+cFmoHz6kJ32GzkyjaXT2Z7gOMT
pgLYPQbQ/kRbfQQH+kbFQnuI7U+MCa6jNwFOMunKieC2cWuwWGM9sIt07fZ3SgErKTGnP+29Oo8U
jgMiV9J4DKEz7EKyb933NVfiXUDxMicaSb8QPqrQ6xwYT8tsX0x4fcJaqaEs84KGr2wXq12XwAEY
hMyXUhQkq3Dn0h1YO03RratuEbOZa5m8oevAB2304fh2LmQZ/B+lz/OxOwIlPpp3UclEj5ndNBxs
vExFNeKSQZIq9oTHFV2XyCyqn7/v9/YsvmXLPvpGX603/ik6vYK4WM8CciCYhkvL/zWDA64GbChD
Kj70KcLnwTyWHuX++CjMft6kcCea+l67PY+mGB+XL8Hs7iFlhg+y8MBXHGxJ7653hDgkoVEXcbYZ
ofexuhqkQYd0TkGK9ddMc6RoxLhBIdvetxghx1Kz8DGwLSzl5vQk+V+cd2FDCJFEKjUjVbTz/hQp
Q0aDdlJeBW7j8lQXPjZRPUowL7MiXdCot/hSAn8oSt4VL5D7COJQg/tvEZ3qCrFMDNLzo8b9AVtN
SpTvG1HEJKf7ixCeV0Ax7FEa60fmUKLc21n4f5LJFSycileeOjwSyKnKmHskEi6g+3apyHgTseYJ
ss7+mLaWyrQvp9AK1Swopi41LRHm5iuTsL0Xa6LnjKuoaZwQWYRuJko27OpfLqzzr8ZrK+hVrGEL
RQIxg/QRnEAJZoGnDmF+pDBIw0fRu4hXFFZ1nZRn56pHclaf/rtabDL+h1TYoswWMFwHNyScEWt2
R36F4ESjYGjpuwwL379eeOsITYKhrUWLxpzT1cFrGVWBX5SiIK47Gk8uAh729W7V+7h8aq9xJbvJ
q98CkAPqLv3D3GyAXLvpJkn/9GjNVJSIgiQfao6/snHSl7xzZrF2oMashGq8+w6kCnq3UqG/Ba3k
+SqySsC0TzxzoKmA77glAD5vCAJHedwO7df/ee2AP4blYLgSPOAVBZgPhpe3ckJ27Xvu2AZ8HBSP
rv5/W8kKMryMlygHwM0N3T+Pv6KQn1fCaCukHJNURyqrXfc5pFw2590fs24VTpjE1URN96QxozmW
Ib9SG90hnqo6cS7NRdSu0VviHQk+AbYX2UCCBzug+xHjdc19tUKJF7Uhdsm5hkldNklB7XKjnvbO
y/50JNtSAdZl1wX6OsAqFiB5FJ/wWsiVBzwdLKBGi2N3B8YeDYkW31lDU1frnP/P0gAPENefsybw
VMcuGNrY2LhKHAUrsQ9BQdaw6/A6sghaUgO7x53YMgfisGAoOCReTObqzNpJPeFfz8JVT6FeRXCc
g4mgjHpEX09F2J84skXseTZxBxSKxe054ha730S9iB3Ys7PLDXmkDdikvutxDiTvBH7N7dl8bxyZ
pUjqWnpaYvEYm0BIZrrJ6NNNQNQSZZeTiI2VO3DnNkXKYwwJu8E6JBpOxTJ3l0wYCveIFBPcrl5O
vC7g2ieatVXPHlRFW2Di7f5d7KXRhtDHY/KYZXLDIvYPMrttEqMfCoSr7Sa/avZjsLb6TdwE7c8x
XKmUbkJZ/7ysnH8cSkL04GTSIdh2JczbSSiRT87ntPAmY54Kfc1lSwbJy3jPdFB/2bAi1kyTJ0iv
ZPvAsrA2f6Pe0XrH+R9oH0AFvNaVMFuO1OKd3sMmZda3Atk2q5DnpamJKanAkuPJA0ysGlfYBvrJ
SfQnBPjsOFL4xF1Y2fmHYyaqUb8ppJSESK06GcSsDUbT101/YVvKMJ04kWYKJWyJvJqudpXYJY/1
f4AgmNtm6VKSgbSHuSWHVUey2WPOa8X2si4wLtWYGJXM5DbOzeI8gacl4hYDv82fH04Nd+0iHqLm
rcYLMFzcOvZXnS3zfWtF79abVXhbfhtesuaPA6c2wATlsliXoIviCsZ90VJuHQjYh0zqhhNKvkAf
tVeSeK8yHePK3I8eDzmsM3wJXqhTyNvRIbggfeMzvjLTEiCEwEzb1jzbajXMBmC80BcnQYUGFuea
wgpiNx1XUZu0a3/EIAJiHPRKLxHk4hsqtgusScUvkhFvaOaFXtntIwdZ4YLOj2U2wjJZlzZqYanC
DwlD8g4nO/IjCXx3zklgLw1PUtm2cxi+48DoQr49dNWI3Vv/brUvDjdZg4zagUYwzp+BXKNJX/Q5
MnMIouapvWzDmM+5/d29OmsqvJ84PrMJ7m6JOO/pqyyu5UCrTfUIF6Rt8baTkyQWHM3uKP3LfYqK
nBOKjQQ0EcTBDV/9TapM9GH1Wp2TbaITTcuIII18Yet3GYZLNrQZ/vUCgdnc8POY4nZlBFkA0WoK
cNTjNYgslIUrXSNGvta77AyL978D7YcuInk80N1Ef1Pa1SDj/9UzBipmkgbHLOuSxNfF0x5y0gJs
l6W2xq1HBWMOFSEI8IOQj87guVH86apgmSH7Jb92B8x8kJEwdLTSrmXQaKsAP06SsiE2NsZyTOAb
B2j+vIwsTG+KlDpfb3QSsdH0Oltg5EB8udeUuL99jnRs1/pWki7ISIVsc5ppgQbbaPH3pORNh4bu
Vz1YgY/RTpnv0bVae9St0Si5RkD6WQJiub2brPuY8HpKTOWAvdTQMHK74xypf/dqNQF/IGEY6pqa
tu2r1DLGI4DBiDpxTShT/z0tY7kAuHGyLG9HnHS4Ikwed070hZP/6QQ4xRdMjzRKzWh/VzHwAFJY
FDOb5igGr4aHy/CZFwoLSvF+03UTc+ySoL1s80w1oSYjOIigDBDA3g0tQ7mp+L5iK6/DCN8pIEqw
5plfTbar84AU8/+qA80q9iISQLcELu6joYItTzWw1FI41VjcmGlM8s4B0sRKuoBicCwwtAIwm3WD
qzCuUW50y9ojJs68UEy7c5kOkO78IHHH/nUvobRBIhyvbsc8i/AtdkL7qsTo9CAUOpvabfOFdxo3
WD57XhB1r6pCBKj5cmnWMZZXuExtDxDBGIXb95mI8LUqT7U9VOwdzrjzxLYI+sNfY0lMzlNgCZZy
tHhHUUap3599c6a3smFAYT7KpcujRQYB9xlbZzqzPRy14L8b89tHWIvNNvri+3yZCAClyCvD8jqU
jwz38WIqL8qf81noGxOfFvS4oMTOO7NAvbgdkTq+EyjL6iSM3oodnbZJV3Xyb6/49ivqfwgr/1YP
GDyhiuRkdlI2nUMml3KNNAW1ndT0nNaQh9WKSVOAqqZatcHisbBCWvSC72HxcUPbg+y+T0ig9aIg
BNgHqCh1W12DDJ7TnqTo/s6lW0Vzk2sBKOXZmivr+bbHgqGfifQxOGJT/t8qgyTZmtiyAoweHU1E
juxkak/VclEsO2nmza3jnNgB0r4/Ewo8EbHZgubVmeuIYD2VY7zKKSzUNBh/KE/Lbd+SyaYISxHH
u3JjrVMaOrdD1lxYPf4BThivLvgQLVGJlOd9F6MbsIr0hJ2H6gZzRI6m8EDs04aF9Jt3EOK7QNMK
tCCSgYkTJJFdkMmtLF8dHeSj/Yapk2stI5FzLkcPZ/lehLjmpI+iCMYzeWbyuACjzUEXei33BEN0
tU0SRCK8akOjJNDGQCXWT3RqLqAu7qJYMtUS3Jz2+vVOxnFXQOeFHQWPpI4wYUn2xrHAU/AzsmfW
yknfsYUH1j/N4Fl/khRhzw4LotZ2Df8D5vX7MAi74zqGPizcQIpYEtsudeVcf3a0aXn4nahZFWvh
RKHMIW4UvgX55+TifL+P+uemEl2b24kxOhdLydaRfldq4ZqoORjzxtYNutYGD7vSEBDhUFK5vYpS
gh7KV+5qI/LUzB1cBJ3E3HTB/o3l1IkOzpq0pfSoriGs99LzzY/b/4Ezbzu9Eihz2dfwpHhFGIx8
X2g1VZG7WdbU4qH3XNdufoZcfynLE5kr27DkEznEt8FFGet9a43FCadiWaUw8RxGQd/NoWWzxhXI
bA1YfLogYkjsp3qOWHyj7boCG/5CUqFZMl/AbMtePi7zZFpaEsxYhyGHJnSmJnh31AnjL1SvXgq/
oEWFlGV7nbQukHTiXnRTldtrq3eGcrKxAXsPCcGYYBTOLEF9fnN7HRVDMv11r4EWxWL5jvuwF5al
IiRWjOxuVAczHdI31Rnu2rebkNNfCZXO2WC8HI7mN03spPVAoUepER1lDWVHfZC1x20j8/+NzIa+
Fdpv9HOEF90oAGbwHF+q1ZQKlks3PBHlE9tPJw6nN7pGmkM8RrayydFBNBMslcUc1K6dcvqAkeVN
7I0DdtIwsoIzrlFxhAzHWKLpKViYsCY2BB12KdtFDJK7okIfdQlqLHBmaGNBnFjBNfD9siirajTB
Zik9eKsVMbOlPSt31fLb3nGiFoJsBvvGfNnlQ6reAX6Cj/u1FArX8o0ZAbehySCtlvXASdW0cLZT
ZZh+MW3jkqNiIEpFdwTQ2g+/8wjjNaPssadsVUXLGCxfTFxmb4gcQNn/XEOeGLZ0V0jn0KVi3zar
u7Dd7ldY6kXTNir1Oad53g0UerVb7xcaRjgJx+soE0+yQWVHmjZXf0QX80+PeGGCqkEYso73QFqI
XC1LRHMtEP/O+h1naJplJ5GzH2v5zqEPTfEg6Q1AzCnST16Fog5tINQnT31fLCjOz7fWRi0tT0aG
ywkfa0d/cmHQ9xkHoBq2un6z3iZHikrXSjsgmbdWtvjTE7TYn1guimiJv6iTL3ix1SXZZw2Lzqun
Rgn7G1kY+EjbxOC7hr6/gGj/f0Tq0PuIvNt/RsAlCAHOfsrEga6cyDIC5m1eljEKZNlxh9hzs3p5
k7kyklRE7pClB1StQgqWfP1oY9Fu8YAhb5Fa3LvwI6xDGVlV+AqMeRtHsSn6rFKl4Y7iu0HWn/4p
TYRpE/YwPPgNurwV6YpFg2DPwAdhHyW4o3W8l1/oHA/4DfsWVhgjtLisEpSvbivj5nP9UcIdwKQj
8atyTTUHWPM9zt449zNVcUgzebjPAan1wro1sWwwWRzSKwq2fS6SJkZ8sbofpJRGAKLlAIKDFa96
RL4Jqg+UOnsE48E1vDTM1AoANnXajVd9K47NfPVC8bIKHl3UbSWH04vAVVqTDW7XW992lyCtucMH
Ehrg0fn2xET/PD5dwcjK+hLxUESEaZCWNulkqc7cOoVn6Z81wOAT+qiv9INjKRT50aBv/9eomUBs
iY6Zf5+wpjQ/nFwx6t16ke59Ckge/1DQTRef6yc8VqLzo1PIYMPplhvIguzOGXyFc2OePs3qps5h
DFVV6HSKQ783RYvji2ZJR17iuGH57i69u8sKqs92Y13TPhvaEGUyimScurRhL/S0b06ObX5Auurb
mfmxPmM/w3bQ3NFAZEHZVtTDu1tBjQQvl/TR018hAZb3Oh1iyOJ40ipsKTqaUOXP8AZQR4jWQIdR
e1/fCX6PM6XeOrfJaVC7MCKWsPMgdg2yiCq9/QnLIc5QeIU824cxLi5SjMVTEkk5ZO3Knn3IRRxe
jBJ9g4fqzN7fodCq4MSz92k248fiFMvHkK6S5mmOvg6Aiio5zQQmklhMZCEdgASlXVZDECWonEGQ
6Xjhkm8HGcpCwU3n3xsQFX27YahQQ4nxjvjMpe10nONALqH7twCEhTI1sVnV7ai/M2QVz4+2D/IU
WTcm/GIdj6qmIrxwDeeJaHz1Alt970z9VRTmh8imzZcE3GGuHx7tQbk1xtfs4us6IraGplMGTzs8
FMAYMAr7Q514hScTZs8PjBuINroYMQn1SczsZ2wW0NWLPPT8YMadm1xap07v48e+3IbpU4EiO9CZ
6RC3ObFUmmPESWMTHSOS+FJSAVOQQXXybRrwSMmOtstd1ngZ1d7SyyuqAhFz8UyHZ9FBW8bzcGdt
pfAY+4dkOWx8K1Jh22ioi/O1NREUfjmu7t2zz+an+ogqPL3dLmDfCNA1fKTQAP/2smiEupSLG26f
PxGq1s41Wd9e0Rl1aMBBgVKdpdGPd9zEjJoIwY5fkc9b7vNfKsv5vR/KRgZh2P+k0UkjwEgipgPX
FzOv95QEw60qSODmFg9LwSEYzL4p0GL4rPHVsmj45ZWdVlEDOZ7+12BfdN38HJaQCuEHHUqSiKLa
m8S7o8ELpBzmNwEQ1n4E4dttax6YtXNACW1JiMEOPpjXZb+sHvYkIQibHYjic9UR6o4iWauB0F8j
Bd1CTzLXDHwegTAXYWVPcpSWhbFhU7zZSxEG0PtyZoyJYG4yndNsLMIhP88GSOH3/YnzjqJSHF+y
AznO/o2eyL0+8C9x31IByXWIgQZL1xEeCKmwigABNeLQeL1Dhn1/RwaQbJmuSd+HE2GacolbWKUa
HPwyfiM44/FHntgF97rPN3NobIdgYCnVNEU62fDCy0DYx/4TsrV1mKw/kPzQMEEX0OvuK7KG0I3P
mbQe638n1Oge5Lc6XD4UgIJBRKqDHTqLZKzuOPtECKnTNgR1ym9jqt6JJpGH+0GaxfzS3R8XO72F
TmpOkXvFbMir6a3Fc9DMLT6hB5qpwRt0Bgcge54YVxmiCx0YPN4ayrMr95AHPoBGDU4QG1ycBX3L
sMWY0BGQ/yQ9kXmuDrzjzvDy24lRkV2YgP9JJEq2mPXM45azhmUZx+aOjyQJHFPEw9vyk/wK5Yks
aFI7J1ZK98jj7bg4A8pejBUJqyafHiYScjY5yPI3R7qGnR0tMZYV/eF/HDVGd0ONWzXKedutdhk6
H1aESeIDNTrYRVSRTAOqDQ+V7tLkTBXXv3QjsN/vCyugolgr3sJ05ks+t45QasKPu+bkTap5vBM6
88qyBN+s+LJdzQqD2ghoCn0IF14BTCINB0hOx6g8Z/P9HEEVmhIi6A4VZIQMqsTwNQIWWI0cRCEl
0CsRPwrl01Hbx8MVMfIPbvvBGTX0KLaL/WUq7yo41GYhmtncqh3gS05TJU44Ue3PjpC+JYcbXbCC
7SrgZWQ9CCutpOhKFWW4i3KoLpwcDkIeYKc1J1aBvK3UkWq8rwo5wKdpa7t1HTX23Z7y/zz+h9F3
5O9BH414XlvLvvfeyioode3BudIiQzL9DFyCZlo/MczO5IA0AF0KFAVy4aGJv9wNH/qiFpwAmjDk
AqmuEr6+j/xAag6nLy5gESQvWa6Y+AP033avWdOgGC7xKzOrstUEJ1EOYsJF6RV7A3WUPOaLwSRy
DW4opjaM0A0YyPEbKgHNFJ/RJ3eEZHVo9nSs/qCdqTIymYJBggfoEBvEnXgPhr24HTF37yyzI2Uw
XLT0iHmEZ7USrxkp/GvrJ8HtzIwG5mLlu3FBH/dkqvUeYz08YowA2fo5yoOHncLvbxXiEI5aEsH1
ktJUqz/Xwdz+2/bEkifGedblNXTWM/3HVwG9YBYt4TIndg1s/sipxaD+uxOYDjSxj5tjU4VXSNBu
HLmIt4apX+QR8H+ZE3uwwJufpQFIYmuuYONTNAOqt1q7rWUYQN/cW7GpTf7ZFMvyJmgHvqcix2/3
bdE5sbsZx3WricqcEP2BPvUc3PcAlvrr5W7YplCDx37VDN8sgUvTK9MSA+8bKGJr65X2/o3InS7e
Fpy03vorYWYVh7vNCR5CKMFEfiWoIxYvyQY8gNXoZsd2ntgqEHLEXbGXMgprnTpAZSraMaN0thkb
wL/CphICq5c/VEySQWJBTEmnkQl+9a6dq97CmIFnJ/hSuFlWp2KAjRnirjS6bV81ACn0z28ffdu9
2C0qJRxf1wEMoLc9dRfqtKtlMMW9mjtAZVnX0yhC/ixEMYXRp6czp5hwwhhII0KwVZwxxkAltRNV
5wUanKytGEzkDyNGSqLWaHwczFyIs8mxTogQX3Ht6PEna2bZv/J9oIPt6eueOQyo9bhezdBLJEH5
04UoaAXIzAzmEoAEOUU0/mMBxFnmqoGg2oQlIYzvNP6MFT/8vNzQIqpLWKokhhQUSP1qAVBDXIsC
D4b31CffvnqYgPk0ZHPTpOaTbKE51HUWB2ABGWTHiGN3IVv229lpVKVoNDT0H7PX22qw0wgUhTFY
mLs8slPVvfgirfw1CeHTIS/RPW+ZYnWU7r+gecivO0+9Uu1IlAsCYsPUCCdVAZAf9f5NM/2suWFS
AZqIus8wFKROij8JVbHPhcUcvIiNE1SJcfUIcVF1vKXm8HKFkOzw+uYY9NXJ+7J+HAqs/QTLgtiU
bTXhHRNbYvp4eYtPKzaCzUYl9C3FRVdfQjP2ZYZJeWVlrJTpIYqz29q7GQtDrSgcydT2xLZfiN8C
67JflUaQy3ovN25+VhiqEw/DrZFWAc0lDwRMtYWQEzifHrXarfGsnfTN8/uCGWa5TWuGQZFBHeQ8
KttbtGpdj+lrhS0RdLBI2b3DSydloJezUbY8qIdQksxJQFNFgflqNfu3PYFevRvnoc+BP7l73gh/
SHWdAbfGoVQzB55nis1sXc2tJxx05R8pQZfcHrH5wlFRaiD1mtUX8Ng2ZIHh7aGxfBV8E6osg13X
zp3acnGTcZErbfk7rpHp7NxlRIl6b0O8IU5q7hme84zuMzCpFaxGoVn32bY8YRuB59xdHt1pyMbU
XisiSgsEnaaW4gBQAFiO429nXL5yxSOsc4fjbNYCQxUorsAWRMLaxDQFXo83MQHjujwncheyoPGX
efO0i2SXkPKd2jrjfoJwd4qCp30vqG1HCRGWh9IvnmfCp0ExWRU88r+fXCNFcwTu0LXwu5JNwm3V
kUAA5jMu+rG9+ROzE38OcwETsiSXtCxtJTorQTflKGG61k6yeEPzjfPMt8sbjHmp0ks6xSzbq2xw
U5hlHY2Cp3WAd7qgHjfwDjeMDPu92x61RiEX6SMe977AD78UQxyV2RWrsDsSlRquwOX88JzgVepO
p9aZt31mXGNplm5JSVe3kNkQmhOHgtzOZfpakqNCYtyfPd+N9TgB8A4FqNg19axA8gw95QuUs3EK
0tu8NvnNydxWaR+uR1J/42XdOtONhxRY4H3ue3L6TE4QG0+FcNZUq+KzP/jQ3ciAzmqMnY87X9T2
ltHcykLO9CHp56s6KkdCenRDua9u37y+SpJK3Au8Z+017rpq8B6e4lh5ruzu6huxeY83Rs6fptlA
l7M9yfHsZ7/IUOP+3EflfhA6/I+/GvC34tyR4BOBRlSxC4mSu72Dj8F/98sJCgHAfsWCCgzxN1nR
6AAMlYXKzGepMQs4Ra49E/9jLSJ2ES9fLVcRJxSXGegc9oEW1iwMGUAyTuFNPri94KtZeJ23IxPa
maEFUMgDtksaekG3zkDJuZdrthUecTlHXquUwpYcmXA8z2J8LpEBo8p3KbhKpRjEeAsZj2DifXYA
j3dC78jgd4xLf+kh3qZTrHxX7EbeVgGNLsSqurubrhFvzH4KI1RyD8uZe+BtvxYRO9F8l2sVGZ4D
tg+mnZ4K8mP4ECyQMkWqaBpkILy5UBXxjJpYOrycPHj+SD9wK/4nPspOzxIe4Wq+C2RqJdpM0rls
AVyq5vLZZW/vHSEhz0anaWD5yRrRcBa+D1n6gXS5ByRVcEuSuEC66ghA02IU2d2ExiOKcBrFY04I
W+pQeCk9ELQbIV9DHcYlJg6tsmfMkIh/7FjGWMXdKu/qQZn9YemNo5brLdSZp3zT79za39sVCx6+
FItKsStFUZzsEr4Xra0sHKyxDFk0EvvJvMr4rji5hTYp+PU311Xlc0FmEUA2c/TySTZ+1RQ5BTsL
HMID9azc098nXehtoJ8z1Z/F1dC9xwtnQnTh5g+WHsFSUdwJB0Bq+uzH1tCuAaaHrWmpvCAKtnTh
7GEc/Aj8Y/1Y9sTHuCrh9Ui2ALycpOTWS4bs2W83zAVYGTV9WiSLbymJHjKJp/3JvP00kXBtBkLO
H/V5R8QdJdo+jK63yV/aHmh2lFQuWN6+SCrTeBJlgFzGNZgH30vc8jAHoI6vDECGNXIcVdacgeyh
0BngxD4D7A/7TyHrWExLZsPYZuVcMT1CjRKMnhHgTFVZdUEItK61MT1I+0oybJA+VnHrJC3SHkk+
7crfXPpK3Sg0cWU5IREcZtPLenA50u1krXfa4z54zKmgTwfbRZmq0IRnzaDScQw780dkMS3lbvp+
c0pMp8jlhWTS0/v1Y+MCB1mIzSQJ0lvhUlvjyFqKqERuvFtgKolMRlnxhYJs/RJsaHObmVJB1fAp
EnkfpoC5uFX2qRyU1EWFhz/odIUo9HjzeVUFKPEp52+jxrOVwayYbPgSypGzkiHphNF4EEwveOZi
Z++vXN9j9kL/9UId7PCk3YQwdsLSdUWHs0aS+SW/YhfylYaTm35K1xeuq9LRK4VkXBx/+kn/bYIl
TPsyyu8sDmVFXI2SjM20njDrnUcSQ7mF8/xPw3Mm89AFbsiiM86b9qkOELmDnDaRkiqps34IB29d
A5I5NxEg1+jN/rTR9GG1qwKVCgEJFutWph0AmDEULg85hlz6Wa+cwqD7looqM0gq5fUUqpJBiKTJ
podkwGfRFs7lR+1Zh3qpse7fXG0R3uRGaav9Yd94Dq5IycdFTHkuMivAVlbIavqIQNmecFdBHV6J
TPzUMze/mdXHXdu7xvODhQlUCIGJBF6X8BaHng6M38BsXTw8YkV6IvmkzaJ7VRxVOLz9oK8qgh++
n5H46+nkOBRQZXgJtRwXkhb84PezOiOd32F/TmcxIBp8g208hShTVokne/fgUWDeTYkgEakYBYjB
/vBu55Jd7PUufrMuaPpfy111e3tT867KP+htYoZ9U+yLW1nFbEY7bz8SEcHRSw7YzmTIE413nq6N
UYOUbg4QN0bxBQex29LZUPRc5/U1LFW6UXglzZBjoe5yzB8VLm9K3CFpTjk1uo+E96xWrcduFLZz
XUlSqddc528zULpPZBtVgCTijtTLULRBDjS4AMS6v8HoGJt00ZEo7WTmJvHYWQmGO6YlcbBFAAVk
lHSLTglL19LV0ynxOJP9KgSbLt6y1GqINrQ3zHRX4ogQwL7iFAj2QQ6oNRyExsp02hlnuZQ8+XAb
k25IJESb7FzDH6rFrtt31DCf0Cxh5n3D8l2zrM+QPI8ztJxBliuk78f7LUl+pD+h2STsQa32VWid
S5evdcwJ2reKApEAdb8HQVhSyfj8XFd6scgyY9mqyvC6xJ06DlCbCBDpifVLhBni66a5+nwQunt4
Qd68/8UTo8PKDdOQLE9MSKovhlRkZLmRfuIbtBPg4/E9ro3TOiXFAT3otoyXgjVfj6zS50toBVtu
kbRd0dTD4OCQShv6ZS+qdZRoWZalwDiSbJp0dPo2Al1rfxlCDU1EkcGEDPRp9pbTHUDKZrvnqQBH
k6Gdio3r6KC80C+CCbW4XwNocNlhtG3I5DiojP6/H3eMLXTt5BxTpgzpQBbRhh+4S1i/If3tybKb
0hJpAzKz12CC3NrdxmoVOqZ2xmdpHBWkh8CaCGo62ax1nSAtHDMlzSCL0NVPtC4QWJfy3CyzIACH
gwH+37MqDg0MzZKUYKNOX0uoWLjy7fD7qjzCd5QaJqZMF/JbzXdZQSFUFtRsh1pZiV55j3Ea5q+e
yXHX8gi29Vds8CvxyMWHspF2k+mkqP1yPYW7XFtmArcwY3FgL7F2HOYavqzipP6mmS/ULALKkYfW
EgiGrAYGHpxD4vWwGQ+TNgWvKQBQp2/v0gpqgZ+qMs/woVFl1a/EuTtGnsL2FoPJUJ2FeFOiOnio
XvvA+2Ys5lVF5SxBCf/Y7pcsfcSRdQTQbGAFySZpOBAszAj0Aoe8jwjG87bRqRoaP2sdZB3WX0SM
EbrB1kogagk10uvC6uKF/MP5yIRmoG/9BSmajNLZVawVzsnZ5trLweLpFU27f/Z6i1PcAEP57M/I
9ymYgtAi1Qu281YWUT2ziUueph+l8ymQ176wLyLZ+MClWPmU8g13bXcxdiRHCPaHpZJ0Mai1zqSN
pbbKxNKSKcI95HHwdxh1PwXFuu7POkeE5qPz0m80WnDen0/feM+mwr10o2v/9XWJATwM31CBz/ef
AukOT/3EO/EWIQ7e70PhGYL0kS5RV7ysj+j6ZsCdikJCro7Ombgf6K6Bf3njvw9gr4SnVLDRxubc
D1GbcGj3S0ISm/e09VOda0XIsKa+c94b16M30T9mXWYq8XrG7xU9KaTHZj+drGnVPLVM+M0NjbMn
eNQqHx5Cv5z+R4C6xWfgbAfnXH1JqTLvrRtSgLFbxk2AYcX88yycYKn8HUUX61dbSMt8alb1oDHo
dMaC4bzj3Ohs55UYV8NdRHNbdFGPr8/V9ZunfeJCtCrU3LsiWcOznim447574AkFXtXmnczIGmnN
vm8Av3E4Vs7q46vbSfMH+wTZtMe70eJIhViSAi7emJRzJiPox00JS19PgXxulnDONsVdZEYGJIcW
HGfeLqk5PeH8zbnlVqHCAoAujET21MW66D09nFy2W4svX9Igds52pBqAXR8F+nI3b6Vt9tiMbqA4
oAeSFh7iW8NAKbiMsoDtByRwY7WQ+VO1PZe9uaMT4ui28UxNZT9WZEe6CzYlySNLactye9PeQAF9
+G/VpyjhD8ECoE4RtxybwGlaC+SCdK+krlg7byK/2FzlmOPKPW9vKadcNKwyDy88cVwjmznujpIq
j4S4NN7pJWj7fRTI/9ouTuLJMgDokKvTGzRwLru86xzZKK3+/9n38k21fG6/dgH3bapNOjJ9LiM7
5Qd9vXYvyxb6Nd0YqwDof6fRkC2LDljJL6e0zd/kR3+QwSO9ZoMyDjlikcI5ijWFxse4EPzQaQrg
xvy66bR27wr7EMTMMNGOUncdi8Zpil4PDRYq0gE03nY+RxAQOVj5vlr0Og/iMlykJxQyk/dSyj0E
Of1nLj7VeXR9OEwzOZjP+JAEPjIqFPxgyMp5reKSxe/tEJF8mhZIB7MsERwvrBGx/vva8QxAVlRG
o6KTrXHXVuYUm8fb7lku2xhxiNVrwq779CYEsriIe4D1k01ylrKfzE9ZXf93X1R75INXGMzjl4Lj
Cqb52JfN3zIJ4wYWG7Zuc8xPRl6p4oJiNlbeMRpR0XFyQYjpqPV0L+g6nUCbVwPccrE8yBOwIkln
lPTSosYto2/IcWMZICB6RzNVPZCTGTI5sbPSz3ZHneJgQ2rHVC6DKkC8TXBqw2zcH2Gq1t9Zmwdg
6SU+CfzarOjXSQN+Lhcqzd/2wG28AFKe9xW/noN2QxXd3YtHyuxLXKpLKBCCMMuxejHGfrYMiCoK
kKGCBroEqEkfu1OJhRzB29e3tIcHCVXIb9xBIdv94AwGDZ/1adaa1S2pYv5m7JXhej5rjOm22AWp
Ieg/FNQvDA+aJDTwj6MmeBUK7KJfSJuvE1sL3ncTaQCrTVBBe5XWYJk17tW/cFGof5eiWjyVRZvf
+CNyBqUZPIwyQ1Gj3dahVMDAUVY/13B5Ql8WOY3Flugnm1ZdZZtlkW9sKRzO5nXpvaRYA4i5yZny
Zt0svO2w2/Y5FH/xVADAHNtAASp51cXtKhyWE8W6govjIojcXKzDDwefpO/PGLKTgts4sLEdQzwO
k/5+GfvtfBQsf9FszdV0kmmVXCrAj05X5gmGDr3KAvPFXiULJ1FHmW6YBAW/hOGCTz/OKvqErS75
ARSKJkKSM/66kahMONZFdLAztMLBvmvSSZBPNLl+DLvZDjb8O5B2Gz0Cu+UIMFWYZJqjI3D2M8Uv
vZF0lBPXYFmIat/6/SJxrFQpGUIeYHDE5gmrsFtuReOgF91jXr7hf7Q07YRLxit0DSOCrtz+jzsm
UNAwIavTWM4pVXMzR9cj3sk40nRd5SkL2f30h3G8UjzkGWRRzFUAcV2/4e8GZaG/YuI/DE7kMDYz
UfjXKnu3XmR/lj8Cm72k1PpUx2tM/I3AFGRtg8Q9OIGnouQUSoskmYT8FHLEyf/HhCrFMxfs9jsg
IkzrFm0MM0lELdBw531uQCUJ6Jg2465QID+X7JC18vUJluFG4m0TR7ueaHyBuOijI2rMLmuvaeyc
U+fsX72Eb/9a891yRkj7NJCp39o5ALwwqikxP5csJctMvYLmHrwBCAVMhuTawKWqPl1lqm+M3sGm
y1f6oZS+5/XbRnT8ht4tfgSjCARmp5apnCbLCt6PdcuM73x+OvRBr8c/K4fjVX5veeXAHv0Mk/eq
pYBDp4WYIOINdA3MUFSS3ym+xXW5lSkQD2YzkQawy6L1ul6QwSXa/QndhiLKXaFQP0Zkftbw9+Kd
BKmkARa6gWIqMboMwgFeepHNrtBJu2X8zMLL8h4rsxpVHsMJUmz4cp/Fq0m3pVcmMxA72JQWm02w
AGp9rfN4jIF+C4GA9IqLEHhixkhOCpwcyh4IV6yqDRItEL2YABUXuIfJKNzH6VoCmOGSwDnE7S4L
8KcMRMqfJozzERschbcJOu2DCKVZVV1DBYzbTioIMGGRkPjRreMp7TQAGDsNex8GBcfvVfWg8Ecg
S6k1MiN3oyntrxq02wjo0RutF5Ask9mGxAV1q2b1uonxd6ytPnAFf2Jr0PqlBPN9z1Hj+6wB9kCV
HvkvbIgbojwqVMnyiPwC5Ibj0cnI5oo07qnahth7G7suYBglr/IrXD7QprfCWVgRWgwGP1d/vmkU
JcGqnbc5c0UdXr/b4O2/jJsHe5bvzB2WxTzHVvD1/WXlEa2zHDxTaAM53h5fYkzlYCFhnvQSHGic
3Ko8tzYwTm6NWzw4BPEYDdoYaVYHKVzNh+pzw47R8XGlA86pTSmBTxD30vXlF4WLhfHhCEEOJJLm
AayFMae+gzyoJaegiIYOn6iFte5pdHotNoGYvL1erXM3MIlOXUnSc9H+/ShzErtknoXEpxn9kiig
t1UxzANXLufEHb6JBHGcqqW76RJSo/mOzsP5moMeFm91yYTNTQQeSg5W85qygzVLGEgE3GHtlkmc
p11FWq4SESDI8S5NPc+/DCkBtNOv+E1reYho9oPbUhuBh5YGpZ8BFpVDPsMRyjsDymiPn+OF/TRa
EDIK/He7DKxdjxcK1pFAK2QSi8D5rYLsOT4kwdFcjXkIezAsg+syMQeT9b48c778HG0QpUiCXU5q
iza2xsmUOB93mNCQRKRi1nn/uqPj24db/d63gh063ztKGYJeAAUT54v79D8yE3Gju/93w6S9wYSS
lljkg8XtwEA8Wj1u6KeHAFpL0/cGuht0HLR62IaGIGC5a9RgW/eLeDmYRN3ie5tUT4XFrInNY7i8
iY5ZEoDEpZDwrFnRdDpm9Ul10C5g52UFCxZO6H4DXkTf1d2V8Ah2XKy2vebClk4eeu5M3iqQdauN
B1ED8BOS5NYft9Y145Iy/gAfO6bkq46rJXuZ5mdwfoOVJpJdOB12QkX1vnUsBtwWBL338n0Vn5ck
meDHmVp4UkCuco+T3ZarYGjzPPKmeQcX5i/o0tzRphL5ZPTv97NGmXI7YXRg76RcoL36DFhiPPee
O64BdfDt+7uX/7pz1DHk4boVFPYCRbls8Lf+6ZkmNtvB2vA8dj+0Wkcq1h/2/I8KS0lZvfK/y6/+
XVyDTB5uU/V2mMULrgsW8gzkheMC+Iq4kf6ecCGc3lEQ0esxDTwhnkD9N/nfDJdCW0D+JEtM6ju1
d358ce1TBt1ibXdMCTfzt1MdXBBistWz3bWgRPVCdHBu/2a1ojsAtDFsDjJvBHPnEBwaLNhJKqJd
MgxyfT4ovBzoW8y5h2Hqwsj30tiubq3Jtiy9Yi3bQHA7ozM/fyymCEqJOahkHAvLYzToOChaSt64
b4DfZEV6ruCZiQ0ilYkvXb0bXtkBBll0XssC0hW3CRnYjK5Dyj2/aOR74N3RZIHKgtysJjgSNBfq
jBganF3FcR1zRjA42imAaHcvfSfLDDLBsZ5vEkCxb4G3ZT43W17VDc6odTCAUMs4foxcACBtxi+i
GAC4WQxlXqJ2HGKn8AZTID6UTyP/UGjoiLQs4PcXPOMmb5h4bIAr4fFI50SFYBxa6y44r92vVCeG
fcOdJ1czzXcHM4sz2mPKjJmrDFKYQnthWfhm2oR4/p1oOhXx82KNAnwuRD7O9jDLZR6KTyiGTm+A
0jVK+smQpm6dHv5YTrnYuPhO7LFS/guvqMNIElU1FpizAXAxUi3qnZdQ/iAgVnef8UFIvOwNdY/8
dLKB5rnzwkFh92EKEGcNpHHwr1tIFt1noBQ4k52hr/7bi5/cZGjoo3H8ZHqcZXeZSBbkaKqoA7qD
JxyKNwHvqEdfyI4Ilys0TvL3b9/LGMUsDhqIX8pmYeydKG+eaOwJRwPTJYBUbl2LlL6R4NuT1+vi
U2D86Uk2etV2aHcY2Uf8fPAVYaHtIWIrulfGj9r02iw2fmKn5igpMDKVoZRA0jRSW04UvKVD/1by
awjr7hTEAq03NnTlcB+RzsLh/ox0Y4aS2Y/1f/ZqCVOkKv2nvh7OpBWZ/ohQAqOTXReOTeQkMfpn
5Ug9myhuq/AJeXCigSRRpAZuRDXsA0uEUTrSNmbhH3cDckkGkcIB0uwJkk7d4FZK24ZZF2VJZA4/
vG3Rl/HxZThyz4fjyRqu17nPSUQ2atYNen3GtonqkzZ+XdnPL0Sw+olzImgnNQz1Ci+UTm3OUvVT
O+ZY0cAb0MoH4SCHG624CPA+s2WEEwWHCI98dGqzAjOfjRFGwes9a1q1zeomKnRVNHPHN+81O+A/
0ipBLDfbYYDP4+sYw27kk4MJwSZEVaAfvCuQZMH53ncOfH+NkB4+2Xr52B+hRPS8PaF+3QNcXMIn
HYtnqYKM6O9pPT34HY1P0v7H0+OH8GDYP1RnyEDKcvGAkBr7IV+0rc59FEpBTUjoy7LOzNLnpHiD
t9XuqNiI71dx6HFM0/ycVRNKW/ul3L1W5CXPSPMrnkXcqYJHtWnJkmu8YEZN3DwThndgIC12X4/0
aAcATHnqsZdC3I4+aszzZ1meUNDerAMiyFs/JTKzsglqfGcc9qHr0c2nhEJxpd3QisuumC21Fdix
UxtykZ9BxR6fC7dSiNkY/mNpidBSht6IRLt8Deo3RwKJcl1wLVkO/A4NI61ZW1Al/e5pt2iOInR0
GksFpIXRMEiCLpMfLNppO1l9Q5dyvMl5anPALym1KicJVCs1NMIVkfNdW4cT94/pCVvxkP4BAntO
TwTlw9yL0maIy/sCPPz2FpWffhyFOtV4E/qh+mXbP8r+L9xnpw9dUY9DhuNm98rKjp6/5Qv0O4VO
iyaSelKhoRGZxgUS+L1jWT0ySGYOdIaw5xPC24bTyeM5GaisBUjJ1L3t2wfEmyTWRf8HEUT78lS7
Uyxk5gpVTDeQbeJlF50zIhebuFporIrjq6zULP8m2je0qslXiG0vjMxdR0C+ABaw4GafnOXs5zct
ZxusZWwFfJq+o6S0gzz+66d7wUk5W1LyK4mcPbuqC/MWHSuDydXL+HXSoP/koV3f8uT6QL2AHWtZ
BCcrJQhjaFQYdG59zusw/yHvTPtRcgchGlKLU3/WBshhJDOzpf/kS4g0PZojZlHRzo9LaR+ApevB
PZlkFZYKuqLtEBGBr6NBaSCe+5U7UIFgydsLqbWFXfS0a6jQJxJL7cd/BBLMqQ9XuUZwn+px0MMc
QnfVusM4WrPeP/095eicLVUIe8vJaZcdviMi/6JU04RmmX+uaZe9UzyBpsLDZALunbqLVf201DBI
elWHtBJzBnS3MVk2okNh9yZsm5t+kx5RO8ronP8rre0iNquR3/zg86rtg+77g3Pddy1tVCOJLXOn
9Q1vtd7buB8BTXQiF4PL/Qdegv+Viut0zphqSJuStB7kIO3LXbeh0+gQcyUhQmtbFAq4Il86DaBv
OAFWFoWCF3+0b6xaIr0KJ0zH8rg2MVWnueC10CQenRHXnOvOgD37Z2pIQFnadHxE/FXl1RiDUetG
VArwCkPq9aKz5uchwKomKd2YUH0WE2Amf0zMJb91L66mJkwCQF/CBpTd7NbV15TkCZ3y9HZKxrp4
ICSkwBxN6WNRsfIhLNu7ohe1ebx8Csbd9zl3vZO/to/5QZHea5IWHnnTund+EGPOoC+Z5KcXJPMU
+AMxrfZzaAaogUgOUHnRl4Q6kMpOwdvbegVA/qd6EJhlxpCxsZLWYN9gp5vJtVZtBww/CJ7xUDQ/
cPyIt15fV01vFxP1/Z7hkd8iUyZizJdzqTwi8xhzR93KljzklZpGE39kvfS4wi4gYjp0NOkrbwVu
uOQrvIFAYqokrHV/cw8UDtTEjP21r8THJAN4/q2gMY1A+TuUW/7GOLC4UBFal1QPsD/tLdOlwDEp
ruf5PNEWMowHPg6AtPWWFHxSqowp6HnFXpLUKG5DfROh93xDlaUofGWio2KMqT5qQ2zbo6x8FXo2
ICoIhirJGxjKPZl+IAA7+ZK/vKNxI/SXczBKa96v76JKLXljQ44MWIlL3Na8fQr10C0rSubI23BX
+IZzcJ7DwtzbPzTqVF1SpVvxk8H7MPw8Roq4uo/c2s+oWgmumM9TxfPHBTzSw/Rl/QQ+VpNv9OlP
brQjWaKcloGMpw+pxKCQqzyAwR/fFZqvpmBD0zRNZcpz4nan5bq783wBFpEFTSvPP5oqOESyKsov
0IftKjdRMmf9+oxEMncmV/foEy/eO21A5IhfC7ffiuiTnrcvOWxqgMdfNEKb8Fdol9rOeQDylEQ6
fIQAqqLq2uaa6yb185MEbBCkvm3MKFBtXeVb/2vs5yuAsQMeg+yk91h7D2WgdzKiBpNgwvMjIBg4
NB78Wzb1h80yoDGxKkjE+hVnWNWUYMnKfD1qCFqpycNHm2VgECyKiMotJeVSH7+zk6ycpOv/2b6M
8mabEPsfFJ+yqHSEjnvaZPue+AdkAzaHMQDgBMktSxw8Y1mokD+s0Zjee5zMq5XlrZNpfwcPH5Sb
eGsyP+83RXJi1jVmbRVXIr6qVUf4c/rxHnD3nF9g1mlTq9XSgybe3ivTFomNryBDIBIgTGqZrJYv
Njwk9kOdW8w199zEsobZSQGlDEuFPOF6nyp7/g85NML809tM+76E0cFQj3DMqq45OQn8hOher4h2
dsMC6Q3PiuTt5QsSu+xEYLjg8iNMY4I/OnC4JTo71ERw+r3/p3pxWRZh2xjKr0wS9c6HKbLG0J4N
goOcYbZ6YR0y7dhVPmnKl6rpj6W6ooUism4TxiXmTyY2nrc05IkpZVm8PibovAcQ2YNRPo1kWjAR
JwqRF7L3eEQan2HhtlByooeNrG/fg9/D5oc7XNc9auO3DI21Axa8u5Zlpru4jM1AKwzhzUjzj9cu
FBf/A7AZxZhi0Z76ZoZgGU9/QpHiycs9U9+E9E2bJHT9soz0VM/4pi/+GTvZugusg6Rcf+bHqDdl
iIivIKvx2lA1SuP5NgdRJI5LqzqCUS/yoEAuRK4iCh+bU5o4en+rDER6gmP89VOkAIG69ZqO1KQd
b0+r8T2uqdHIw/0hhOie/DrMo2YenZhe5z3JUGa5bWExaJKYsWyfXtMhZ0hq3E4F0If0yt2PJmxI
4kJfBoONgwomLclxp4oEdjFgM9YIkd6F76d0HP26Bw3zulbHhTXpcTdwo9wOUS6/bWebWl+Xrw6y
4zwfWiiCQ8Ad5QwrR1EedrOsWyR34diR9v8905wfDljfR8J2j6v2ulXcc5BGzjtEVvxlxKFh77gN
vs6PNJA0BIlR5JehBkyTnmL4pD9NUpTL6TQP78qeLvSBMcF/km7RpWCIi9hgvpwzcXBznBaQ8UN0
J+/WiqEwfwj6VSg+K6xIwUdX4IKimg9mP63NsgPHyG0w3OrUhDCgtnU/JxvxshHWqH5yj2Q+Ta3e
9NFq/jNmZ1UU3O2UxZ89erfom9XlY+Evi//ESzXFqBbmwD8ua8sxhetA6oltiA6dsxNep18SqZhJ
3TTL9KGwtloEpTFrlE4poWdoA6mklPif0P9XfDHgJMgCVMMIz22RaD25aKoHeLP5CRlT3I7AR6AN
WTAgV9ahP9fODAm3fDQSMKYWaxMVaNUcJ3WZ9N1pi2kveHcmWvlrzTFYXDBXZ41labTIUhBUnFLo
6hisW4Fon3lFAePS1oefSj66MUQ1Kj2aoPeJmyltlaG2SpN4BdESZeo1/McdBZiHBHc3k6Hq0/af
kF69k8OK7jbcp5KtIGC37Me91CUv9ve/VNgDFZaXfxBiy0hT0iye+GAX4gDBE/iTajk6WdorckRi
/vTwIjqLIllrAnspuy0KiF9sWnL6/PSJBtaqAd7evG2nejJMith4cE74QLy0t59Dw3PQ5nzvIrGJ
JQgNUm9Q35jp/Jyu7ibizP1wKGOGa+i5YCeu0HjYy4W67/HJ4LwJgtK7H2QJvkXLx7wIsSlGVqLa
nwn5Mk5e01nDCOlf+KUpR6gYMq4yx40gPCGwvdaod2A/M+nux5RGNz9csy8mQraGtDXefvKi9u9w
YG/zzdNQHok4ydwVCLcfJaaLkqxpXJ7BwLHMVGchosyowG1TUs/SiQ7peTRIsbZHl65eFyU540Sn
a1F5jCsb1xjMdDcX/Riup1OANihcAAnEISD2KVsf6P1nuVp33Hb8V+pzaVVw4xCdUIkdx6QeKakv
MdSLHAjnSHuMRjMV/UV8+G3lVZ/3EKMwAO5ShfyUP7XC8XOQm/VMPaL2qLUIpPT62hhMV9p3r9Wb
RdNiQ5Vqkgqg6aekVPyjf1kyuMOJ31YAj+AZxAqeidlKU3fM7WCPZDz4AygHMyG7CMvVYjGLldkZ
97pjC8BvN5zfQe9Kft5cO8vLki0HcIRnIVAZoGMSH0x5YAT63AxoelMGXi4kIzetfZmD3gkqFPcG
dtKjDd6CU0jNhrgoCwe7M3rGhIxzORu7WLNh3MqLAiC3j6RD4Pngf8lgD8gj4KNh+Lev0pG9KqnW
IpyXHykgy5y9dYv78CxOzEGHskNROkFnDxq4KBWZ+xwjtYuXZahn9+pRBAXcEZiOQApv13erg8KT
xuzGLQuuKr79sb+HVIxxRDqjHRk1Kzdts0MKXYpOndCuwPDq5VTdm4V4t7GxSqrLkK8GviS0N9b4
fN5fiCISKSXygWw4gdD2iJAGZ0joa18fCiUQ+0VrHirDYsvCGd485cwVqNlOKWoAp6acz2diA4OM
6Ed42NJciJYFd1mOaM5NZIF7zQnVfDB7Mf8C9Yt9ylO7wwKhEexCSbTbhZ8/oetIV5vq8eXHILvo
+oQe6FU5YL7e06yWehmJH8Me0NIW5QSmES1MHXx7PClhMwdKFmUnknviIsGQLXqIiJshTnGC26YE
zFqnmq5EQT4JasMq1SEUwv0/pCcJAYrqY1QbhXzuoFWF094uhN0JmeuBbbkdyMPVS1jal/ODiYbD
uj3cZK+MEX1PFhJDMVksBdfdNBgADGg4FQxnkxKhxgvbDubOeEZCt/Qx7zmovlZ3UIzxqsj5v05C
9IMeectHh1fi0caphkI22mjyuKeGEr3XB2YOruW3PqkwJ8DSJLHofOs2BCllnfZU2QEWcJyv79Tu
l5prvqQv15xgrbKPYTXGtXcN1gLTLVzRM4H6JRD/5cVdGKkbLv/PyrgT6jggg3pskJNUFzRFq7Jb
hNXhZ+WZf8jrVlOohxkHVNarCFQlQ+slYIUaraX+3MoeR4kpuXiBHh7MohDbtpmzI4Z1vSmmIW6o
LvtSDDuCZlWbfH8ujA3b64iajKb0zdUBoAYP64yvoW9fFYbRCRbq0cxEb31iXh1qjZIgmtcgV6st
E6v498kELnPZlRTAva/1JL1cjBX7K9QYd1OVEqb9cvjAQYhC6Id4RX8DTFI6VydHuBP1lyr08NN8
lY5tXoApZDREwsZ8MCg4qg31cJOhIxp8ZsPjoUJp+A6SNvW3SVmciV7CDgZcVqzii0fpcFU58kpZ
qOntGkgbK1JYtYniI6diihwBnbaXc1w47xdTQGpjB3M+tFVQrAC1IwLH7RohaxRi1j3g+BIphbC9
pa5ooJnbFOpxJBsy2YeIPP6BCGGGqr90z0oCSWA5yNLc3PI3iWCEN+4n0gNS58ceu6h+H2ENRQPj
/GIXttGrbIIoWsaeCb0gvscKG2BEeMoBssmFT1OlN0sS7PbR6+kKYvA8EZekILp/hsbxSWva24zR
5QTruOoE1HagKOUDnny89coE2m17iIts/l3AePkc8P8aKUOcoCBjvu07kc9XEamZ8yqJi9pePUya
7op37+KlMoD56+Q/qMD7zmKMzabGVHJxUrT6v2nV8aveE7bSMAxw5l4Aee96LFbGeiWl87+XVxL4
l9hWXNTerC6M6rVP8K/ln0uVlQ5X4txcj+QkySL4hgK6Q0k8BM9FCcA1gtZunciHTO6hR9M7DAQy
xRJpDlnPIZANG8gfZUO/K9Usjz9+GeXzYLazQCoV49jZbdnJlTn1hcdb+id7e7pJXN0v3Uoaixpq
9bTqPiJd4JoO3fZwa6o0kd9cdulS/kd50PowjpuuAJ50HeZXnfJ+6h9rQhp66AfXk+TMgEvhY1Dd
DloEb0rSG7z6AYHjayddO3IOyT4aqR7B+cUvYbTYrEkqyLK2FpqicoBsV42d94nLJHP5T9nLPYcg
QcFe5vYIF/NVdzDFIE1rlV+RXHIPKW32rIcNvDvjuOgH45ZP8g0SYmHGOEAjnZlGmBybjYdQDwW7
mnjTWSH1eH9jg4M2Vb8Sd0YlE5CFTmtEYnzod6NLSy8An/HCSszZqiuXFdjIoFCQU/Fubw3TS2ba
xDxZPOuldX/yKyIxba8urA8qVMYfN64iFmKA7qGCrRllbtQwHLW6vvyG2GHot+7F+wySV7vIPDN+
QNcMz4fVgYhoTJVS1iiHWoK+q9y8tcj8nJaFUzL3qMYjflwyldLH2Cpa1CUZjl6j7uvIIep3Xuvh
MThldiAFfLO+rLIX7GgkLuDOYnl/24q/g5xx2q6o58Ja5oiYtmDbOkNi+N03YNAsHXZuOtmSI1WP
wvnz4wcNfSPJ1hq4VCY/VOJl9QgRDtLLY95WDXsrcuvN5CUG6M4ExuMWpesx8+LdoxqoUrYYbO5W
t76dmCMT5RQ/vfCyY799EcRKlo87X/xDZchxwj/zfvSpc7ZUVLA/KTwpBMUwkB5besq3i071GSem
Lxd5fruLpcXMgNYFI6IvNDHMFhUYHWxMxMupTk7B3WwxFVbYw9dIFekME33MqC9ZIrJtMMihHdEJ
I0zBP1R1B5In9MyfGRXTrI5M1YbVTcDhiDQ7Bo3NoTymAJZdbK3QjIw6WXFL23J8JDKPtWgk2HPN
0FAXH73jKmFkGg3zakZSPM1MRMoMInE/zwyIrm4v08PDfA+c66ehjdO4Dxhfm6RVZksZYJojbruA
1aOFnNhBktmzksIvXs3bzOVAGBF+MG0LmvowoisWRe4mBEiwSnf4HgYljzwuSh4Rz9G9H4Q7rX8C
0V87CLH+1hMTYYGEvs90gdAF+VTpZOis0DNFFmcaf95J7VznEGgUF60vg+S7mBI1W7zRSpIJJ86l
gvNe4UlbuesJEMoa5tLD9Qli/0g72Uzp7HdvLwUswcfJaAWjrqQR599FlxWTnzEx5uPQxcrcduul
+w5rLU4lKKk7/nNv/NSnXGXUlTW/vViC9UPb3nZhpRjjIGKnEPLJdLzSpWF3fi3qCL/hJhI8ODOK
qKt/s/GlCC5PXw+Xot89MrDBA1siHgJH1S+z8S8diSxcO5ZUP1K7TnxsiGn3I6yRxwzSNN9q2cX0
i7hLywjmKMLHvqx6aGhXkvpg3K0DRD4UddCyIxo8MMbkmlQ+TqzAVTv+SMluJJXadiamEGyXv7UH
Sa5s/mZgvBJL5noYcJ5EdfmrAmQwdQeo9VFxy6muiQMkKhZIbPBvJEGg5dae02DMmJ5E0If9lHc9
wX3GbK20saGOoH8jGm0TFdrQpm7ehQnP1iTOChL0XdA6i395n7RF//byu6u3ULUor32r7wsx/wEn
ez2IO2XBzCgGxZfwUPeo9iFbZgBNB37MSeMs43hKazve/ifCcbMYEU8t9UXKcrfzNoXS24Nnl8QI
Hf7zkY9mFv8JEyvRQwclGDN30KLGT0dZfC3xZfJZmRxVvO7RJuTqWetZFK2Lv1C42dgQZi+SUFLj
SQmudTjXlcnrqTWwrN5rl2wqocKHHh2uQeHV/3QFmwcz+gEvIcuy9a6psSSuhR51kOoyD1uhGb44
ZM/JnfvDVHdpsLynxPeGjedqqtVq57n5rcKbLjcNP37RV/gni5OO+drRtFkSDL2S1whOirmtXGS5
jsHQUW2hD0nzjbeJ3U+2rNtFfZlkLvWYzL3l9lfaVXKrF6+g50fsbmKoxCxmEbo5CNMNKmvnTyYZ
zCiE1w4Phj75AiOQtBaR00Ue8sKN8LcF92CJ1+4U7w4bAnHooNV3Jvz+H7SqeF0S12LiCtpHFC6l
vx4xUfBfSa0F0eTh3RPOKakFVIoJp/w2j+zYqw8dSkkqRw5Ln+dnl2B0ghbMqYY9gK62ltzyvdrF
zqeGDanIDCueW0/9+7xYZ6qLWj0kZ0mkZIkOGnCru7SqPgAhR6ez6sxu9YVXQur5v+qt/Q4CRQ4/
yEZEKCE4KrQhM28Pl7K9wUXi5Dndos9J5D1vwdd8G3sJ0PgCyYUeFuaPd6TADxEo/b1KLSvyq594
ohmPUE+Sgfkjo0xhR/h+RHwXX72QnRUQmTzcn8rIovjU2vGvEgowEhk2cgneNB65f3zALpqDQThl
fDldPjhDWn/Kcs1BXNygmneO2GRuZ1aqUqVxk4MjdnTCn0ZtHjlhQDqxHnrgoCl9AgUY2paVaOYl
gl4E3d/HiP+K+XLn3ljkp0s76y+GawV1MkBk5vsOHRbsbFZBpqGbR/auAodZqw7nGSYCvhjbWKhV
CGdiKG4o/4uTuEucKufIXleXCu0hfNpORH/SYe2XG0/7Q9OH8xVwa/LYQ9ZEhpTJsWHv2caibE7R
6TIouTrs5jkvVFGM08DI9GkJtT/WbQnlrr52+cWmqIH9xu809AlVS6JVP5HnOApVBal9qFLimiNM
xMgJ4Y5Az/DVbJr338C680fmGJcyNMdljebgRwyFN46sSrG6kaE69vtl+1y+8d1lY8gvVTviCrLa
eRHOubcwk/3mpA6rS875mUMA+Zx2AsQLEXyDI1m67WbO0TPL09hwTTTefSr5nz3JzcgOVeJ6Nxc5
4EZKXCmSpglfQB3VBlhYUXKmqYqSTamsZ/SMAyPUdG+/j4Er8N2gq/HpTCI+81A0hqto8qNIw/KD
/9QxdT0PA5eeN8yK7WXk7Dfs2fUA4UuB7Ezha8oq3czs7mmul3nCnSWx4g/vHNfhYXMgY0+3Kvpx
QG9UK3N/fNlTa8g3gDYeknYTmebsO8zMoluwByJ5FOhl7o8yoqC221sX7jc3gYePYPWrbfkMU+lz
nhOJajuHnQrk6HflNpWqV32JMpdJeZeCtEhDjjSpKbf3pDVBEaKYmplyaXHUpuqvKcSoYYgKrjwt
RsABLV5lyyL0HCtuZYOCg/gsv6yz0taaL1iJWvNXXhYygb5IahBDM8UDjO4P/ykvTFZ8gDCLPjPb
mRTEf2JDuu/l0wceIpzbuJImwGJ/oUb2j9TluVmxqS5hf28HQkOwpHbTSL+KmSkFl4YqrolgfvCA
UGGyPxa27cMuSkr7WpI7aL9pGrFMnlzhMqUhZFZdZKyWCYFRlDlXcd8yBqX6wmtJGEuIaqFvAwia
EBUSg2j7FstledvmAApwXCez1B5YAv7HP+E5s2hrSLwAumWxTDKDdOI0b8udOv8rJN1dxNA1StCt
2jK3/O4Vml7gyOgDHvbeZjCWvD5sMKXDB9L10nfDzaZNKKlFu+60J0aSXgnctGLG3op46Q9U+njW
CotdYjwDsBxx/P5IH4eiALYzdrfRWE5vrWCQkKAYZjZMPsK46G0OD7WSM65TiZA+thhnyJww3ETJ
FfkpBCeht1k2UqBPbwYb7Y33b/ostufNyGr0AiVRVq32qLVV+ZIbTlwJbceVo0hOm6awA4CxsKuR
l9kZBN8n/r4DGiHmMyiwQxS0O5K7+7dScuwDtTY9H068OR7gpPmp4uSrUSjUuLnMmQMpEqVaM7wy
Ff3nU1cNsTP3pjcGr7NQJWBxGF6OWxOSCO2rgjg9FT+5mlJUTi0xONHWHNDqIKTcEMS22eyTG4px
FcQGIUsB3XpGuq+gBu9BwqVwABSe/9rFxusJiQ6MH8klXmn+JIpmaMBzh/djApusgtxRDARHr6eK
gzeP5nO/TbbeTkGtcbDe8JQbGPaNaOtlxGk833Jsj/mZrv0aXHpXEEjMiBDEJ3P/dtX4zYG5f87F
FO7FHONXMTGUA5bAGeUzSLd+MQD97MdQH80FDvzcKOSN2Ci4j2HtOl2o6jZX0IZsfgTcAFvTo577
wN0jWyyghcdlKFtGP4gpD+k4r7nNTWZoNJAZr/N8a/9mgpvOawwMegubT4GOocO6r4mfFR4/JoBT
lhPfnEr/e1WGRY59LSBnLUDHkpHaps7I/l/13x16HI5iA0vJzksddrw/TEwxot+pvEACmLV7++8M
nJYA33fbfQUUjINTRPYkZg3K2gqjDh5UMHH+hJ7lbvzGpb5vC1MwjVCt9eHR+9s49QUCNIjv1os1
3Nr+HH/9h5kKRTpSy/7mVq+cB5SdFBMC4PlpxCRJgrpg6HCKZ7AN8R2sw3KQgDEFn/f86pnSsiD/
EQhXWL8RbkDcUgaFr/Bn4kLadsT3SdZUv2PIESw7VRChuj1qRGVsfd7r6jPZf/nqyaE6I/YApipX
A3zvEqgdNFD6YfYXy9A9GUZNPkwg8WhrVifQTZyhNFwMU67ZREE/1lGUrgxpvQKPyfU1MKx+ubEg
jcD2w3hV9b28bm2zKYnH7PsJzfhVVm+aWkBnrmplsJKG5SOi9DJP10YRP4b5eo1qya9aAfhi4zDq
kjx71tXUdoMkqTY+w+Y8IHSGCp48urTJiWYjPBKxRb1eBiH6NH2ZM12BylYrhq5uSSwtmUeX7oCt
Z9l8OcnFu+CsXXGyMfGgojKIjdp1XcaoDNfk3plxL9o48FYbSpMul2PvAyqSxXiMe9w3iBZXnU2s
C+TcmbCP8AtVs0OUG8Y8pzAGTtT2wtU0YrsBoP4wUS0yM6IZYeY6kEqJwJolAs6ruQNKIiySTE/d
qv3B3BArL3N4bZN9EA19WYvqYnpj6ba+CRZPJS/wMBPjeIv5p3G+PAguU4zQQW9jbzlin8h/Hk0K
V7NPLe2yzyW9nLbuFy8TRo9QhlvVEPkZrivWzAbfCsFC5v2TKXUYmAqvR3zRSddkgB1iIy98COWl
IrHriXB0z4jsQmFkMDNj65QgFb2CZaXbKwrgOLUFgPeYaCN5fBjElaRoMZJxg03gw/WLAdishLrr
bQF4LdrcAKSatzHHqnvjN4f0xggCduhIA2fr5MLcE5sOV4qgHNAJmx5YjP4EATn0X7AVpHdwK6Hk
3B/C88wAMCibrYXjeRfLBunhgA8q5w/4Y8RRuNCsO3dXxsrf9xjNGwXK/rLaNMZX+kbPs1CMXk6e
A1izx+fowOSaOUFrNortpb+McERp1De50pMbY9ReRwp+pprDxnJiSElAhlLLI0RxKTn1qzz5Wr9j
duVpq7EvE7nKoeFxvWR+B+QsKIADeJRBDt3LKrrJmAxkZhmkH+Y0ZaRaJE6LYhNVxYjpAEkGUnAn
vCzvhJv42Tf265G09MISULcmPlK/p47o0KrOhsGBO9aiI3toEfpzXT/AhRJ6p99E9yb1dhOHa/5i
o/uEB3jvygtgq5AyvQe8dI7Ie2Tq1VOnZUocQOHyBrMlOQUhWdU4/xAd/ZkfL7/4eh1jt55jl0pa
IhuGczfRFyRdJ0YWK3SbjSrao7wvP1YCBVrjh54NcU5s50qZFDBnxLElWxS7jyBInnu77moeg2fs
IfpLP/2g2NhIPujEdRBT8sdJ9I1MMUBIaZ5IBTttId3bB+02gIxFHcTsNlsmaI1iAChOwOcnKyvk
+uj8cJrBkf+Z6DgskgJMSGD8mmJ+1tKEYqhjyVqMNKo7Dk6LQgzUKU95+xmOfGjSBrL7occHw31g
Tl7SztRLNsMPn3MWRahKS1L/CElB2FDssEnNsYxdE84uV6fcVAbNGxONwgEdY0yW1KJYQIbkBMfV
Rh5IPH8OHUtXxP+y98ha/gpEjIHip1sAlniqXPtRmDdNMXbvh6HE8+g2orw9JkyuFPGvHQgcele+
7YnZ5P8rxguDy496Q9JMIV+pkcFL0/GAqD+1san1UdQeqQzJHLG4k1g80hweNUF6IQcd0bNV29dH
lH3pGjOqNzsvxzkLYmMseBPBVIjfIMQQ29L1gsVbJukfWZAEpKbUQhMr6FA8EPzOBS42VHCv01+z
As/43C0f9DoKhIYCsGKfvB00dJT+h9MqYtv7F518wEZkRA99xei9ZOoZByrav9Ty5er4UdpXFsZ2
246TzuPpK+tUKtEqM17YSD8fOfFTRPrQt61VIS4owgV+Se3ICJ7OndBdBuSookIBUSW0s3xGrZUj
lfM2o17HlaTEPQzFwr5BePGVbQJ10An3RWVAfu7ZfLszAkrhVTSnavMbl7TdLMAxixszedHAbvc1
IXa+H0EgGHU0vrE+2u164WsidMGfygkoXaTlKe2SnY3t9MjzexR8ImyiDvl7Ke/H276FlQ3Th89y
3LuR7EbHxAHroMScJQAYGzZJA98PB7RJ414+LHC0ToEPLOFRMaUI8zECIjUqVYCkjeZZRRvZhKjh
k3KEW1n1g4szl24p4cZoxJFNnSqtL2ELXyCJom6KvtAGJNaz1KCPI4nfNlINQs0sJjIKo8eEBGhK
K8urzxKczanICTtoZYQdkv/xC8ICJvuVLWfpxcGBceghu8+XpnZDefMjhjAtsXbYW9xwlDQ0X5mP
snW/Z1HpCKEEThlt4u4UhDcLT+bS70ukVtDm8dYx7LxO3vjpuJ3Lp+HQ1oCLNL4yh70QvixEhCzB
YQhnK6vGIMadSDMW3IgwIkTnOZIR1pnED8v8z3ozqtiad5a42dj+A7JGpQDdgpprIYIhoi+bytzc
24oPV4hxJ0EIRwGsMTmI6dvzcBsTN0Hq2r05q5xTVBHZCu4cvnqDPjR+yZsR2e6NJQ2PFPO8eI1e
VsYwNHszgnnT4mhRVe2mv5eq/1aM0wGyLrvLL31HUCikbqrZr5cN1M2IubfmlDbdrteF317hHDxF
zCfELZhH1DjSe6HqS5yMZTgsY282agh9ftSc6aOWfpV/yXFAcCvZfgOfk+E57T6l0Sn/tUMGmWzJ
pr95C8vrcj/Wsx/muOP60zY8wlqGBtiHmKbjO1DoP2Cj+QXO8kGB0sVnNZ9upMZppLoQAo/kSXhR
7pQJgY1TodqoQq8g/zHMzQJdao59dN1IBZ5u+bu0Po3hVoWTuuP5ZEyiUKI9IE82lD+/iz1oOCve
sgGqSXBgHhKPHxdKcTvi4k4E+AsWX1w4auI7TuUEhFH1N029V/lEAmCjvk1734Cc67sXs6JKgSFB
4WBBv75A3ruNX83VIA40NQa7WRWsjYdEUjXib+Ug0YTMW1IjXFRYURVitiuQ2as8Szo4k3F+XaVv
n3iD2u/hYJYvaOiw3EEN8JyRZwEky6kB2Uap7DIijkNWD8CEOx1oaTSJ1z3vsMu2BJQMTmb7Veb9
ShoSgYf38cBxfEKjDltVTqk8Qt4KtVxaVIWfi0GjNxoPL/QqQjJuV55heAz96pjWTXrJlQBx9tUz
AjufUrV/dKxw74lA34kP7MMHwoklFwMNm7u5oyH3CBlxJafe7pZOh7bm5Gy4d/lchDiSVCRo5Q2N
vfVniK3vLCJuRPDX6MQ1kIrySpEnRmyoQ1xN8hfw4bKi2ejkfZrcgZgrGg+NP0dxtSH0Na3QRiFC
v2tTNSJifdhAaToivJeOTNM3NrYxXDePziX3cavo9nAEDzek8LqHV3En6/YxBgQezdLd9kwNKAmn
3FKQ35+bXpi4SsnwTedNN3jiPh2P+XH8cNPmS+zkGVbiyMOjvlP62PQ6rJMFAaS9e1Gbjd143Ms3
HszUGSnh3UlCJ2RChD1AEBrsqcahoPjgFN0ekCO/1GCdl9soVpyS9frL5tO5N+apx2bx9i/avWHE
06e1Nc4JVzZICBOLCak7b5EL81JKOBuUtwpAR6bXTbZTaH5yRxgl2cy1u+i/HvHwBWaoe1KBd3/a
4cFOHtTyrumyyGhbAgJA0tevTJ0FFww4ECOixWZD+ZNBruEQFcurmoQ6nRyzhrnuiJY3Lut3J1oH
fPtmqOLZaxfuLC/LNeakeA+waLzRJN25JXZCXwghkrgMTnkNM1RAyrGoYSss9kXaYrlylQ1AYgPu
a7br90S5FG3B6UfIh35uziIceeZh5deuHzsYoIz1BfuCF+uljwD17G3PIaZ3tL/aw7jqzp/wq+N1
Ng7yFGUpSFzeBITmvAHGc58xVif0XlGKolbC8pDAATVWomFYLtpiJTIQ1l3+BzQBVslkiHaE+9ti
ko41zDdi6b6H0UgytvbzFM0xDqxrjVdnDXJuKaRGkVzHu4BtLHd7nVLN4mG2bP6DsK2siMLlreUb
rMnmI/L01mAgLSpN0Kd0Px9cx5Bv5T2csi1t+Nv/msQ5IjGIAZlHXzBEphkojaZz/1qafusHd0aH
W0AH2G43YasC/q8959BF7wtxTbNN+bILcCzRnWE8H/YHM8ymxVQZlPI6TVO3hzU7Dmgj/OJ3/yfO
swOUae9/5kKpAX1S6her41Osfj3Gw/Z44x+vP7sn1tGj7cSeDWbIdgxsJ3An5ojtYFKCuKzarTRZ
FxsD/9Uq1GBRodblU5KfYMqh+lPH+AOLJUtxLOHDd49/fr22z/iIsz3BxORiMY9ZyoG44U3Up4PY
WgmvAX+p0VkbWkeIaH7/BqhrDV/UMkRxttkjKATEYVHgc4m7XQOKM9DOw6CFfWvuIaBgGYSktyo3
GhbgIoggBcIycLFezn+nsl/ixJjFEmyVH0N2WOP5VRAGcgoS0tDJZZ128e1XeH4N2EJx+3NbZ4Dq
r0oevBlCMwpWy93E1rZtkeNrZQ7TccjWhXKPtUwIOgpMy9KcdNWbVGaYcJQuyfwFgl9VH6gWpiMx
AYcyDytHg4zY1jK/dfcetQvSoKi7MgyVsH5IkCRg+fkCihKGcJqSIJDQ5/j3fnKKLpnVzhDemap7
1GppeTmLUWYHN74P7zIxgs47PvRHA5X9EPFiewS8gijrlxEazffnOZ4T/wzuCiEPAsG9DEDi+W9N
MsrnofLhSWfBDfAS8Y2WGA8DSKA89vLLcjjCVerOGHB9ZW13/x6CnxSmJXYkgh9Vfh/mGNODdOEV
EUyxx6f/WQcHBHrzP/hmC1xtzUs8c3EoaznELnbbPaVxWUbYcUc2alIiE+0MmQ9oG5s+sLvmAoEg
4S9wg9G27nytcyoJxaUT4ZI+2Xtgd5dmp+oKixcrhdtqCTXwBfJVTI7Xhi7PgWkLcaaGtPkoHqEz
kOCVPOOoMtqkT7nqYZzsP/WZlWVPlZkRSM7QWZqa3rExq6CHlsNguINX1e30W9GDQA0r2qPCrUR7
pKo6F+W6kkoGxOL9uJPYMdxk9mWk5Amo0SVJzqPjPjZ2xsGREaI6EgJr5/KzVQtYOyJy+u+x9NCI
SVzkvS0ZZwDwgWKpZ1zufsfpEBqbb57aPxJfUDnTMY6mclic6GOTuMyQV836VHmEV4Ra7EpcvoUJ
QbAB18WVwS1zd5CD0gDphdqZeQQbjyemaAhb62NbzzW8hu9WWmknCp61s/aZ3Uk1WUqVmI6Z6XnP
XcQ6XOwEhhjYpPV6NjlN2hZ9Ch5u9FTPcGQ+Op0yBEp0AqN2CyKmzMrqXle4XE7uO1AQVcGn/NZz
+lEsjbKveT92FevTgcJ+I560D/vB4xEmnp6/KY10l4B1mDmCsCp6tS1yEPKAvw7eYFxJuGpPVAMd
uqfYoqZSxAGSImJSx9490jNa9D9s7x8qPvAolq9PqeYFfntdaZpI28tmybeNlwWOcLxuhXRxH+Pk
TczqcgU18dSnCu5zmXSU8M9Uvrqeg6Uu7CfoT94nlf8hgvf4aOIRcmjgvRohlqe3liov1FHX/B8l
VZpYD9oXCQ931ELIq/KOmdl738x/cMnxKzp8INp/J4+OUMLvnI1uR1yvePPr6bUWdKUltyA0Wjbz
qniincHLuXOxU7GKiF5E+ZGjg8aD4a9AjGL3QD8PgNkHBrA0nIZMpM3u6dpMfqqMZL+IGW+Hl1uZ
LrG/EBZcp0UEFQwTFwmqEY23KfQnt97Bv9vodk7IKwNDuPOwF4Tgw1KV/3gABwcDcJdA8aa0GCNc
XNUd7ynRG4uWNaNo1ois+eQg2FE6VF/W9EeqKZxRxGJb2SCB9+TPp5LfAllu6TrTMy59ZJD0htzc
gTgzHVfOzXAbB6dp8mu+q2eAUblDC0q8q5V07WjOp99X9gJtenlltPyvqCYYcEtmkflr/p2qh3N9
JwGbW1IwwBco89iZAkLuNdSYt98ulwN81h8A/XdoYwY3Svxy35FnlDqKSCzpQ2v5Q8NbGojOyBsj
+A24QIVMDmviRAKILsMSU3z5L/I+ZZh5Zxb5lRvKpfseAtbsx0o8gpA1R0XZ+Oqi98lgsRHUhERw
0q4t2dRhUAS4D43PoQXwx5kLt5PqtjaIXSP/bsHnomOQlEQezTNbS1v30cW0swl0NYph/qEaJPGl
kV/S1cDaYED9I9y7MFEhRDk4Q6EBh6sTWA0pSEQzvc3btpQLXIFSChx2GXexsNa4g9I6d/5FHCtU
H53KMrwvSEhtoj2Z6iW9xm1VLYjVvJKJfn9QSSjjDfq/lCP2BUIyf0i4MVDH6gmDXRgEmVAEgiy8
x5CWWB+qOZVIIwuriQqKAosMzOiNmA5PF4jLK1LnJEguuQhQ8f5iqtRXTEz0CUsjAfokHT7BQDVn
eomtmmoVsOuhQQ9M2jGyj37irdomT9rJHKkAFjp0rH+jmcvUXr2NYPE131PnIvoLvzUIAjUlWjkQ
6hfCoP8YN8wwx24mowAM09gySdwACK1TX5gEWGlODUR7yU45R3weGxtjjk1NF6m75X5bOs08WhpZ
ZfXRGMeVNI7lxMfE7k8Ye8scDd3sWp7nJTtl8WS3xeTiQu54aX8xTP4M4/KCUyGnskGAZl6RgXx4
X39HmTIi8FpTfDCQ+87/umRGipADN3hNUkD090Lx3nPehr4JEpah+HL7yFFvLxNIK0BSQQwBQ1OT
5/8hXBSNmbraMTE651w4GBp3QoVDawteENpyaVpRdfQavkBh5gt3Cyubz8boZ+hOPcPyBAF+W9XD
AzsRLFH3IdR3tjqU/EzKqxDpVgTbUKONlyMpnIWDv7Owm0rV+0wm+bcZjYVz877pGrayJm7diBx4
+T1PRrIIdcPut0/mBM9RbKuK8fpO/hWPrJAdua+NdpsapjGHT9kp+adaq4TEm0Q6YoAOEvHnJ8ey
sFm6hmnY1aRHgS7VRrUv1olwCtEp1pFN4yxTz/5gUPjz2mgxB7Lt+m+WwA/YK17xx+Cu6tp5Sszp
DzDPuoyz2fv9gzuym3Tr7AFm50bIrh+EMX0jma5T/GNqrDyuyJrXQNooRQXic3hFgR2TkkS9iigd
8mKA7rPY0WEm6u+kKlLcA2epcJZ7RYmLcDENo5oLbBYcpgGP/AiSEzQ7noTwbwrAgKHf04JA8Nvo
M5pBpzkr/rmr/dXqPkDPFXemvu3RRr1R6xzOx/0ODaNDpVGOYMiWiosfAZnsWLErsOiOd2brSvzj
z0xqeBrfUV00f3mCZpDEbjk38/q/o2zoHmOPllswiCyW6kvS81EDfvVmCQ7+0F54eYBC5WymaKE7
X1UscQvtWsxWhWGINtlxzNDqpZjjt3K3UlV548pdeWimQSJakhBlc9yI5XW69j5zTRD5Fsn7Ut8l
mPrOjdxELicKAuhcW5idlWRxz7P7ZabDNU8MdDeSPict20DqucVNoNPtBG+geKCBRTNLj95wXx2/
bZIJlKFuMV4YvRjrWoqdK+/YohzHS8n1HqNkw/JwxEmkTkCHzFZfjHoDNErwuoBkSO/WH2cdqcei
RzTH8PmPDRzEWiJ1Ik+JzGRKvs4EqZsYtq1KILZF+V69cjjx81+3Z8/FcsV+9THvPDIglfVRzacJ
JPGbfio7o3CheGzy1/wWKK5whCGwOnfWXsD9SEtAjQ9K05YKaRu6tZMY7AahRt5khwkXHO3SmU8+
EPzune+xuacpMg3+ACt5YodJRKe2Eg8HwKokMkKwyGIJ3IIdR1rvXTuEg62jhIT3Ae/6UjkHhWI/
ZDnSCqtCN6/sIGHB9wg3jv+L50adefaPQP6S8ya4toIa46pj1GyNmhYUbvN4l4ONKy39FfXvvYsN
/0XccRV69EdykNOlKNpJbr/SBN4Wb7tjwub6EuextrDUxc30DGJgnpiGx5XGQg6yDS4C+lKhZqN+
DztwNHh0ZrUTOUEzSmS1HlbHBgBGeIKp/3Ii36SjQegv0ny2UexlVhCZbch6u7A/WYi7d1Oy4uzG
wrP9WMO8uo5q08RjgWXj7QcusZ7O+wE6ArhIxUlJLOiNQ/Qq0E5kyaP3yxLMvYSaaBUTZ2sVjhEB
shEU9mqJFoZib6h+ORn/vGuXIl/lN1PIvckeCInOnIHnYobZfgLT1A3dABs0hl3kOCt89fXoBdl0
ODIM4W04rcI50V9WCoVSqdAYS6GZEfCKr6Kw1fKtX+ioHKLCpWm/9YobCdGd6NiSCLvcmoehztEA
K81688olAA364ZgVqwlAAI0/6KzpSVjN+zHZ7hyMTxN7CzKILw3WbuXfU2MbNFxrF7Zn3K+NFwJK
ey9SzmTHIGfM/VKRXQcVqrHa0j6KWqDhDrrjOPA2hJdJaG8CPB9IE+qSPtNhXqP0muOl3beXHhQK
WAaXkvh49HB2lMGKdiS7ERNPnvlsNjg7z6ye9QXcZ+P1iy1yogLp2LRH/Ms7+Bxl9jLePhC7uG2F
XvprLKS90oTyEc46Ob3SXoLxkpd4BT3OZhUUVhiYclgZb+/7kyO/XoPuS108Pp3+mHVYxXUXMJ0J
HqsdZihmK4tq9nAHqjOWx8ipgpJ7W8h3j5x3mxTgxQCItuRzEG+1W1/coGP9vbgIOGwI/VcAmJYK
PW2RwA/6LZfVMrF4tg/paIq2tugcBpkRg/6Uf/an1w6F08hoR3tGqSB/4pU5fMLiHUx6N57QTLR/
18DJEs7OdcSlFjMl4AU/BQdqypiyUhdaK1s/sYSH9PkGfFSKop1WGhGhwTE4N1TXn2qmDHi4M/GG
mcm2GxenxawN3GBhFZNL9PBPPuRTgs1KI1JkOOfTWbmGbEhUj/BTWHI+WVB07IJ/dtDOwH9fOepR
u/1nhIaoQeRAzk433qALrQg2Gq7gzfycF3SBgpBH5mCB8/1GIjsFS+e2dj2M0t6Lhy7svpvnJSmh
dm+s4XiWFI9Xq89jT2JIPIT9Az0ZFhkwdi45V30VJAGzIm+BBXoO6qgXmPXIC0tAcdN9Y46JJDHD
aHnnZOoAhUR4j4NSm1dVQXlZtF+f8vxJru2wVD3o7qCTfLvLeBASuPuXd+fNy4TDZ+VIZBNmwyIP
HlsTamBHcFQF+vSQDnfqhc1dQENXXpBXkPmlE02LlUpYYGcQQHm2cYEHRh8uNxnAVAM2cuiDq8wV
xs/54BX3Zh4K5Lmi1SE8eGN+Jxj4nDTO/9w2DdB0adersmxq8rnoPXvNl+LeeG34eFsfcLOc/363
2JXJBlULpfcfd8FrvyJKP8RWryCLG2japxMkKiMrwjBaI9QLbP5DRMMB4dS/EhhcmL+GaTTT61Ek
bkngxdYWGOwFNZhwSx2bGH1xQHsJd6Bgi/HmTbtOlwvNQj6RafjL4XAt78h2fBxIsmtlDNCcPPYL
zA6tTPawjmlpLTGlXlwXw1xOTIDVmaAndDUdHa3XCFCzA9EQdJy4BVKBByjmwjiMiZC3nY0NDsYJ
yHvo05xJFGpfhlfQZTZ2tG5PtCKHuRE7qiNJGTwX1CYpXxtO8SMZgimFjyBpnwlYqIq0tp5MxJfC
ejF3NAeErj9gx4FQgW9LBVtBQrmHsZaBCRGVEb1vJLk1e3NakUIIVk18PufzkBougjv+0gTBGpNs
ODumXIvAC6rWh/O7cpNkwSFvjIXlPEKn4Ksv6TTGMNGYP4OcC3IJT4FX7DkyNsxwXfkL/mV1Mppi
usVHAEbuCS3QvcX29mkZxX+45v6SadKDnGcQMpJwLEzPtdzK6X0ZAQ7EkkrbcgaLFlAtQe8Wa2iM
7JJ+jshwQUF5AjChXDwPIkCXY8HtL7J/TnmoiXnd8Jtv0CaufMerKW5g2D2TS2l+PD/VfMOn45lC
BN8G7SwHa54gvQ6yaXkTfcm2MV7Yd28wy4jCPggouAxeM5PdmoR58A1phBTvkOLacI5h5F/tMXU1
mw4fGmr+4W/2Qbzuha4JdqyrmfsWFjSBHDMeZgVUfIIf6MGt0yJVBZva8aJXbNu98Pf6Hm7BCK+0
opYBGGbh9/RQ0m1KRl+oM5ZwFloHdX1cvAoCEH9JUzWM1c5dlYIG/4YdmULoEA5Y0pjoKQk+QaxA
dT/im+kso5gyRdve6fR0yyHL2m1pyAyNUzztyJyGF5IrIOHSTyWuDGHBQhiprq8gf9mGA+eV7ThS
ucRx7vtrF2P1f/3CM9gFszy9SryEmuv+mKUFOrxkHLbyFgeuny28EOm/U7beJS4yfD+KGTKnVbfM
dgDBtZyXhT3V29+p/4VrvVkZ8e2MOPI1Hcj8p45xoPz1VB32WE4r2cZxwF5BewaUee3MDznOUjpd
Ym8DKdSHkO1CcJEPIXGeofsBFRneE5OVCQIPoj+cgoECjndBCYOBVh9i1CRIFUN2DtfcGtTl27Vp
dfj8jjXWDdF0nxdU3K2KG80Q4gbY9k4YGDlrHlpyf4MeC5PrGeIdkRyUmU9frGWXAGSxEdjOWVgs
hroqrMFxiTEZZJBMHb1W5JAJ9/tNyMCZJfXdb+P7toojD7GCaV/3o2TlzD1jmAidoaOkJ3xAAsn6
9eFte2/J/JuxlAg6T5YEIh7qRQfu+wG+QQZQdb89HpW85X39m8mBKv68zry3YvAwiReUZXHpcdz0
xCu05mjXQJ6/sCTpzCuj51SK7W6+L74nnOb6YRVfD48rBsiYQrjgWPthmTdExHc0x9dL/J10gWXK
0DNboU5ej66PrTVxU+y69TL28GV0n6UHGQYo7Sruy49LUrfITZoI5Su7KuZLxThosMHU6u+XTftz
cSDqhmFSzmHcdQQ/9P06M1vy32rnBFyq2Mp0D4AuI3jbNpaQeuQwQsL1hCTECKxHRXksYP3EeLqx
nETiZBmROCjy/tjkyC1iO0oR/phDp1fqZ+QuCkbAcAAtdieMcRuYZl0bDfdxXW9FcXPRD7rnv9Bx
KO71rhTbXUgcL98upTWHhy2IbTm2E+xChjgM2POMywV8UBzlvLUDE34ViOQS6fpyc3vlbWlpbmE+
O9wZBOZ7guTk8wFwdqdLHt/qcBXUGlR9jczNGP6ZmCjQubwLseSBgBxRpN4ZBdwg7bKONKeYXJFl
oK5IuxT9EI7va+KsLr4XhCEYOrxxn+dkuBAGPB6ooeAQsockhMqUtgHjG1bVzrmO+R3fRG1/MrEC
VXCJACwhdZNGFni65n7nRXayokrH8EImY+KUisQEzYBHTT6qPzsyqdiGQK43VyEGwKhKWTdH88oo
IZMIjnkVSbKguw+HQtjfLj09EB/lFuiLg9aMrTMHgILahD+xG9BxLBnAvExn+NEstnETrU4OzrZ5
/IV4jdKhJ7n0NdmMHylJRHEP9LyYXEaHUlkaI/JKsaRuTtSiaPYm2/J1etfhwZgBP4DmOUxLBUuZ
JzHnt3wzkVx+HGp4GYoJxWjGHQTNSuAzT4sAs23+EKdy0Uw5Y77XFwZWZPSJPrPIkPfAFXAp0vQ0
8SzOskR9AtVRo15ubXQdIUV/CVN4PPDX19cZiKidsNpHQ7XLIM+zwK7QqHq1js0G6FVxywpvI/aq
n3+SWeQs6BbPM/Y0+Dcm9qP7DHcw8I+aWwDSDyEbveWi32CyBvMv7hVv54atiTG1Y4iFg/6rxvNO
99p1uLqIwN6IbpYmtoigZ20r7lK+/AAoP7av86Crwz8nAnuF77RMqwU7qO+wsA2JMSTVjYQlpi1v
J6MrKI/UlqrOsCc6wJ0RYLZa/nnDZlBJIOnvHqY2iOlU29rQjrwWje/pWrA47e/HuFZQk2/COO2T
nMChjdKdT/C9q31YEu8ca58HJ0iQKC2fhQmoz6Y+4fExWwaSbvsCkLZ+x3wOPn041n8vhpQuUSyt
U1KIGhFLzv+TlfW+TpX7kIlaywU6fCDPO5ESWto4+8SOkVaoS7nQcQWwxgUysAgbD6KyM2DgE5r+
AA6O2Kw9a7J7XyrCl4vfdM461GzoPOPmM6niLmZ4/n64Dz+4a83k057nXNVyckYgYXvMhSUorWuS
wJm6gtAcmRJdvdu75cmmm4S5Ac2YCGW4PkR67B58W+d8TTmlKkQFY5AWoIZKzqFID33WMuebdS38
9igpy9KyKqpnLMhv/3G+1qp+Cxa+QLWDxldUM41Y2u8Yul1EW/zGyi+JewGepWKNVgBBLJgG2VKW
uOdzhagWrroK1ZzLS4xrRJzoGOVku8YL66ncYa2xYrANRKdaZG5CtuHvGeD7rzY/4Mw/b6MkkIdI
XCjxkbMhAv1R55nTnAWOvJMsjFP6DJ8NgKvlR/qHZBaLvwqEtnAIxWj+HTVkbzx7bXBYQDH+Se1S
/lk7FkiSac1Lw4nQEpKfiVoJG9UFmoAsvJ7eGeRuwoCvPzUjuIgWJIk54LCWw8fW6UAny54/ACA9
/yAzfhi5vp7l/VqYj8PMTZ+6t0PQVV9SX90+odJY79qF580PrdsJUR9XbgBKloCmh/HXQQV9y7xH
H7XM0j0Vn/LTEWffCkN+T2PPhZ++CCCjVQ6GoELyULev0REUdi6arD8w4NOZslHWQ0+rDcQDARVc
zC1Ro7xRX58UHaape9pKUUx/eBvbcL5gqaxz5DpysB9nWplamT2GI4mqbKk/O5aAovAgrleHMEmZ
eDKWZA54jkC2ozUB9bMuJHjs1NosYS9Tk3IqpQNErXaSXWYrA0aZdX+RgV8cGB3wXTd5ACqRfqi6
OEHJa6z/MGT19jp/POteYTE2vK/QQAKLJFaVcqZ4bvqw1I19DFbkrUbB0yUMTwbnJWu7vt28vBK+
ilUKr2yhl/wwrjfrZe4bPXilgk56My6vhhvdbL9A+o8jkhEZ0iDsQzcKYG9gyi6L8uepdSamN6bd
CFROONmXH77o7XSpkuBXUefo1wxZOnJb4LMLv6Q42F4YAbMF8MwEHgA357GxcjW6aIc6R4iwfnID
ke64W47XQ/hu0BhOJRhDrrAFoOdWJEeBsiF2M2ztFKrxtywOMnSJ0apDYbX3ProI7NlVA5ASKP57
+ME0qenJ35lpzdFQiNsHNo7A+/ax7OXYgbQgRwJD6mrjbNTttL/GvZ0vTQL8809byfhsCGL73piL
MaFEj1LGpm4CDTL2CRSjhWhPHWnLJr34Cqey30fwawMzSNyelHZZg2nPQGogUPiOC1b3KD6UaBkk
7CqpQ4ZAjnM+mQ7JUQVTJhbvXL+NSb1xsVDPLI6bKCUWTdlNDl1/CvyyVNvGyaxYe63B+L7mCvdL
LniiDjW84UdUQrMDN45EY+FKVtPyZ1IMfn+iB5KDoT0t2TBVV1HqVYvYpEt06tDGfcGM6apuMyOZ
sfboe9ozMNBcMIVAsH6wMlDkK1EFeCNGxk3qmZhpFbwyqsIFbiFMD6LGWk0rGsXWYkzOJXeglLqa
hEqwRlevWvU594csSH7I5MZwDEASAb2PokPqC4A67zZ0RZjsz0deDRTyxbkRWP1Zka9suuV4KeTN
M665dxdelzPuo9VvxMgPgcnBF3pilCd9nt8BA2iw38JWhewI8yUBLEkOMVs37247P9IzTVFdckXI
6vR+RwE1UOLj5uoXRz8sdwDT9B6KBkBgRNVSNpkZtUjc9oqsDCTfbHvLIYgjuGGqn1ncQarjZcoy
Znr/F7RSHKj1gh1forklQG7lIfGTI8C5YkwufhDfXzTxdsgINaVnib0RsXrhuyZpuMLf8VTEoP2V
qn0RpLXG971q1N+HY4N5BPb2RqfUslg05ECF4HQe8O37uAYLV24vHE4S5vIKv25l22cWGllIzWCR
fl91MAUCMO5b4RXGi1vkw/3a/YHW43/KCSCasBsG9KtFfTTyvuR0kC8hpy1KhcPnRsEkfUcztARu
Tf+kqhaEf0VHScdy1xjkWslYDSDNiYAPj2JDHiEZCUczl37KW4Q0zFfntIhedrclr9vhMeC83erE
gd0G3Z9bRYAN2h/J7c/jIZDHYN9jizD/xT8jrUmaKGCwwPNybHGfFLGbu2+fnGxXgvToI5WXES3L
9Hev/w+VVGE/z+zLb4LBsq+7mZH+9Eh5Hf89bRoJlh0G0qemwaefuACbHPj+5v+jj6XXdGQWrg7w
Y4XBB5EIXFMotBZNOYiPTQTAGmiEWzjDtstoUUPQimbhXZtb2K0kDlmA3C2jG+CXAMydItnbBaJc
7UMr64+E9BZJnoxeGrvkh1nmKcUoAxlrIf1Rq4iiL3RPQ02yjipeVcmkUFFcujsGxl4V82Od59D/
Quvv5xSX2OLfcu6LHlvhIvNhiAm2TexwuX/p8q3SRV1x0cREHoVAr3VkcYaU0GOq3wieoTWxTnSa
tcwOo2MZ3NUrv/HVIRX0EO4Y5l/B4cQIOLxeytr6QX5Pyvmxb+Jrk5Tj3J7XDf8iGzIHULr5iy9i
vbWwhkkWpznM5Z72ICOcoiv354aDmiC7hNqO0U/st6nyGxTxnQvsu1mbgA7yO8hBhY4cwIZjk+mZ
Qt2pmqxDxaZtzoFNe05U59DRfUD+ob3nlvY77dO54HQaIsFv/NfxM1oGdxtADCfYf5qOEdbcaGPG
Yy8HmWrPb4u9sFSDW2lr7hvLtkCcgPNZ5v86aosaXQWcM6aTJBlvkMa+U2cwxy8V1zwLHCQUCAdw
w2ENec+Cp2n2E/wHF9bWXGHeBSOoj94kJV4L2vCX+rMYK7LlKB+cIdRVhsjxAxO397oF/6SnQoMH
+aHMGt/b9WaX9WWFwKxHk7nOpnaCT3OwG270mxt06WwDTekiNuOYH02GQdjLJTrZ8RVuBxSwBfdO
/uHM5gVJ8oHCzVh1rtHDL5Jz4W4jMLX+dk6w9wpjsRypMk7Slu0u4P6stApTjVj6MhG239SqsXkQ
RIaBi9ca5cKR+/7XcZh0sq5Q0UeQFXct3g741910iHLrL/5yAVmdpqgAHxfp9USWtuDRR12QcFyy
I6nQsZZ62Ofjzh9v9iggUfdQPTqXwyFE0qlvxNVZEhLPSYAfIcZAsxeI6v+TW07hpEpYxw172pGd
oEP91EZ/YW6GriiBe8Uq+7ok4+T3Iplvr99ntAnxxLvh0KIrV+KKnuBNqXfm1Kgrwz+6k/D02BkA
JeJeFyaKwIi4/r/3/5CbPr/FshwWEq8fpdjrPtQkEsFohFoWCVDPeQ8+dmU0ho3zM6EnTQNcG/HY
MbLFEQllOtn2uSlez4I3kMlX+VMWhpuUYwPyyhzdQsRx2FpUcHZMHxK7tFj+MGjQM+3x857aKtEN
W6+3pgRfq+itObxDMMIEOQQ0ReX7N+o3PlK4sgUhfLjETI1Q7uLr7k+mNPZIW6caejVzitCEMu2n
OrRPCC88xiX/vpBJ3ZI9EbJ2suvKGmbXK++oonuTH+TaZcOINRQNV7pGNZjGV4M2oBOarx75Az/Z
VZWhgGoJikhPtGuorMHFhhq45J3C88WVlZ9ayiV60AxP6eUiYJkCTPhL4g+G6Npj5dM7Oe1O19kS
4GUy0XLtEbYJB6DBSWf3yW4+1UCYARWuDir1zDXEcJ4CcMgveuyVx05PF/BWOPqiJ8JWuPVVURX5
KdGgA8gCYDphtHQjy7IFj75QB+lgP4Zr6OkEFMzUiIHJWXchxSvsgNiSrbv8R/B0rnBufU5S2QhT
La6VzFnU/k2IuNQ9a/BvS47aUEoin4c2i+VuK9XwLILhijIOe0q2++MB525G7BSN88KzTodSTDGd
CrIPogZ9H8h/iMCwYP2HL65AFOyedQr3yzpYLRbwAlIqwZT7qYcIyisyNh0L9INRjx66yY6r/Hu5
So94bdt34gZ5gRXbRw2x8oKDsRuPGx5rzRp4C6ucmOV1/dHK3JoPi8ufEj/Vo8h09biP9XxMLyaT
EvD3gEDtt+W8XfLP9u01ybAafry6E9ZglJmCoGsb0yVZd/DouwTm6WDCNeyE4IPS7al4wrlunrca
GEVAcmkeV1mU0ZEKzrCwxrEazKJI6CVjj+AQ0beR4vUJcFelJr8gxS8y/xeRbnJXhf0x8Z+Ya8Ny
0lFH8PqJpyfHmofkr6rcQbswTGXq6o4AFV9CtHFVxxG72fR72z3iQHHq4d81+2wNub9ankw1VlbD
YLY42xn74k2nPxTer9zIpUdEx6IvpqVNLtcfJkr8YO8Znb9xug2DdJBzYoZdORzw+FMJUMf5BInD
VhXfWrAwnLHUTgxfY1rqWlAjfxSQazzCI7gSEo2hAljX3oSQWmktw3EqVj9RGauhf2zA6SFqpG1v
vA31RnzRwbBPkamrH65O4/J7prJDljKudmhdRsIakesxOLOxe5+hWiNU8QlZvF1+jmISJwMMbgGF
9VOlKQEIuQ+ktuP89UdWIZ4RAh5xsxeAOOIEFHlHVWH856S9BteeGuT2zwTJwcqwj9YVInNx2tiq
dd6pKQppq5TZYGOrngOPvLu67Zdr4oGQ1T9wYcONLI1UodtO1Cs2366DfZaIa/qcoMjd2Cz760Bb
+wxo+UMqT6Dczy+TmquxAguEvXAUgK0mqkzwQuKqwXNO6uCYIHi8FiNIbOyY4CMt0RiRKYzBGco+
Gth1VjgEkonOqzz2Q1ELO4CBeFWnApiNmDb8YLsERHRzy/dLekw1g3qao+OVO+U3UWcUDwIeHGUG
bJ45V1nSgm5MYc2hI+fxHEbT18LjUoo/dW1fmasnBw8CtTqBZWhQy+3OiyIoFClxDVvcUFgOPWhG
0zWPhx7GA0Ct9QXtb/mWRuXmcjO4Tmi4Hrv5mtmC68dlPNUk/0owm5l8ypKnmLaJMu4ANGnysyRz
OiE5QPaHOwerNG42Rx8wJuqQbh+eYBn6NHJQJxUJLzu20DXfeDQf99W7pMMtThagN+5RIS7T6Xe3
FTl3+aCWdMGJKjFDFhYdOo6VUVy/ohIkPeejc/wyDHUYW4y2G3d3Pn4mPi74EDtple0/FYNGR7sX
nuWOrJQ2+6R80GLBokd2OAqHOwhh0voXG6lOjtCTXHCTbS9eKinCRvrM1vrFA7JASUFfkx08Nnes
4dV90EC0fqP1D1ESmEQQvoY1ijHUVE53hNCWRuoIuDRZNwa9FRGLsZpWC3VPvaqK2kKdaOr8MDe1
2lRgTirNYEYn7uLkV7VWBIIKlfCbgEaLqac7SRIrzp4vx+kkiK+lA5yQsXcmvFrEPygSA7w2gjgD
vtQ1WBSmMw0VG6IMXHOgmWZRxFdkWaMOUiJaSVVL6akK5g1SZjuOyS0klD+sNRyxyXxw55IbP1tO
p9SVAIMYLB8c6b6iTNgwfxrdVbaZMFEK/FVJZNEUrlgn4Tzz8X7/leEPKnIZc+0R42nATo6GnnC3
1TofPrjoHNrSDUTDOQ6YyHPC3p3XPhZi2MvnQPt8u3+GLyfwoTjvErwoplzPP3tC+J1rL8kMh21x
H0DfcUoXYLCKb4WYAU5jO6KZSOCHkxkjQ2sOdJccoLRpmTn7EywznJ3kkXv7LtGaQkgAGma8hPpL
u1yRf5YFniLh6eYErgfzuaXRnSNttNLZSVpBXbeeQWDOgbDpAIkp4t4bstwUvJTDAiKK4k3T6TZf
Ny3DZxwXhD4HvYNPf/+NUn2QZAAyGSH2nM1fBAEhsBazK4fNahdLNDVneWsSW74dLPVL23b9IbHJ
qZSQY2n26CLP/pYcJdPAwCl6mY++o1TpQv7eDn/S/AMkpBASWKE/Z3TuEqhK6S26Gq6A3Vji/Vbg
PXOuXl4bKmMHHlDI693U2AVYxKZSY43qHNctDBo1QuNzZohZoZaHC8qdJ/WPTFURDtLyzRHE+Fh+
s2bnb95vjqjf+BszDSEepU4IxTD7Gf4eYgtCtsGnGB3n8611hgUl1rW8dzWz/GBEcMsWi2TEDFSc
vmvCWjeueD8Z9coMPY3YZ5aGP7eTkW0JtpQk3AgI59XqvipxtcJDVboyRNnBCg+nQFllDaoZRO9q
IXLQ3RTXWmwhe83DnQjaKjMv0EFB6v+2raAKX5J3GPOWmlL8rneUR2KFCGxehBTItrcJEePvQWQz
bNY2WsSffrvqrHaJEB7EyF/RiI4GDkBeiucB+ptJ+X6rgd5cO+ChucI9BI6++2uqhsl3ITSJzeXV
7agp8Hv20FBBWDI7eI0EA5CH0nWnHJE4qxWENOStTrad2hthoeud6//yAUk/3PRWtIrKeMk57cnM
QCU7M+VGZtN7pN8amyNjyLhkEgjSIGM8hFyatdf+qWgg82te+qvRelg/cLmzlUIHGqnotvzFyWy1
6NU1tSzYElMdTfF+OBWu+NsUrAjp0RHhzEA06wc20bmfXy9MlzDGvCEwSYBbyJXptuFUA8m4CLyO
F+tXuBg+hOTdZ8tEyYR6hSK6jC6EwSciHkg95qwZhWg6iwnnEAuwmmDLORTcCqOQ1YZjL/f6m3+B
YaKwVlzpu96DV5JBmkN+IRCflM72GhxNIQ9c0MZrWoTD+ZPB2Dg3WDRMGvHqBt2gkNC/vFwO1qvv
fA8r6s2TGvvpjNayzIUWcH/I88MvGHX4IOLX4LzfeS2/2JlRjqU2q9GZ/5oITB8l+nQHbBRHG7+A
swIkH7kEp5aMcPxtyA6iZDm3VpPLKLxbxTp8sXf8lSUOwQ6V4/s93tDbAYaYhyRsMJGbreCIeULz
pv9vJOGaWFa4cYX8GeOxT7eZ1jElKGds946NqNtVH4br1yQEaCK8qgqF3brH5cGDobcodvfflGZA
MQUCfq0bQR+CqCzoAP7kxaem4dsw8qeOeZPxup0Nx0ItxsRpl+QOjo6Y2n6tDoqgbye5BQOXAI9x
zIsSsDdlaDpcQme5yjJHfgvmbbofstZnbFX7JzYVg5ISkTFeBtXbWQZYCLmL9Kyov9bKfa30ts/W
Gf62EJ+snQWhkeEO3CRT35P7vOfjrarkZuBNw0moV+17W/YlSWGIoS8WBtCanOwVXQA9PB3ipwm/
0qGnRbSGwRa5z0YdiQm4UHw5RJAl7bQrW8osi+CWJj87tJsDPzEh1oro3znhyDYOCwr0t2//RO5N
eRdE7tgcevZnKy3K2No1St+ekszB1yTdYOFNfy/3gzLonV2Ddq3iXsmsAPzusE1yJdYOISkBNH6J
L+vtKUF8WAM3gEJC6GbFd99l2q7Wyk57O1l07rHM5Ds+OaoZ8ZrzPXA2yYmEujXT0M2LcQAMBac0
XVdhp3zSIgUOd/jKWv4ThGNrpyKJl8vPJC+/ugAjKl1tYa8hd+CxsQWFY+O/Z/9kALLM6tR3bQFv
rDdYKbX/SqTjeQZTVivUAhfnfz/6WZmyiXXiwNJyMt9mvMasx1EWR/cWEiOjhZM9b9AUaRv2zVpj
qnAXOMy6y1363qzIaJP9BNyD54N4YiajxJCUwPC0w1xBO/WIOf7Q9CXgFtcalZcTtn8K0WvVvKYz
y9yj9ZZC/Fn4RcRcrZjualt5a1EaNUooI6H5LL+/aSLSISQeQUcotizXt8n+AdYt8ggcaLn61uQm
sUxB0BmUq3tzUcaTEnP8+wxwxDlkTeE/AaoZKl6Og+cxhqSROomfIBrmD9yqn6jBrHv9ECQAcI13
l63654qyEXuWOs7gfw0PnNUhb/SAntzz4KlsHcws0NC3L7aLQsrhFzn9zeBQ+kpw9B7KvZxxwwe4
xpRAdLMXYtbmJjNvDqsYA63hfCU2qCerM8chLqcq/suCxkqCcjiGzxs7kZtG0axskG3dDQve+Zsp
8Xj6Dyjx0cdg1Xx4cYNVfYIn9TM5Zt4n/ogoAeMxE6nryrs4aPx8DPTZvPZfdwguX7V9TMrPrqo8
du8MuOzcIsX+B/NpCbo58B/IclpdZMfBR22nLv2pSwrVoICrm8w36HcEbtZgWqIfc5ht5BIAIQlb
DdMgGtEvWmfjxAjYC+psJMJEuZpM+spn+J02rHKmYd09ywoE90wQRSKnFYd/qGWLALrzdtsGF0IF
MAfOJWqDkzMOL5nUsJ1dTO5SoBc4zXmax0cAly8gxJ8mZ3OE5WDqS+KO8Ss2ctN5GryaRgG5AcpL
jvRZf5fbV/p90Wf1x5skg4AxW6MFEAUTSTLP8Y/3KZSQszVBdEyGKK1BAwwfU4IZnBxAwr19Qfg3
kukGqeozhGLDVuQF8iALMjjwPuTdWJpdAbjUB1niMtCxq679CN+S7ls1ZLI6gZjyhcvqthaUPc36
CYcjqXS6Xo9aTxq3POSGRjYDXBIOQhAcZaEuUyZeNw3zcHvB4KpTTIUvAtHYIFFMrhNNY9yPvma6
5l4Tm1t+SBXYGlZdAl9J7rjv/TvvNVIU0mEi9PckyREaLt8xQ/R2i13WO4ipapOkObGVRVz5WHTW
Hv+ojjkgZon8xaEBdzaEEe4uJfakTRDyr5KYksz74AuKTuu5rrggPAHCVVOfPnKUoaOEMa29sGDy
iplVVhtNf1S+LZjhkClKDSl8q+KnBkhYXLv0iymsaCqM6TYWuk1MugMCUkgKTC15H7JEL9ium6Gt
6Lqe0Mt6Dbl2f/6tl+W+t1QFtEhMLVa1FSgpUXC3OSwRGIyLERdNWxl76Ed50ju+scGPa+KPkN/U
SuUfzlGakGgqW363mXhWwfTe49GF/shMK5la1eWWdPKmEYOInUnEBoDv31XhlDNLe0cTOXPMxdcb
e9C7c/+oEmeBab/8UEjcz8ZJLKb+XW6KbsG0C3np+HmBRujiadyU5WvvMVc2YAsNm0suKZjZcBL7
ZNreq2pyP9pAFjhl9ccfEMRoHncHgmFU6IUoGjTnFzF9R7SP6uyRN0Nfkaa37DLQbhQtixksj0b9
pXN4bf1BgLc1rVFvzQ0lRUZSCiEamMMsdwm70rXW9HmJD/eLGSvT9jBXPb/VmSAShZKf/3c0bxRS
sajQSmbOgxeif1AQXgk1srIavXXAHMrhFkJYLiKNyg5PZRY+WxNbDwn7mkNQ2LZJZjsEgqLODO2f
js2+ebMWT7ANDmZ2G5tFwln4JTm1tNGhHHleKq9UcRmZQV73V7v+AoKsJAOUdwaJmdGuB/na+nE9
L+3M5bshNNknLFdpa2S+6zA1AvtcA1L46GcCq+Tw7fd+kTEvqSGRLP3Eb/qI+gbACHbUQ39N4uOq
WJr7ywPqnMMKjlvztPcAd/ivo1TEPSAbq8DDgUZ8Hx75vtwQgxKBrN2D7NeWxa+x9MDsTxiLXG3l
t1VQwzIh365zlZ+BVpJ0km8xUFcELDSgqLMYAV78e1A6xuIvb/UxetYvX+h5JMNIrDd/Vsw3zbNW
lHC1BAbHuvZAeHmf7pHF3gAatO08YIi0M+Qa1vy/hFujS3ZI1tqsIl5brgsKGQ1q6T9A9EbNenlv
hW0cnBoVo6JjdZjIuEsR5ieA2XHw98xfHdHjPRF7qDWCpDvueEp3QuYgLbQT1upuKfWD/ptoS85f
ouBIxwLfzwmhIhb9WR89iMgGB++Tk02U7m+yfvthEh8jFN003HYv4AAgVOsgiZvGdFgpuZgFS06V
R9qnedF4fVl+j31q+ofoF4H4KPtdC2iLfDjE7oVHoeAvGMfZRw6/0mTQrM5hTFB3uZGTHY36/h/2
EnWdEoNCPPF6W08ryJrCDepaLlMySdvwhkAcuDdWjNgAuFnfqOaVtHmwYstIS+x/0moknkDjd6mk
lds6rxLEgiIIPps5P/0Dy7FPZNyg3innV2JIQ7cOaoz/QQnc0WZhCO+mvxO7XuLu70IJixxeA/h0
1jg6Ijq1dt58lYTLK40J2zj7xAt7JGbavCKsJjtRy1q+pd2ja2OlmBnBrHrK52w1iwBfDvMishNP
0krcWFztLwMdod9bnkXnjVcrAEirNSErM8A6MScT3VdTeYcX01t9xtf7XzGG1wNKRHvm9VpogheX
fUB8+rsc2vi0fAbXWFoCqbfDDpqPZdyE31cIYbD1ozO/0WesSbIirF0Vv5Y7cAKXDBGnNL4UoyTC
DxIRAeYCfA2BkknYj9zHId3nNUa+QywW0xsnxKSSy47HaI4ho/vekwfP+ph11/zlkeu9S9a18az4
3lZc/sLeEJEqwBbiU6A1anpmoVcFRpeLB+WP61NYyQBhmxkteYz3zfZT0bOsLzvPExIdTGantSKN
SdKXnujczjAMcE2xozPd2CeCzuq+3YQaJwAERSm5ub3M3Fa+5DFtTVDraS/K+R4G2Sn/5Yk59dE5
Gu8qXUp1kAB/qc7Hy5GIkwQkxxmpVOnATRDeGeeCsosqbI6cY8zpho7R3WFreXEK9WduKMAQpDoW
YTBfImwpqXc2FmGUwPI+P5mdeAtMyivRdO8zWCqA1Uis1P/qhhITBErQ6DohLgL5xOUOwykJAnc+
h5Ws2cv8cneJ7dCvov0dZUpsf+shUCBF6CF85HFtXyckS0bIgD7DAQ12uZGNjPZMoiR8yns5eicT
NZ7QKxEbz04vmaNAZKWV3lU3jw8mS+QGdACZAceR4ecYOhg2xcPVXk4Cp/oJ9/aJttTd3bG7YfLA
rPyPkEa+JUEFPzxFYtd0jZHBIzEQyeO3AnqAH57BrpQDANGt5MH5tx6ahmWKsiNlUdwGyrtQkz7V
nvqdh7FdZv5u03yPGrhnTaPkhYJMsDpw98eWslkZxhh4Qd245PiMJGPjXotpgILqrQUKbOtWaRcU
m5tRRXnu4K87j3ZZ1HnsyJEoKdNSju+X95UKDGse4vS4fjvrnBhGnmRq4RIe+4qOscGG9r+/InGv
ulJhnADj7qaM/JFnf2GM2YSEfjF/Mw9rCjvX99iZmZqPol7Tsx6V+JUM56naE6mxslAu1CDFDT6S
8DKy/blKCm7SybzXFCthAMOqb/jIZKHxYi5emaZactmMeyt3m6vjZ3RX9Vh23FvcSOwcOcrpX8tU
LNCu40WbslY3XCjxVOFW8HI2FTsy/wgsD4qph5+z6fp1q+JTy8LMiC+2q+Kw3iUjxa1UiIliH0MH
URXm6lYWSIsjwxVFlL3ZcaoUPpQCPd9Fu2shbBiEz62DpRBW4h+qZF+619Ze+xR8kVferXBvjJse
WNIUNaKUNA1Z3ZNw3uDOZjEztF1rRRUQ+oJStUZCWMUakIsbaH3Eo8MFOem1ILFbLoaEXmd70goJ
i/gJjOmp5Rwn6K0AyXTb/6kpdRJLelB1hR0hUqv0P7ifEViZENZyQn8lJVjxln75Uc8+OWo0orDe
4zh4SX2CAYSaFM5jna0cGBWKyM9xsXBZF7QS0PVZye54eSvqSoyHQehPXDvSEeUNe29HrMYwJQFr
SJeauLXb6W/jjhQ14QI4AIGycwyd/cSec3kiYQx0BlKy64crz+lWfsSUZBe6VAVJFR1R6KtSUyUT
08zdoa5FPB7Oc3OWDF1piHxz7W2M1DZQAlFQCDtNhLeoqtyGsDzZ2dhqJwkNyMYoYUP0Tc1uZEV5
4DUOyIzvVZijQ552BdQaN+/DjDrOePVWUdpiyLJ9PLwYW6FdPV9gO6aWunR4/XnqqpwH3s61Xey9
X/OgpDg5WVo2iB8hCPh724TrWpzBWtE8OffT4F+bAQmllvelq25G0uQQEQKNScmdLRLKzsksMekV
mE9dMY0pqF/zmi+BDBwAzn+oua9ZHMX91fL56DuvXsfxxYm+O0I+7IPaWTR7pr0Y8ICpiVjZrBay
c7b/qEm5vaMJwdCo5+sQViNHlL10G2wCU8o5SZpdP3OrLuoNNMZ9ez5MvzpezCyOiObOdAjLdjhV
Q6nJzc/7r8iBhfTtjahQ50GJ7Pn+czhGgjbOsKQ0K4eF1XTPjYEu7nM057ZwsYgpP0YloeeVidoN
zRj35ni3xXfAvTLCqkJCIV2yCiq2w3s5EMZVPI2qt/AR/g/Aw9R62wim0JjPQBG47PyCgXwvuXe+
Cyg1tyCB7Z7ZB0Lz4aIA1y3x/L0GJwEnhTCwRNjsUKhKhi5wXdFRt3yitPYPy5x2/J8fGuyavVx/
seoLTSlEMiBtiS3qJeNKZf7okVG/bZqjUg850Cq5lQMIpfEZhjNSeQBvils+Fv2QlT+S1ESpLUi7
Kt7N7T2JnQMbysABivnXRqOnL+HiM8yRWW5Zdyx4SEP1xulz8ybagAWVnBMVMGsWJ1LBSZCH1ibL
YfgIK2GhhWlmp9w2sCCZAkEpcTx8bslyRG0UMYLQroUa7ihgD5umeMJGKHSJnsWqFuHc2Ji0UpQ8
xA2u6ZSZJBZXNbzHFbzluwYtTINtYtHIFviggGrXPaedilnuSeOPWKK5H7aKtYBktfiVE6LM70E0
1/Ypyggw3XD41KsS+lAJnV48Ity3cg4t0Jo8D3Oxm08SkyoQOgIuSlvSXzwapjGNkNivpmQvczO8
p8YlatTWiGsaRpCd2Vaeh7BTpKwuioHJLyGMCvyR4VglwUkyUMS+aYl1TqxZc3PF3sqQxfTOakuF
kpIKlzZYTT1KyIxqtlUd/Vu3rmMS5EEp7kEnWTOFc6TspR8dXbDpAg/whw8ZS+ipWomo3pFplbQj
cGzORVxo3RvhXpBcKZ81h4EMznUdC2dYG6uBsmdQXfRdQQMxvr8aCEzAAbKcZw0783qIxFwdjpzs
mFKu2jYGTuakprczp2+PZypPdaEBSqlXMU5w6x2r+wx1pIdS+tF7oipAR6ZGotY2OopE31zxAtPY
lNVWTd6AFmB6QY+ZbxJOOECKraOTINhtoIxGJ8yW75vJDmRwzm4uRA2LS18Kl2KoAO14h9Fk4DUN
lqildC3S1u0cguyI79Tz7C17BydClGDNg2aNPq85f02yeaG1JkYQ7z0ojJMyPLeEaeNEw37imZwW
CNxHXKNhrWpCvJBGw34gNihaxMkKTSQm9JXrtcKE8IJxDTmAVuiLa9vIG43TJzbP+geUPQFiUfJF
kxE9BiRPdgIRifn4cXZG4HirbwJAqxtEdNSsSkbZZ9zZQn7XrK3XnQZ58AQODENojX3fFV7jDS5u
73zjy1imncxY85Lz8W1P0IdxYi4hacIq+y4TPAm2KqrQwhySRFyt4YTvgEpZpQR2Ri16yzmg+NiV
rTgMFzwSUh6HggANGn25eL7G/PnYxRPcie4bO71hWupea/U8/FGfX3b/jTGkatpoXEW2CIXXfYxj
+NthUXnR411pUGIo+K93QOFgb2Foa55OS/AngH8i6U8mm598tLqi3vA7PatY8YuNjzmMnjng/+Vl
RshB4bIMIiFsRfMLKVtNrKxAS73bB93uUtzB/7E+8W8O43cX98HOFIRsJSpmwa8HX6AjrTMpm8kk
VN6Miy/ASz2QSM8n/edwUXd8KDJWBiDwQ11p+PLBPx+4y4q1XB7VIu63ueYCi0xElpg9f0EqE1or
pQ1oq79hNsmaFsY9EX0ZMzisJ2/IbnzgUpVLxnR7do9ff1InsXQ4+BzniRL1B6/EgZVdfW3g9h4M
oa1YOA0C3LLUmWd8HneQhGLtqzJdPu46gbBr/BC65ariQBMRNk1d9yNH7u8r1ab46XPYcchf13Wx
nFAXqv91hwM1Atp3cTTLOxQpELDBBQ/SNbL+6HVzVkJ6OX6rxxvYMXd5ACyCvwZCuQGvp20quOF+
IuiW6eAxXhhwsCddRWTgDc45JvwIy4JM0b+roanUKJzndbgCVCUJF3usAO+nr3KsUNgnZnJxPwQq
kSG1uySL6Jz4LdICDd6QEq/VxpBZhPN5n2OtAu1tb+uHNdhFIGrIaBJWaC0vgBgHF6GOweX5AvuD
S60QntUbRbVQCkEqnxQSVlGfClDg893RNVxVdgXHjiScRK6kbDnmwmtx2QHtMBoeg4Yro/XmtlzZ
wRtQJ6us9In0G4hFg4+8OhbeZ7LOnlfHSgkUa8TSEHcYvTyVzIIViFkca2nVtbDsfF+yOzzH4oi+
WYz+NLlrvK3KTP5XlGHSXe1PMmE+tyEj5Y+wtQZBMTFYLVPy0R+mVIabNA0rIZ/b/VZ14aN1cPu/
GBm6ES9wrHoE2d8g4RKTpTHgj9Z0PjnYWVcCjKtUpYA+uzfNQsitm6HBIgH7qB5kP/xqdQhCJcKi
qCt7xs027KS722vNqT34kzohbovfT3Qgvb+AdWmT7RhXXi1GDYrsN5dfhGel0so+jOmMEgFPikVf
RCB90a2DdNfBqtBJaiCX2qAegLCdSKMOtMZ36RPfe5NybLyGaTW6c2JZx4ooNuNf9LoU4AyYr7vo
VWd6tmUi7eM4Gb5mP9vAsOzp6qO1h3ks4Ts/dxXHoaAg1Mz/rRca+gILkqdyiSPhHyke7Wruvtxd
Q832RfzH0ZkJtuVD8EDMRlcDgXFuzVG5JfbUH5jbRvuGdJsI6UWyxJ75/bRDjLq0zH+/f7/ncMw1
7y4tYE+J2op0JbsK6TXCspUVpyw+5NAKyLIhJqAs66ca/ZONZbIiIMDLvwq+HqMrmWEacquVM6P3
bJw1M1vgUOi+fLlIkqeFjMIewvCYdbMzWn/Udyw6D7/6aZ7704P9rE4poH8eGT6CYV1uVz5MpwQN
SaHJwDg6cnjM9LrZY0Frjdn9JaDuUMyxFdT5kNWESkYza0iEX2DXWmpTC5NZV531RkkDGTGc7SsA
OTc1yU6mNCIquWcYBBilaazWh1Kc7Hhvk3ZC2IyqK8CZ92XF6gJMsKtUY5Y0liuP2Y4CBVPNChxk
olTsyWgexPceGCVnwMbrq9lA5fB0s0A4oYLVC4+RCiyTxwJGh7QK4Rqxb9Q8O4qrfMQypNIq7rn6
k64X+4ldITIcvbG7dgT/uyxhL61OjI72gzpN6J17abmLqBPsDoOSMnodeQG6gQHfWDpDU7Ev/auO
7bii+BkxB5uexRIiWsZwKJChcq0d0+R+yqn5h/O31tRuA9ItpCUXQ9+niL8TIen9+ZLvlmTRQkQG
kE2fUQcoCCFC9ZiXM2UoKTg4vvZt5VfPt+ZyAvUU8LdWhHuNAmxLcCygbRb/QpCDNR6tss7vj6x3
pv73cGNH1Xbi9BBmcizHdy51vtCSRa1M+29oztrf/Pnz5/r3NiNJnp0uJIamAv+/80pJW/auBSK1
cS8jdvnxr/AYu/HnLZnoKajgJsXcxSU0N4DKGYzWV418yGMORySZqJoexMCqsodPBVifH5R7pnCX
ZJvFf8yNjNKxena37iXHWtxwN3Osgr6Chbv0PJEJ5VG+mLuCFGsrIOoVN5KnVCh0Q9sQ949FiPhe
+nAZGaZokQ+fe5qHMhdbhybgy56E6pFJn71YgFJi2D6de3AFgB2T9HD0Wp6mz/eK/PN2SRKBOg4L
cRyu+RBjzARoO0sserfztsEz8FDixYmIOutCCj+m+Egzqud1C70FlS62YIpkjwElJe3lSN7M33v5
dvzj0hZvm+war8eEBl2IYjmwvfgCUOCWID1Bv2tGvfI+ntApPVHh6NJGoJaJ/fKW10YmPYrUPTjC
QBCWV7df3QMS3q4G5PoBLkXonWB5NBbI2qNVFNw3iNBbr+Vl8sWpXmKYnl64F+JKTpBTL/iK19FY
HfMNaAeku1moAQMDB/n9AvEtEQuOFKYaYli3dVRqnty1nCsScmgPhlK1fCapV1QD1kefDgHZx9bU
iIBzl5YpvzuxsTGanNMzvDNdleIOGgWrxVlgL6w6SLG6MoVn5MkrcD+ijTI9oHKP0R/fkTa01T3u
Q+yeZAFOTG7r3f5qYqt5ov9oaxskSM3oF2KUulNsfGDyK3xlblQPw0w8W+MDuurB8ItE1NqaNqGP
FgRU9AUlXfpfTRLqEdY9YgDIIBIk0QyZNsRpO3SGfKjjZY5v/ZW9OT3X7EvngMbHi2WY/O8y2XAD
r5BIjH7gATpDnrMGb+70o43qa/NLH9ndBA+FwMArr+ZQJIx+7h1L8p8xH2TM5ZnXylrK38USWjtx
7PJEwycqV996Ny3hkx27ISdTKempeqULrnEfXjERXpxxMCzDAS+gX6YW9fr/s+09jqLWbNilO06w
EpK+FYxyF9eBxopCBSvVpvCBB5DtfqYCf8hkBtcOwf4WIfiv77F5wA0xZzJcG3ztWIBXXxN9gmh2
2upwQhFigi6mRWJW+Bh6a56UzfrKhHK+qGFpbR1e2WWTIvqDhbUdNpStepQ5rXoQyl0RdeshNo7h
zH3hSSB7KqlfP5uNjevNwNNGxq9/Pc4AeMeC6J5pp1QBeEmEtZmj4XWWJvVHf3uh2z2mh90BPFT4
mu9kviLA95iHXk2qpS8/31DVQamxm5MYQ7HuTULTkWsJblyEQGRZL2ErgD12DrfCyEAsg5PM6sur
rIod8w4n+oPBeFUHJI34h5qqj2a65nRwtE/n5G5VkY++ZkGFxGuwfQquIGAIvLXyTFoxCY6q3jp9
0uZfp2AY7+X71iM8KmGCKrvC4rBfk2S/esPqPMoHulXpyT41fc7Tqw90Y1GFHTI86A6avavts6iK
vdDDvcLKgpRmvSsv0rPt39mDmPr0e1QsI6F6UxiPKAhxtiM9jTBhEx92JS9y1JaJoJbnG/cu5ZM0
+G0Wi8UcvEg4vflStBZVDY0r6KLsNrHEJ3lVaTd2KkOwzjPxv8qCkxmpCR/QUT6shpoduhepUZTW
Zw9NC32ZJT+9Vj1m9DN3R24y7oPBy/c+VvAHcITXOhE69d1NqlIBd6uW5HUPcbb1DSXzkg+m11al
TvNHkbImphmn3nVebfIMLtWFOGaIcseUmjrins375SM4cI+hB9veI6kxyKwBkQQe7wnZi+sXWqZM
JzTiEEM4i1F6U6z6LTDwRPl/CbvKlCbYVO3fKsIuFLt/33G+Dh9qFShnlQDSZJNxKjIjJBWL/3G8
IEeMVXvHOpHY5yqDR8VA1oRbpof0qgwbCXaZEMvWJbHOzqxd/U/G3QvEyad3jXabdZuIRNb+j1hu
xpLrOrS2Qjz4RuB7cLpDQqoc/8zyzgDFovfMz5+/7wqBCCKRMKJ+TZq2/ZrrQHDonuoA+NKEfE9u
dQ5p+Bq+n6jEzz8d4B6Rd65iOGOzsc6A9eKC40PAxv7y8CYM46d7VAXW3lzQc3Ax62kq58MXYEUo
L68PrdyGdw6QGBJe61qTpuY8mTaPs7+YRy5yE1DX9eRbVXd09oPET9USa0UAghVuSYxPAzufKL0B
Ll9qzoP9AxXvRPs2+6VjAjoJ6ITRZOTbVLinBscC8XKYhMDFB4iHgHTpMu2CVTvCUsd+dgqD8bSW
pQ5KQOhrJYJKd5aiUa5DitGflrchyNnZ66xig03+T4uYbqT0afWBQzgD3yMmNmnvUG+e6AviLE+A
8qUEWF9dvnHvPD77eGmftFUeTwzWrK2d9MDZABuSlMpggkPE1+Tv0m4xBpjnBqQB0VjUvqQD7pUI
jJ/J2qpBAPl0G4hRTi2Fw3l/a80gblGsgeWmJ8Jy3Ob01AJSrE22v1GRH8zd1bGYEpvx22ZbgJWj
DKz0S3I28/FsBdBM853knxWWK605lWg7okZm+bN9Ex+2xX6koI8RMKG7kYVCCZmfsM7nGbYO4fNM
eDf4dgBSKcBtQOrfjmXhff/zuhfs4jYAVEIaaqGj4hRh/Q5sRNblyKaqG5n/jXkUdSSi7vQrhwx5
G2pvM4UyPxU3wogr8rb072T1sX0lhQw1egj5jdEsAROnM8qq8PT+Bs+Lw07w4lF7jagjzKe9Hcgr
8/7gcD2zbXsP3aSS9V32Bfw39vMrDb2OMbdZ6NUX8VNROi2pL4+tiLZK2KFWbogZ5Jhsfnx0QULM
jD5ra6IUoeqFSIrHnMo47JQS00ws5mDR5lnoVYHcuZnIN1g1Gd4Y98CJ8BD15vOxM4/mP3kgCX66
d9pJSi3IMFu5vEtSiO1uSlWnaZzxJgTIzqNFxHrtktkZ7aJprNAhtgBJo4N3DFpHYyGLjW1ggj/a
eujDP0UgGLX8tUV/7ixzKILrRIy0oh7cBqNwPVRUq7bW2xfnrgCNTdH6/RV/jgZwL38rI4ssfR1F
q4f6A+/+F2J5uWukSqC/eSwVPQGkRkyR+x4VAsPLIbAYYor+r74xr0VX9GC3akXU7W3T7FlX1A1M
TlujfzhyMEuZz6WQhISgzGsmU+5EKdSN5qKrBI7BsmFS+zykbiTuKstBAqExKm4HsqFe0eNJTfnl
D4be4+WJGvEUP20Bl1Mgr2hKDLOOicTAo1lcEcuagMWnWUoCAGkkK59CN6oTebPmQTKY1tW7SwiJ
miZvnZu9SI7QEUEyj3UcpVBnP0nWSv9d5QdimE037MYBEFnXNLZLmWkF7hR5KYSKQZHs1eqnpuna
nzVKlhAsfEfw0/4nuAtYr/fB3/1RmRt7FalzRnKW2UA64MKB8S5kV3KZtlazkgi4go8EjcD4/bck
DAJ297flvUh8cZjjRoSuwAFDEHSS/8pmI4GK+T8Ja1F6HsHfAIzzkaFc9uxTxLPhU0SS00soww2A
RfO5R0Q3C4OWOmMAl8mm7jeNrGdhpTnv8Uq8rYQ0JlYj2v3M5DxqzaMx6XSS1qQ+hx0ehocVJeMC
kKjGRyqI7qKonw18vaMb0F3mn4Alcj0t2s5A4gMe9qrXAT58F9hsPW4GM/b0V6VEWLZ/N+ymcB8m
r/xstVfylsnXlr/Dw/8WBJzkK8B12jFLuACWyBziT5uEUGsrNolz1ftnYNNVZW3HC+HAK9cx6spW
qNo4rzDfL32H435To9oreTCfyeQcfb9c/Z7iqtjEIARP/PMlWXv/YFj0NA3LbiVgoZ0NWSj5w2wU
pY0qx8HNoNVrXA/e5B0JdYxiZCElrCkdu8FH51XAOF1SRh5xAQ17JwWvVafQBkXvIVam+rT3voJp
Zjsr8qnCiGYf4IIvi5zE8YwjItIBn56MZA9x+JWIc/bH8/A4Gd9czLnsi9BUTfTwF1v6oNX1QxxE
1amscEj26vMRl4M2ECwCYVGNvNCDYj+CGZuer4xP5XV7D1StdB1Zi7YLGf3CfUHzkcheGnUw7FAS
d5oRvU9WKaluxeg24fw8Awyyv+YOjZZ1hIhJNHO3fg4aFErmIAzEjZgWRdu06Exl/kWnF+EUqZPm
QCINkX5CAFx26b7d8rOelJ0j6x/DMxWLgssfpYiaK17S70PuJ6JI/3gyT12U0B0Fsd4+1bRlqXM7
h4cmkejUjAtwwxoO8JNKyAwsnaCd2kWNNzjoCCMVAm5PWvOQtqJzSEpU9m2MYoo6PwoML+ZhBnDt
E5wz4sc8752FkSW1QmV2i2+UqAq3TrIxV9UiuZb0wUNQm9WTjeHpNftpr6NJz0i4vovP0NrPXjqB
g+ZWmHCmdBRvlYDcnU2K0GRxAmOYvfWmJcqr2lNcoPXG0XwdGwlzv+TU0dXPSgoALjeesHjeXZuJ
07RzsmwMrZEGGI5g+8b/J6d6CszkMRkLcN60Y6AHMPorXBBkNudnEA0byopU3mkpQSJTXb6I+1qz
yVFdn3hYdzRdMBzv0+vfYEllMvIVN+DzYjGPotBNImTYfjUyzItUQGgnppgk9v7rgrlI00bdMVDi
UjD778XP7HpG+7qkrJB1/thI3vyyF8RUbt02u7OpMs8mWUlga8pMuYNPQSrtKZPGPTQxhTY3gO7W
3LmH0YNv6KsZd9aVSIZphSo0NTWPfBWIPW8BVAllSQwukw61PRYJIMdYz1d+7G9nxIY+/AzmAuxV
3iCaKISVt4YcTPVrnKnanOfOBhfgL9daw1JnqTTylTe/21TCa3QGySJnbAOnSp2eRvjHUuwvurrl
wRsPUIG0ZfEiBy2cno40/Teiy83BOG9WzJ8KB/e8H7LvfcpdN9wS8XaondXXOEbH2yy4P5eraNpu
kvUPmPOG5gcGDE3fa1Uw01PvfXXpmrGXKMgA/T+mG9Q1gka21k1aEwt6v5fF+UUtm5dE0yYJDWJN
agVSlAw2RgrEzUP2JSsm0o8Ir4bud95HY0oUXEeAAP0TSoKLVDHWY9lM1qEGHc1oJSp3dgHmDcWX
/QAsiMJp39AvZT0Uhyz2Gt4gwf9kA8ASpF2FMmfYJ9ZhB1bSgzUjb0GHHLkht8whQ5OrexteHV0C
UPoAXHPb4CTmgIUyEkAM6j6MQQdnPMpacDGcBL2Aort8huNO8Amd/Fm+i0a9cC1ZUYdBKJwwyd22
yPBgsHktpbQM903PuzyLxL2Ia6jsXfNdDhMbjNTUDFpsknq9pkAi6WbROa9iKirBrz83K6gsoOuH
LjxUqxAkTpIfWf4CDYY9umVyC0Wy5PfA5yLl0dTdc0JwYszEzSOnd2zhmULa797cATHOVyrnSZN6
Qhv//EGbPrQCBI+cWffYkry6y/x/iaHSXFvyZan/HoUH4mLPWMra7nkQ2+sr4tsD97oRuTbojhpN
99qdfBpf0sw6zqwnbjvBNYR9EsI3gvnNtyi5U6iOorenFGfqOPwx2JjAsyh80ARv70IWBzH1XujY
TI5/emGCrUX5Xrf8RC70R/EK3QPwMRFIVDHju4rv02H2KGy1WylgN/ZEgeD0kvP2y4dZ3SUIHn/X
fqkMQ9izI9IMrCPQG9ASB6DMaGalGMGxXzQAm4MULLvzNLMJdOqpzGVnbQfgQxYjpzhpnEgiWxO3
ltST57um+lGf/gnY7JBzwNiZxfkTU830p8klGaPzrXiz8xXCWyY9s2UqwFmnSGiyhFOrlfMqMDJZ
tB5BwzNadCH9R4vgNPyvP2H5ujcizbGjtAFvOyKhDW2RRcIXZerg/ghaYi/dtr2iaxiohV5PqsNF
7vJG4i9L0+he1+ORL2kIe5a3Pq9iU31wZsGHgESWlFoIHI+J+zcUsGvhy5hizghYlP1fpKFrVCyP
Iy+kI3z+T6eAIx48akdsJP589QYP4Xt8boO+Z9rDcEHWVqm7ZAo37uAhE3en+iZnwSNP43euQNhk
jvc0gd9K0lNF7gI5JYjTHQogVuQsoazoua3WvqKWa6ns2/w+DPmMnoujn8qQJQkOdm3K/QV7jTyU
BAq9RNpxdpfSFkM+ANwGlhFfIp8zcfI4ZqgP1C+C/eoUEnrGUe9vB0210RxrHqLroL2zifP9oLTX
c/gtkY+7TlbiE+S59+GRgIv/C/BG/Er9U+lSXnZR3Ht6jFDDHV6rZ3wqqG44zFXXJ58Al1finhUK
8QMTVF5hN/sIzNk161aB+FoZNLEQYvlh9MkUiq6VkZRvjCb3hpOLkhacFFiTEJMMAFpb0aPskdNe
xxe7cfquyEyfH9ZAxqNwH4nxPIPsGuUaAIU5qxBtu8jQUBeiHpW7ryMtxGPjrvNX5AjaB7NcJSD0
p33+Y2VgHFUz9rGUOsUjH86xXYgxSTZtr6mD/v8Xxcmp6akmhNllsvaKAlZqHKndWoDMJcoOe9PY
r0mz++vMMxdvQJYtGMDkWd6M4YiSUJM8ZIkoB0EeqO0544E+LViFDt39CoIR1SopTeWPo0bRW5dg
NESnvy6UNcKVanDPXxZTmPYfBsfvXSXBCRv1Npy+qHjHv/OH3YzhepyK78+PmXCRiCbAFSdc1mFK
0rZ7ll6FSIe4jVdzEmhWpW4HkmhbELfPq08dvR19sY5uvpnVSmGXChsgKG0zNu4T3tjQElM4cJ9J
aJe1RH+jJwPWDei1lJyz0Y4xGfvuFjz8NwpWL1VLRvbMAYn5h2w1shlzR+NJaqHzmiIFp5uIu0DX
M+8N0ipaFbFHHyQtsIPM/zHRBFzu3dXdVOogOeYjeBD63TBNAQI4AwFe4BZXmVnkrSXCHAtliRpH
6OPwDkH3oDDpPtR4rn+uzSr1Y7ktGzaTvjHm3o3x5MZNJes7I/qFwI8bdkbLme+IjbnMz+WiSh76
RgQmJcvaqHz7vIFvYlvq1votv5ZoUf/TZl0XsYuF0dlSKYKBlPaBewpOUc462HHPQBSMZZjhdjqP
GLGfTJsbXrs0XSBmcrPIlL8bHldJu1Oi8NvtNUYWwMsghJLR1OW7KHis+Rv+HZdIhHxFm+X4m33K
w5Tfv0z7CUamuQj9X92mArLHuanKjA1X3ZAsOeEGNWePlphuSx7hIVdleXUPYmd3vs+GuxPvbkAb
u+5SN4w5PAcLhryX/0jpcFOWFrBkqs8Wu7kFptSJoinYvDHQXXKntizpUGM7F7KQwVtEHZLz4YDd
gdu2am2pwuJfxXJGvF5q3Jc4Bx5ylOlt35irssOE10Ew5fexoxPSt3pw8KMm+p5i4+Jf/LSVfu8U
49VQN0PWwqswebfOwnJbR7KcWlKHjaZDI/MRPJOC7qYlHFHrPIGoRZZMlCSyGsBMmgNQ2sO7PXNN
AcbgszBed6/lHaUBQ5+SIQ00Vj5zbweAQweiNoo8A+we8RNXD03rjG3ZYWtvnTjYY7panu4z1jat
SCVODU0nx474OTstXPeZFR0TPRrDp1KzhUFlcU7pkhpX3YGcyBosXRf18STFotzuiPWukDmU8Ve5
g8WC0TdCSLSI3NTiVYsLAtY6QwWwHR2DHRGjDdKRCCQhDuTrC4hhr2AeGRtND+SKfRk84AmK+k0R
JPVP2SnYc+9bdGffQ0C/ZhO4xdstJD+3/y9cyi4Op11RxBRMtkglT1pzFRaw3dMnbGU59opFTJ9i
INaDjcCrkguKz6ixm02akqDNJw7Bl97E+PsdtvuMhk4sKWEZ2uZ4SPAnQXFNhMDWH95qMauIer2g
qBQQA7h2oWoVFW8KexDG4TURxNNOhrGi0HcHng92diZoOBYgK2kAb7mA93rSQyqPkgXOMzNH0+I5
Rg0v+QTP1MZw0fqnVhQaZW/7fO+0qkaUL4w7t7G2onMyFFTulUqoVguw+sJTtedAmUrPObivRC09
yCGGFhWiH6/+ZalfZ176dLEAprYsy+ZYT3V9mHb2Tvn8eVlyMKOsiuFXpLR0WOoYK9ng47QkP2ZX
Hbf80i3N+T2U9R8CHCCXrVkGnLi1f7j3GJYDaBTgR/akt+7W2fZBlA/v+BpwFZ0TC5Ncg0uMAdRK
04dbGXP6AVUoFIojLchPOh4ep9T6mTuF3YI12O5a1AMmZQSb4YE9NHM6ZtmlHqRAhqmI27bIuvmt
f0N5N19OPeANECmMoyaVWc03Lhs+tgucTwLVC1NTOgsNguD98+hqWyZrwJuvdjBvUOCQqzmDYwQw
JLLTSgmmO7JholSeQmN2NSihAEX7I/9gd/n1guOdcG1RrN4cul/5ihAuSjivvgIJDoCfsM0zleHt
pUaN6gdXFibiw1aimZuVt4Bd1cT0enOzXVgm5fx/DdRNgjytdeD8QWglI7nxCRudGN4S/K/ktC7I
0waSzXCcHbYEuiJiY10QLRDrDosBPSyAMK3ch1BxmveZNNQVCzyJjiucyZKJCCR/hM2HtlAiVJQx
iBXp0QIkp3Q5uA+OghtXKFq+N4RrLNYu8rtq5G3ceBKTEZ9XjheCQhwICmX1QFXaR+KGc1qjIgt8
q9MaxGK6J4DCKJkkrZrwjapdenquTZhed3IV3xUaSw5n4ecf2cDqDMK02kYDCUE2elqGjZdXnIdL
7SvBkMOWYftDxzLXVQA3h6rsUkwhBZn0sf+9o76+g4MVmLfQfafmkbnn6+j4oH9d3Tkg/BF4sfJb
eACSxWfvBrtWx7zwmIdzdoA+GEnDCbnxwNUDbwgJFvMW9MM5K7Vy2DfsBNPNtak4M0IV9LU9EJhY
FmSqRwz/2cmmylGCc8JIH4I4yCnII7V71O8xk6SSI+csCmguycEx6GyrIcmVUR4d6jSuzFhQvNGp
T9H2zt0OTFQrZTmnuT5wpP0YHjnKggLwZlL4jYfVDJbhYX8q6qhElSUWwImgQkhxnLc821UWRWW9
AUSr1xl/w20LuTSQY42GsHdTDT43y8devGFCA3zW1F8RBoWHRrysjBseqSkSMN7DP1UnTwk5dhU7
7Q6xPrm1b5XXYrFvylH5BXeOnvPrSJ2/4F7rD3MraTYA2ajxhz/DAzRIbXmJUmnd0jmqHoZLzV+D
4sNR1yXVW5hepSOkQcOdixCVwUMkAyLyXc45xX8wR0S5aeE8Ftc3KhkgOcPzjRtCUdJIRsj8X76G
hOhwHY0jWPgNP02iKZ5gGtT36/WIFoPzIJ9SdOinXwXl4heeUrHhnM19cwCfF5yv78izSl+Ft50W
EMWyobrxfv49Ahv0w6phkwsb7nQucM3RETqXvn0jwZS2YILQk0SVyvwy5k2IYvNlJr95gHP68cv6
1RZX+tmLC1oqdeUQ9nR9kLVwmdcfU0D8BoFKRyU+igXB+OfoU0BtwSZvqBOqLSG0AmGkWo/twYyK
6+/5E5y3VCSI8IxwNINBqfqpFNRDUxizR5B4trWDetkIIWbtI/DWkYcxILEN7kF0kVeN9jl8pBJ5
XXUYrIBW3N8lrA+RHGgLIQwxC5Qygu8ecxMmaQqwEZBN2zeIiIMlRGP1QDH7xjOeDt8wZD/AujTM
Uf/sWFdlHOzf9m/uj+LV1Sm4MQKaPKBNTjCkujviUxjr5q9Y+loJPqZduMof8pLB+5W+VqaDLU2L
SnKFU6ojOeZn7Ei4AgJ9qjyAk1OREAxPwWay79cBgJGMS4ahb99LwwQdTCX/XEQ9+n8TJSQgD0Ft
jUbRdLByfzaPDhbfkbfTvaQFAQb/iBfLqBlEmlP5ptSIGT9SKBe3LpqWeFr4Tfiv1OoESM0hMNlx
YMSEQU8Vt4ghlBGYadIOS27GpY5U8gprdOaqolBoHagqgRFJ9KQsUPVsWlNh2XSZc9K8dXObYfz7
XYHfW3l2IUYbeLic8R+fv6yxyKpnqqVdGGYNc0K04MLZBtZq9T7uNJViJbBPOlVgS5hGvsqaqI9x
z9kR3obGWQ8+i9F5OTKwYNqhWbSP7k1kBVj7+ps23+bhBVtuADTH1refWwZKidgbyL7nWh96HlW/
V21qV13j20pszPxgpKfvja424zGlxJMnkVZC3HkhUjfEaJ8m9KE6YJfD6QL4+Oyfrs8V3pR7y+WB
DgTrSpCvzXONFz0PKQENuMIAZWQqcvXnEtS8LD2YlEi828YzZ/7cPhMnvXdQaE0gZC5KENkECiOS
YW2AFUTqiT3ix3BHJIJgzbuMzPDnHddn/mf10C9d2oiquSqihq7qJbc8mkjYb3E0HNdPohOLq3kx
Sb+eu5oDMbvq5gmCN0J46zJIgLK+HrBm0aa7mbW67u9VVVGdVcBK1l0aHii4OIwPtWL18oIcAymq
J7H17Suig5tO/v03v0sFm3OvQI5kDyqm4d/FgxWgdKGBBUcndgX+Q8JwTbqcThWfrP7El/hb3+RY
7UqpWyrTo8laA0Ze8fmCDDWVbKVsFf1UHHU/N8Loy4kO8dOY1OBA1DQb2ZVn4aI9YAbo1Xvl1aHU
ZiaO7aHs+I3MFB1JZrUueF8nVXhvNSxsAU/r2dJ+9gBiFfhyRdDTnXspp81h6nqspdROR/TcieeY
AYlurNWGoMEoTj1GXI92h4//gAelKhvDYSrejdmLaCXOb8+DAcop5Om7Aak7u+tf9OlIvoDog5PG
J5X1IxXl02xhsojIxejnwfXOLaX+oodZ7eASxMyvo7tIGJjAi5eLDU7O+I1WjkJKT7hUfgpHD7Rq
UPdxlYlLIM2MnFBHn/n4+1ZpAAqv9AvjBJwzV0DLaEfcXj9D3/rM2Hh9aBl1qRCidPVcVIRkvmko
10HvipXiN+oxw6SOWdkWb2T61zjhrx/jTBmHGCM9nBavrjZvwLSIz3zPmzRY+RJ7dSE6qjhAVUhE
P9fIVRHSxWd0OVhBp7/iK+2Twj8sZMaNQV9MrRDgvsUM0xmt2G84oBmrTE8wxUMAoVHHuy6wPHQy
AkKWs7G+/b1iDTqBZ21OZnu9AY6gE1jMMyOcpKNpRy9ecV/aEi1oWme5QYvqrQkR7y/wdCRxtk7k
ks0xGD8ZexVdXBPVOGqXPCCcVGzU+D76OvjYmV4hvgL8OKDhaYKe0q77y0sgVIJ+Dr78ViBInkQN
9NkFGsRexPFHcgS+SQyTL4zdy5jsedzlcaV26EUDm1gicW8VftkcEtBew52vIEaL8Q6Tq8Yq+is7
PrJrOazYmST6kpEI7V3QUQkM9qS4Nl/sO2T72XGmgR9BilhYnmqFKNJDNdezOsbdMtHzyunrYjGo
LN0uIQEev/4AdTfIrN7dWck7RNCfHhcxRalrJdmv5VqDSB62KGSaxDpPWjGroqfyYODLiSYXP2YV
8gyn50rG+GV/IrgdJR7bYcNNmoC+Pw2nIoWABEUDkkeYlRuL7YaPHjHDAvqMVKkWSpxJ/MREMLxb
PVwqp2QugdleNGWBL0OOmWelIjvLNWUr3zMsCVg8G9IlSDUkg6kPgjIk5ZYIvgXrzOyWUAE6iNg/
h6NOlEYwn5+Ea4ljxm1wTeu7HukNz1qi3XD3rxsZsm7tEAVtYfNq9YZabpYx1g6gDlpO8ZMAgeOQ
+42Sva+ehFOnoVn/v1qu+gAxLIXW2bUtowobITuvvbgOhKMcCTSVK8NAdgoey+hWXPFu0Wntpw9F
Vk3opGx1ZL7aRNmBFBaHBDi23b5LPtSkbyvmzFCltB8X1ug9XntsWK0Bhv+orZgRPD8UGDvbJ2ji
+coB0gLgl6nZ8Bmy7SgJXFq3odsvXDXxD06OpBkNDDN99wxAcsDsPUJk9KmTr5BIRLKy80lHv9hV
4KaPuGAotOYwb3grHV3TDkrXi5JfCie+5uhlZA4TPjH/8yA7hK25GLtT8b5FNMRIz+DGIqbUHc6L
tKqDfDHpBRNxSAg9K0bqS+lnIKOGcWUkZ7r83QdDmhnrI4n1Lp6neX7FuI+0Z8WE4TBg9Ka8sVe9
1nEheF9PWjmQaeRZzNpVxr7Mt1YpZukkSXq9Abd9DsA4Ha8Xp8mr19yKxIzAXvscfmaaiJANdrC+
7AK6jXQjNleXsXwXBPRYWabkRluDlpnc1hsSNvbIP6IORzpK4uSfnwV8j4Bkxu/4PfiWMPZ7GCz+
H0p/mIJGp7whNFr9p1V2dXIN8Q7JPh1Mytt36k3y72pyB6VM3ihUKyyW2CpKmlVyg2fuLyeO/JHm
WC0k83TqZ2FD+qgERvHQh2X79aaBw2Nj7rqSGrTj8M/fozUmg+CNrR34hpi5LDuXhQohEZyAyDQC
X6/knopVw/ybjk7OUaDdMsIpu+sjnMXRRXxPHGtlRQviE2yxe05TfEmv1UCfQtJEOMrsXKAjx+Pg
LDK1cyBzNxJXIDx+1JotGtmCFPoneNa3EswApovx7xh1Z/SlgPODXdV0G0Mv+YIlFhDjbZA/eIKT
fvJuGU88sIjUjPQnNnkCvG5lFPWvL8P2lgdwDzOIPivlkUYBlrulhSW1olt24XNiEqyiri6Sgmij
PVqEXtk7t8noCU9mqq6tMzNLavZ/gq7vVeah67QYmPE6dWuEFvBWaUO/AC0TFbiVqdwSZ6cUihZY
Gs23bPMjQgNonk/U/XLV/oY8dTI3y0edyO4HnSuGGl5U286SjtgKCGnpjvnFoyYL8CHlK5BDLqkg
rO/W3VsWicWg8+CRFPbOQHvH0ETAWtLd2noabEyPlobhfmD3AJOE5OY7iDSfT/UQRPHapSC5iCPK
aryx7I18/YYmXFXFio4IB5g7gt7jHXiWEA5nLw2ZyNLXfSzYe4MhoA/TNnGBmzrh6gzRuQCtEf39
LRUxTdK/fikkAR7wXgOKW2osB5daZ2WpEH8q9jF+EcIexhWZirYAnOVyO3J3HDUoRcBdOxnaLuTC
FsaBqR1q7Pgk3uRtogaBoLeNdJYIhJd3exNFQv1ZBAjpSBUJ2mI5JEd88/RV540tHG6I0XTWrzHp
qdmLrMmCMh2hsmuMoD+gW+bHEEpOuB6GrlmJCkkeNdAMXWUmi9xdLhgIwcqBttZKW2JTLCoHoRvr
p9uczYXgR7Ymwc8Y2yuDZF23TEMPsWosXWvyUN11twxdwtDzq3Ydg9Xr8WclzmdBSSOki5ySyteI
R569AK53xRG1bU2begAoh4AI6BDwI3DR0imMRM924Tj501i6D0s23ZrzG0lAlOrZLTjyDUg7oa8y
qNkp5nb6CzpGjF7EZ3r8dbcYXm+e9WiPTZLFlzmZGnY6ddMSPxHvDakmVntbO8US9q5VT+lH8iTg
aJ9vFZN0YK0fYu6KSAhkIM4F4WOsfZuuxwu5orC36S0ThQsQNE/CyAXIqbWYtRY7EqEeutNfrTA8
tMTi+grXZpLhla6yLnX2tGj0Ejg0PR1Xnf0Bs2V/u2uok/rHfKujrUH9wGmr9wkjLe6OIJZBwVm7
SfMbRWKyDIEohdqHC9lEj27xPV8Q87xUlvHoZGcBGHtfmviR3TleM15p+P56ugtIXfGunZZ68Ncz
WX/1yX2YxQjJs21h/RiLv8NzZpH5knCtpAN8d80WcmK55ZbmaUBD5q7ic6QTdhu2dQwmW66lJkdD
jkxU0jQnlUBcv+E+PiEHc/ZTzDCd76Jgkgxqhgk0gi+TriPYLTWDc/1X/Az/F9XE7M2/0FrnzAeb
/uMdil1ZfTjNhc0lMCb0/n36YDjW7Z4kktHUcFEvvaCUCRgDQHJ5y1/VFZCEI2+TsQDFItslikCw
ezsLJSSgUzSRCyl1Zrxvo4a7SlsOnRM25v2IY8OcXZcb/VS7Jny+1vaUjuN1jPrIfhjlgCmzsnez
TlNrY/cGYSF8y8ukVNGJ/n/6Y/MmnkJHAP9+kMhdgBdp1odJfPgOxEkefm3l+HkU8gn1LcmvbY8z
/yNkk7VjfdKfgZcvlnK/mHJeoC4GbLRsVlecZlheQgIvYWnmalIT3bbcwDhhFl5dw5B64oJNXodc
Vk6xYnurB573PXeAyLCnC79pq19M36n4iuBnj7FabtznAufCZSt1i3R4Au5nYl1sYwE1rmzQw/G0
lofFv6Ptu/l+0RqlEGnT6E9up7tJP3Nb6n+uogr1n1FlPx7aQCZMKrSTdd8++ijr6697sCgAI0Bk
ZEFDt1PtKao1iRM9WLKFwuGXNGi64RNkOlfCLHt5rehW9xZQ8nxcFcBM0TDYVxuGzBaRwEIQ9mVV
6dZbvILmQOPXyaihred4DRQ38rlSX3m2P6c587PK2ajB/Motq1HdOa7BOuqeuqs826bmz84OHB+P
Bh4DAjxiaq0Yi7IX7DrWmg8S2WNX99IaIvpD9G8yR2bAUP7PR6+rMwQNjk12MOzpLxCgnNx7rFHM
M1wxuqKtJeTh+lDMv0dnR6eGbI9bVYnaa+oLYD3YxuhQ4KPxhiHp/MmzC0d1HQdWGFvjNHfl6uNI
LXYx3+y9lTk/S1i3K/b3UIH2l8HVJgPbQh+9kqoxQYYFDrtw0ovIYbFq/8HnEyEwrJHfyO1q/Y5m
9HgsDmXM28jCWn/czy7q12rOa9nXdMq1XCL+kmwzYKIn/ezz6NA5G6/QtQ38d9dAVPRjwtMDHrSH
jnMOi8NLFQmb+i57LtbNgC1KlteVcKwjz5o8x/YybutXTdmjXipZtVOuHctNUjDj2LEIxnmNjDfh
IOTIJkBWdpLnseE6pL64T4bS5ShuhN2mxJRqeQmk0sE5cwA3ufasgqiY513da0fuDjnLf3ymGrML
e39sgSf0b6NUxvv36bWHNrknyPMwAPShJ0bXzTNIcNs1sbJg+JgYCIbH1IuDArkXSxFw5S4gyVJv
IE2PfBjDJHf9T88r+bUNrymycIYPB3n/lrLSpxLhPVoC96FC6oY4hsFNPXlKmEbxqqmFh64ppysE
9E87WGnTg+zvjX8gKPKDa2OZc6PdQnwVyL14c8bUylOaHJNNgoyD+FHXQdXpu7nHO7+31pJc1f9z
+5zyd7dhr9uDPY5CqRdF8mAMsV9ErIWH7QRxPXyuYFwxQgBCWlF/8mIlQd6oholS3a5blQQOF2hc
UApc9ZwD1UHxEjmFAfpNg5cG5xxm3jf1I7dzNfqHjjRyhVXNxUR00sISzEwLVuAvT5nKhOGzRDfe
CFRoLBFJedeIE7reDwy2Lm5Pwh9iLbLLtbQmQzSXpnyy/OXVWz6kdoB2wG2ALirQUk4CG4gkhv0j
dMFarJkH46kY/rG1TWN8s3G0/yBu6Tk9b6znhdM4IUHuZNFHel4x7ZG8aburDmhiOUM87wVu+KLe
J6KkqSco+zF8H9marVgvRBTNg8RjmW3HSbwPVqT0l+zlbsi6ZH9/LXKBsEbujgi5mHdrDWQ3A45d
sFb5+BNEcbmvXm3gKofRd6lICD1/HqvcF4e14EfD+B+awG3fhkLNt/5IsaCaCw4wLS/d+NY9HUfZ
XQ+MMEeYi/kvFEKs+5CQlC0KbC87Nxzi1TplH9HbpBz1lW2dZkf09C8v8V4Da0Ehuk+SRRovpBt8
Ehd5VO17K0tc0pXLWMxtL/LmTkMXU0tLXC+TL6jk83fQ3JaztyEcGArdYLm+O5tHhcb8C15scoFC
F9BeMOfkctVh8dg8/EZeKOfSMTxprvN3+3iPhzfZ3yONkX/j/H5Yo+X5KoURwxf2+7rVkxkUkZt3
OupDNzeR3H8P19q4tSnvgcy7qPzJfxGvYN7L5zHHlpId+vbbgRoA1He3r42uFpEf3hITEAgeZgE4
iY06KCX0ng6zGsON4sAh2lP1H5PBcM5fUvsNCBnZS96+aC9z8HTxd/96FiXGeepDl2XSb5tOU+0R
lFWw2hhOWHyOIkOeZgB4YECDgPtxdWmmmDMm8HVRQDLbgz3h1AaX9D5X9QGl0UYYdCrL0ou/Aknj
SsI+fzL9yQhksTPQb0YVlTcsGPSuGDk5ZSrz6EJwlyr8M8J/YkeT8/DmZeIP3vR6KEhSLVJLksQ6
qB7GpCL3z5j7CQmn1xmCZS4OrdfDgCFQ1Yf8pykNvGONFv274TxohMF+ijnBXo3zkTeErE3DR7JC
rPbor5EmgQDleR84nBq1rf9Q5Xtk5RRv6xTtZTzqjZCZm5NstqQteYPwZsxI9m7LgwJIkoWoQRyP
nn8nsHLO2zzHMjbHbiBv+O6ommVQRCs3UoHLiMNMED42UwI3I4Ao+94TpmMoV5lWSudmNf54C9Bo
eatqrqUOvHE8GKEceuRrtiWVMqunH3/dHffM6F0BTFduKH58EjojWw9PPlJNv7N9wk3TfWpPDzEo
rePNU86K4F7rnp5Xy5JDEDdnkD2sV9Q3qgb1phZ2EIAvFcS3p2oAxrnJO6gjlMbkVIMHppa9QfDn
WAGlcRJ7wx8PGEcfYMD7z1uR1ShFTK71fd/eJiY51fMvtxbLG8MS/lyu1zT8ry5jGuFdKYCYiePB
084f8G5wPu3cWXI487da+KPVYnHEswb/XRjh5h8yr6Cls02VGF3oWf3Aa+/5O9M6hdB8QtTxkg2N
plDNEaH3sl3gUwDz7wTxVKUzAVja0W5FAZ50Q2WuTzzZ3mSE0n8iBvYrU/Lsrp5aHdARq2ZOp8yX
cMk1/a+COASG/PuNREgbDzQQjIu/GhpC9b31NG4ZaQL+IDfsS9z8wE0mK+2FDPDS6RSQecmns7T0
yIdXW7J6/sPNCo5R9z4o/rUD0JjLHRL2yxf0q0iKuDCqLpy5xVWKeYjhlebvDOve/FQ0STEnSns8
AT8LWH3fmmfW4ODaA6stH180Rrgjp/KOkmobBlBQiC6yBT/o4FoZKKuPnLzChbsgQrAbPG7VaoOq
vaBgBaPU+B3N94H5naCbRlTTMXHsL++6slYbm6df/6fkgvSKZF+YRjYQFH08ySb1QhTSCtDfASXv
XsAOwSfzu2GqHWcycjzJQC4RWgiHSu3hm+ywCyOA9QWTpwjjRvTjHAt+qlfrax5IXq9HgIE58/5c
GmZg+/T6ZZXLxksKJE/novVVeXeKfwYffG7PtJ8C8DSICe4EHbzqtAZUL0ABrsNIQovzvDgEvZSx
+HTASabBPEAZK/tfMxcT9jUMko8P5uMZ+/24NPmfmjrwsgQNWYncX8qfg6wTDsqBc8Ue97/GqSp7
mjI/W4HtXd4Q5VpwnNNI0J3OkUSqmd1GdgtcfO78M/161RXDbyHRBV7YZuA6dh7pWKQy5821Af5d
zU+xEXgGqGhenmyCQeddLnErw6GPtLyH1i0+/N8iebwuBzDI9fmZtg0pbYDoqr9ZRlK4ZBRCxZjM
8xng2vfsyMMtTikb9ioMcAayJ1tipn1jxr7rgQbGnmE+RmOibcqR6ZXj7R/S+1mXq2/MxlNSXsqo
xMjJoNY2y7zvM/IUIJl3cX0QtOYLN0DPKbQUVtOdqzjsOqboDyNNf8m2GU1RijvPODOjQSO5CYvB
KbrDT5jcwsXAAiG9zSyqJMil6FiuEUC1O7SBpAWKqBI6Bjwg7UZph/aIbk+MVy9AhkJRs8Ol3Vbv
kwhHaTN5RroMdIQyMbt5bDaztMcgkPUu9oGfQOeYE89Olo+IyghrHbfU/CVMjVArYsNYc4eIVqf9
1vgl05oVYGlANbpYa2+ItGB7sAloNJ08fzu4vDEUgBzRubTQLAus7thHvC+53fva5gGiY6R5XOjy
wnXXGhUDWIBWMupiHcjh24f2fu22mZ/orUmjRPUFHvO9qq5pxf9G/pveGuUPUXMa2Vj45NPg4SyI
SwZdrZTCse9/OZwazMxA+ahJfYDgbTS+URB3AN+YUFd9vLR/vVpYm5fJE/MfMIT5q127l1OvLW5n
G/REIdYE6/qHL4D3NFYZcxXweKt+QPmnuKtOib1nlX3h/gkpSgGHSzyHPpAD0Y6UucJlY/ky/JfB
7QbwGWTekzfhcrJ3M8q1UK7s4utL8hHZhJ65W/UHtwQkBekqE++GPhD01BbfXls6S3g7ajDhyEeY
n+6tLYkyUEhdb7YfSFhDb2AG5acCecGVpoy16qAC3AqqhYpwyjbTNTiqFlDW8SYLUUnW/VzlGaoZ
0FFUHQaMg8X+tXGEIj4WGpSdRzaU77ufBoq1lEfuH9bD2ap2/NDl+bfDn208AiZnPbHtz+UF56kU
1XnRhYbIqaPd+/MJUvPUe4pl1fq5M051Ecf5xRgfWHE2UUgwD/pGjCi/vycr+9aSkDdCNJu2eL6N
YrWJHXaK3TTr/DvEiMsoCxrNrAV+VnljellUYKEDWmLughXpIBXp6p9LxOUBbwQ9IZnFQ3JQwMNe
rQ7x23YHqeGtyjlwmkQ7S+gYulDzzipGMvrDij9L9ZNqhxWbpd1iAB49HCGVo+Xhc9GIvh0VbQ7c
804t/rSTp6c0rkVbrS6NqyrzJdU3EahKMtXdaMFclJboYY4L0zRBlV+aCt+tpSZdBljOVkTC7CVy
rXSC1A7E2pDGzNTX/jSp9918CYy+2XQLYI9ZcoVrjEQQnZHR4sEehfJNFZvzB2pJoKE7g5d1yS9W
O9f6cW3TPrvHm4H698ECAAx8b+2akVLjuPwHkzdwBB0ZgI3kZOSs1SCBLHcYUMicgIUr0vIqBqsL
agSeG4OjpkJRfm6WU4Xe4yuA0oC/e2tXsDu11U+V6km359mUt7tLjdUSZU8Sya+vWNBwcPY3fhYC
a2gBIM44iPFk+KtkGxvmyNRflpXLp18UJS4f18eAkzddqeKyzTzjrrwlE0A1ZYfxyYzejDhnXwD4
6gYZgGCIwFXJH1bbHZ/w2qee3R3y+T/nS2OojR5sQRLCONQqhFPxllw3ERXlwXrWIaCq/d4AvgdN
lmN1G0yrB4DScT4hWva8/mcHSfXb3fE+wpEiCaReAQstq7DfkccRmTVed/xjH1GucSOoieaCRMwW
HxlUe6x7sbdqvL8n3oLeNXOgEUbK7ntqWlA298kaxcdxgKVAtK09Kdc46xvzqoU4vUe12aT/pcfb
6e4bVdjxIB6NThmbzXBU46Kxuy2eWuatYWnYRNk2iF95bcQq0dYhGHXz1CzoRZ+Jvke+BO6zmoH1
mmydY8TrJ74UfVTZ9qyncPLgMFzPWK/y7R3mLkkc55zRopyWe8N9mik6WGzlrCZ8W+2Z/0lgxDhl
rJ0N4e0ndTj/1B2yV4zp4zD+wEyqn2RXzzsPNujR1Bovxk7kyp+nvTN/7HreYx/o/uH5iuIndru+
1ocmD2hBs12PQSykQaVmhUGU8kHhElj1vZ4ozOIX4Sl6KsDrtbrZuO4fTV2bdnGgoKvlCc1gcjOu
qrfzhax+4grkU8XKEEoyikuQ5/IzG8qUlK9iSwyEPgE9OSHcT63YpdAFUCJCkIgqp43pnYy6m0Jb
aXdjLBN+NrbkhY1kdq7AZDKuf6p+u4U/ANW2asXGnvhDOD08Hd90/45RMPw+Mc3bfe72USASQ1k5
jnSh6C6AbPyTkhoCcERW0qwK08d9jhykYkTqbsDUkctD9ElKhsHYmDxk6bveiMTOHamVqnUSjJSB
hiCdAfxmxfTQSxb/OC1W3iaDhKJZZdQbOU+Iw2d4effFVQS/OzzOc+WKKlwXJqUNUOPCnKkW7dU3
W05Wqw858TNyEIQ88F/xvmB5NF2phpuTEYUCtjs9/VuGNKSywGE703rhnfgk5bAf1BpTEVazNPDE
Ife8nFioxik6QWpMQLpoG5WwI4NT+hRG1MXj8N97VObPM5gleAg6ogRxjrudhI1l/2XxdJ9gV99U
hM6hWcBKBkoH+79/bBUBkDpKoc5d5J4JMnYqFvdXnISvUyIdSAYeoUQwraLZ/snKf0LubrtiKV9V
oNhWztJUc+etxD6XlQFDunzwBoufc3og8DW5ZCcazDUZBx8fN1AWp08DAe6LQQLPWGIcuOhaq08x
B/kyOCzWQEXoaooJNcBv4voKswHddJ989D8YuAd1Pr1cyEQQr+9U4iG+anVAa2AcOm79XqbFw3VN
JOORUQciysEJG00FsBnL1ccz5ejEGgVLhclig3sTz0jjtxfsJsebIYAaPfqffdD5REmoEc3jL2KF
Yk6SyyzN0jPWjo5kdhYzPkTmJQ0tW8AnRUWskhkhyi4CQ+vfAR5+/vT+dZFO741+yZ7vVDRN2HsT
I2vy/eH1/m62qDqbXs3hAxR7JdD1+IPYP4zZMok6Uc2MWsuhgM1/DZ1EHagHAZIydr93fLy9UaoR
IiFaz5s+K6V5zXhld7XO9wtal0HSIADNDkuBNX0c3Ar5kIRVQAhoRxPKdrekEyqLnral22x82SIQ
vgbAzCthIkZ5V5TSVRKr45nVsQMwFCd0k/FyBdr6iqob46GhcqDynwRlrhQ8hFO227vzrvvbIOxq
r9wxoyIR+a9cCKagXKK/cpo5O2RaUaepq/jQB5nTclkAqMUr8wcD97f+8D4aOBeWDoky3Yy5y7N8
xPKwCUWir1r+FilPmZCyfBUokncQSLQ5BphRfYZbp6mT8CdAU/+xkeV6FbmhxYQ/t9JQXKf8o5RY
ZaaZbQ/h0JJ2RHuqcU/mNC2bTqzmi5l30X97t8GKEmgyk2PCaGzSTqdKI+iqPDsjYB0XfbKhuiYB
4TngNBLpMA/4sXYzwnVmUaNvndEzHm5W2HgC9XIYSdHtt7NWusDSYYf71FdEZfWw0mlpZOfe5OGT
GkzMF0mwVT05bl0ObBstLFyiy1lr0aUGq1/2WeriKKv/aBlrO3Twk/6geZdkh+luOOCy2El3kc6I
kgyUGXKIWsbzLwjbuZnNdVGDdEbABJ8VOjwBX7264mgOU8NU1fYr+Q+uud5ZpOTcL/R2Sbb59PZE
MgtfkMB0raaCFVLwyLRok+hmgUGCO/ar4Atj7cu5zCsLQccmfcXtDzYWQ12dGRqMChdgjVbDkV8o
xGSHH6JjfsVSYk+O/WUy8C9zynLzQMgKslGJu/vmUpgLADl+UNNACbdu0AzfHxiMVFSBALkyiZdc
7j2XQNQeuPoqvaKvIyfqD2VNzhQFz0+mTnaX9iYrKkKHCSXiPSH+GqourKujVD5aMlWqWoyY9+I9
sW/2Dhbyg+zbavg0BoUCNTrhs7usgH2xiDZFjQldKzI94QVUTAXbfoICFgB4yk+a8B5cwDgC+ARe
6PkBFQRXT+qh64BrM8vm/pJBugc6BaRO9kHwThKwWgL2d/Vo+e0dps+bdXdzgT0EUYzxjBBGvK9S
WdiyBAZsYDgwRWqwwnu6U6ZXuBjez7XGoFX2DoezSYve4gQqoFAX1JhziObw1V0aUFGO01DcNJTS
yZDdV86VDlo8hdk31uCSwPTxuCrrXr9ZxHEnxfolF+JhcOgrBqExN3VinV9/gzRq/+eenmQ1ZdTB
LBCMsgvtvs3QDVT7nZ4MAruzuto3LfAeMDCSQwq70TRFAVS31NtqAPokbRblYx2QSYI+/h/QBMYF
hPpipVZZNPLGBYTDMwsv25NhcLXB1FROrs6QcYG3g28d3F5mlajTg4T4xARVgxvzD9nY71rcmeaV
0jeOQbF2Zsnw5Mhf028YCqQ0B+asMt5pKEl4IQYTmk/+aSuZ2iVX/Ybm7KSPvmiQsFB3hYGa3Hru
T/HU92TWv8ZdIP/2RrgQwDThv+yEjkDQIKSfH4Yyr1C7OjK0qdLWEi+smtJ2CJLAHVKmHABSYzHt
VZnK6WuqGcXeO+AH+xqAjf5ZAeKBGjd2KNgiIqPYJ4fVdLZTLmu776b1kwtvwHalWBl4lOKfDJyH
WLdKm7oPp37B2cVBmn5fmXEbzabCYoYMeWGsKlp2kBj9iNAGiVL2AgY1KiUx80An4UvyLBdPpAqD
OS57Um4nDkacMdaFWXVf6xUClSM0DpYHVX0R1I0crB9+PrX7H7k1OL6l+1HVTo1WAvwXfPGFwq+O
xf65cpDXYsTMufOn9JZfLz58Z1Wgf9AbVhz3sUVh0tH3cmDSVx8a7zAd/FzFAaRs23MJms/b/H76
Rek5x7Z0VmxQrRWUqMF+ICRyk8ssG/VehjkiLMSDo2idOM+YBrmPF0aZ10S6z9lUJMabD33oSJ+i
BRC58XhH86QrjFbgR4HHIBcdloq5Dh42J550jiUcGlL3jj+MXsM3PBz3UinvZxTN1hPEf/U4uSoy
2PH+PLxcTFP+BiIIYSQeJ6KwAD+xGjWucTx5e2YttjbOCJ/OE4YQ6wUkWidaFiCbITK+zgcG5dw9
Er6BkAbPrcKm9ij3VNxlF69EFA+PRzFdb1PQs0g2sA/BXrPp/paoZG0Wi6Y6hVp/EI+WRtsQUtap
Zb/biXHQK4v9WKW19YoqCHK3yHaeMPUzuhAljDVX3ybp2jHI3viLXVfG1W6iwLbQxR9iiVIlQWiy
buTbIen1rk+BWV+Ckv8CxAQTn4ycn9POzkth8Ejq4PJwPt3ejR9kHG2qtRfTDXp2CN+3L6I2XGSd
R6FWY/WYe1gcI5gQnS7Pmd3bA73CVEcsa6GY0WkVKWRiLtVTb2/L+fvAUNGQBUHNgE3eD2gsM7Yh
BEXGtGq2fnRUfjJZmUNiOO3+JESFruvxSdpU0sll/nbvAzgPlQOxCBmTwxTnzE7qoIn6EdDlPe9T
md5wfeROhAgPronxIQ9uBlKpyS4H4VYWBF8baw9reGEJk4TlIvmshw2DBwqJEeIOVV8LJEWYVinD
zpNGq3O7ZO2wvdbuWvZaE/2q9NH0Rmy3xKpxLNCL+IZ2gJNk6ZzLnoSyeM6bNCysAo2Moi4iz/Me
2ePsuVhBp8DR7cnyV5uWg44NxUf3RZZxgSamshqO4rpaaxnY6MPmbGqVHoJwyD+b5BIxDiw2SSr1
1joWbPCPd4n5TTIh6U86UB/yv91zHUgSADeLwQSoTGoQFfzcNiUI8iOBVw+2BqmaMhdb/EBVtjRi
UnHmQcROZppfy4ED8o26aG2RdG8so0PyfkktvHFI0MzofxhkjteF1cgw28VtYF9ipVcT44BGwmyK
BLQQcoNsSSA4QEj3lP+FRJVuJcA6r+iYE51KLQWP9abXRx1JUESY48ssMjCE0WFN5uqLK36G96EN
NE7gDGz4SNjkKZ8S05gV3MqIifoAXdh4RMC5Ww9zS2lyqBWGCj7onNq1DTg5CjQ/dUxwYEZI5Kc9
GwhsqXU+WfZpmksu/6784DWNdgFEDg2axu2uyuVlIQw4l3O+bDmMZKLOZnWsTWMUCndwV4rlo8wu
z+IuntH9K9glm08mxbw3Od3whhicWasyulHJb96nODucPUplcrZ65s0vzGn7pdblyehrw+Rx9vZ8
ulz0gTGKceJGHo1CTiysBE7AO9n8kAKOqIPfWVjRv8U8kXsAcY0a+uEZNkh65orL/JjPXrmi5zKc
+z2x6/oNMgy7jWtl7WRqTBiqzAmULAErnqMpL0fWc6+gIaVHhsw86OAfuVrvNfqTzvsbox3ifuxX
/DqcWXGqmt7LUfvDCHDp+exveZN3lsYQuC1UbGkLTSedqku/SDEjIX8FDxFRoamyt8g4OkrMLuZ1
6jvsCJyz2ifDiQOGLDA8tML83crS+so4hjyjvReQkmogzyaPS17VHby0Oox1Nicd4vhAk2leoFZY
+HeuIefHU3RJuZ/MjOnQJ3GIz2qubE+WWpp3qfmJe6vmvMkrYYB8QaXRS/B0ISbqXE16VsxXciuD
XZ1L+Y7BnNbabb5R3qzcy5nsRqzFgJTfMb6CNhNaa4sfH7Sf+mmZgjthYajPGM+WUjsrpB8Ps0yN
6kW64IWtO2veiTiMi99j/JaWZAYg2ev0q7Qo5zpSdChaHLnQdouueWE48cazT1epzOOv/WZyXRVd
1y7QJHQnbwU0PiXtSzGBZtwISn6fTtRGoUqm5faOHRfDhaPspa0aMjzulikG2i706GZYEUKOZLih
ffZZ9MKlI4n6KAV9VqIeJjM2o+KH8k18MspcxmEttlCWUK0THLiU5/hNlh5tTxHVIiIO7Zzdn8ub
gm0iR3nsHkacNxoA5Rvp6WDhFFOszU2Ln6XLRG7DY4niTZkC/nTqbo7DyvcL64AukS7wI9gyRWHa
Sq75GpFSLb4FsiGJOIOLa0Bl0sLtEyRe9UBpsM8ibvkIbW8t7D2fD9bNESUzVuNuea81/agErfRm
tmU/Bc3X1ckEdP5VWcRnDvSblDKbtTyrTkUp4rRVTagiXUsXEXUbycmpJP4nrPdulpcL+S4syHk1
uGX8G7x4rCHc1JSPtF9K7wpQDWd7NViKbruOR1vIuQR+kyfb7v5RRGZ39rO4H7Uq09O3rkvqxCtT
+n7b00VhmpDCutEAvhZ/p0FnqKFKTBuAQkGQ/zwbGu8aUw/33Lpq4D7P441j5qDhqLj00NFFFkFw
PkTN0024/KLjMFqTLzRD8oFlLwIROwTfQKrvB/AvFOGrciST3b7gPApRB78EuxFaRTEd/1wRZyhF
AwKEiwWhR8gxJ/JhMBh78AsDR2PfOD/Atl0vB1e6w4WiQoqVlyv3rzHeyjXAelrREmTDa4+AFP5G
LzRmhMM6SMhRVguw+U3CSnjnRgjxxULCqwS79rdvNqpY0S/xDzI2Gx/JITzSKVmfinD85VniOD53
zaZTMGEFepQqBiIbjTyw8z70UEiihXN2LyIxQSJAn+SCYfN0lmlk19w6rRqpqhUZszg/0Ot/Vuis
qkTFbCScVnj3+DZHq/INzUmd+qvYDc25ulvyMcj81fNzHINs09sqytopjeXmBgwyZwROJBUeeQYZ
YKLEEBsx0K1KHUIRbgIBSLETZU0YAiqmg8napFySzx0GYpnqOjt704U31r+SPBZf+AWa9o7WTnng
qZURpGHrEGDLx+MmbXxzzKjWkQKx/OwN/nP1n0marAkXZGkLC0jupsPj8S8M4ZbgvopXsTKHXAHU
EFkjGYfROoyx4xjscpa8Py6ZM9ZaX2nuVrxfviOveC2Mi0jUEioemvkUjzGVkX2X7aZjLf86jDxD
MgTAZnMmL7Qnc3m/30fp6LlD2Ku5ykLwMZnVun4yGnSncOr+v9g2BNC59h5A77Kz86gVZpkgI1YW
jV+hasyTRncZWLNPpaU0cXhmne4zcUeXa5wvvwq/iztn+aIKpnM19x34jfS9Ixdl95Un+2Tq14f4
YvdbT2J2WO65K5u2lfDKO28YHebra8XUFS6c08b+NFwRhFKBnzN1lMcFIGKf35lPRD02A+ZGShSM
XsVCU+LarsLItkOa+2fkBrxP8WJK8gQtjaqKHQwH9DhbUZpOhjCdP3uHTDQNAUso/hV10nadS9zt
44v8pphK8HzsdlmN8OVH3bkZdDLFJRnkpJiIzR+Ppb0sBgS8oYEr4lRkToTeR/f2tz81DwwbVZpr
XV07WxnNS5Eah4v5d7HQLeNxXWOquWuM46HyfBlnaUZNbus4nxpjS75q/8UjXFnCI59k1yvlpA5w
Osuj8/nbjSUzfDRDoFCqM/qOxMy9kS9YbvQxB1xYGAVDHcuzp5WyHc98V7KCG7d6bgpbd5TFCjac
cgaYmEZdnmysCGR5kO9mqctQljB5oaecsEbCDOoXUu3gVV1sedTB2e8N1GSPNRPzHz/mRwKMRA/N
Yc2hedPcHiyWCfKsvl+piuCiF3YPMO5YZ7xoXtwC4XpFLdBdpCOyKgyH6aAUw68PPBHWQKJgq8l9
OZRAqruYjXSduixiaeeopzm5g2jzuLiMY1a4O8gSUkqRsNMFiD2QsYcaoljvs+WjHAvS4jYMlkrz
RcQB7Sn0MDwXN8neyai/k6BNl2sCQvI77nwK1xbL1hQXjzkAX9rL0iWh4oMFxa8NRPr4/WA5WW+C
bp62jARmGvbC7xJdn5GlbEUxBIZCV/Bp/4nCtdoJ8YpUAxi818sDH4YJMp7qRnxP+GWmrDyptZdt
CAG3zSFx6xv6/kG75cwwbBiI3JCdMy/zXXVDN6tjOLDfXD0Lta5lquAmYobGql1dtEpuSFPcVIub
f5RIDsZhokBBdgDkeG39oQ76D/4nWPF9WCSvaOQ97qrj9y/bm4JqLcQd+1vo0L7kiIrQvHKWeErF
sj1u4R06NgaPn3R1l6b0UOd3RpSuE6/aLf0OYv2KCHxYW3WWBWYnqjGrUUb8yQSFcf8pkCVctDNb
2PdP/ur8e4k//WGuXeGHjn3Izes41GOYntNc0kM0heOhdCUTXIoIr3WHNFwRnvcGrkepdRIH+ON/
z6t56fIyeCnoeC6MRUjJHESDAb4kKKVUAibIAtTxbggFH71sGuQVQTh1qQZTYgQOfVI1zdnJrfWS
Lt3Go0pT4tBYairDI8E4on/vV784iNTSIbEV8ZSOMH7CsdHf6m/aStZRfntof3s68x+WJEJJbgEK
/CY6REgPnU3V91b5giSqzFpLNY0SzEXLb4Iq2miV2uh7Z7zGali6B95/r6UonQF7tIWGOwCMFsir
7wX3qP39zvuKC+0aqbMkyDROFM65MyY6l4mCXXTVwpoFdrDMNFzQ07fcGxTMw9Jo7fdhgXEes8R6
S41LWcEN7NJVW41v63j/b9IQSodQoV4qOImkb4B6QO+0PeBVZuNPLElWIvkGlKEBK3fdpPeMnPhb
KXJxzSeOUG4KqXqBoK0xDDlLTYfqlF0vVn8YKu7gzd9i/tW33gFJDQStstRUv+K7Rw3As39O1kZe
+3mHfJFZaE5LFlsoHJsJm9bKf/nZH96wLMnyB5rpIA8inEOWFcXZppmLI2qk4X2D7Qrn7s4+MMfX
dv89BT7EcmUtzzJ9qQBcrNjMPYC+zcovKx0IS3LV7850IFqGkYsEXIlh9YpbYYk1vFjA/KKh7wNp
siQbR6Y/XkVKmUnc3sG8Ohy7XJUkCInFKSFY7rWk9br7MaC3M3WZqHfT7QnnUZQ/gsqCcJxiZxrc
A9FhvDh8auX4JYN3qp/SpBr6+/R9yiO9iy36ViWSbzz8C63Z2zTJPxM4Zqvnc3sYXqXoW9fZWqlZ
xcdePG3b7mPX2ed+8WX8eHFg9dcsimxa1/fpG1dv53WCa6m3MT9VU4dmNrDKa5H8fMAaxcxyhuhj
ZFbZlPKspirNRqjf/few03okZW+m2dmGv9BKnjp0RoGlz8eaGZOtukkzRBcwtdl6EMNWbHRqX9Jo
kMk7cgGx8q5vSVIJEkA9yyquKlahXS2A7hO02o5yaFNF076gY2JOyv4dZOv+81MqKxWSibHPexcn
kuEyEhEdZsjSkT5nyarZmutjy551CmluLDe7SQnYPp9hxrr/O8BP3K1ChDgLWwr5N6oO+aYlKK/W
qOOq2/t/qb6NN5/2Q3WAAsU9FPswtAIuJtUF957lhqZxzuGTlPjobVfF0I9uSJrHW943H6K8Ec9v
lVEMjOaEximLZaq8w0hBq/NBPKQkoeJOq856IDjXPTivFZoWFlF13ap3lwajC9IW4+wkYgfDCOIC
5MTo5qpp0YnvcHfLCb2IJ/Avk6PdeQxOncmUrMG3k6BFrPcQjGFH3H1wMmTDNlBv17xxHfVSiwTl
RKm1v/lHjp70poikKxrgufnDnp0EdPrsPczwo5B7CPYOE1uEdWkAQq7Q6ROHl5O5TaIwEIwgNBEh
htGaYEJqf8QofeD85Gs2ZtZHEXrGb23ZFjHn3UmEhEPkJMEejW2j8xs44t0nSzjhT3BoGmthaCmx
KURG0VKfh5rTq4Eh+RFzrHOubrtr2cqPwczJ81BIdHXRWk0yT3i4nRFhgneDDcBHY7PvLVA5rDIN
lRDqFloEiaMRXDrsLqGHiG4Z6BW4SlNsRW1N0bYB5wHgjfgqXq3Q0It0By03/wGxfxwcqxWwnTKm
9XL747bEybiOiHQB7DFsha8ja16J3lRCLSPkf3NHVgWdosJ3VrifK7FjZvXYJRkWX5aQ4cLogcY1
A1op3wXQyG3nbIGflIs75RbczENc7X9R+3qutSIFcABl1Jtqg1xMJ/r5adNSFRZfu4fnUaB4DsIh
AsXz9NZNQ9NwOq1hYEv2Qbkb4poXH+TiKQtDjk7qH899CE0Ty6Nw7/Nxe29X07M3QBuIrdQiyNzG
ODznAg2e+CIIZqrdtEtsMZHKkU96qB/0R3gCLtQ8LHBwMZhgAim5JDN2RO/Cw3ObvzAi48qnweEf
DvCQ5HbuNlLBqJCMEaLIsMiILPO/ng/pGlQKYaiZbuuazhmCdHJVcpgDxrfkjjECzrxGw5ecT7Bh
NgmkNdV5Ieh6XnI0/f6d7rvCotFPXhTTyc4Pr14GvWj9DSTxpz9vLnxDJsWrqCjX54kzfECzVnMT
yrh1Nf6bo7ccuO1RKxCfUZwqGGELC8HE4sBxXrdlSL9CGlrgG+FIyBvCBrsa/boNheAtdNFcSunY
HWlpH3BzhfR+Z8jJNp0c355yTMjVYBj/b34z6WNw+okFGZwB8WU2LsiuQUiJBj5oTySw7KsWXZIW
I5XyQtI0Ou565QuElvGPDu/OMqU+fHNYF3XW4B+LhQ8RwIEIFFw+NDPsefrFVo9KyIefe1HgK1TL
Ba6z3Cbinyx/OrXXRbpPVyHYXmNJENmvorxKDakmvScd1W1Nn4Yu1WQ/O/xwpTZmeGF5rA68Z0rQ
r4UK3LXI2R2qcImmneyihY6GouoMXA2mi7GbiZTT0mtJ3UFTseX4Urjz4CyMwiG20h4YkCN2OeQf
MnVyHCYccePriAbHDFEOWbyqXdqixWt7OaB5jhRXV9xhWJSe971b1GYVXKNsMbzcWFr8DR8rtTF3
3DKu1GCwm1KO8U0DhDGSKKGynkiF+OQ/UHop0ByHYoqldrLUNZ3bC2SAW5gVE/bUh9yCh6I4TLNy
mdFCekJJ2YkdaOn0KLttbQmQYEvGwAcpls/HdajhsjzPa9fkgsWdPWnaW+aqHF7Q22pxR42xe6o7
7z3FLtgaDIDMUQBHpAM7K2YsBBHOZIylL7dKpMHdSCtTn1mKMXh237N4zXGg86k61XIJPFyELv7r
sRTgImsBg6AmgJCSyprVqyYHw6vb452XKpstVuOEYVZ8HQk3OTMuAY4ZwlYs+9pCWXGh3Rw+JKMW
wywvRx/FovvzZcqMh7i4oZU0GT6I1FCUVi4R7Sh+yWy/ba5EvjL7pWCioX8bfTc/MgfTNSqfgV5l
Gb/p0vspX1dWcxVIWILSzDaFlxC8Y2ss/2e+L0v1wQjk+y/wd+d+TQmagJsUbEyeZV75kE1+SjWg
rHHeuIz78+h6Ht14615UdkR/DJi7jAMlTg/8eOEwyr5xacbZk7iav56I/gJDJb90hEz8Cz0xpuwN
KMeXXzNCM+yYssBe8ihXziHRQXbXeB5cgwTXYofyNEwfTb1gbFqtCSLQfgGWBWl74LM9RY3dAvLb
zBXEsrZxC5ngmuNFcgYg1QfB6sPQRSTDfMTihL1u2/yxcXw5GzWXmYkpqNjppbNbjcSa5AlGZBm+
Xa6DXytTJrDiAfyY4CfZEP3OcEs0m7GHbQwfk3ZXzZ2sDIpl7RB5QrRf79nn46VsDIB7vX00LuYu
DsTrbFqPI3rWNKXmuSJdGKjfEnv8vQjq0YlazTx+Fi+ddu+8N5FmH0fbkY34nzrP5pGOYCtgnuYo
nVUZYCErFuAIKK3aD0zZKNxmeSZxNdDXn8xvDYFxu+x/94HxwFk/EfQN537UYwpM6wLyN/j2Qhro
VjDl3skAP0d5czDsBiqbiCIFXYCewsfgmtIJ/Ic6vnrKP/jYwQ4933+lpOpyVEn3irF+xcgzBa00
kwVkwE17qce8iSKLg7wEeRsB1/+W2Rne/2IZNK7jO8K46l/FCVAT/v3p60QOanBVFcfxczhFxhxZ
URoWIgZxIhBPmlhaVOzYa9OW0gzLPRWHwd7Uie1F5P7YpT8fUfX3EW2WOfdIHrtaaeRqTNL0Ygdj
aPWMoo+TDCG5wfeSbzALkuTZ/qurobLB4QJbHRTE3E9JWYQNRt1TZf4xhRjgv9gl6Dwe+q8ZyTvg
tSM/a2dtyKL7qFGAXyzlstqqkuO1uA6uicABySSkYLFSDiox39Bn41Eg+DAGmXcUqRyEcu3KbuEj
q3WB8ueBV6klr6J7Bm2QV8QpQ6AsWN8ndvHzjK/cH8h5Dsw5aoVas0AXXVLQD2NmqR95RKkb1LQZ
atqLt+SmgcePt/1Cw/Jj9aZ81DO/xkfDICtkSen+IH+qAnv9USVWqY3CXliH8oT3sOHGTxH3PHEL
JGzu8tJNAAD5eJTAE5F9TykW2ml7LgKKJ0kzzN+c5Rp1ip+1mFRKTW0RT+zSbrY7Rbpz0hK4N+Bp
fOM2tyOVSaH9XS9SaSKNp++ambZQNPKbBcx5MOwIVeNQ2636NojzvjjWXEGAOZbarPyrWopkomdf
ObdBxHltArGd8ajxfjPcJQbUEZgYCKrFhH4MCvPC/oVabLq6kFoFN2svar6uCj3RIppN2rkdhvkx
Nm3d56wTaxivEe99w3q2aBqDZtYRFt0EMS0VqVCotn6+qeGWOKp7KEBzBsAZyDvHe2bB/I4GhKMP
jX5+XJl1Y8CePF3f/Jf0eiod7U4lE8F9NEsMxJ+LnEDGyXgbnyn57ie1N+TobLKQXzKMXP6rAvwL
/i745+QLfCo071zipYp6sFarKzeMudalLJUu0FdF6c4F/QmI2cVLJcY66SX8G3rdneBLB+AJhrZz
udEDTZLdZCeeGwMF4Zl+MzFLnGUTr5lCGQTPuaBfzs14XnH5KUug//PH3U4GHVcnR1LS4C8doKdH
6Kv8EvqbU6B4GtDy7unL6Fa0fYVqKbbbZtoSu8AJ5JFEC+1TLr7jSup/MGCgruO+IGJRADWs5Ezf
N+ErSlgptyNVb+bza+F5szXsH8HoU5+Q5Z55B0znlSFFe3zGmKwKeEqqmgc3+W9d48vcUZr1NPA8
qZlSKhvdRxYwN67PeRkJ+rkJI2S8ZDjcwjEuGg9dTfRhgzb8DlgYxRcALlS33nuNhAQGqRuBwF76
K7bIyRd/H5alRkNr9tF3c4B36YhP5lMwT8dNTehhL2LTmnYDuUF7CC5sZ1sbx7esPxYk/yTPeFXr
G/7GjzYwZpaek7Ga+fjcOV666sIDZDdVOfQAu/1nnA/7ZYukS2x/H9GnqdM99McloRjH3CzXmaO3
N7k2++sa81qt9gvnI0UbBJlhreBSuoVdVlmfSzo23mZg0rXdKJOspSUiMOSl1F9uY9bHfZg0/dpZ
EnTwxdC9VO7QVC/VwNKyF7Hwx27MtK0UdEgZBjAwVpRQ7xxmyYXhlNaZk/SeSjhz3trCGFXocCBG
RhYpi2bDc5F/MTg8g7SxgKfYHqP9+6zQAc9pSfxUgY4Jvkf0XjOCYxSL05ZrtoOmXMP2lwmP5GPt
noXMQHQb+D+NwOEBUmcAqRB4rL2pysKnlogU3XjHS3AOHafKxyYv5WnW+S7HdOCfYgQvLoxWHQgQ
3EE0scfBUmm88hMREwMQlzBd/ok4GspuyuiuWT2qKpfqqoOIZpUlkmSccGTbaYyTWuZRpx5C85hd
tTBbKl9Yyf47G2ADPCpQTqNStewwOQH4vOCSzp6op7ay0f9GvfVjPlab1UIzP/IOY3zA0kbaSqYc
JtRA8vH93jdSSQzZL3KPeaJjItk+HPXz4rhv8moXrGnPOZ10nAmwMmET5rRcYDxptkv02jDlXp4I
SsXa/DSeUci7JAzlKVstbqFH/3XQ6rCojs8E6ept65folo+fk6jF8LhWVd7Wq3jN9FmnnJBW8cVB
1z54e2fK4Y1O1vQjGWmxYW3LTpk0ocT0M16eleHjK2FrYkb0/edZBWTO6fr8Be6OqLKzvLgB5tAP
LMLRj7UbJQmCYIJagNBVrEU8JhCKNPme0zchzb1Bkg5eQb6Cq9m9jSHig6dQRZL5QoRj9AyjBu72
JDUoWJ8wBIQlrvopN/he/XT+Ja0A0vx2rZ5KIywa7D7BKJGN7OeXvVWzAiG6mlu7Wb1yHCDqMRF3
zM9sdgki8/D/WVQw+Ym5J3wIAgJcFef9lwrojTLxaLieuckwIlGVabD8GKiewvl6N2BS4AQpC1QW
Fod+xIZs2GmkQ83pVvyjY3yHEWoaIT6FecePm1XF65uiilYTLONyqrjDumztuqeYAjTcia84RnGG
CiokCzSQfvO6MrAVaaa1UbQ+mmYY+QnNVINJbAbavWwjVvqIXMPDnqXz/rxXbsfUoWavJeLG/CN5
z5kxkawDkT7ziEb+U+GPt31PmuVAlr+eeB/tZmDHSEYwaTu4L/D/2JgI2QV5gtsWuT6tWDWgtMu0
Et2k9H7Z5I3uclAqD4oxth6L/nOCciwXzsReTRjpoXF9jmCeSCiKHau8x73124UhTfZtNLlQuta1
kslVf92dwNJwrXIg31QAP/TmqFQTJioULPxEa79NRMDNFQ0XCBfVsXLN2t1kSEIpNlxPfVKowVLN
nkapSW/C5Q+yofNpdgEKYhABPWbWch6ROQqIgrfULUqy+0kH4t+Sv/CCHZUWsmnPGfnHI3xoGkU5
VKmuXQIFi0PGF+qmEpzprA5MhBW28v0I8kz53mG5LVMy+bdX4Syq9IUbADQn5JckU+FCsd+kfmTv
qq7SiiQnYvwZg7Bi6xEvsBkjrP3E35DtqiO9B4uCtUq6jHrOQa2cyohzpzVBkV8HepwaU/Jg1mvr
Gnm5xYkAC1V1wfgSjfEKWFlVujoELNyT1b4W5T/kqExEWbfycXRhxfjN/PLLv1DynROImsFLXEA+
Z25PH3H0JBL6hUjhDfDTI3M6PjlEiZHB1lQjUXOy7+Rb5skNVdLPkeVw4Ab4AcZqnd4bnNMOCzlL
598wf9OpoGuVw7mK4caBA59gFnmf3orVxEvHNzVCUk8VFLWkudX3/7Yv0GkNBy/vpC4j/PQFdObQ
4Gor2tgdCSv57qKKKkjmkN1mOoGp/4F8OT4wELbDB9Ew8G/GF3v9Eo9wFUK7XtisoaQRXVy4gdSW
ZQJ5MU54meFdH2PPa0WQ1od/wbYy/gmvnlMBaGwKzprKqGcB3B9uzhAB0Z2jK7j/f5WA7oBYc6XM
lN6+9Mdf7fLhMboqSp6hwOiybtghjLrS8kuzmnfGZ0F1HOPXxWV1Zb1sdafgQFMhOoBX6WtoT16l
PCBILJ8tdQ6cuEwoR3PYLYT+5h1KZDDkwz7KZWkEhibxGY8ww7pE7PrkqszLRox3lQt0lWkghRYa
9Us5Jsb+nU52AxIWb/ZpdT9lVGGTekX6SCPO97XAujo0Jd4oqrVKbC3xKfnB/RXovuuoLSBa5OxC
8zHVY6TElTGcTng8eyZEvR3tsNfPRLQTDeX6oGUp3rjRE6DdNAVs+cJjE+L1dAE97mV5OHkVIO2Y
tUYlYGbZHh/coC+lzGB2wNnVZ64D+yXJvBF8RddE2sC+EbzrYf53MEbZSUh09Z+/NFkRfdx5Qmrj
CUFcalqMMQc4YUb1cmkOziZSRqHROK3X5XeHhwqppArxoajUy4n5+62n+z+L0KmYE2i8y7CkjYxP
DauF4CWiw2gIZpD1R39Uh0UlM0DPkRIWDiad7xY4RNV0M3LGQ82xkPXfA3C/fJSOk54zHiWvyEdt
kR+IhJD9IhES63ZkltzuiP53OKnBIE33l1EIBSWT3TAcdaMxRG02znBLgA56+oqvcakhJao/rMSm
1XdW3uXWPLdo1r2PJwukOMdouf3/HRWEc16tCelji5WmoSbQx25Ny94wsX5aqqkkgyqsiOdHW14/
4IlPviGyFuFsfoI/I1EMpQtrOE0nHW+osgRvzUjFC4Niw+bxm7Ov1N39U9BmwikKyo5U2ho/+qCr
QyAS0Cp4pIRjb+osU/zdf5wbEApfeGsdC7DO6UJP7RjV7ZAGZLMeFPoqgJErMZ9D3v7rWO4O/zeJ
HPjp3u2fjl8d6DxYu+MngIeEZNYCZRtGnpPP3IH7HItsKytl4ootCbI2eVpw+JhZXpN6X9Ep08eJ
VRKO9dbwkl5XbMlCHtqOL7yeG1CWT8m9vlgekTC4MJORIhKQfFXdEs9XWzwZjQK5LldwKk7CL6PR
ivMR5ZLVnWDjKtszsjByzEHErGxY1fcCz2fjRaVQPwlpHyC1ovWaF1D6bx73vPfhUCOeetzUSgrt
uA4VGEiRV1FU3e8QlIT116kyfSOuJoNHrDtzZviOTGq3UvfyaI5PpbPZoA9s
`protect end_protected
