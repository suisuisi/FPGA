`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SxRiU5m3pRlAj5USwN3/QbFDi4wilQqKO5HiDmatjeskQ3ASrppIMNzHebfOzJXggUkFx2grguxg
0sk56Y3shA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tDykn+grM71Uu6e/yG446Uw+MIRlJpkLtrdfnM0lIGJvwYwUGUBRWRjR0Fu97VJ+XtFbbcajOR1F
lMkALcaxLV0AJvU4rDGEtsfpfTdT7VxwqIAsu5TJjPXAu/htb8eQfs+L2dJYQukKr/VfSAEZp1fq
HdKV8mXQOAmRFXzIdaI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XAJbIXtfmqQCbpKYtCW5y3044wa2G2Ol6okqYj/SRYk1KN7apSKLZZSMWgXZUUlXrFflPIkF7lRu
1v5Xa+TpaHKQKZNyYXYy8PMlIxegoXYfTxv5GRiQBfUxo23CZk7xa/RfSmeyZgiaLZDm2bNRBNjE
xRmDHy25FHPLhoeUjWxVOUZHeMh0c8QrT53gWUXgWwarZBBb5fPX4v6KmuswMd7smsszZ86fSMmw
9fpgt/uwoGhjYzGKA+sDbJRW4iAlsPpN2MkNoWqC5s/fs3SHuDrhOQoZZHAQVXH4EoZ5GXUt/sWT
4dQdV/imVmQUDzY3by9kI2fbQd0/0Tj0Hy0QCw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QzCn8QEWZVTrUxxYiyrjKl9zw1wjN4NR+bv5bJ/BmvCr+Yy2iFWkJ5OekWoGNLnaIHOsJ9mHrA3E
j10hKtlDyY0gUWjeck2k/i3uD7Q6EvwCDdedv5VajCQApRsGUvEzhPfLN2wn6qW+1Mt3v5vTQe9j
VXMQ6PiUlzQqUzbHv2n9ttmq9eYBjCyU5Wo6Z2Jp7XOttnPsuhrH3x/nFDjMUVu+oGPfey1UYL/v
apD7IFJJZAMCQgytTBubteBbnIKi6mxZ7AVJW2BEBTnB3b3c68Fmz9/tbV6vud0eVVrzNFTd9v0s
nR7t4H1hYDIHryA0jk4FIV42ljvHmOI3QKGctg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GLcP/n4mWm1qYeOuuTpKAvi4/zAHcTZGJJZtPGPLpHlb4H2Bioti95h0M/sj/LEI9YHkywLDirrv
+rwuj04PZNmYNaRw0ceYbooM1yCfoWE081jVo/jtkzz9t2B8R/nVZYVN2G5ZJxMO7zjHmsyr2iAA
qz1yLpRPJcK7kkMgUVI62SArjenSFzyEpGnlliJ4CRvMBqbmAlCZpjzQb68CdhrkHx9bzUBRf969
2U7g4qtxK29js0QycuSrvObcQTfL3Wy+gjogTH8tgpZlDuabJeT8rD1bL6qsNYPh1T6QtcdEMMyr
LiLak/fN0x9buXBwajOt32bP594Ve+MyhF4SHg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
s/CgA8pmJooH2onxypWzsGR+ZsBvu4lPjfkQ6fYr9Cx1Xiu62IFhsI6UXMTcIt1hmydVGFt4Ke/P
2A+RdI0QInW9Oq9cNlDI3bq6ay4E8GTMp4MdhRV7hKUQf160W1hmo4oUoXe6zb3te133scTO9RqA
8InhaH8k3Cngy7l8/Uw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LUmj+7O7n525DnQi1mE9ra5fU1tGjqZxtrERBm8GCTMCWk88CKw3dDxwo0NpBIE2dnr/Qe9MUCOh
BqyaZF2Y0ZZqWv11A0huWoJ8aDGdbRty9sLwm0SiUJhgykOmmqxNDfK9+aXGIoyXz8NwLyRpRseJ
YVnuwwaTNC6ePvQDZqt+Nz460+FWex1A5GjCYiq0uqIbAbae+HPTNJtbYIpIGYy0xzYDubwaPpgk
vABhPZqH19XWfTwJr6uQvu69if8+6rs6fvmty0RdVkIgebxdGIuJk8vla33HfNkzIMMT3QOgJf6D
abLkC2J98bSHIi9DwqIqLbiX26O+uAJpwdUiAg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
YG9f56rCLqVBn19yhVHwuk2ifXtp3n98/y4arE4UR9aSfHOdYTbqcfLsCwfx3c2GjHzefaFIPEUP
ABlXbC8OTOq8EIPHhF6STcVFm8A51Zq77XI6pJEoBlpdQ+5Z2K6GOQp3Q+XSH7m1FauR9+GHxfaB
ijoBQSUnrIhl4kMDHTTO/xYVCdPPd4CJcYcasMP3yhuSGCxxhs8SM76ulb0q9OEK3MTUQdgxn8vB
gZikgHcTqLf9sTjY6zBXv+BRDyy9y6JjWB1wPHvip6cxliXh38b1VX6Y08q4TYxVLvbV3IYOUS6W
CFE/cJM2QcM+CP1XJ+PjDObYvc/UGKjnFipfkUiRdJoAuZAXdOdsWK5oe5x1Ovvf/oG9H6hMSVOn
b2IAOhRsLa4yDkPQcrkAWdw1/EE82rNYNpjo04SCnVAifZBgRJ8AZm6NI0OUjfsJFzHkckvMrHGq
h+TxYUSLQ1IUFMMYddzeb7hXhOCSAoui2n7fbuVj0xkcBvd9wRBT0KqKQJR4Kfvc+q68Sg2UiUu6
HrNrPh8wG63LwwVfzKrbT7eP6Tgn7zG+vhK/JH8Ag6cBidvdzv2Pj7a3zfEiPTdKumPTCjuzdACm
BuT8wt+iQRR2373e05T51NBKip80Or7hVZM2RJAWWpxK+NKcaXJnhQ28PQ9oKCCXLDt+b1tZYy9X
eGAIqqqCRw4j0NieIj1gltRl3REAhj7v81kaA6sMRw2U0CObufe2RRRYJy5lyGrVnire8EIabYRD
Ujw6XQdOx28C+mvcB4EEMgHANc4BpotkxQA9APAnxjD/LqydoyWDpTO6ttdOSElj4t7TTxB+AfgC
WO2UbPN1fDBIHhg2ktJYtVu7y4fkDps4Dm1NY1DRcOmjYKjsRgXpO5Q2MZSUciOEsXZ3/Qdwl0YC
fKo3OkqYQYMcLk5EixAlz7tdVQAOSz/waPULTHS0rvE1idSzpKOruKJLknpVsn/TYoxDrkbwbX1Q
OWw7GAq4oPrGCvM2XwEOYNOEUw0SI4NDpDw58FV+oWoVY44DEdqKsoGSVgcYGLx3AwZ2WZcOd8Nx
B0508QvZCuvs2xmx5Kj34I3cQyiTQlRHccAbhrbRUoCKCiOYwWyDo6VnP/30sFY5ZXR4+DuOSkBr
5T3VImFRFu1xtCupntlse/Ck/2LnFDzkjEgMMpO+SKXlaKCzOk+LPo7KEAfJ2oWsAzzbWqbk9owJ
n8BdGKqjdu/pihuN05EOJyyTnE72Jj1AKXjajJNZBgfZBifbb/uVvNwkuUXvylDLeV+GI9bCQG0C
8Bs19KPSdZS7V541TX0E9tuTyq+gNTgo3EVubUVg2DOUW14BZb71lYFl9XQ1flNMnlvRmpg7j09g
5uinl9NdVvGrS3ccnYT6Rl0GaGe2B4Y/qFPFRRyn1XiXgE88OnnnNqTtexNOI81caUdx1zM+6Iw1
SKcc5XL7OAcsXGnYvzVgmFHjByUZfVRt7l2ooKMCUq3HruIR6emvfVsfcyDRX2rpLc5nXrOume2k
xO7jpIdYqv/i3lYard6tNRXwe+MClhWezBLdzichL7ZrL7DLjn4OIlvtYQA0o6HV+WykVgXSPv0G
+523PwwtSmrQXzYptwbXawES86N4fYQVjjuTTC9iw/6j/V5fVlpaVo01WV/nOcWukElN71UBunYA
1Uk6/HDikI1dAPjWJL7sHaVPF6jqUwYnccBPcU5/8oXHLRn+ntcj8rP6nH8FpBIoJQZLIskSo18t
OkU7UcOAN3CAKWA/tpUryWDQaRu15e//f6751seNSdH0mm4hPgYl/QKQbVUzklJLd5czWiMdDMOS
sUJrfrkctYELfxtQ5JQmTKye0qbkvNWGkE08w8MsQmoAOEYYCxqcKdzSorLmZUidf8skD5maW3/L
Uxlh4nTCBXdriMfIJhTv++eKlH/ylGJ0HpkgadG9Ur6q26Dk22RSoZYbp8d2o4VNjT3LL19O1yjf
3Y4NWP2j4Sh4BubmClWWUJ3PqyiFUaBFjoDP8UTS9IKRMcu3bbiy6V2BiC63ZbK4KVJQbec9dmg3
RGUqiIjeFI7pZcTRZDqAZYCBJi6E2ZKj6I1WGrOzEpC6hFPQ6o4d1Co+4oVvIgm1oBUzmz/Hhkh6
1YP81dtPK6T8UtbriA1ft2qcsTK6mDN7VMFg9krR8zuKPP6Bdoi1KWYD9OsrileBDt7Dl+5pgReE
2A4i/ycsTZfLXQfoJJ+g4z2EWQO8T08E8aclKpS86zk/TdmrCO7v32sp2DZtysxp8iq+sZvj4kYq
NdkwBHXEU60+sIVZ+awnYtqAMr4jPPjRI9HRfiZawAarIl2SkV9pnSAVS4CVhZdYZeg8YG670bUb
kVrhWuGaVFJF4Eu7h9IjvrugjnP/FoyVibXCdCe/5TvMCePbny2KEJKUpeEsNs6VK548+t5QfjMX
PNpgMu6nIlogIuqeqOm7SvFSBtsY+ykGDOciVqaxwJux2obcm26TQAdkP3QTN4wbmYqvN0TwQ29v
Rq8uWNplxx6UM0bRGpiEmNA88joiNM32N6APXMxCL5ZakNp2WfJYA71AUiVromMWAqAsn2O2HWzm
30zoYqW/UhN8yFNZ3+cSofOHXlSI/KPpUqoR04eXWQZjkygETnigIT1U2FuvFDvBU3/w91wGZK3S
8DhgCYGUxp7ejz2sw57ka1UBeqpdWcKiY+930zwVIfEa3ypHUcrEtvqDf2DGwU+TLhdaStg2VuHC
CfYjx1v3gi8/TpW7hPNbQy/W5F6Yg4szr+QaIj65pUuJFIb3dyMtpQP/TDaaTU7oALJilf43VXmi
LQ4YQb2t7PGkwjYXjOpS1G4MNvtngC5oHfRTaxHERU6puy5wx94GafWoP9Z5a07Tbv4irc3ZHPss
YGtM9pv1HZ5JhRTcJ5ApefqXS2xOe/OPcwETfwjmZjCyLBV4COvmV1hvkcKrVVJAxCfGaseymUxy
dQly3IsInMrTnEnYF9bz8rqQ/UMVQ+HD8IL+1+jsy1qs68/Jl6NoYkfsXbkPmdShn5ZhwBc9GGAJ
TZbnhKM1jhtp/BFY2YjDef4owQzDxbOYJNAFOWGExzMgYO+n7CGCBffbQw5pE9J2eSBZjJz/qtrz
DDbGU/9QzDKwIqIUxmMCAtIOaWkeNaI5lsGOmHMhdYguVtYeiJLyfEUhMkcLS0NVXF8KfKz5mpcG
Ln6ock2Dwqqh2cyuLskKMUpWMthgqc00KvFKOCs0uatQewyijidD0vpz3ELK9zth8s9/ajgWzfdC
3VYHIpxCZOTeH3nYW54EAKkJ1TNYQzqYo7ov5SLqRTosNoCd0T2UGzliIU7AGqACjfNuSSasDZ/y
+OvIi1C7WKvuc/p47iioR9Da2esEJlBfoATm8bzM76nAvynpgte+KbHeXu3enn6O8UQnWd7NraFy
zDHMApsU6TKHIK8iOwh5v8aLpMcSTqyAd5mB2oM1kOJTR1Bmrpbr2MW8ZiWN7dPB7an/H9mIWNQT
ipiwwO8WhfFSz4uscH03QxZMXkpzwuljN+LICRuNsgeGn4Wd8TpuyB7JyHVEkR3b8ZVvrXH+Kx30
5sxNbpCjBZF0ndLtcL4KkDfZW5DbmJC2qOwPazhAG3M+cBCT7BLNxvpr+0FyPAFcF6QyvGLwwvDg
0aXy0c83MW2euPD3iXMgM3J22BI5QOdP/hoevvCDuBD+RODt1my2FfWm93kHLUM+4oK8DGRKLQly
7JE93qiaak1DQFc1LVCZsc801BB+FtULNMYtiu5TpVsJair/nnYBzX2DrATm2WqV4K074oHdxVd2
oICyihwtJNB+uSm/RzIYM7qE+FMyjAG/jzVa0RTXN+lCIgDJ1sDPU7nKA3MsjixDxXVEQ2/t/qfr
JqpdLz5Oi527e5W7Kygm+hd8hWDfLO+GRas83hZAXCHy+F+YgZPIm4RlxA4ONIab5SeuxgAVS5wM
NMlV8IXgD8RBGmmf9KZmJFoJ1XEqvu2KRaJs4YIUvrK7E1YRUBuGwDM3XGJ4h/8R+q5GfOlF4Tur
fDZvzXLK55xSsVdJGgb6tXhoAAgXFPFhEG6nbo7TzlHuXlurY6T+J+dqauZhTQ61Oyy5/7LcZY9T
DtPa8ox0dYL5hP5T+tW5dvlDHG74ub+xKOJSfcid/5kZ263zNhe8LtFwsmj83Fr4Ipye2/b2OHxd
ULFdV7uvSXO3PcnsbUMjEZS0bAGpPVgn5EQzJfuIQBJ+HNOX42wsAzSZeWACFxi4YqcRJDK3+D3K
Vz98i8rDRWjL2GbpETTfMsgCEuxb1gNZ3JbGr0yaX3Hvdbilftux1L5o1L892EykOGYdH0QhSxPJ
F/35kfWh83B5R3P5vKly7o8wwZtZplf1uuddI5YClj6majWnBynmIn3G0Vb/NgeeqjLqxd0kzsEm
3CYrRtNQCzCxcCDpfuyJFfUiBbXizRcMMW3JZMIAPWwSeLNgUwO0P3KYCVC7EAquLlhqbFoQDvqH
AVwlwvvOlEuISd+uO+Ryld/N9317cAOiSyufwCI8wZJC0muxZq5IepMz1F9SSCSJvu/JDysRGRvp
AiL16IFZH+2i9zs4tgTAAj1LZnn6gMn2QIBfLCPsE3ESTH0NkyCSZDbeaJ/ndqHmG3x1SMnZrm6g
GfyuO/fYULzjjxmB6T97VPDdNn4E2TLjotWz7GgwOlOwjkkMfh5qzl7qeEfHS/W5dvuRgqr7L+qQ
abRURFMPjREISeLSb2Qk0t7V6jVN5eXjMUpvQo12TRTUKonLgf/0KXXF0VUNxWrWfJ1//U25z5YS
OqLgRqXmQfXtY17owoUoVIwqzN4ziZ/m/lcEG2GExi1dphgtUmVaud8H7YVAY/AMdKtbao3JYiKr
3Tv0MxSQ3BXEmKsu8rTxryVXWOpxnKBpHBXrzWC3zcgrHx6SyFRNRvaK2RZxP8TV9Ub1NrPPrQO0
3cYT/D+md4gOl16TIzO5Po8EFMBkhZKmuVincdMQ9A+u9bBfcxvdUfEuyxUhzhfS8MHEazdYZK9x
C9AlW9HlLMlIwpwd1elT+5e9nlsl2xpK+GzHpW4C0ClQipxQ6k3/VCyZpHUTKQ3ojdpUfpzuVtFk
p5SjjWHfjmyRYjV+t4vvv36nuzeRlF3N5xLFfcGitTmCosSsZuH/ejovCgmMKLeDRx7zERr8ThH4
li5mecVDJzr97G0OL+vpY1IIUuxx4t0T9lGIEmf5+cZuJuV+HSDjnlXf2Tq25V1IwtpAJQ66IJtR
ckkT+T6/O7QNQhRruOBUnjhFUK4ThEXRpNG+YgXgs+MHJPEZ4/5kUXnmH7ryHXckI4zkqH92974a
uiV15wkciTSbtPqyHS2riI9FK1RfiyRiEbutOHay3c29JhBJqwNPLvyCBRbUKvsMHTI6YqL7Phhi
RMLnBa2bspxP0uxDZaKm4hEJ2fFRFIbIFFb4p3XfCnQYg/qp97eZ/XmCnrYbixB5cIB1119oWisd
hp58rqK1BkwE0eXB0GV970wY8CCwxWchfCzjmegYdL7YuXfp9WvRoZC1i1Epe9VsDFG93WpYA/hp
mMv5tMotnF3SHbhqBZ8rWcvPCXmngojhlCtbZOoMoIwQgjLt4TCEEeHJgnzHzybSH5zt6WZhKzhY
nh6qvg9WBOqVS7K413r9vnyM3gvdq0BVgiDRiPHZIHJZN/IBAmPlmL1gTGVNRiaDhKngHHqd555k
eeNhWyr+SktfgHicl/1t3vCnbmAtFEqfLHrB/pMYpxubOriD50tqMjkMvEeWjmTbKL7KA9tXgxPM
kF3gMulNQj/Aak/q6JiNrghKgitwFOQcvaKyG2iIVYm9PmILMY9jw777n4STzbfKF+6YEYc5lfeC
vH9ocVNTdWFwp70VTJBu5qqIi4+pPAmOAAunX7nwSPjHuF6LqO7eUTEP92/bSXd1sbNfOaI7CvgO
97rGzBUbpE/sYuHlcYRIzQ7gbyd1xlCXCcU6If+d9h7TMGMIJDx6crZ77vM2V2vVUUs5XPX8FDTk
W7i6i0IXlU2+BkHG9W+iQq3K2aoujN9xYUZ0gEGutwMHnIcG7lA/rEpOIyQO7Pe9tZGo8JnvDOXG
hLNS9SVyYBEI3TKqwCjkmGzob2Gj9AfF+yqmwjp76rokn64It+/+NkQ85z/eqbytADoQjJTEuAsU
nwAx9IFJACeLLNjUp+hpP4l27DzPHKxuHsKayj6CMCWKGCoPKlCLCkt5WhOzHiFUj2kdV4o8FtL/
HotkbFPJYSVOjKYiW3z7Q7fNhzosrcS/M/lsMDMYVPnMKwM3kARRJ8OdrvamhdaiZpbaGVnwSqJy
4Jf93pbxki+jKS+KnOJBA2WME0HbOAAIr1jq+VJG3tIPkRvmLAncwZCYyS+qEUzO9D5GGvtFn4XZ
ME5lloQFD+/ScJ6VhRLwCX38swS4tA31cYeWVBwBv04O6RVSpSiOsD9NKTMmXaKHtN02JWdJswDN
krnzp8hlJclPBht6NCPZGsbYbbCuv3tjK4WoJmIUVqwNcT1Tre0WbCuNUuhAzKqNYd1izN5PTOa8
qp4Nf+Zf9Re7eBQYGvL3P9mgmPl2gIbrp4b9mTXuPwN/C4223uF/o2R9NlEJB5HjuaiQM+F/VsBA
6B0X7mJgUgRodS4xS9WSriAiieAnOb/6Ra2uobDLFwTXk2QvkGcLtPFN+QvGxG5dVqqt18sMgnF6
xoFGlM+74vIcVpSRhJPtCSYcAlk1L9Ej1bTHePgDkrQ56apgNI9lVWU3/3Y6PcLN22JKPcp8Aisv
UiTMokp7eC40fFwdbTn4R0+Y326FIYPu9w8KWC+982oNM98dIlh/JvAkqn2OVl0cMYhb9SpXfwBH
9vg1UGnvqapklLVCy7r+avCtib/6ExvvVPNAfwz/FI9ViMHSGkM6qsto3nC81TnbQPbOzd5XbGuG
S7h7MUd8am8cTAQfx1hrSppA/CC42FU310TPkeBcZRR6tAIXgGNSZpmB1ZVAO+lHjwA2lKpWQqxH
UCjsZHKj/Bh2gLHZAmeJJJl/4TUJ0m2r/W8KypGYWDze+DSWrASf4uNFxIO9wbEwmfJaxG79MnbQ
pK4p13jZLA8bwrQkfw71wzivM/4H6kThqWMtxgez4che3BSiOcWOEwSV7In9bexe4NSbHbj0xxJr
KvoPaSSpNfhq5p3zq8E881wCjbnmDFBRthmIlyRR2aFZb+Y3AgAwupW5DluV/U+i2ps55AYqmdFv
mTtB6hFja7gwI6qRWdNIbb5uyqu4gAiTpZngt3w5eCkAArN80UMwNRjtFiUbR5uwB6hTkbV3/rPJ
hHM9B5iB9rCdwEAKmiboKd5XeUI15/X0b2see24Kbu1bwUl5f2PzDkV0Lo5NwkPlKBYoYC4DjJF3
ilOZ2tdL3K5rvSjC42z/RXVZ4rWXDOrp58dFm3vp0he/Em+wSoXflnXhhCEAZTgHH+p23VfDuKIL
C2eOw2Kd03pbyZO4xakHcM2DSzfBEH0OQ1RwRtygBgIME/pBioHz3NlpHywo8E1B8taiwf219LNS
Out67uwLb73xEORNM0fOrKqr/87TIkBKrrNQKE0OluiTRC7s5nD4RyB2b9yx5izdWH2ZrA1ZRHO+
BgVe2nYt66LUetXf9/3XB4UpbNZLnOm9v+MzQxq0MKmPwNE0svsTTJF5/s9+LPHZ1HeLwkCxoIeF
zWR4XWFqWPReRlL7Wkj8R+1dh+SIxgz1tZgco6ypfX8clscjn/a3BOrpYRzOjbZmvhwW1dVJ1Khz
0n9lrR8aTz8QdlcUn04BPeIQPeCAXMMfkRr0SZCYK2hIrq20S+G261TEK2GOKb+CHA19JoFUgnvj
ph714uRWj1pqc0DEapyVZvjNOFhE6Ihb6g1wQwj2F6g6p1JijYoTaU0mrwkK9F3iDFw02piOLbjt
5JrvtY2I0Dy7anvsCOeyFHy5kKz0YsGnsg3pyxlfFO8yIUES5AUyvmY7a1S05XwvX6COODhUPxsC
LleOzERVHK4J/c1TUiCO9eNtR4rgFYctpaVHE7CdTZp4RT2IRDjUyC7shr5hUt/EH+xdVEEupMNX
kqbNi27VBj01jFADiT8WFezO9ucUFlV9fGDPMVEyBUmFKH5qJHa9BtEoxAAGs3lg6MrQZRKF3Bdo
iEOQGGg/BBiVCheR5Sz2oCjvoxcuxVjdQB1ipxJNWu89A6rw1EekhMXqgWb6jj6U/UqHd53i7PYW
/WP++3rw/zj/qksG3ZYrJMD+r1wpJdqegfsHS1BJ+yoNk6C/8URfLZ8iyfj3f3iy0a74sI6hu2p3
NWD+WOBhgoondZ4k0GfBIyP4/4gG9wbbDvN4LJe/4cwp9t4OobcwlT5lvVP1V5dykKcRt3p95HSI
OBkyaCOXzngq27e9+HNRgNye9Wg1G94fdSgraEWk13eM/GOk432a89SaEMo9BmzAN8XpCKI0N3+8
Pez9TTPSTkDkUPbGnjgFG4R9zeL7Uv6aHa/HH7dt/joYrl95l1rfqXOQ1xxSSyrOhxaXOTEFmnLP
m74EmoLPfLnsdByyzHOrFHC3LwYEYp9l0NIO0OlEpQXO5A+S9cvnfGIj3h8lPVrAPaWVHwKAYVhk
5FXDjmaNvYiw5+OYpquOd/eQj0FkFps8LOlR1TYi6iV+4OAkQivN4QmMaUJyvoMLRym2HzX4MHWF
afe2iLp0uH9Qo31CWHyA8Rkft4p3nHXusHcWWSrAC4Blic1ttLhao1GKJqMyk5JblF9ksf0uuWVB
usxOXJ08X/v5PKJXVhY2HycnNSF6wgkhQi/JqrZeitvB+wr1slJ01YV5LahPwSHZzrbZRDNTL5kU
2VtOarcL86mz7h2rzk7xPqKIDFIZ1d6GOGy6NNokOuxkhnDB65lMpKFsMTaTj24vBSZBz2JAYhMX
H6Xby129SaWUaHTAUwqweWUuszqJy8fh2oE8zDv4yRWBB5SLxUoFO6dLv1e9Zm8dKZSNbw2+Ahfx
EYy5EcUWPVvZs2QVPHoigW+7KlG0PQTdAoJKPAFgePQxjkGNFXaEPvKyZB9AHk6q5wze06R4SOXE
QocNewqV8IqQC1TWECpxB2KmTA9Ma+pcvPlIadiEwF4H7Efq8WFr4CSCTLW1gDWl4Ye5cg/XgEou
uRqFhsoXSVzpTsXGLNK2LzVe/iR1EJ4fGJ+BoEp6t2gYXAtPdXjI9nqNaEUvUuhZ/pN7u2CyPEZQ
XnFkXdStLF13xUMp4uHALIKl6dwbB65nICa4oju9uk9tIDotUZ37NIIC+XFvYHWLxeJGsy5BJUQ5
hvmMsc80PxVKcoWOBViZSiScATI1eN9PTHQuvkTnwzxRdIPs3USQ6w60LwSvip6GnuAbSw57h5lO
mWoK2txm3MtwWMtifDSgGbsSyTNT3gyLjGiT65FsEAS+w+GURXrlX2wneU9GuPGBnKRFKKML4tKi
+bEPhuJomdrSy1Xhg9xE1LrdWDSyF6Ib65QDVYSmdVOlvduJsbX8xdWQ7XRwnLi3DKOXgJ3XzH3S
4bypDQASlNrgNsylRSOqZc9uHtdCpD5hLzZuxfrk7A8tx3fAC3LT3kZeLf34O3+3KgZbtK5rRZKd
UqLQOZ7XhQs0VB+IMi1C5ObZM71eynqtSbv0cbd4uk5QVx/ZCRpr0UFTfNW6pi9J8e7if/fr26wX
nDXQ4xDIQqr+d+YJb5p80P8UAxpW8swaRBRwgq4xueuQzbgoSBFUja9WlbmE28KgGct+UB5d62xf
1x5WfRiorIreD0LYg9+hPOj7oGmuBuXEXDlCXa3xrvNMaQxCntqoGYCGTY8Oik+OQ0bNNFCLVUn4
/mkPF/saj43bmSEXbGrWBxJKGZIPbsLdIZMXRWJtPPJtvpoTt1e+xg9jyoOCQNWtWrZj/y9KXpFw
QyS6WaA0kjZzuBbD2VBMzCrUu5R/TGZk6EqJvXZzKZ7ShPHEHfqquX3agNF8Qkg/tVPIfAHjwiaF
sFs9Vv41QruT1byc4yQUjxU4V2zWusXYzw2NYieoQ5aE5mxaRlGBcLP+nht0ZCNFfvMwvDCh/RSB
myn60m6TiS9ibsSB81DYijl94IaMNqJRe+HnvB7GiXKlBMBe7un6avfI0etZYFiKwtIgLWXH5dNK
+yYUqWp+VuKQ9dpOPOhSVPShh2/UyLlaTtGJZatlinWeKEXHbLBBXMxHH4JuwIDdLB92iBaKY/gB
oDmHu3a6OrSFZKy78ZQY6it+ucm1S/ENKjqqOkT741QoxRTgJc/YlW8GW0sVuBMM+HQnZ2FhZtj0
ySIbl3hyX/FvoP+jFAG1mLRHaym9bmA51wzoKsORI9xmoYQKKDMHAO9MZnizHLuV2BCVrjzz9Mc3
xS1Ct04CjNxVrKlvbWaTc8uEmTyqqS2q3Mdy0pbfvRZV7wyDeugmiGci8ZYGNkr0BWpQtbHXrtOw
JYoIqW3cP6sFvKOj6HzcRuu6K/b4XCxsIK6+TCUxZ7eNZG2xGGNSLBAdpkJZ9hXxoYE22wtNje94
mEdX5Nwc4rHzdhN0nefT2/vgx+yo75K68engmMmkAh+pOV/Qk8pQ/H2WcHARmbClL6sk1PVCKt7H
PNsV3r0d3SpRICG7z4Xw3UwtR7vI/xU5D8sum+h9My/4q/mGomZz3YMybrLHAD6PfdHqnTLYM2Sz
8r8ur5QCr3w4lTfmLVFJoKExZf3ukT0CKd6Q4IQsmpriIF/T1pMQqqMi56FY8+EIzaMIqFvob+Bv
eJrPD2yeRBDZCciE7Re2c08Vu919Cw0vwJN52ALm+Rm+NdLmx1t0APs1b5Zc3gEsQq4rVMLmgIPL
8MfOkcY02s0EWwNATl0RsZ3MVY7CKr1EyrP5mb5COlPTyrNY+DMOEW/3N245iPSm4wg3wG6FeHCk
4sDA2oqlFKmWUQeOep6aryPCgENBti1i5466nHKOkwOcScsRgrQDxClUTfOg+PhmKhsNG4yJspY2
7B/UyCrisD5VVyI1A2wGo1sszdhz2QJJYDIreYkUfa+jkOBxN3r9VTb7CI+1bn+2Ox2aTwWGbfUM
KhZ3ayz/OHDzU8aWwI82daekMo6b+r1shu0l/cgQqjZ6PvQa0F5nCn1J6NWzamwc8268foD52tf4
FcXwRFMqyOV1yxz2XPwsat/eMHIeVgzrbQWb+vAZWc08ScptS8dDHAVPwp7QKhyyrI08+85/vE4O
WUjyHdO/AakHCG7+VqXtbOdQ/FcTwKG1lkvstpZf/a1Cy7k9lU1E2/WGJAFwIEEqAuOVn11scY2S
1NbXME5Sq/HCEVjHW4POzlIsoZXVygo91CKinf2bHPGYjyxiPt8R+pgykZkJothBLj9RmQfxG6N3
Xoy1M9Vqg2s/8DhOA7yxIaBFUfyFcx95QVKMr5yChR/hN0gOLSNZybAVaY+ax+SZXx+FQzN344QH
Vxp5TpbFbXRbp9daLPSTyb3LX/PUZX7oQGWB2awZ3IWnSEKm/664+nhx2wfAgjJH/mVj6tnz3hjF
n9sAOFRfPoLc9dp2g83EKJWR4r+qIiHnnrs41bOCiU2BPx5Je/+/4wGK/rN5oOoAYizA8rZIFpYp
bhYfKuzH7b0vRoJFmw7GAY1qvVfWgp9Do2T0gLLpV+4LBlkECLWs+krTr2Ok6JgCRoCjm+9ajh1t
wz/UpjRrrg9VHElP/iB0m+8SUti9MNDUfuAVUmLNn6RV+IbrcHTzCWJ6oWRnvNSksTx9VGUUJX2A
XqEUQv47MTriu+HWzxbYUytLSiIPMd12sXAjfvoi7lDEUoq8I1/ueWYGTj6GEA4TTUL6WVPtp0zQ
8skrnKe98BxIU4+DgzXH4l93cZa11XkRyM5YEfOre+8VCRHNl7TwK9eez3B0LbvkUC5xXeYRCQOh
qGsJGJUZoAsF+/qiyCcRaX1ltB8FlXBZ0U/DWgvie5/AoIgCZW/pncqheWZhP/9mkKGJ98CNftwm
ZFBNcQACmqzF0OM5N5pmhIdEh1shgoCWEsN/aRQlzlQ31IeKVlwmF/F6kjl+K5vuXVi1o2YkBaOI
Rl4zym5h9fm/jCUITdAHG4qcIQEyt8iA3cTjra6Ew4+QKBPnqOf0GTnd5VqlxwzoVm+8CU/hWyAb
o/UACIKEurlG+VbdisSzosa68hPeQNtanuCE0GtxIzfpgf6ZV4V76iNkxZuV+/MPoBps5fN3yE81
KoFJTkGcc6Ob7jOUP+fHbg5+8Va/o9LEX2ZxTLgp4b7+/cIgVIBA64Y5wQp55nHu7bysLC8v26oG
3ih0MgOekTRm24SE5cw1w5JyNwIOUYXfNpR3jOvX4WFPQQPioClk6wpqgWS9xCJnUMwOJaQao0pX
t38JEo5yf77u6kq2UonUil3u50q6z6Th6r0akGU1bi+O0BaG5eU9/UhBOKJ6lm0kROk6KkAAHgyE
hF7M8coLtS3dk+q++hb+cBO9RbrVIkniERRNx1YRgdtJhcPsk4Cvs+ENsN5JwFEed2qMMtpx/sLF
HGs72Nd+qXymAbigj7eBo8al9JX44b23Y9TpqkqfW4XGdJyA2DlE7ooT9Y6hSiuy35i2nY8NzHQ2
hya/EkHN5kVgwW67PtFkROSQxrfRAHOLpAl4Zzc/LqqqhV4CZKoBb3GqoSu/wWBY+o93YEy7/DoZ
qTDDGGeWlsv1nIXQoomDrM1h0VZYf0DHXEKQ6LqSGs4gThpqOdRkedNvqqLMIo9JRac0rioFAibx
WwupG77Km4xuH/B60sihTwkv8aEvZoiT7xM31Z4H7pjjoPr0nRyZ/g1+dbAyCS4zXHYkuykUu1Au
8QPXHY38tGavGlksFx/RZf0tzhHo8FxDvMq7YdQX8XmFrZTkhKaH9Pfyb7w8g8Gkx4eV79z3dYJX
1Oh/W5gA4WrGUWIphpXSecn88lSra0bVGstU+PbUTq1TTxs5rhx4IJhsJPBokULM6yTDdqjK7eyx
WbPam6Y7DCn1B46e6ywp6ohsBMjwJlb9KC/CJO9rc1IvDOb9WD+b6mO2XWh5IgWwgoFypLC9VPqj
BV4XOYmrHWqybDcCfif2ejWWbHFnuHX1zJ4S/bcNrQidC1oKfZSDdbpe8wYs69UtMMCvxLSwi1Lv
5wxMoyrzUM7NKMj5cmPpafvPG3ah8J1+lZF5Q5/mN56yOXsBW5AWbKpg+vV0VsBWYgfUhKKYMS7N
deHV64ShowIpoytGHTyumy0eBkgsDmO2Wwq4nHQaRn5WR5VlUTijZb7QzsLyZfwridhSMC8V8dew
uyBWxJ6i1Vwmx6J9Mnkh5/zibts3Yh1M+VageJ3GVuf6v1E2JPvjEoHPfepcu+l38H1D4Iu0KUyD
sHVREhGa+NgOHS5Rn2sdP5SzqnQ+rn9SyjO9C48LbwBLKZqjeqnE4NJ7SlJEUdNYxzqzxPLTIr8Y
/hRJzfz1zRTlViaWBAk5ZYlp77082Qb6fsS/qvxSENDpkpzDhLH5haiHojv9L68yh318NhX4K+Q9
UHZ9yCCdJCaMj7WAzVcAm78WMNGolw7fHJEaggw66mO9LGVKtELlJ7txDFmUIpw+Jq10ZR5Ylwz4
huHIB/CG4X+fcydt4+4TQx5uzlnYi+FmJmtKpkvK1kgizic38diIi9M3HXZ7hXLO4wY8jQA/S4pK
aHYufDEU8fZFVeLeEv2gU/11Y3yWMZ4NThHG/qPl8JxQJuz7ZvTUG1rH/jQ1mo25zSqcUE1QCrFB
ilSzJ4ynCMa83SF4dbbdky60kiBoUS7A+HIjNEVfFsHN3SB/Pw1ST04UUTHVqsztDXmsyxR6DxqT
594DzrL0YbRNVke4qkYvc/Eq0XuGj3GAYchfjmRaMYH2+NFG5FnV/ILu9h6/hVVpi4OHMiM9SlUW
KxHJNd/yaxDFKEnqA5z8sdtNIXswx8iJQjZjCnGciDdkcG0tAaV/uqH0Vm/6JWZDvXkwWYT87mzJ
V11b+S1wbF/uGUMwvGPYtlNSX/8n5cg3Vjojl1jTzTGudqXZkNUWk88snte7XDnFZxejhD94o46g
dnh1dlaZcmeendSqd5TWdHQb8SXrJYPYGLmeKex8T11aWAYzVopivRoN6DSoA3vzD5W2Bt2GRsxi
Alt3QdtBVzQdOyLc62PCNDQzleuzrm00VD4sMMxpbH2ebUB0RwCuLzMjFXFbHfyu+y95NNvPDGir
ODoFSKqh/REegm3Ir4cIOQUwkyPWJk/OCOgemIqnMPZqrSfX/0WvldK3v3fOtJsx5PjTapnF1ONp
UEJMrRm2/GBlwYQGUpYqJLsDZ4SJhJcwzxCBWpFkKnZYzqPk0VQJvnBPQ3D7alKQMf5PCMH8IWsP
N0aqs9xGOm9I/xnH6hh+m46UmPYd2nEfyrpABfHY1oLjZMLxyrRRZNLgJhwcWE1reTXBfVq2mRmp
IxVhmJkEkcnp0VCUBujrPelh4CQxc27m9mZicQTII8OY9Ec0p5gbGQIBsKuvAL6lob/oh5BnmeXP
FtXVeTlb4haT/ZxrU+MQaDFvSqmy8lWMj+2fa/B1ZiTOuOczdtTLPwRZmVpKRrGw5qRkeBZe2dZh
ZyK/wk7JBHPZMgHR0vCEmGDptm3WBYIMksoJCGuur0I9cHPG9UdU9i+arLfU/L7pbjevB60ULPyq
PHSPMn0kqtdpqB5oljousp3q+c2rlwX/dXf5SkIkk5ZU7pQtM3+Xu8tlmV3eNx4Lizq54+58NF+n
kJPAEdYb16tmD4G1dq0GmCqFARCJ92OPQqW78OobNMq3wQ2gKBqGkEoUt4rw1FAzv0xlYX8M9w2H
DcQQRy9qWqpRs4ib5fY2chD6jTJ594bWhIeqiGvWSpdnV4gcGbkQVkxNk5KBW8Zw3qzYprg6QmAR
oK+VvZzRjk/Hni+Fmp8Yw6b/+rD1yDy6QDWkEpSpPRXMpo9wEdcQlYP1iKCGfFiGZPQiSHPFhfYn
wE9fNrrY7J3zmzNqCn0d67CAuOuZy1+rxsgMk0mddT+kLJm+UyNHhh86F7nPlhhdRfYtcQaYXmt2
lrekfTuY55SoenZxmYzi2nE9DbUZ0toVJcofXrYsHB0FoLLodOyK5ZxyCfsEa8ttXb/6KaE7vjpL
BCkzwKfMZpAM6nwVlMmtsG3N0SKkawL1qQ8gKmifVkutx/B3ZnXfFUcnu8hDKIcM4j5cb55n5pyu
10ptwjxYPBVGMQ58rpaT8UV0pliTK9cVmVh5OEigyT1qc4HoYRXurkfL8YJhIdw8u2cMy1Cygx2b
B7ju5PwAbPmAuloxex6EtIzY9aU2ktETIkyJ+9V/aHwtSuAWn5M6A1Vcuy7yhk5x1oVmFWoV5SWa
5vLBWKMZxUlqenWO+sfn6RQqk0pZ8LnDI4e9daWpsxmpHsxodmTokYgUPeOGf5Hn8+7bWNDKtxfq
8of1y0fUwS5SbuLZj8y4zzEW4ctXL+nnzpmdRLgRb3UnwgRW0HKxZjNup8FyMW4wlNRBVTOyGovD
IIBCnY75C/Ae2/ipc4RBedm9MW/iS1YejydlLPY6aqTRTr9xOy6gQfbWQbb0kqyeHJEAojc/azGh
CqZSrseObJRrR7KVTdDfuGEKHpA7sLbvLTm/5npEYRkumfJhE8UCxVi39cpVM9dpFjjTxz2AHq0y
8hv8axSIr/731NUcujgPf/GJAz2rUIorPmL2LkfIYJoJVRrh6Tbi21OhCvadPrHmAf43ceyDQ+Fi
+CIuzh+LzGK2/0BMx+tTl6z3PTjw1bILXry2wEQldMs2O+gOWT0QCOFZHYy6sXp05uG6Z9cRwm1+
tI0BHHcaeU9o6UCFM8XRJCQ0AsAoxfmkpfyXRoPdPGGL0YZnroe4Qe1MRhIi9nb2ljm6wS7cRRU5
CZ7uu2RrCFPoWSTNMdpDjT80ElTFSeXOMusP+15PHBm1hpswC0UP/1J/3Tre1eUBqhtj6LUxc9zS
V5fFieoapAO9ztfGdHlLsBk8RQULYiXjmdvwfBnecyUp75eXsYMYQVulBXAQnKviv6z6VnvoISUd
LG5IRD6y6n0LPdvT4ML0+E877HKN0a504+tolan6GmU1zIYB2u/YtuD5sEFqSCgFg265qNY/LUHq
sumob9tVB9h/81ngh1MIm23cRyWIHNChYGO9eGni9o3fhRoifoBr3S4fW4sHyGyzXaNlIu9ETJMH
tGPARpugrOj7BfsQ3BOpRaq+HlRE71eH6lc8i4NaCk+V+6BERrMcriwyWwXayfDm4HgfwAdOjCv8
wmjqFK+Kziw5Ra79evhBbs+YV/I0AX2aWez10Hf9P0qPkB4AXA1XPFi8+efnXzL/Rp/Za+T37ZIj
8qYfcIoHm7sn4b5+GDAZIKBJfHMEN5y8jrIwCY9X7F9hJuRLwNbLoMshx2EqCgstbgiRfbF3/hzf
yQu/fTQqEe/xxmrM9v/VUrlp+QLLr150/w2eAIzUmoM0K+h5gcN7PYsfYdbGYB/IaFdIg2Yb3jsm
T8dfchqaor0qEIhYTYh7E+yjYDAMoMenf2iD+6+fBMKRwLiOwvYklgTCBLmfRpS2w0homqjRPy2E
kjUa5xJlatnjLUvqVGRktxneesKLEGwLSk/2uE/VjFFulqobulvaIp2PPMAx/RKAvYUxsY5+ZhYb
VkshACHGT0jq7JqOBtm657qq1aXz2RwqM5WmI4b8dOssqpbpvi7D4hg0GMQ8TZxiiCHYv0ioaqWH
G+ReSFekLX/7YvevEvBfGRGB5cZrLRYetnexSUow00CK1Mow8u+WCTmGRq3ApuURTCgLLGfwV6Kw
OW8IqiySR5Omf3p3AMuXBKaPVmI2Ob2qj9ejkq7g6u7X08P8NjDddXuOpnKXGpVEPpagWOyaFjgL
RV4ArGrCVJSiYHHeTxdK4t5REjjaxohzRPBhTxdwYYNxmsgc3VLQq6MdP9KMdQltWi2VixzKThlE
hsRzzj29EqObveroBpzG60yZe8TN+9p4UJhb7XZCK0v5rmXZP0cf61FOijtaVSWmQCC0hp9qED6q
Ef0+JIqO22z4fqNrOy34bLI88s52mh1Gk3FlMkEDuW9dwFgF4wPFbiZEM+Q6ERcZV0c0/UWAwrNh
u4Aa+L/2vogef++Rv5JVewVpbyZC5O+E3QJZXnAg3Ek/3YRspbonTajohY08LDiFDUd0IxTlqFG9
GUMW4neNqlSgsCao2Lbi24bWI2hBkYI4AMj0CiMpSVX3VAIL5YzNFFJCLEnXc1+qnwHHAkwHjzRU
gHY+oV1YsO8GPnhCYV7rTgH7Q1kxRwupiMIT9YuLYnDyXedFNtVTbrAsrY//jo9VkJDDeA9l60Wv
B0JAXEAlUtGwmz4EFBa1vtVr7CHjT//Rv+Oik5Snzm+sg/ICs/7+S27tHMx4cIFgwv9/wqbyTbPg
aWv4HS1ps3Z0LuJTiKJmaPmdhneyYpjDz3e2ix6q2Jt08ibBHanYD0LBZC0Kvae784eebKQewX5n
/6SrNUJN9E6iCq48la2/DRF21bCx2WcLAKcI6jiHAuHSZVh+XHyLXqtgi0U1156IHNqst/H/yDF1
PTeIkKbeXTYhE/mu2MZEckm20A/4iSLhIi2M2j7PXYNbVq8jL6Esx7V4d05bsZKjwbMZIKIfLkJB
64pH/YC/+kAAVgo7chYaQqe4HkpSepOxX2/nQzdBv7Ql/93C/4zKdtFWiSnglXKbrrHpKGsW87P5
oEyGqaO3THhNHfOL4Dr9Dm6Q8SwOnAt3EAw0dMuPbZFBq1KgVSplCrSV5061eo1QnynKa5Fgbdcm
K4yh56Fyv/gvg1tv/Preyqb7Ebl1V1Lh4n6MGn6erbLIRgDF/HYVv6ruCXWjbQIGnDF0EtMBPIo1
uxtnfAREYJT5kDfuBugcUo7EdNkgWll5ODOdZF3JOGquhnsN/V43OMz2vTCuLFvOJCxhnvRaREcz
QSWIgFur635Vwp1oP85mmG4op8ortSUVu4Ad7HqcJ+UgahgzE3rv8wh2uvW0NRoOxmr4jnwnIoC+
dYbXuIYxEbQ15HGL2brCngJxhaVSt68NcUxKfSICPfF80tRx0NhYxBLa8mvnHJIqv6sJJ31QJ+6z
W2I9y8Up5taEEwJkVzhhPyXYBvXQ3OKWD/+QxfuSI9llP2sFLSuYakvrfqTHe/oVcgN02eO2MmXd
EzD/Db8OMYWXEOhmtRxyJcxkqRFCcWtep1jALd4esNev8F+r1H0P8Pu27u2vaRrjfTIcZxJHiXn1
Ws5nwphWjs21a7PBDKuhyEO414gyjZ9CH3v0I9vtD1Hy0IxliFE0gliB2razl4cPOXuH4rbio1uj
p9yTDhNATem0uUlsuTUTrgNyoJhBQyI+Oi74Zy2ldci4B1pseisKRM2eqVcKV8H7EeMHX+iwhdMs
ydVFT8y8iok/rvu2fMiInkGTbBn649Zc3YtDaTZZjBKzCTn9Q+2azKMekSgTkDa+jiU2e2l8wViw
t+HZ3DcS9afFvrtiZl61ITcPI17FR+8TBu0xTDTgVVMCyP4V5vb9fWKx7/dAroF6ra7H9fcmj6mW
XLNUD5o/OP1O0A15TutlTWMvJ0wJkDA7D4KgtkJVop6yantmQLUfWMZOkYw7MWPqdapuJYerm95u
l2yfXPWs3FEeo90GOUkPpA1kQ3ni15SNGWwo4UQ9TDeyQezf8XmOKbConJtAh1KAbv9NyY6QdZM0
WVS5ymHYFB0+emShIH9YEPgUAkLKNybMHsKa7nh8b55v7bjufOinxi+FXetgHJYPY7hGy2Qi/blF
6/zn5Fq06QuELAVn7M88lfViRQWDZgzwhBawkJJMXHLO6uC5jQmF+SzWmCz2jbGY95tXtLHtX4au
j1hUonhDjby51pKL9niRyg2gRgqecWdLr+T00lCw3W/xSBDD6BRomM8YYf6sY3YecupvgJ2m75bv
JIb0XrqobdTjgAHrN/8lWyFT6ExFv0JOb7o0eyQ47vLu4nROPlqc1gUrAmBspM9Ae1DDXB+W57gM
Dfsih9ifEPgcQ/qqGr+EqVaCzMFNXgycNEUM41m1T4rlO5zI3/hVJjxstVr+oX1FnNnrlLOPeYgM
RoPZg1AhQKFhi2oCXWK/rpSrD9WgePfeXhZCcrqlCuNvgGTofVpGOzlgWFA38Ql1xKVe2hXBpTJ4
h7vQnqWeUBF91KTem/l3mCUBIgJ2pRV6PNETrPcDTt/M8+t8mXUP0SzgX/aMXoUwDSnsiv9oM/se
/CTlbZV+1oFok6i727AEnHgi0JqXPgSLAiIHfZAZpIco0cvgS71zWLxK3uoubfbNODf4wcBqATi2
hsoFCq9iSPyTGFn5xVxfYZIEKQsn4gdEOSMkjk4+bq5ew/PUSLsXTVnzuleIlAcwrMX2xtI3z56x
cT1AQIirUxn1Abb2vW2oXjV06SGtwq5D1YjMRxHc4PmZWWT7lKaOd9bjjZrV4V12lsvo2+vtwQMs
HldanV2JdeuqlFbkwzW+peymFB4QJRPTbWUyltSaZ8JVyVrO83OhC1WuqB5N1X19EWf5DH7/QOyJ
NKjKuFivVEVn+pkxIsnTRvlcJ+tP4B6zWUQPcnbcca+EQpv2DCwMf+/1Ttr0bWilWYdMD66uSruM
ydWwDO7auu33QncYu0kbA8DIfll+D0EPgbFfZexS3CB0eQ8Ufgwun+fPUCMZb8vBnmqaHp+hm8yS
BKCKp/NFub18c5lI8wFtjljF1QONPphrCzMKn44WN2eam2f8GQMfKM0sKIH26DeMJOoku9byO1go
cPdGpJS3fVpbnsfftbGe3+qNauiVh3ujIENZbz/X6MZ25EnDzyy+hhsWn+zhWwbd6QQH+TaVvbTg
sdBsxlM7KHAx9bZBZBs9PZJhpQTYkcmltYfXJsi8MKAJJmfZMS3Ke+utrz7XzvPli3uQ7BX4y8Wy
gXRg1w4vGX+hF6Rl8S14bTA6nSkrrGJD26X+HLgCMYLxnzdYOeS7P6i79swElEF2ekL1TzsBIVZ5
SyCgPhFL924aE1PJwp3bYjq1n+ykSZ4D8mRjAf36eJkEoTHqFRMkISd5Z95NXjYmHl3eqoroAPp1
3YhMJxbVbtsZkPBOfw0+oohsgjcHdMTcDY9wRrqlwW65ILcU4cnFXfzj/5WTshDtnqq/gBgc/+kO
bSYgVZ1pRKlqbFaAJn0F8Q+i+oq+f70EhL4Pqhe6HZgUs0uGiEE4qAY19Fhrw6AIGKpzRZOG5cTf
gvQP/oXJYZwMJA4klXBZIx9QF1I6DW4M6EiYorgMOcYTqkmn87lKOEIK/T1bqcYZHUEyzgtENfRa
EmAe945Wvfzqb7lBjrcU4skVgg3dvkAGHAF9OS/rMVhgdJQWKUmWsBZP5d4eWwoPppfy/DX6IGNJ
2zh4lyG3+kuTt9gVxXqCBzLq1MvVg26zApzrBIlkGxUazl5maThRdYoLjuGJAuQmTtVKkM1bP0V/
V0cRlrNOiZsaSq+ABXcUVX65GT98lk9O+S9HgBM8KxgrprgwGbQQK99l2QnK+2+1sHkx1kg+hv5G
8PycpzjdmnL73jikmy8jAJbBw1TZvubBu83+eHTTloC2Tqsm5zo4ddn3XKxi2krZRpm9XVaOw+cG
12H9LAcYEFbHUgt7+OW6E0GGPUq56XOUOxQGZaqEPwZMrBBI7codCrIO4qRV37MjXXkmIGz4/Ldl
8H5x5aICuuten+1eDNLC1ra0ZDTBLRVKcbEmYwYz/DLxKRluLpWq28KPOOIhwZm6Gs5QqX3654D4
QDHQR71RbraU1t/0t352FSYeVPg80EgUT4uoO1AhkFIS4gpVhWJHZFSpnwHGuRR6O6sGU+pQXMNk
zfYHRBUxkNqKtLvkdBlTqgS5ggL2SddsZszOCtyT3gjXCJtSGwE7ZFZPYkhMZPy1OhFjoofw/Lxa
gLlXpPMF6zNCIfafaTxzT0rg8YDBka6IGAucznUYqwilH2DZwg33IwaXK/Qyo6ququ6DLCWTO090
8jXWIzE2B4ChLql0iOcQZEhkQzO5wPTJ1LY6OOGUFdHpSOSg/aV32Ae7GmA3o8k0ZEvWYgF4Vpp2
fCY+wwc8MvIqy2QgZySCFAiZF4ZVBtSlbNxRaOKUQkFj4t/UECqHNZ2Aq8CRKC7y9C83UJQK3aB4
2HUZ3IpfYd2g75pQDfPH4TLXqB+0RWE5mVZ5G9N/BMTSYGJTBRDeWyUNxRe/GKTbBQfTjEa0ZZZc
pR6DhhhFRyObO9Lm/rvBbZk0yuB50pLDsQE6mvL+YgCif47QP6O7WC5mZFp5yb79aWfZ/aw2si51
fHCwBaiW5ML6t4NaC2sWL0hXHj07CQTg+ZtuYm+h/r2zecJxYE4M1juzqCj8yTOSGtBofTRzs7K+
WxTCGuI1WW6bLrzNLXztBc7CCe6bAhJ5A0hc4sIoJmOPKg7caVfeRTFGSkrYkk/k0LoEUUBamm09
Ab728zc0WNf1tZloapFiJ9js1uE5vQmDrUu0/UTgc6O2cVE6UF/7cGGPCPSu0uayjbQmXcHgCHlN
N7nlUshWndYSp3ISBPpKHiGlCt4MDII5hiiKL+apgK2E8BWeyFI6QnWrglmHE8ktYFL9R/bsZpp9
Ipjpah0tnaS0uLFy2zd8d5NhkkqXBjClE2TZJyWZcZp6Rt8c5Pxeg/opRViJRFM9A+L2XFDWepjj
xpZZldCElq+6rtIjv4TeXa3FnLM+bQW/1KkkxUZriThfx19wnQXBBim8gTnYtVmUf6MkdygeR2wK
IFytzBOfePRK2YozTpFlJ+h0v2D38R1Qsl2Hjf+yesvcTql7J/3khgwxInZQymFmGZgOCwbGug/9
RR1ok7FQ3HcGa2+f9mnUWmrlm9QjPnRJ+HeOBhIQRAjWl4oVqFXDjxjZyrNlVtrQZa/FIMnNC/dF
I1edoqZWbm9/VCK6EPXnQYH4e2IqhIEKyIYBxqctTgMKcSjzSxKO6Ayhna/SablbvRZbJBfLwzHf
p01vwb/6ywPKw3IsAPm6iLIoTLn9lsHl+VtrCupqcwbFjYINcUDVQfaAgAobN7/zSaiHfFKvyfbl
ciyMTTkhfkssOZN6h03E/zMlV+p+gO6I1xU4LdmMv9TuIT9Yg8Kl45G8LYZmM6Kj8b51Vn5aytw/
ws+98qjBBZXCO/ZjdVkZ0DdQA3ujzCtPC7/8bGor6lfnpcflYao65CzOyc0hczSqJYSEOy6GJNMq
thrrXUiT+oHzqIPyL95Zk97m7pXmtheXqeXdxUQPbtyPl3aZxUG3FUB3w/lGMX4v1Kf14l21hcry
zYTcVwo4HzoVt9plKEUKByMAVG/+gcxKrbusdYJufXwmnUsFPZRYz7F4kTmmlnrsOFMfn8wmdTg9
Wh/ZycbHUnyqHsMRY638Nh4HC0esWv3U5rpbqCa6lAmiKqmdxwyLBCEnLHxO1ARdaDhNVK45d4ro
TxiGWL6OuECkRL8flp6sWCmGhjJKT2NAgpdkzcV97fkMau2U9KEdLfUCyA6EWQTZkoOAp4MxoCAn
+0jOOfQ43ETzmAYBCXqy/1q4pvrVp/UCsIfNu2qA74alRbXz9Dc6l6VotF2M2HDoVlUJcJI8nmzV
hQ0oVQtnZ6tj8OCmr3YPp7K/4q+YAComjABSGBEvSDpfF4TU8cpSUe+BGNfAxooCAGbd432GAfdL
vC6WaZ9thIOhgisigVcitNFGe4EC7+pf27dbz4O4khhBX5EREJ7vDhFbkoYrHsbx+csWW3/O2pbd
k/bqNsPaCVp40H1WAZ2lxHJ445HboT0rZNNf1Dj9Iwedo9ztWSO+11F0dheGxYk614tZrEa8sNQ/
jI6anEaY9qBRgal+EPb6V/CZMhfoUAK6f5DYg+m302qY8O/4vx2ivvp0FyA/VCKOlLgs3IyO/gSp
UItGMlyOxqd0DNAR5Eb1Gxn5cezW/lvfttoPqSpXT26RcOrMzuAMxhmOWPAtqoh5zjyUe5mc/Bh2
aLDa8Bpw6H6mBodIjv8ELzfodCd8Yfjy8TvEVkS6WVJGfFP4D8Hw68n95v5olhOwseebrIRM8A78
uRdzh+pmRkxClHwu1hzTlLRlvcX6FCRyC41Pk5Jvr3prhq56hvLRmaojcHI90mj0LIi6eVH171nz
lJsuCyAZsljU/gzx4WJFTTDvEyj9nwZ1ufqOdDzrvfxOnw0LuaTlOX9tuLtwUFGiqxS12B5t4XQT
k50WD3K0M6SU69goHiDRJhR4dV+QMr+YEWznG+97rDfgJAw/saUSnD0cxEyU8TPFPB1KbH/op64+
U4kRLwV2b5qqraMnFaID0naN2SrmIs5c48zSQc3ckTYHryRn1qtZ/1OQ0p8xgCAzmBT9otAuxVMZ
lI+XURYmC1Bzns+hUGLfpTsl887KNK71rSwXOu4iv5gAG7e+i3bPpypyfqPke2+9HM0GwdMOzJK+
QyWmuJr+zNDa1A4aRhSHgLAf/Un3sXGax3rvKBdypkHPTO5XBe0RCDYIwINY264XIKY3M05gmThk
0tXu0JM+FRFDlFijDxLzUHBG3g8WgclwdfYqcdSqQLziyggTEvrvslXmlCiKuJEicQPJAEfJszBc
zSaQVXiXh7a/MbFe9Rk7Yh0Xp1lodPHpXqicDjNNyr1QJ+mCBWZWG7z8Zr3yF2UfVJIWymGaQRm7
PwIbaieR0q/l9NqZW2rPHwDGn6NCTubSGDkyATgGR24ddZm7HpPI8oIsGlLM6NZoXr7GXTwMxs1y
Gmhv7l+1AGya3O3+ZbJQ3/cZHeIL+79SXw0FjUaKEv1QwQ8qSOGAHQi4UcUMdVacI/0g54s2eJ1e
eDl7UHajUOmlzE4334RONvU9Y6aorRqiNuGdOaxZUhR94zxQ8VFy3/9z9nYzRfnyApXwWZysQlsX
hQM5WBnABfMQ6IcuyS+zt2NzICMsR7rtGTt/Fgvc69EuxPKjw67sEZhPVH8i22n0k6N7xmO5sGw/
cN4joVpPRsKOl2dewckFIOPU4Bl05HhrXZWgqkrCtfzEM7ekJHW4zlayOs9MKT/sh5Gu30Vkt1VA
vw5HdlhAT2RzeUH0whE2ia0BVJQIFzOzmI2rTOt8UXRBd/xyLD8BgRAD0IhDEzWvc8l4MRswyrbH
KVpqIUA5TccIe71iNT4P0VAKkASV9i2QXevCF1VfXWQ2SSc6xxoyaNrhp8l1FuRgeQdjqQibYP75
8Md9wS7EUGD6xCP+MXTsYWL9MO/hf92LA3kI5VQtRB6920GxVx0ZAqq1WIBOcUGkOyfCsyvh4qqx
Tj8BLSq/bPmrP3u8ae/jb74FxmrT0GaKQywgr2fP+FimGNKHCedi3qJeE5BK2eqweJHFy8klkmrP
rc7ieqC5YyspNy8ccm9GMG1pIEMdgXyzJfQh/xH6jETilmcWuKdumELqEWN8PADY6QC46TTN7tbX
TteXDwsDZXLc+fS733JrbXRr7lcJjIxGEFOcLLpEZW4UiiiX5AY0j7Z0NdiaOxw5J2e9Tz8l90vt
LE6zJt5I9KfnsUxvVcquDyTqud2mMGAnDSAsVNRPt570PlpqwhdHLM7bQ5dKDNwgsCkyq7pHzjn/
EALjcxaf63VkjBe9bPmDTHXx9Gh96OkMVMGh1KiVy1OKChAAou8orr08JSMIVeI+PXpL/X6lvY31
/bC47M0qUe0VQVisRiiod7uuU3ZeqdxGKB4Qiu4VZNhwr8QSBiuYR0IbtfhWOmt1EcHm5agqFyUZ
Dewe0MEI+V8UizEcGyAk9R5qgRsm0r1ruEsSfFEIaubiaIfZ1WpWIn7PpYiON8OWbhOP7F/M5KxO
8ESJ5PsZKG1tcMrkKvAqdt+P12y2PMY8LF5DZZycVC0exR5uAAG7PTcJubko3m/nOAu1Bg3DNUiA
KkOjtWjnl7bEkdO7DZJCw7GmiWZf+7IOCjngKa8OgDO7zQk3H1+c+A8QgfnNpajdjEPP+CCJYBQc
HxrUoKrbaipgL5O2DYFSSqNW9Nn5gQqzudkj4m58hnf9d2wRa04EB7fi+4FcBrthVeY+aawc1+Qx
QsOsYdMRJnj7cpDM2ghsedWKCYnTCb2DodPTgnALSBW6rzXezdOnocgtktjf9qHyLJ+pCrKfB9Zc
SjLBnl2F3GBxe7R0dqA/rdaVDIZ5Xtikq40+KqLzN4Xm8bXuOYTOUN4h8Hrvf8kmte9a7St4Sty2
nHNZ2wEaPiYHJz83hS9U/GwNSzp5OQqn0cuBaphmUKvZKWOjwFWwx71Oeto36OE3OXoldO/D2OSA
35wsADgowEST72zC9DIzphQSk6wC5YG3N5TDaQ48S1mplXdnLicnAP8cZ++dq+vuF2hGZXmDe8FW
rgjTqq6VDA4VwBKm6Hk4Al9bGFj67qLohNBHRZUghqYFXBrxqA5uZG9/psCUfj+7RZFW5NrPzJtu
rtS5MlEZXU8l7FIg/HSdTYa9AlBBcTJ4FP+JPIPBrvnRgRVr69K8vuO+78DUifDYsBZ9FdpsIqfd
lHX1b1ldk1WC8zsZpzOX87y58MZAXcZ/t1n7US1lE6EW5CGtLp/BdxP7aknfWoY6MxRrO498BQF9
DvBVPP2GYJySJZzFBf7SX4crfCsJ3tIjzV8llzml3JIHbBC5nbnAQbv+G0y8+0FJ2GW0PtkQyNU5
/WVYSlzYOGHKZeuzqIjRa7M5YjZouA6fn/eTuCqddnm1bJh9u2VOxVmnQVXVJR0EtTB+j7JcKchn
2UWqv/lQJjGYx0V2/SdrHnOayc0WLVDDlfr6FNctsYDCX0Lo2QJms2pxP44eaX/o4mic7zuaumwh
teyU00hM+B0pvss/1bZf3JCHmg1591D2vcB5E2YwN1VPGIQsXAZ+veedN01Cmv5Q5v59pysu50q/
GXVsQWI8IckPGdPA9JCaOpffptUYE6fegywZHmSaNqTGp9g523elpQUHcwza0Ih40wRx0m7eVSSp
lLf30ofjtHXwxU5eqLNOy6LAEe6xS4iXCl8KwH2auM5phi6fBP8RF7xMnBWmEPLmziZ1+A+XKg8u
z1dgXg4ZymuTTn0YaGOF5lVdXj+3Sy5s3Hap4O/1XWwtOnm5TSAGNzYTtNOzyYAho9p/i4km6Lyf
PkX0ynEYojn9Ms2f/b7WQkf1e6zYY4RWPyGWZhtDBLIi9n4vHZ0+v6aLbOPay0L6GwTwDcqJSxm9
5NjVyXJM2Tih0Zq87ddgY9gB0b+QLB4F+gWJBR4eiMhILQuiewZoMEI9BByr+nuhxLuwbt/HBvoC
ZwZkRieYlVa0l0jwiCI0oNiSfOHw/kZ687t5lrYPBLAgFFGeWRtdiOcLjzteZygxjH4JoCQbYcUu
8gxOp8UzB4Gnd3eVVVNbd0kTRfMM5FGUu/dY0ZCAFrDb9LzWy3iFvo9KWBMwOeHvB7TaRYIJeBl1
IOQHPG0t3Yb4oCvqXDnOWxARcDvBdV5YYu8Ubo9A/+ceHj3XpjsOuaie/JD/cPjQldFORlOrbT0C
uJ+cJi+mJO2XcGK/miPuTkLQb7ZIJh10pa6czqvjKWH9mrPArhlgD9Y4Sqy8N3FKK8PVPwD/q/FX
kLxOLIx9FhtIegZjVMG2gRYNmojxRc1et77d0OlMfcklWNCCrZpfB89V2S+XrFgOpMEhZ4XsqW0F
q4H0zZCuqXib0Y9ukMZKVYo75nGcKPU0QDZHNSNU2WaRu2cpF4tplWv0s6SFw8WSG+ulWrzjA7iB
CweV6T7Xn7SoSLoiTZ10H/UGTGyR6TYkTL+UbzScpQIcJSNnEOBY4Gay1yTb6qEcZV/SO9ULKDRl
LC2h38/NO9nyCMJpjKDkHOZdx269h4WNfDS2qze/PsdkA0qRwPZidHDnJcEXn9SW7rmJXn235EZG
dRp+9f3r9gfJSh6CQmXD35NtkiDsSJpW1+WExUo/ZwPqo10W7lkqdFaPWqR4jV4lqUF0omahpQn4
l+a8/NH63gN+kZkHKP7HyGuROm8pFOkz1p+Lfbm/HWIfyXe/xe5Plf5f9vcpFeT8MGCUQhR3EnXU
dR9Ki3zH5hKAo8x8MPrXDWhyZ5KG7X5Jv6MSMXyNu1G3I+sWWmw5r9YLGJUhXzFTQwKgER1ub3cd
fekSdueRS7mEs2OmvszsfGu3WBw3HE4x/JiHya7I3AWNy5Bror0FnEpGJ5Nh4zGt7ZvhsrT+eJD8
qZVk5kob5EjB/0+G96KG2DK2g2CTCCNcTurrp/nyo3qxp7UiBkIS2R9z43Z/0sE13qVJLv6Hoqwp
Egf8MGXuKfgCm1MEVJaiNTnx8Q71aGFUk9xAELglRuhSZVuZUQOIy7YKaEn2hVHnEHigMCcSiDvr
aly5AQ5D2Zb3Mgsk/vzQkh/PsQm8Hg7f52MkTnrvdMVyT6swmx/jrBizzXSpyJJRyiVtYE8EJra1
jwoGITLEHUQg98cWAXpgiPw0u2kDu2nb/NIFDJ9Lj+Ndi0oLJq6ULSPhYQCv/NOUdJJ3pgHnvXgT
KotB0ykVO04q3SPkT9TEblPGqk/rlDW8HLMZAFAcaFzUexNQi611V+f57+sDlqi1FXRD84Ur7I/U
lJbBGmqlBIHgv3T03Wc2dNAH9QkdunpeM/YS3Pld+rpeGMQ2RxzDa79IyqOuASrTdQgGw0pto6tA
rs3rrFnPt6L3+pr7TBWLA7Gvo7wU6sH+vN6B4Um63KmUJ5fXuAmqJRnRNbIrC/C5u/qI9I47BziE
y4JPBtql22Ey7WO3N1JR66H3PdgfHowPeneRW2Wc3WDo3RQVlc5/bMd8TryfsffutQ04YnZ/lKZZ
5wSlbB50yiiTamuKaZdxczwZeex+RXSsjonPsrci3YTFJcTQTgpyHkjINOjBzboeISXG4pza7QyH
8cWunANLgUoDvCC0cyIHp3bIskhDGx9byVqMU23aiL3M7d6VYXQiMJy3LZvQL7I5TDhEBkx/yWGB
XztDbitdjya9cwkPKTJOQQag6VFPc741P5KArmVN+rCm1wXoAbNN3lwio16CfJmz4wttmZucnFbk
bQdv+fYuxgM5rZ1ZMnRqCuI8CwZCr1dIdvXfdyTTUsktFhNueq9mkIeExlzJBV3DGYyI3ZfbNokY
wcxiSn1t0kT1rf0XkMKGEs59YB4AX6nA8IVCLhHcLwqGtIObcQ4H4zd67Q1awmGy8yGzxk5ZOD91
ixiPetljy2FSvVqicFWBK17rdheBNmkFzoDdmxOcyE5fIXXtEsMJUcLpfw21QuQyvQvwjTwfag3f
urAjmExZbAwPBJ27tRLgAHYSrFupx2dsNPsmdjKYUmP3FjdGcJ8OcZ4b6njTwnQgNqgqdBHZVsMd
PkW6JRZzTTSOhaB8LCeGwBtdZChV5+jmBJplCTbIgmRp2ZY/TioFkzU0CsdYU6VHiacN7boSKl93
E1heFUm4Wm+1dOQv4mOfijm+Ink8j8zoAt4pnBVicfhsiu/+5DBNgf0bocA4zgwRoiz0j2WeukgO
HboGx7zPHoA9QmUTE1EfwVp6Lu6vm6KY12OLS2c0DOZLGvqEW7HN51S0UITLjFy8d3j3pTJJmj0f
6T/IuyOKg1pcbcY0sQlYO1YSKwDW34gKt72Y58sv7woFq+kvRm6pv5bJ8/KEyZa1qSYtrQTplrOI
hMxEcpn1vv8OsYUHSdE8acGyk5Td7tWZSeVbJhQ7sin/B81KaWDUNl6MC1MS3IyKMXPSxoKxvCCR
On8aKE+m3SawsWYYfc2iqevWudNZh9wOAxxTRbnukvi4aJPj4Fh1JbGhLZ6KNAr19Am3xQhB7WY0
CNPl1EWAoTeg6/oMpkWmaxbRyw/LIr331gbMXbR4yPHWjwT4JLPsWd76npCBAc56FU+29/yoS1kF
Y0U5UsSkeUZjyHOkgzsbj2lwZEC/jPuY08ENbd+LVPdmr0MNxeRZXlw1GvWhCJhTlw6+aSRJlNTp
YOk3LC6qh213fL+F0yzwTi+WLx9cjrQBm+fMgvxNTO9lGmM9zuZn8QLy6d7LvcImxukxtejv4YBJ
32etaYA/g3o7QuBF2yfokV35PLk1tylffYvlJ6kr8r5FadKwMc/WK3AbI37neLVVk20NGmOvDvci
PfpRxqBProxe5sPReGGc9+MnmP2vkkDjKCdvffgp64/CXbdMU9ETulNRSG0Pq4Zo2jOI7HLB3Zzh
G4i89Bhp63ywk3XvT94WPrWlvhpLqi/LZb/vupCsj6+bkA/t3uOqWsmUS2ETtu75CtUl6/Va/nPy
b8aJs+9sKYb3wYQUtp5lrEudawLn24JHDNsddr2nV1vEMv1BzlwawwSDDUg6b/+JauB+pVIkrtHw
uQBb6T6jklTJa5NO/Zmfu+ksUf0MovXxaHFTl1axNM1yq9crE8cMdsyj6/pomu2RbfPeMJbAN2Wh
gaH7+BUTow3kB84DVidisyqXbw5f2r+ozD0BCWFxK3ip3BnsqAqzUv2+CD+pcbzNrf77KRWPtDx2
8QQQmjtDOL5VPLr5Y1pOAST7nxTkTZQ5GhMJ2I4TJciN7OiCmqy8syNED3T6KrT9IxZDKq+MvjBh
pHE9fyADbJ1w1LOnBqTjQfV21nwnYXKpsPUbi5WQ+dbn9RifhtiJmM+PdExct48hjtLZgSXSZVtq
aeQ5xqsuvg1DAyPOOwdHScM/6RFG8nWv9CfGrtpJ+09z89sxLBENSy6hhbY669SppwD9pfjdndMi
7hDv4WLO366ZJGGv8bvX1appbUZCz4j4vbPd9WGG7wDcH6JbD8Ishk4it+Z3u1xRw3r/eswpfyg8
vmNE7cjEKJiLjHTXFuq7c3J/TIFlvuzL+eehMfMduf/eaLOvJXIQAZd0RerBbQhgEi7mT9TgBQWJ
tnlQf4TTNfzPJIUV3ve/9lIa0VpD6H2hcIOq+4/gIIxBjwhvvmHbYll7GrdvrKa6/f1DmcbF/6/7
Bb0Y0xLA9v2LjT4vWcqsnFzJUceLUf+RftDTYFOdxbyvvbYWTAt6iCgcNNzBW/VjgJpDP2AfYZtg
JMQR6t6ATRXK3AXM7SNjt3jEfz4i3I0fBXdSGKL6t9VHglAp76RDlwn2aVSItHz+QFCMQ044+tgF
RLXEfoYXYYJv7tEJKTEyhdPEUD3STbLSlftIWibQ67rqGJnH3q1P0ELlpM2kn3OyxVgKllGcwXVs
DErA0XutSz5dmWYYlUXWfSrylOYpIMUU1KnfgAmEAtq/uptgy2sRp2D2xPLz4VLalR8C4XcDHvWf
zOXb5PxvP0+prvqBfEpV7BjrMUbt8qEk/rXHkFxQnTo0L2GLuJdtrEozHVqgqXDmtUaYAmnN/9rh
5PIGDNNO93Rb94RNugg+Y+h7XAt8UV08DycDlEhCdFTLkTgyd25bhMc+u0AQVutO35gpxneYyNo/
Wg4BaQ0OHAYJ/buwdORVaL6OyVz81G99zAaE/6uYLomBJfPQPRAyVo/D9Rt/sWQsD7WYcM+pcSW2
jIkSHrpos9zpFpLkaPHatL0+9J4cVTrpcfKF/t/2yCPZv2OlZOMsAry0RK26oWT4csmhEKPLBgD1
OZEi/fPPX05Vs5RttfMPReB7K2GDj7qTq0RyB7MJuCdTmpBXaIrRkzYrVGhRdT+vd2p6mCo89f7w
hzGNTb9p67rgfOCX3zk5/Do2h7uWeZEQRZ8SB05jCPVkw6X7HQyRSatAc2Cl2ts+pPQ6VUjHfpHN
C0//FMBnYj7qIJUSJtX2THY1xkK6moD6IsvYqHQL6nbuV+0psaOnnPNIUbnu1fOi5FddBd++kXFz
tobNfR1f04yUX72ABQ+93xTsPSnCmglTsP/4BXKfR6jGr3uNUOQj0yj3Hn/xYzO2UDyjVyCgOXpU
o844KY9QbilNJX0PNxOPAZb3TkV5Q8OP7SWefyRtAa/hWzd0s8ByQRXByT97tF92IzwnwF4Kx9Jc
pLcDMPtwx/AMm7+2f8ZLRLfzjsqqq/uhInqheCSG/F8XzXO2h94o68EM2yxXBqmXXwBy1e93mHLt
Q+dcEuAnV8ThGl6/4uzaHZibngB6p5LfR0h0vM8tnybu5GlVYC51Xley0tjXNR+qQE2mdB7MRJJm
rvv3tcskhgyl7fElgZcSOw3v5AVx01WRwoTipImHkCtk2x5tw6SeFI9x3TLHdKc2S7Jg9EKCC7l7
7UPgSaU1bW57xdxMGBwDdlkrmQNoHdEYwNdegCntjj2CQ9GXaZtB5zoK8mC2Xo9tlTp4HRB8/lAV
2cSr4Fsc7nvXgg+j7G/arcEzHUDo5roUzutILBE+O5YBlTrZBreYJAAJl8uTy1FbrpMK3bcnuZwJ
rVJfwxwa8EcmunSsu5hNHQkkt0jZc5vqD/mUJuF0Rgop69FRYctIUm6hE6I8I7bRjz8WpukC343F
8wairkgm6ikgX5TnIXeeFX4amevJnOjLTNdlhYTwJZGp3EcHoypx+MQbJZGXN2phofQcxar1hkoq
v5d7LNMI5WqAvJE9hiXZsRUlmI4WYk92BxKYQavIcrA7fUgmIHt2XzAc4TyHdmNghxbrujG0Z09W
mG2DdEeeEBWV24mFymc3FqGqQLN4JKH96aMoA9C9cimmvS8Sb0OY2n4/EqDBZLhgk2FmC2feHRmQ
YmEagmOMmZ5ksJ2L3BBAy+0Os4vHNWeF2TE7cxfZ0kOt144+wtdNMoSuVFRZEJIT08hJEWu0aPf8
7ADAhYca8RITFvhERiiWVZ9oWgqVnVmxcq+3c64Nrt98gHb573M4I/BLeK8xsN8OUfgw2seCivcx
3OAEeeVLHwjT0zac3pys13HhGdgbOerh6dwh60Rj6nkN8I5Al42UiuI8yLlRYmUShNtV8CwWoh8C
vTCWHCh5OlYBCKqKzUQLrnpy/Z7da1hKYH2B5XxdJPQGfHoSldN1TZeIYYGoUtbrB9Ohko0i1iND
qsQQ3+aLdswZpi0FqOq3fqZuDgaXJimBftM1+kQcYf2SK6nnYF74BAtQJsCKNmO9vCR9bsPvmo2P
vLstD0NaKEyOZ3KAf1DTDaIa0WZxumGbPgtFmz1GdNpgnVe1BWuj5MQ867UwaUwmCKCnyIcL+UTh
G0OF9Wg9dGdqcodgxzMvCdC/T9gk9+XY4kKGOPuw5UyDC+EjLt6FTfn+sbIrTsWOYSfBLHWp71rT
QEr/LiwC9dZ7J7CkhlfzAt89gtP7G+QriH64FXN98IFIzQyoWJUyy89W94hTFxj9xLzxRPh738Fg
OSRCJaHNE6TYjhyr3lp5ko1cabzAzcwBnDmY90UY2ibQrLuew2uSzcFPZH9mkYPB3B1TAg63NN0H
XuodZk+wxR4aT5Nvu4+LXLjWScJ1RFpdjbz2HKmGNop8W+oa8B4JC+7rTisHq8PTs+UBApmj02/m
POoxeWZIJ15LO2fo7HyBEm7Dj8FSoN09P8Ufpmxb524ue+stc/AXreD7GuJEkTgaTwx55mP/yHVy
DT2AmKfSpIgX6fiUpN0+S5L43hFSDtg2kl+nIS7XDiop/qeRgUcqFdqnzO4h/ZHUU6/0V+zzjFpH
C0BPz06nl6ytd5NhXLb8lAW5sh9dNWH28jlk7YUuZLlRryYEPSgXLVsCda2J+fAyw+4gr9cj7mv6
7LCJhDaPPI2+4CFN/k+dEjUtt16HQEbdJ34lFlYiUZaIBMsnG+S1YFiu+QYgRzmt0I+bcf6UfW4t
FMQ1nwxfk1sVaFmNahv3PvvnCXJc72lJ4Z3SqRZXA5xKvW+xflaYZxTe0mHPGllNOEiNpsaZrcqs
vzjdVsi+zVePBejlNP8onfqd28qPzdSZqpdMHjCU/HhDUHAVck3l91/zq3SgP7RZWeTFy+a4KthS
ZmPjMY/NCXS3WvaQNTD8n/6JkDnT4PLwsxVCQaKuX6QFxYL1gznf/Qcz6kq5WyIdziNicHqpHeqh
Blcx8MPLYtuKq8IxWothzseNRd9MbMzJRBnfqtbxkK28VT8QIuHe+DD2Jxo47x56rT+SanFwb1GL
QjfKrVBXK4zQDuoZbLeak/oSM8SzsSjhAy/DyyDDCQd27/Q5Btm6WL1UikBwJbAqZ+g1UDX96HR7
adT5i4hYHzl+reE0VxmPQ0lHmNNPeXNsFLD16QDhhC0Uji0bMemMGoqG+ta6HMQKzjhy2fk/TSxs
bGDHu43jsizaO97X9ZtNBA2JJGrQE0hpCETrVB1tT2FnCWaLE/TyMVGBrKd4LybVuPSZ89Ce/wIR
mTjxvRTqLUak26WRz8N0hHfPFFQRMc2p1HNxeOqNhJppt+V67WRCOZV5A8sgNRK7iK9LN9lZF0u7
rq/x7eSJg6yHlbHqFKODkjILXCHWXqzQwbPlanDw16ce8POeTd7iJNdeBIegWIn0hz3D93MUHTbR
EFgy0/tbyO58uHZqloYf3zkWYHDcS4AmqY3yt4/7Sk50Nnk8ameM7qUgL5LaALlwM82xaRH4YgmR
LV4gQboVL0jdSdPUdv56j3J+n76wfhy9CxyZe7s+0C+fz7U3LsoNdSTYIxpus/s9ClOQ1CZlkDEO
3FCTkD+9DY8hVGM0Cnmdle0mkNPvVahBzfEWtAXX2JGldL6lvWgN0MhICICp6SVJAWPd0qWEjQ0y
b5Rx4oS5IdKrbnP2VmmaMUsIsZ9FUPF4oZ4T6IM5QafgFaPydUnJmoBDY9NyfyXE/O2AZU32wsBS
RPz/doT+mj0eo2UODIinzoMzLaW2SjvVfzftTXxmk0IGKEmXW1tQX9/ckJmrtVIs220hZrOLWDIH
JHBGPPYc3f6ACSL/33RxzUDMp7uRe+fkww0v3WM4y2vhv33E61gPaq4m7SfhZmoXAvToP2gmC/LL
kfTaM4XCBelJffIdhsjsiXvvlBaCyTsFOYpnAlPsxfWco6wlGa/CCbllVxp9QgE95ud5LAPJ6APE
tDy+DFppZ5JlOHsfMsYvwp//l8Xlw1f2P5opg78tkN4aUMef0AYt/Lc/OST53+wyThkVvPgxWwVE
pO5f0GLjCI5lJGHRd4SVxJe4LeonFkzHY0VmwJvLjoMftiJrPJSJGOJJHXKXgwbcRZ/K+z7w7rbF
PyrqF2SLufHykG3gbVJDOHCPz4FBXdydEJB/Bmad1TVE38Wu4YZMwMYZlEQ0+haAMQ/I3rsjFm/t
4ZI2MzSzt9GkZosxoFVQMZ+NFORUoVFuWNkE/Mq71AGHkSKPUluuY526u8CS5IUngpvzzqulCd0M
TLEnvjoC63nmA3x3yAZwwFYaDuzYgqXDAIUn6MmDXt97/gb/u1UB49mYq/WByw+uvSECUW1hTU68
3Jy6KernAdL2OtrtRDCPz2ifk/2Y7FmsT0Qz+0FdGKO3wf0eBihAbgf+1NA7tr3AaYcaPZ+3xUML
6KTxaBAzZ42TPcwfdIs6WfTNfGoXFphdCTNJ8zBSI45TvOcU4vQgq/sY4gO3tsNcjpoikJ+qXIz5
nGTHPbi9jP1JQi6Y9unYOl4hpQW/7Kv37q7Towq7gPp6Dn/PM7nk3aHgMW0uB1aTzucu8HtJdtwc
nsyVRMnI898IFbUin7deg3oTvwxfoHpcC+j3b65japP+SymqDFWqxtt/cz37tDKsuTWHFNyLEzGY
ilUPplBNXIEMZLYAb80j02TzmHJq+UbS/Hh5pcVSPWgVC6dr4UP2AmyobqftI6ONSCtu3teEk45z
tW80YolzXwV90Hu6qVuf3WvwWP4apOQ8ciRJvRUnz1yzVQ7MTNBkh7rmg71geu9YJUGuwh9pIuUY
HQ+4koVPo1tbUZtEOmyMtZupCyJjVfIZot24T47FMQqdvkyOYXoHL2W/ovs4P49te1pUKEjUBHgJ
tuJVLrT0sE+o9oBWQe9DQkYucvS0DE9MlTDIiWrJOXeHp8c1wJGEC0Y0ciksXEgj0+1ql0w465zH
w1wNdmpsA9FlgH3J9QkeT0P5y0MVtpfshyFjMI9pW3KWSEnuz1FC1S2mWNvpSla9/oEDH6V/K+nB
mn2RECZSlYR8j4ML/6WS6wi8ezp6bhnD+CfwXvAFTsalTHXMaFpUyqAf8Eg93h7S0gb3JnqQJKt1
RQAURQlnVEREi7ypHcN0w832xPwyEp64MpK0ZnhWlLX25jPk1CPaiq2zj8Yi+kPoOiGo7NtbmrNC
3o0KF50D5oRAuvh5lzmyNv4qyVt50G+CN55DcBfVS4Lh7Z3rsO86sMgygA2jlfJUi8dqKKeDoO6P
eUI+Lf39oxGpgrgvyhhMIfNimXfR/F8GyPFHca/iQ/XrBsyICePafTUpzkaplhOop2XtaympX+gW
PaC3OZ4o79WrYgC/d5Xu/V7WRo7O7jnpg8k0+QXz6rtd3OQcuRQlgHWDi/R0iYSB8chXyDlD3zKd
GP6sVf1oLUlU6Z6DpTQQoEsBRSpFLrjBMyvqBrhu465P+HijDgqxxcI0QWCRxrNNwhErdZbQowBT
YfhCithOxyeRVUAi4/Zd/jUnfJTG3jawYXKcNocb6z1wiuIPiXsFoO4nRrfW1XZrpot7CzPy1IiA
5vUvd5v+MWJWBbjAqnj1SNzOBaZmyxo4PoKaDf50B11gSxZh1LZORQDzoIbHlX+oJyb21Q/7mzva
vt6SaMpttrmI+7lFhPy05RtX1i4jTRzpo29LKvEuWgQLV2GrgakENGhyFNSrjV4m/fIgMQxlXjpt
ZRcjfLcijy44+gEyiVvT4sTmLsyJl4721Y12TLmZRX+tOXkHiP39abK+/BtZss+cHQl0slpNGu1/
C9mdYQUy6pdpqYRQCfzSTP+CM1PS3Z3Adw9og8gLAfmn8HVJ3BncWk692xdAYQDaFMqetP6z7FV+
ddR2Y8Crz16WCrWnGIgqn2C5VRnXgRqmDs/1saK34d4tkLEFQETEiDZlyOfsTvHdmvEXv9QcUADb
3v0/+HfI1NAmbKc8YsNUV1BhzxrHrel6aoHnLAax3lEzLKrIrx+5u+Dh6h3bTWXGbhaxKskRF2eP
evqYQqQPqNJAsG5wxEQXgJYTObvbaPM+28Kme6vGVnMlaJdpEN2042y/dP0QTQS3muP+UBTXhgZk
Gyyc4zdDJbvnAdR+uU6GCmUymhgKILK0C9iMfkwylrDUevBBGVTjsscLU8A9kuffiQPVdQLRsFbM
WCDNMJ+Gst8yjsYcevtXXnzSOc/o/qSuC7vvEpajvg92W7xoEHhoB+xwfkve6E8mIFiMAggkjbIO
VBvW4GL2TQP8TaISFaCh7XVmrh5x7vKzduvzLq6+iKKHDu3c66We0X+0Oa9TL4sreFZJRMWJTjXA
5E0MdxfP55lqVUu1cIQftkMInI6LGsB22Sa2CjuVHbh9fM3tFL3o80EYGrlUDjB9cFDTWnJWjtAz
1nKvseiYpWekTjmnN5KC1DIAcoFxw2kOgc2zUUoiMOTBIWkQ6Hw2OvrINZGqxWRMLJbmcHh9oKFu
fFvqK9VMuroSbfxdVpCciFfb6N3Rp4jdZwElbgFY9VJxi8mBChjHJOpuZ3rMyd4NdjVDZxuEHAbX
osW+TPMkjWTJg5636/BUGDbYnMrIp7tVw5vUAxmObZIJAefHLBrdh8iOVoCR9ZMderjEu2jljY19
k9U/ZWWDeQN1s3te9I7aQeQZUt1zeWRIkJa9yW598oO8gggI/krAlHkRgTQ0dVzIO56GwPWuXt0r
/jeYBEBSSxvYoLyeAypayfByfQK+LnzUqsuFBGd3NfdlyeEWxEWhrUG8lQSfLKDS33isvMKNEdRP
aaDuaPtCVsoRiQQ+O72tEJ7w86zDWUn83tq89CTOWpxtP5FNypvc9klb1yM6q49DNAlqP39tSY1T
MygaHudf49UAQ0UIreSM7hxfMFMeynDIWEMPoUlbSmwun24HUw6/StJljd1Er8QJRC/ZD/ZtF2GO
ehcz/CXO5JiIhbpwcH+X2kRf4MYtRvgxyU1pD7rVU+/rBKbq2BDRRGOc9Sais13UUz9ekje4Pl+U
GxpzLhl9nZWKZLSIfXxyijj/7TRYjxQJeq+J4WzcbWVbmlHOsA7+8eu24OluQENOmo75p6fHwd6C
jWTGBKLq9F8OUfuebkDSsjm7HlBhRDOpbE0TyfM5HVBfKizeZ7J37WKklIqMJrbWf/RE9ii+auu2
UhX6lehBHtDNpmEW1UqvHUNaX6Vfy+M5vxhnu3wbcv4vtn5A0aIU0+4+fcDGiMlyXwG9FptF9WCA
uEPKsNzkh/1W15w+IvsdLSJuQ836eX3ck9dRWHVqJIf6giARt+9qzXmulUXUq0Vdv4mLwmh2WscE
zGZOYp2RZ3I0/gzX5W68lrdSSZREdSPdKYrRsHl99uyy+GIoATrgjXPYU5s+9JbEtxnjpn3MKakX
44G6fDIMwFfafIF7aldl8CQ+YgaQ7jXJTtyv/jM88HMGhIOtfWTL2KcrrzepiX0vWKYYpKtE7l3k
Pdu1BuZLPoxsGmUE7iWPZFN58GFK5Z3IY0fYynr+Gw0X8pkzk+rpcjJ9jkqFv52XcSlXBBLONAqI
nvn8dbiyVqFTVl7RCaNJMUnVrLKDSo2N2SXJReqVqugbQnSWZO7APVFnxW7pAvzKvd+JTfHms1In
Vt7a72yU8FS3EvkD/oAzaKwLofuel57tk0tbi8xN0ohjlpN2oIKJZE943+ZQeYezyUl5UU/yYJY1
pqeh/XfZI1XfIvhPPxrOguxr0oXDsByto/6bEg8YJOTQxbUE2+de6wuokABJEZkhpO7+u9F/+H0O
A3QK3q581CiF6w3r/oQpe7wiOev40bMH4IX7g0m8guGa0JZsMpZzbYmpIIHDh/Y77AP/cM4nDODe
dkPXuYSw4XgTtMOULGGXrgaUaOoof8ZrElSBzj9irsImsJtYbh/s6aXtqeYCydA3o1gUh7Qw9L0s
66U2cPxBfrzu9fhw/DdY1EjqmsMVUqCcF7xLDuOgOY36gAugVzYDj1+V9bsXBXEsd8NFgSSQM0c8
RN4XSuwr9DjDP2quTNU7fWXGJ7PIZIh+UAqgWysPBTfBf5eWBMlSKOcYK+iEkrUMqfW8eixAK/7/
bDB8kbGEw6J/MktbqN/WEtuay7A8Xy4Dq4wQLqb4OCIbhNNJb+6azliaOMAWIIE+gIque+L4Lxu8
iYqxwCP2hSwQiimxLIsVh2jrCVzvPMMDpMxM2/e1pmcifKoW7ofAoO3a+rA/p0R3ZjbB4U9ozjUK
QJ9b2HJn7g2m7aCgAE8hmX0QY3amzIUgF1BQUuvuWSg2zHiQubewHr3mnr1ykZ6hu5oUvgGLC1OF
rXH3YAQP2Vd9cIR30hVpIeuuFx1z7uFUYTMzJIPgJEIlbIl35c1HC9NJ+v0Df8x2+rwJO9R21tU7
79QjQsyl7qMrOQksAK4q2BGAQXS0jZ17K/GZhb8nJG9pc4WBU+HNvNJhGrtvBRuzArPZ5yyIjRlg
Vgdh2uCNwdQFMmocFP41d0lXHOUqh/KcVPfZ1yn6jkMpT2NV8FLaJpi0YeRBiAQbWSn+YBVQHWke
xysyk6B26saEttpzql0k+44zZuSEmGmrL743RMisVPfx20S8cfq3JFSa0TZYNSRN5tbsj5U/FmM+
M0ApcJa2MI0f+WMxS4qzcUNfqHWBjFLFkjaGZxMUtuPMcI1mpay0LXsjy9RniXXHRXFZlY9due7Q
vQraWD4jdXG+acxKUkd9o26/eMIdi1haVdr90EwFMeSXcYKHWTtlBSk6N4RVJjRFFKm6mHvXYCld
Oiju6Rp/Rfbis/vY+G3QM6ic37M6i4g/t06gTw7ZD7Ysvk8sOShQcfJhIEvvuZ41gxYuyGlnmASK
Ydo4zUKZmuNXiW/056bvn/76nVLL6Pv942uJsYhBjFFNMifP151SRm9vCsNwoFVBTrNVnjBhu4uH
LNw7Yd3eFvtnj/6fJtt/4wHyIpbFaW5r+HKrH2pn2IIrZ5m+mmB8kcwWoLL6yz7MEp1JYrYtaeqd
VD3VTrmgxSAMcjcniCA6ZRos52XiSNC9j3qGDDJrWKtxsrwKB7Iirt4eyYgZgoy7MeivMLBPS8co
McoZ/7Dy14btG6YpGE3gOUhTnSRAHIVSXd4SB1khMBsz2ibmWKcRWi8YuO9lunIqOyMqpsRcxhjj
1ctxFzxHvcRdqNsM/F1cqBtBAKjMv1CjaMLEWWGd+1+KgcdyMNDKLSr7u6Xlj2fzTVfRN6pxrErz
WLNlthM/OLH5LDLLHBaQCgOf1GCaZzcU8pqodklHadn6S+U6qPtwGFbhQv6dq72LZ1QwZr+K+2Am
y+to+Fn3UsYZjt7UElFiP8GP8Jgz8FzdOFdL5KOEL9uQgQGWfrE/SuHTSjzC9M9GJA8VSuv2522u
gasFlpXQj9c/WJ2mljPloLxGN3xT/qOKLUr2HqxLtuNRZEi9UoNpoBdldoL+m+XQENsNL5mzINIU
GYojIucuiWTrWAa63bVm11n1WWUVnQDmgHMTx4yen7jC/ULKvME/6qZsHJ9gb+1IpTzsSy6CKQAr
JnlNBGPDr55Ufsq8IU3Am5QZGPkJkVBIPjcW+VzzbJTb37cQzAOQI0p3176i8k2R6RCM+POMQaj+
mCtvFMa2byAzcFNjqCrYDPwBbC1trobPUi3h1p8DF59OP3+z5/KY/pp1sbKNKLaU3eJqhcsFIguS
VOrWPrxsHQHveYvObF8/8RSe5XR512I/ppTaAQ4fEePnGO2PEmHcjoGeWGUSvIZvnNHXGgDtKfpx
c/zWhfRjO+F0KMb63HJKy8Fodl00b1K847q4ExSVcDb3dpkT2/Mst5Be3+oDEpIrO9DpEil7CdF5
qRMYtNw2HNtIBq2+mQ793nulHPFzkElnFMlMN7dRc/l/L/x4sdqzF1thq8GbfgIvm2l8TtPVLBX8
5Q0X3+zx7VkDAQbZ9NFyT0MTR936Nq9oMStO+Lbk28I0K/WmPiv4dP38md0urfj9u6XPq6ZbMaXh
xO8/WjcgRDc4VIaDLWzOlnU/y8PNliakTp2R+vCXmRS1B87Erz2PQGUpICboQZVVGjCk1NPzNKNh
x6yV6z+wdxlvhNYdGNNyZwoY3U8QtFkOTjOBvTlAOB/SnOZMjkTY93kMMNOu5VpvQhf7p2pLzEaO
k7IqqHCTUuh0il8W6uGibET/xlZ3hwGjvMUQIsrtdwOcNqLA5z5vZE1JF/u4AG4e7jx7MkpTBFZ0
+K+h6O/DoOFN7EYIOOkaWxXTO7Ve43c9jsU9rqnvAxEvRus5xO2F86S57iQhESM3U4ombDK9BeC+
0gotPksu3thMEuHEHB5S+gkyGgnZLDCdXnrdU+5YdBErKhdj0KjGEl9OD+NAugFFynxOgsAjtw6q
I9K3y03IOez27FJjwlEYgSOk1hr+/693zPGFvxNBAwS/uhUNSIzaLBorksaJlNrZdvKdNWVAdTuf
u9l5LrDx8iHAiVcNGowRjeK+oH1yGN0FnmKMOkOsx2ktR8bP1Er4i1lCL8aKE93OynYgyQG0w4FP
OMVqN5aLzhrvjmE3wo2Bc+Gurm3svVGdMPZu901oawZ1C9hd0XpI0zwC4uQpTeC/+PUaa4O++Yf0
xZ2+M7jWdEV6ebP5ue9KtxCPNzw7yRY4ni+SWhyI3yGWLTtVKQZA1uEtTjiNylzA+mz8b5idR/Xe
zsTNnXnEfm+jMlznwuvIXRQTR3BMtqj3bI0xQL4QRv2/69wIaT9k30JjkzQxyjslvBRu5bdIPl/N
z7MWjUWsbusxJc3cUO5N8Dtuu/YPn8OHcW/+sw3HG9rNDms8Yq915FE1+JcB/1yvuEOu1FGCTg9c
VzMKQOIhLwGQKNzVjLk9nzZqz/Td9LrItNPVKYTpBRsGcw4x2HC7SosO2z9LiIJR7CBzkzlQPsTT
pwnq8fMbK76XHRbXHmbArnhDh4PSGCtNRaK5LPnrv76brb14sKZvyBJPB6m19YB8Ujv/NP/cB7fT
YZR0HIBz3mrJhJiKl28wekqr5ad0mmvjp3Agi1NCrbgCrjeMComXdorNhfYyQYe+vWbenXgCiX40
jo+HptbSVy4VI5mpD4Nseb0j8iUONsCV8uWBzEgLyZP3dOyEDJeXdx+qAvC6kVG2Bh0esXbxWZDS
0qj7zQ7X9DaOp9FNxsMhTr8NasFM7sxTwFamOWtSvc9obpI4xQ5C39Pt1P5PzGr2CdEiXXoIUC//
C6cpbtS6kLj9Dp6dtM/HQgyKRhtMSUsw71BtJy3WI+j1dzPXMibxQx/EQ+tatlyUBopKMtXaFc9y
WXTlJSdrYkc62AsQG7GE9wmTOH8Ftk/mzxbqSUbnyp6Fr5mdcp4U4EwQHKTCVghbX0q49BUFTmKq
+OlymCq8ZBkEynWjtDMb66ofAZksgzBr4vTFYcn2CHscF3OevE6WDosNILuA6ER00Y0vvVXpFJ2d
VnTuYO1BobK2NDPWzpHbrCsD3dZ5L+ejkj8YtG6mvDyGlyOScFf8vGAfl2/4M6d0WinCpyeQTYMd
4DbcyMRIc9bI2Ro6cxl8udajVdASU0jC4HmUMZuY9hzwnbPMST/jSPCKp1gUQb19fLUdCU9eK0Md
XQZ3nQytKCdnLCoRqCTC8c9X1XL7fot6ASfN2L6W1CkGOtBTP2IHehQzoPz7qrgzthjp3j5ArG/j
inIs5cbACxLe2CMBzz5ZB/HQD4SDKFnXZ0vP395Qw74SFydRw8t+/sQ9nBWcj2BQy+OxCc4a+Dr3
QQQU2gLfVd+DvsE8wMIuv++ARS/aWCE0VEDD1o3BSWrYwWfXDJ+0KHNOfmd3RzNetRq1gowaBhBD
7nAuzO5uFBjalJ46Unm80jpKaL/MLS15+nX51KwKrMR81Agez3AI5pWgTQ98SweO0RwbVRcEFCwA
PcTqF/5cKnH0oSzqLMmHBcD0XrY5gIkFy5is7xsesfGj9SLVe7JyWGqFs0Abt6zDftUnD9j1r4uq
5vTi+Jo1ervj5DKs8yeE0cgJVJ3uF2rPN3c8UNabqIbysSkUNXxU942lEMcWBKqcZxyn4DEOjpGi
eZSS+Klfqefn3t/RXgBMTwlfp4VORnx4YEeVCNsA+XtcG/cwmNxCfF95M645qgemQhc92xDZNd2c
1/kQqh/OYn51lhcCiZZWf2fsb3m/oK0fjPQEsT+yZT5hwE0F17gx6pyKNyXFoBHRPxzCaEYzZ84W
AdnIay8jJttH+Q2ESrg3EhRGX0X7QqVobflA8a1/cy9SdjRZrWRzTLo63s89fY0I+sGRd6H9iFxw
THoxYE5W0B0+v+E4izAX+FAGSEUNX9LPaszM+sC62lqtdqSMQyv7pmx4LRx5f4PxlkUH3MrMU+DJ
2gIdtGnE2XdhqVjEdR3htIalbM8gY/58woX3a8edQIFfF8BHg6vtG7hoO1Y6Xbsk5X4/4jRuTuPC
+Dkxx0bvm2imdRlSjwJHTh4fCvXJYn8wkSoaAUPuDSb1NKufrnrcM6RkFZkJ0WMw60Yw8RmWHWtN
WQVaBIW23aODMbvr9UNN5yUIlU4DCa6siNIFcjynOatHznX36p9o4DcaicJwD9P9cNl8xlQXY+Uk
nXMFpDs2QCQ4L/353cgphLqDm4PQM80K6HJKHXR+a20/QhkvflO6OWdGPFikkX22dmGcW2ZDPekG
K2FsynxgcPOsh8wZ/KHcdB5cCf/JGQyKqeIGBG1atkwhqn+msMYYCFPGi3ad7A91DcavBcnnBo4O
0I6Cn/Sm38tnrS9EkCi5rPpFiFCnQCDbQoKIBo5mqE1E0wqBUAmJ75ZtQc+V67rMtjBgeC6m0HGV
WjR1JBa5erjOGsDKZ3bdIHmucaS5/p0cc/3FOdYOIgpB96YGJ9a2EcN0xiUlO8oRTJ4lcGXdmGm7
rk2xjvzMgvntZ9ezdjhBDOE+C+9OcrCsn6ykUEeQep6LMwRMJnHnxY5OjdJaDnxHSeo0tGQ2lz22
GOWwbkATM3js8wYqnCCthZ6LoECUMQ0fKFIwqDrMSg1oH4FJOIWCtx6cuWE4+TtN2IF3LBPSHUNj
CP497+/+7c7OockEF6XX2iTQeDQR9v/toJ5PTlO0m2JXf/kG/WulTDZjmawLSf/qkdtajtNAl5En
lN0hMSjdas8bvZEeDYiT5ceY1RcqNLdTJ2vfEaAz4dHuFgfUnBFBFMJzHhJFKFQ9JTv+njiOTXdn
mk51XLcHig5juS6tAlAbvKdhpgMqkHVRrUAl1tI48XI5MdirSruWjXJWa7f8f7yMcEK0LZYKCBgX
hFUKOp2CPO8NyYFnn04l+0pQVtK3dKwPvQqGbWcDvI+Z7ZTUgWm1cgMCpwX/GjFFowIIC0hS/iCU
5DkOG0JkGUlUw4l5F30ruS+gcYgUGO6E9VIkJM1BtryTvvZaqY1ik5wxJD/PD2thiS8enCqPlDCA
nKhmMLsy3EytjM9gSdOrRj16NHqI/7ZqWyrGqqTLQnppUJcwkMd1pCiOa2i3oaSMpJPRfkFmhGk5
tpmnBrmvOif5BVLOkhAsIsPdRNtdkyyr3FCA/CwT0TNouANtBZtNqfUNIx3RPfr5D1h7r2LPEcjB
mFzPwQ6EfhyTX/wGxEO64374Ck1JRNAzbGJcHdYC23QgXHu6P5zSmW4c9gDE+Y9w99FW0OMEQNz/
8XSOItqTw/OkiSdYBy4fVMCc4iW0RJvcronZ4lUBwWVUjfbhwN4EcsfAcUzsXvwSRhFubtlx34G6
73DHveW5L6sNt13x+haIrfT64DcEJJ9ePUoNb5ckf2PaaUPCeV9yEfE6YJVwB5R0J2yiy92bg3md
a+uXM6BInehHBjmhVWdoigmNq3mFkfsJpByiznkDpBqV2oSEaKUiArgllexeIXlHLOUArASyuy3Y
2OevItNse16dO6DPb2bsvZpUctk58diCl4DkkU6F3i635J7QCguA1ae8xwkRTBWGE5yj722aloaj
UdHuI5GSNufbW/ok7AGIYhVSM+I7j/MG7px1HdjGqdM9CQsdAdR/SciMooGHAal3/z5hi0d77kUq
AAVBgKLBo2swlaMIw57zMZrlmAJMT2iARMpVRTq6/NWyvn/nnolzAFDa1yzTf/rWF7QzVvnAzpam
U/gZq+xI9e0Qw+mk6L5ClS/jbdQNcnnL61uqyc1+LguhFf1j7XI56LgU+eYqMMiFs1vhATzFHKlg
zXKxAGloRiUYWldBaRFpVRtnq/VCjTOp+9Gg+WTGU1iNfwhAg/vuwAK2VjYQ+6Yhduw5/aoqYLhD
cW6PWLEPSVcSh03BVmvj8KSdW+C0T/OY0y3+M+5LB9f4mv4QgP0m3o9KT8yz/I2WHj4IJJh2MwcU
gxFy/gN/zzybl4m43NrTOM30X/pNWvvyiYQs5b2e8EQJeoUWCzHxvxmciqelw2XFmlQjV2GJ51zQ
Prf6Qh0mewQFSG73KEqfHwwPQG1NXzzkklbxo+6xL6WgHPphvNaCiqKcj//pZPrdB4u/t4jWPHsx
ELOrfA4fbkD6zDcgW+GMvYqFSBQZHXUxF+C/VP/y9CCaeBSwKzrgLcNPWBT9rmMiFryrZaJFsgXM
kLFSfWeoS9cRItRd/np2KjTSPmdL0Dbk59grNTMVoqh6+3uZB5vT4ZXSBcDdV1ZqduJzhDT7d0t4
k7HN5FqvJMLEUt+baLQKIQmGYXCnf7AZPZCTIsYzZ1I8vN/kakO826D5oix7zM3a2JSl7vH3kk3p
RiuZ7iO/7DyGWKM8zStaCR0z1WIQIYOXGxnjjyT/lXB/NqYT1+6j97rpp7rycA3185nEXNubSENi
1JcDtf2DzQpqQOrAPr/f3HEiQNgWfI0B9c3eKsXXlTkdkpqPb+kbhzpojbxq+PAfHXfVT8Zh8YAR
XxOO9+EDywL7YFjA1nsXyn1OELGOwMbvasoLvr7BAAdZXBxZyMuXuyZNDvQmKkvv4/aOio7S69Ck
FCcwutANyorD+1mwvC4XS3eRCkSEBGEhZhsf2RDrWhVjIznY8s8mr7XlVlpyCPx3BTPIniR1/UvT
0OLlA5+yCBKKSXAoI8k8wFpUGimjIrmxmoq0mz5wxXdFwYv9K+XZPWIXx3ZGz+Efr5wZrSnbbpFl
0ibsrKpGg2gjnBzyWdrjhMFz4abKcdhTahiZV69+vmp1FzE4SB0fYxwuu6/gli0RqUkjAMNTEjva
KJ62iLu1NrKRqQt/9JGQi75pBUTJHkSljFwXYsvcEIJZvaJjGlYftcsnZt9ff3bkqrfOYS1e6pAx
g9qdsPXfnZrRYD/UmfyUUajBIpkIxJQfb8FKOWycu2j4qrIA1UE2wvr9udHnLYOcYWvJPlX8TE2F
i6MXTzO3TbUBMvblAsj7RBtpQeJEssLK6HkRcro5ojpT9n7DMS/dMTlZsTMTNFd7g+qQFGe3IkSz
4BahhEC3a9Vg51/D/6MZKsyF8WKOkcU8Yej88yhDmaXRolEmVMIg1WaoROXTQCvv5t83VhdY3nkJ
lVngP7AkTj8zZ59OHM2oUHlGjJ81byJG4aikmghblLSg7PsK5RFsCaKGp7Oa8ogzzaa/wKMx62tX
CFROogmaz1W9YuwI/SmgyimtBycxddQcmWjI6WzJYiKjOZcji1fqpLf9Fbt2EyWd/6cDsk99pVlB
X0jKrAnkXQLHyTCYaupLMROCl+/goe6u6vf1Acn+7r6MSP0ZXHMsV+TuOppDDME00oefGqq0rzvJ
LrJM+Fx+bNO5NNCdsrmWr9jQ15ciz+s1BvF/u6A8jbBFMrYAQPMOXSn/IQKcuCJjWBeY/K3fQ0LO
CAY9SBaoT1MtWPzPc2xBdI1g1v+z8GQJ92Ibq960jVWWhdi0DG7zo/sqiMfNv/BLTGnKo4aS/qLb
C6qTM/afM7QaQcMt+kDsIj2x44O4CgMbwN6u2OrD+3oDmtEvNN/hHzCSa6LX31+68W5CaMhKDNxN
AhSMQ2CKXqspfRY9GUI07S2ZvbOTIYjeMSn4ax2gSYAdnR6TwZhqioqaYfujIFsuHkiyI9xTH5Nl
b84F6jRxoJbH2vmp9eb78hj5PgMar+CstmfZjm8bfCzIn5hMUOf1fAi1QDzQAEErB6arz3h8LIBL
gDRWaSzAli4dly87TRG8Iv3TlEFCN20OHlhWUsvRjdXL+hbnW6xDFgdZlgkkZ5tsLVGGNFSiDIox
Fa2TAYFC6w4fJ68VPaFeW08h98RW7bUuOrcbf6KseyfnspYi78dmG+p9h1vd8glXRKFLR+tXdL5p
MiQsxhLJRUR6rlzPYJWKr2AkDJE4ufeX8ESEw2WcJJ+eVWjuSnpL5m2vDKngzPvKkAbgRNmIvgWh
2gMXB+LB1rZxSHB5rss1uk/nVjnj05KCLuMxxMfTm+7og9aPECmgCJgN1Lrrjj0CkNC9GF4Au6mB
4KZZeZXUDZJQuBDJrURzsG6kKojM1MGQQsQH0ZVp9buj7wuUv3Xf1ZWTkGn97dOg0YgnYEwmvkAX
FekUBFJGRGaCSlgrhNHCII7Ot0fbdeaGSmmy3GZIGt/wyCgPj6Z3cQ4yhLVtsRYjFTbTCieKGNR7
2ZhuSb874yvYPjN8ijk4BulePudQHSfUC31sbu8NYeavZj5rouLgEbHbWrBfhlMOzJLgpchBIJIg
O7Tf3xHyxuwQJSYH/O8gCliXgKT/fD4/xX0SR1hNs/+q9BjtcvC9LymlPambhXII/4UnS0Y8MN+o
K2TtCrSDJ7RpIPxQ7aRdiPKCrXJyOuKg65C/5q4LPr+b3M1fHsd5itRj7o41t/SB32AFdnJ20auV
ig9y2Ttt9HPl/ijV1YGjZU81596Khn7pB6nkDc5kzBhTBS3hdBXPKyMzAPP4+ggWZsphic+p6H0p
2GurANTdggn6iDEGfXqPmHXX+GLDa0GvOteV19i33uaLD9H/gJKYeBfyNH3ys6k7h+FWB1RIgJGg
9BfxZVzwHX855M5A0q5i4OC3M3zxaSIJ9WmC6CbYOEO5BjOYmGy6WvThEoD11c1gp21l3QHhYx+R
XK+TyuhaI6xXWAtMMm1c2UqfFbMIEg4aVATWVW0p2eaPys6T24/PaTb+G5EuD4QmLEc1FaDOYBqg
oRIL5HrHgXFTffREUIHLVJdE28G8+ygNLbE2ImFMKas4bn+CD1PQA4ZQpkXNVgkKcbmVi32JWUm/
cTCJsGvtqEPnoO6byxIN9EM9iKxkjhRrHh9gHki9z23vF1S3ea1Fu0oM+LUyZ9kT4M9A2pAlYhYA
D5Ro/RrnpFnUmMLxopBPvHd33Wsli/moP1Gj7FboWXHxKrbj4z0huwYGLbf2QbRgR7suT98E7OJ9
zPFIX1cH09DbFJTTs34DQL85d0CBgqmZu/baZBAFoy9nK2q0TBs4azYmH2iM/R9sZKfZYSeUoTtU
2aaRShyF8J3jad6dyYtS4HfTWk7G8v+sOCgOcSRZ/uAX4EaMqFhp/WFOR7GxUKotqpCBl8b99JYC
hsWGv6C3a5mNHgwZB2u1L/pANt6nu/oD7VZJSHIirQ4kmdiVbSYIFIxMXD7YO3DP4eUELFEnjGlH
3ep0z1mMmmSwXLE1U4t/nwouQaCjIvKqEK+vCDlgWpCV1UiWjCPs+TTYH8kgiGrv4FqdRGuleKT0
1NP3Yd1kBNESh9o9wzW45NYLuOfJ8y73zUzKi+0xCFEJtw6PtrLgobHWKwWDDaZKPh3GdMnKkFwa
NLzQj9pqvMGWPvI4Z++CUEbBhaejhgO0sxFBLDNV2/6zfZ/0Q2GVX2oQHEVnTsbXSQUE2bHtQIEA
1Hwa5j0B29UZyvOxKCIh2BcYOrxk0NCdZhJy8YYBpIqQakmOG2EvKT2+jGZplOfixXLhrfW0J/bq
xmHFokOJEJliPcoFBvrFmRUN/uQhNZZPZzJr1cIBWwgdh8yQZpztaAeG83T0iWDrTyeQ8DdoYp/1
Bjsz7w0UctfNNZ2OetH0eBuWCNomOtEMmLGyuAYMN3Rzk4YN7px1j/g6/dE5P7bUK9aKqyuwqPY9
boKjW/Q1JK+CPJaVlogDf66rBo2UDWSMhlj6HiFHmC4BysHzfJONQyy5zJ2TAnb1uujkuWQnbUHI
S8EYZ072ivZtuU/IwQTZ8n46vBv05AsKMTdYbfUMOO9r/byl742CUnyduVfziZe4tAYr6S/Wxnci
Lvj97GqyAtvmzvfcRWwFKXDFhY84ki88mpCOT9zwnwzK8n+W0Hw+mfA1gavzGp9WC73efCjTou2W
X6qeTfqaQ9ZF4a82bRJslen1Pij6/6B9gyeF9hpzc6Oa0zfolIzcHLb+2BScgbkFVjuJy3lCso++
nRV/OueycEthkQ+BYwOaw0NyVCg0Jgbes5CdZjc8QQaulNngifArn1VCwAfcCkYOvt6oMsWqoRty
Fgg9GA2FhuP8gu1d30txttrio+sMF8dwGd3iOTbDxcQoxs4cUsDXYD1Ay2qmTK1WSeV5yFsft1+x
ENzw4QZXswAfIGhFsHk2p/nvYA6EoPTAvmLFvMDllG6wR1Ik7AJVdNSQx/aEI1k096xlHxTncDL8
uCiKuStDNE7+kDJvQR2lcNNsjCOMwqqoruOVqibVowKweQl3fT9876Eena2ROuxM8cnfZHxcy3c4
2M3r1snEsdXTUg909y0wG/UAu2olqvF65BmbaMURcoVEs0BxLpW3fdJGfo2GI3Nfo0iZDtdB65vF
J121MkVwAdY5XVmLEn8X95qLI245Ffz8SYpJcJQJdcxATOgn12qH5FrlYmWPzR9BJ69v7mysTpO9
Xall6tC0F/SHxrMQilcfhy7WQVaYqPTZFEBfaL4oKm/CCkGeubAQ8w0hL463esf4Xr4FLigMmVdu
s4RVp8KyyWEvdtJYou+wIzEiQEf4Pa2Lbpa4WDozd17pqTEWrhLt6vvdty/ZF+acFltyfYbBEhUW
VTxU6OYI7Cv/cvIOCYa853/L2hszbIvVcwnCFuYecvJGvJ/jmFwN58YTWw7T9BZj6Pc0v0CyQA48
Gem1QPA1JyZdCFY51iY9bD1AXOtWNmyi/gDsoweoxhGEma41ZvGA/oyjILOz9Nd8kQ+ydRZMXbK6
8won9ZJ602DyeZ1WYwNhsvdPnbROwllWhEA54l7T+kly9az7L0VavUhRpyjxTjUb+/yTKH9t3z8U
XJM86hX0HGPCP7LW9O4lotOC7B1AxScEt1/16KgASlrqMKmLU59YOb3nhwuvKnJv8y4OXxRRex7e
p7bdfLq66/EgPq9G2YYjnuo6tOtlxWR5BCBnu9t4fotuVYkEXiNX4ZCUNY63tUJ/aZv2Uid4/Yuo
absb6BLZoz6/CBSnu00QEF3/DBpqLfkNP6w9adcFVKNsKT/cRW3AzaD7C9TP5poBYPouWi23Ejhg
IjwG++EYQ8ToaIYAPAnq9HQYMPmjDIpNyGwnJb1kr2tkntSumZO4P89TMiKFLAc9+L3E21zl4Mtu
8e458n7Cas8Clz8cll5rHMIyizbIEC2T6O03bDddKYOzffqlq5X3iXYT/rHkqnIu8kY6MyL2Xllu
KhePjzr9S47gMKrUsygpIcLLWPYhxG8jVA8SK5JPeeCxqviZUrFyDq/h/vmQErpMLipkBEDVsGWR
fFCTCdYd+4a9+fxwCq2JKh7gB+GZZ+/Wzp9i+lWoUz1C3n9KezCylbuhACRNdcG2uN4HGkXZbav9
drDWFAeaS//8Hh+HZZi8R5kGDHxw9wgyZLfz68y3+CXpKha9ausTDz7Gu4VNrOUw98R6wwB+xUJi
MV8zBQUcGeOP05k753lKi6L6lYSSZrx6zRB0wEWx80sucHgg9NPKLAOIvkxYZl6m8aP/GBfkTXHi
2RT95uIbayohDxMUF0xGzS0YYzHrZNviydJCfL3fZMQ8Q0PRO+elnBcDW2XEPB6BZz4NR410Bjp5
1crxMzSQMBE4dojFJfFXFxI8a6jBJmVU136mrunfM3Ii1ITgAzUHjt/fFERm3eh3pOVU4LgVyWn2
Jm20h+Ov2kwLhcHDSDowkEZEZu0PnJ0Rc8uhyTK5ML2e4JORsaFl38a+N2JlCMWlBUV79gBks5kw
PNy8V+DgOehikYfJBQy9XCbo19kIEki+pX7iVOr9bg/j7N9kxAmpiR/RULtcdZ3graHpfmTkQEFQ
siAZg1Z6d5G6MYLt8cOFUgjlP6Ac2OR17O1/Bm/vlx+HurlNrAXPa3y3vYy3sXuz9iwmjMQrTJiR
lCMlq4P9RRR/xSroyyWs4W42dGgaRx5Fxw6v91zmoPWDBs/qCD8EATAOR0H0oNKFvPL2uVGB071J
TKpPjFhSYmNfUZzUQj9Co8WqbeRUnw/5QSU8yaRqLVijIrsfsOmrM7J7XzOvvqNATn8fEfG6I5Q2
8mUoMw0iHmqd+SNAzaSSQRs6NVXL1v0HeoUaDC+0lFET0HHzAVYqIrnwfGC6NQeu7WZECEYj8lbW
h0uR16p4dicUQi4uBZXP2J2SkBaUiX7pwYeqGTIEQrEd/f3D4kQ0wUGt6Q1XdlRgdD0wXYyb0GOH
AXrsGZyZly9uYMBNdIQlkZKvqVAAovF+GkNHzRvDNnUBOE/VFSKFjGTT65paS3X6iCqOjaqwIwYl
9ZvCpWiT4rkwFRMEds6TsM2bP96JRjxStX9xQoHxEu7fvJ8Lga7MS/TRVqM1hQLsUbFCF9vr5LSv
5n0oFlseJjiRVXsST+NY6Gbe/RZiGHWHgmB7al8SK/39QlagzStqv2CAXzG7NPfmwZWKmD2PwEAU
dCGX4OG3aEKZ9vnenTcuXlDHG0ZkHqey0k2sa2RFiArLkvscMalcGq7Loyz4BXIAZGlqm/l61gJg
+NLOL1XSfImuEWDEIxsJzqM+GMMiOVlLcfcnOI+lziaFSV5nqy1CS8dLNsh7YKUDg+Nwv+dpET7G
fIfXjQg7SxGXsdrSzXJzujIeLoAZHhOZnDkdCgsalz4IZqpXfqgeNba6HDfAUyRIGpy4ChZo+D7Q
GtDMOqkJRBR5ScP6O5k0KcsFmEz6tiG1kfNiofUwXW7nC44P8+eUuulk+aHEu6RVwVAh1bzHr1eX
9fg6LZajAiY7tkvempnVwjfm875wSt1MwGntz9X9YfKrM1u/CQ2K0ShLVJOfogwYtalbx8brlE6g
5oWxDBRJJMwlzBeCuFVkQJ3DTxQP/mHDlL3qGoZn0+ZkAcBbaoIc+SPxorQdy1D3URBd0wByYXpj
zfpXAeeKXNP2JIrR1iKfLFCx8074sX/CknR0h40TDGk235mHhvIpy15pi+Fk6UEceSKSn8RHzexu
IVAm1cJwA0Y2tWORwbnZ9qlaM+/9X0KCU8/cUaK96iKWcXwPBrpUxTyd+lrG7HyiU6s/JtU7QrKw
oaPu0hX0teAIzkTFA5NiLSdeWvV/5mTHaXNXGEZDQMNwT9VLDnSDhzzIswcLgPxLEUZZX0VOxS2f
LcBdhh6eu5+/qkY9QGyfl0e0UQx2+2txpN2BmUvJekwDqsv1KLYH86uOp++mlRiOMjgBksvtKQww
QAmDIHx3k2WNPC26hRb++1lDdOEqoHBYCZPn0opR+NNzFrXlWZMWSjwxDwDE8l7V0CNXrCDW+sHD
YBrgV1XWnaDDIV1jn7PCiqNVa51ehavycq1Tp0vRV1srZdUD+wqiCuIQwleCKt/4yOcctGf7YcZA
WVD/NX4VWSHMEtiCvRgdWmR3blMlsGNM2uytzyvDDhMK/fiBH34einXv/okhjLZJNk9iRIPiyKtp
onxn5PGTj0b6bT7K4mjYBaNk8bXao94KEh+w+vkeGSskw4DKphbR21on3h3M78t2z3U8vrHGErQe
M8oTW9mrdBLgfSk0XTBfFgdkCgZ0EzU8O84qbjEGbQAhcJvpBbO3U7pE4pcLJIu8rhLRsbfto3u0
50avLshGUkpRt7pzP9colRGwvRu776BMMGLhGGbQPd88DkOPQY0wCabrcIUV2UZYb8U9ScI5pJlI
y91e5LeWM/3QUs0rk5xLjMw7nVSruNymcpyWQ+doh34KIUrxepYFhZ+7X1AZUqr5GjhYo6aOi4KO
+/I+NaFk1/lcZJtIa72yCHZrXmExsm+AFNP8/lOiA4BIXBLkj9xr3nCRijyyNxJsTzFEKtsUYhkZ
HoCIPN46ApXQO5VgKuP+m1nHgdXQzEVL0occYVoTWrUHdO2wmS4WBXK80Krt35OrSvgtOSR4Vbnq
r0HkLiKnU/xdropxQ7mcJJvGcz9zXnig5jxpsAFpNG8bygzkhGS+oXbyNqHfEX6zmTT5sz6pL16w
noME6vtmPJeWz8JttZmhR/h2c3/Tp1wzMdxOGG+tZqpbGCXBQqBkTLecb5VNey6mDByhbH3GZe5R
e3xlni2/YGlXEbsxrgS5AwCyjLeU04cMgPIFq55TgHs3pHcoTcPezW3bIv3bhdvswZlOwf1z250N
7AhOtSibnvysT+jNu6YDSreqDOUwyPSPeg52WG/yWwl7TOW3y+SnWOqOj/eAEFLDcU2OPHftepFo
1oKEYKwT/yrrKWrE55xzs0TouPLfED1pKqONzKVRid8McI20HcEQ4lWIfS3joATB4kg9FgovxLdz
pnXK0Ovo+xfaxvlTYvaUinHkhSt+UwVRASmBbOjPXA4BrmrBxNOfVVU/G+ysF5f8pKLR+9ngrF9K
GLRdi+x3mepPjDkl2IiXaR1EZXPZBDmAH5nRRKIZf3zb07a8om7OqIA+APfMUoGWDZJazuORK7ZT
gsG/uBOfnxMPRiGBFXEAN/lRr5nwWviowT/AeyBKXasY0p/gIEzippc7oMtQLrdIAX0A2bUADWfs
KyykvV1iZS46WpNRQpWUwaZizxuTuYrgugoxjAJcoDudElQ9769ZTthhxO0h4DWHVJbHDFq4v2tY
WkC7I7BAmIXDXzSPKLqtCjct5lBWwA3nLPWNgQX4JFngd3ZFLtsrSlVJkSE3PwH7QlRAcZ2amh/M
ImcJrWwAyHAD+rWhVIfZLneZZUiWNUsYiSAWEnqFpMreJ468N/+lGnVhEsr22ynxF/xYp+rPfj27
/qeU8xnka6vOQj81/XVjKg4uXbActcexFRVqfvaDPe2rctPVGznkupkWIE42rdgNZmkmgpHqS6YI
Uzfex/TzHISWblC8WUaz+TKdXwQNLbhhRksQpgP/BwP/QmWZcF4g7ABywbqk+TA3KMka0GMQaUyg
1BaniQWb3W/tu8qTpiJX3oyoH6MeRXKiwA0nrki8bPR9fv5S4EpqdhoUa3gn2tfY2bjLK1PkWKXv
/rf9FSLD+l4JfD/WTkHr0iLmNV+nL76DN20dvXBh8n9uIxx/j8Rprs2iBjBGx1sKrJOID+8H9jKd
pJQTeMV2z8jT9pUOzMD9JdIBxtciRzqeY6gL1oem4K1qYr/p8qiuL0kvZ1cTJOYKZz2JmqQZpaUU
Xe+f3J9KWuS11hlqXc/8qGSVCAaDA9r6EJeq+/YzDOz4ebnXAfxwqMbUfnLAeXMSIpYutHA1EVHq
Qz+V4wZlS41LEseW7Hnp36HAvDFqDLmf95dKsjvSTwVX+Qf5dVXzPoBGf/Dwx65C/bviyv8uaw8V
PLb6XsUsgotqFdkFO/ARBhc1vpXT4aPkQHFGYfSckzjnoLq46Vr4aeqXr0aDfEim8YQJScJG/kA+
Sdkiz3A42DbZ4DGHJzMg5vgaOmyxtLjvFepFoc64Mo1vUPjSZbQ87XrWhljYYYCrWOtMVMLMXV0T
pnfxO94ufbWiv+go7Q1c9aA5hkbhY+M9gCmz1cfJTqo5ucy203eBc6xRjTY2jKVDp+CjCqPBg4mA
RQj4yjaYQu4g2pu7DaExr02wjMFFy86piETPKkJ4SxzAN+COi+Paj6NEJJFXhEOgReiYGqvvPFkl
DU2lrOIhZ0mPx5kymLlc86L021/erKwmewkRQNXDr21eER04xsW4Dr6UBTWYmdFw5gS7rNjcjS4H
xJxG6xoHqrGKKvR/7axDWbex/EiwFootJS1wbL3tm5i/K2OkdyKumBnDww8k2yOHkA30plw3QXD1
M9elo1HJrsiG3qzTfk+S8IbaJ09juWJLB4yBZHSFGbULXVKKz/Rf92j4TuaLUtC/pFT4N8z03x54
GjrCQdodQelRMFofrOt56AMT3AJ0Ullpb49dRRc6lj8Y0EM+rY8z3qJS66u7gBJ4DiAVWbZWA9NK
Zohj9LJOVOlKZL6uv1vBPosqTmD9jUf3CkwL1Bc8N/wjF+R12/5UWv5sGKx5/OSjRBudK9BJC4Em
xQH1Tqh2bCemqBakxFr0whQaOal6DTi7XhWCS5g+mJ+3ZBi+5t4FGFQSotRTZrZp0HZMqSekCX8t
hJYHhvn0/CLuYz0+4KAhpy/5Oj53/haWO7kokO5nYk5rirSLGj0EvQvo2NUeEkhSJIBF+ptt0qU3
F5zB9SHfRY/15rK6SUsZbQGMDyHw2LIP+yCzVq5nmp6inuSnCbx4vtGuU+o1+5i+vTbBx3nO4m1F
zW7jU3Hd8HRxMmm+B8csCYp9PglLrggN4PDB+XhcYqlY8/bWEsiBkrGHSRl9/3SSCAzEL1sK1lGE
+NeXpJar70uk2rba/cRF2sNPf6ZmbfqvyWofH0lyWDrZV8oJGGDQfTp9FuMqK+vbksQrgrMYVRcI
Rui9o2AC7YPYrOTJgS0/1y73QSrtQkFFG5WuQbKHw3MCLUxykjgnSwU3nNvbmndX/hNPgN/bWMu8
4dktB8m4zEhlnREvGHtJS65AqRGEALnCiGdQJ8Djxd5OOrRw8NPMtdlmrJQZfIPAbIRvHc0FLciT
YjXFT+JuFDRfRO15Ag4MmjsLBnzqjcT886OhGYVh6E2WdsWrxfA+iMhrteQylBMjzofbd3MDc1YU
3n83WnaO1hbsvjpged7FXwPSWoxpQIiOlJzcbs/bZXPu3hUdHjDNMATijNUdgkubbhDhMJAkAoRy
wWtQDRWo7BMbCBjEC28QwGdeWP4VHRwGlDqOFfPdartgMM+tIrUm3JmAE8MT+6qALt1HEi10Y0lJ
sw4Ex0ly41N7qGFi3re7IySzzfhqi689goNs5bdof5MsF7I2F9QQmNUKamnd0mHnIAIrmKVzjM/M
h/BEtwMh0X6tNS2rTh17dSQzRYEr9/aLeAu1HF37DhWdrXbbTPjJuHUxWePzMqPU+XQNK3DDNEPD
UMCohavCE3zFSixkA466VoUFjlxMYy6l/VYSVYU07ftVI0UnagId1ppkHjs9bZrwx0bDE29AI+wu
ce72N6uJ6MVHYR6vQGkVvF6SV4iKXIaH6bgTybMoV5/kaqkKjCiwDrfk9mCyXSsuLr9U805hTwUc
YqQp+Ir3jre/5GxVO4TjNLtz5X549npdSjw20LxEBBv+D2PWRaI3L0ZnTwQ8O7BQv8ISTFc4lrvn
eBKVjJOMFrVmSs0KFuijt8S1jC+kql9pfHtPx66ix45Rt7Q2k6Tr6eWUc7T3bjNrR/tBRKM5FEAs
81kO53VN3QsZuM6W37yDmGc9klCFcU2EqzoeQvsfldxGnQheGS/QAir7raopDpaRWTtZB3HwYryq
GmWwJTgR/dJ9RXtXkpvwmfv0GPrlD9jqYtucxh0KAogNvZgXO77aXdl/FfBKz8YM4dr5S64v8iOi
fZPXaCVSxY+SBO8rm/oLnuRHsUZxNo8TiGh/6bjZkfVf88Tb3PiTkkOgaoI0SwA5tbOjHrEAKo3J
UlKBZAt/Ai4CP+MDrepjE9CVLOAT0uhFUs5+WzQonLKRXUStYZZ5G8uypnoNSDKiDcIBNTKn1b6F
2sg8lXNxP/zpUX1L+/15tbyGgogZ0xgKsjmt93byMlVjBPzpfu+d8B5wtA+Bz+FryvCrBnWXdD/A
Cpl0BpttYgQYXZXO8+X3rWZT9+H4OsfLskfkFthocMjF1ZSv6R6M7QYRGO6TjhDf1f/WFvvvOO8Y
jpWKBZrZdOyaO8CJlpS5U7xAuR2GzIFSFKeR+bALsriXtX9aTMUbg+HQ1gtzMC5DDOnrWwxsydHG
PB765aWwwircN+QiT+Qs7D9bdYqKfsR1Pd2ID+o3E8iVFDaHlWNphcbBRYToRN3XuW4eJFWfE1WX
B8knxwQb/4xprBR1ILXgtLYISWzkZajwxa9tCGuZWkdXLJVONdnh74hBHwEgRJM5G6mbp0gM/2FK
8UTQNx0q3HeZ50zXfU1n0QfCcegU1kGF3MvzYdV7K8cABYO7plwwIGn9icS1Zhi/jtIHUzIWjV9h
YUhdVZ7ydBMF8RLa+hUpealx6hnuHehVGxRW6iRhnIS0FPoc/asOesTOWWZ1mOl8jUAssiu5+stx
tU39uYeSdR2xK+CqKBjlWAJjS0de/SbihApRvfOayr/OL0KyQOOLEaS2OvFQ4L/9h6JdOyftmb/b
VUSAjZ//xeYjQzVO5OGN4UbzbXQDk/F4dSfhGBPiu++ctZAy6561mcPObG55nWVrpdInpYXECI6l
AVH0Z1X4jY529PnUcolynzKAm5b2UxIfD0ONcDmzpZ3RxUFYKVepwatMDc+AhsuAhsQfw0Azy3kz
lWPQzCcWgBtMvGDyO6iJgQ+x8av6E87nZbjWKlIXY9NNatqhHjGyFoWgJVm/AKW+x2ZZga1kfTKy
HDfhYOaFRLBcUrJdGrpb/TszuudLzNT4+//+5JiXDqLTCVbeO47e2/FxZMwTVs0s6IlsoCgUyCSK
hC87Rucyy8OQMjL3yQTyNeE6D/7u7DByS38kuHRJOWbKsFGKLb61HlPbLGlBOjQD74wYZdes4nI3
RBpiCsRQEkIYTw61ju7urh6ay5eSmyHlX2TVHYR07wFWOEfV3FLb4o4lPVS9eA5WVrPE1ENT5eZa
SXrg3MD6icXHO4ZeP7pj+8cmo4B2KHsQXUgFeQo7oAI2DvsoCi5z/2s4XUQ01IISSlq9c9jUN2cM
S1/brXZ51JuApRXMJRNFvuEDZpeuFccLDXQeTPdKVM9gvPZsgJ5zup9PPJeQkfSzVjTE8uAEDGrd
8UF9MF8Ol4SAMNIL5G4+/9D+Cal5ZT49A7xYM0txbjHPx3jz12mL/dAgp16w2mj4IXXpV3/5laF6
Y7sk33SambvI11b78HZCy67iSoDROwCsnjHPS8gQpKNfLscr1Ms2mG83V36H8t3/8laTwYqSwZOQ
tv4DftkdaZXup685DAjS1QcwSNmvcx95YkSmp9ujvNYz0tcjeDH/xIpV1SmtjXLrwTZmy9DXjUw+
RVItiwq3U8NXl3tC0k8RN4PAm+prL1cB/rXTo2QQjICngceb/cIGxbpYoXM/psx5ULytIBgjhDyU
dS1P55qhqxEWzdY6oUyFozWoaivpn1rfTy3pwq9u89Z8fGTlWltDgz70Q9sWxKhe+qQ37cU1Xxuw
8rjHs4QhNs1UEYzMlt3vru/1rK1TLcaj8gxJBrODpNT5tFPoC1cwd3OgFveNprX5jwU35TGo3ZE4
lY2pi/DKIguZOD3y0x5ufWE4ui3kogflI7NMMR6uV2NS5d+tBEn2it9TWS4iUge/x557MqYZOjcE
lC4VspjuzTQZ0tK4Wy/ktqzp7W7zCexmNdMSy99eFGICKt8J2JV8sysYpXFEYU0cNOq5wbMil3jp
mEWY33j7FyPiDgJ+KQPnXX2LuaLl6YCsbMiHlOW89y4fekrLKwrIkGFEblS1O+PWitMt24bq5pdT
6diV07zSu8dxxKS71uGEHCfxLHBxSjJ/ZpZKPQvpgKdANTCICaa1AMz6HmF7y63+DlDV8+wIuE+B
/ZgOzdlHtj6KgT9lliRn8l9Vz5FrIPz3pbL2JIXk7e5HlXK4QsWEKB7umQRA7V0LrgMIvq9q9dB1
vLcyYS5JsR4g/A6LjvTYwgkoj3Y/D28w0afaCLXfG0rvAyN2AVzhuW8IuR+FX01SffHqdEsfMTo2
YRZN7Nsmf36QZK61nL7yRsvLwIuyR5mCBs4B6gwKc+Awfk3kTqXcXP1J1fiabfOWoJLVNUyMsb/r
Q5OehzYrC733pcstpuPhufa9lw4bG22d2g3ky6LDrphORFAoM7H0r4DSQMcdhXv3nu9W+jmj+MWk
oUpHwcBx8TQ2I607Yz1e7+wQPel7yX8qN75l5jgVqctcAi0WG30BBaOZg8fTha7eiKyD/qgyU+do
uR9THLLfp9eoNiu5RPc8rR98gII29KIbIc/bIYQHrIXuTJGMA56GHohaJ38mgA7ukjykDoQ8Tot5
qKy/sigrlX05JgosvSYmPx7w2X18Mo0iTznoKEMO2LwCddVB4EhUORxVrOQNi2xOzvn+pHmfoW65
lySxWagE2X5qiIboQE0dJRk52DOyA7DV0M4rqZ0vUi138Ol7ANhEmXoTJ8gRM5EoSJOkdlMzEc5K
lEGqfrqDBS5KtW5xD8QrYh/SBod2SL+j4ZAzSn8bC+fxk7S/O01iGYM8Yf5kakEc6wmpiZx3A09z
b2vGb+AoHoy5as4eW00aYGhUS/A0MLfMnjyMh3+8NgKi6BCqrj2aGULk5GvoxIKEz0F8/vcLJkz9
SnOZxw3/BiNEEr6D14borvQ51qJ/R8hcKMA1IWVaJqtai+1iS6nCCfD5VfmOytgA1R9EDEQ6bFom
i4boiMoboFoOtwblgSunpdAKbgM+KlbPXn0PmYFxOf3FiGjL6Y6REoL/yFrmUvT/RFpRMWSulIcq
kS8f5PG4FnbGQncOG4z6t/MiwOM0g5VNdH2UL0oO1vUow2q+KVpmuc4PcLFQT4rr+LJwl9tRnC+g
23kvDPdKTZ0eM2Rh4QYWxaa0IjgWleW5k/Ja8dHP08vaKyixuasGPv8J/a+FP421GRF/xchO7Tip
TnECUvktFB1K5IuxjqYdaK/QCsCUbKqTDtz13ca6EptMex9j4AxiFmBO6bV1mW6AqWk0mYhOlG42
+f+uMaqDPSReRXdyaHY0/lvFpQa4RG0il5sUZcKaW/27DLtmzKl6q+5Drvwk0Yzl8Okc2k3YDr/v
MSOS3SO/FiOMYq5QufCIx7+81sUdlWCn09a0dSlHK17pIXbTQuJMQZuK0yGZOvgKbgXcXCVX9THx
XKHTEF17twMelpjMgyXCVvWSygpkNMhaq2WT2zs2zJJsR02mkGWN2MTlogoIUe0G/vKFeA+Wz9Os
yXllyXbTFabVNKqa6W21SLV7hv+pBbXlpI4D1e+ogNSuRKAuX9GxyEr8XtLzHGusqO4ZqAGukJS2
TVREtli9l8NV0sI5WanRmPimBXFN/Gq048lHAy4GJ9fJXwkffIp38LJs+Ob6kC0mVvLPhzuD5FN4
idG2DsC+KBVX4Nh4sMT4pI/PwW2umaXSFVj3VSoa0VliJBBu9KQZac31hfAOL1bIcsnkTyyvh+UY
fo8WIru9fNhmD/2axECnFhtBw7ecCISbX7RMaHgRmebJKL3Vg117PPxgbGGwTt73+aITVEchbrrb
40CYNaEXNn134edNEtVeLYvh9yGIq0+bQ6ItLVLiCfK+jEsV58tlXTE38XRFokUJH+YGP+o84NkN
JtMykmVKV1DP89ZEuVSwJ6DnS22GEtTsXESFhVa7KE6dj52HzUCqu+DLZREBMMLijwrsxNBZP87i
NEUmXx7UcahdQJW+h92Nj7RBKwvaj/m2563k+yPhHR9Kq1Hcc+ErFVOjSy5M0rx1hp3fIN70L3uQ
rovoGS2TUxtjNQwPVPyA5UD2B7CxW8JXHRGb9DnmZDHIgkTU9/nugbVW+r5ktOBPbfb/d854tk8L
/eF/Ei8gvaQw4Oi4DqHZsrfw2tswam5toz7TKIZWGdqRwqOfXSIRV3h4zAiTprag7DWyrX51FFQM
Qi+w0V5IuCRBVAd4XQix8ydYJ11Wh4MIRz9Cytd76cBAiNctu4a9axRqT42jsSH/cD0sFAdm8hv1
x1j4Djj5p/7XcAKTXnPIKUoWoe5a1CGEo3pRffvE6w9tKWLk1TC92Rbquk2PIThgS8ABXjdvrNbQ
hab2/ZLEnb1AFaueyNWdp+X0+Zrf4YoUqyaK1nC2A/GC9W8omaV2UlLT8UnkBDY0EG0V+7SW/l6Y
dkGhWkKx4RAwFrJpDZxeDy4eJ8kTGKRgCra2vYnsikUYclgHIlT/a6HQtDS72CIaZ41nbg/A15FK
Xfb7M53L7puu+3v/QLNFWLl/xTHWL3Qg0YrOR5b0XUFQuCV//otey/YTaSbvcIUzmuKzQACZZRMA
IOOt2N1xhs+8d/p5xTHbDcE71TzVN3YmotuOPu+zgO9kImJ2ABwrDaMEZnzMww/JcgqfJf/zt7H6
5KcpU48z5jii21w6nTCjxRcal/PuujhJ5UExqcctDR+quvDZaIMMjZwhkYmh6Gml6Mosh63v8hIN
GDEYFV+BWIelchYcd5otuZfmbpCH4FNBLsPIqyQ+fGEYP2Qyl3wNp/S273Amli0MTfm10R4a3Hqp
fuRWtUVBNX5GI/3hTw9Cp7RKMrmxBV5QtpOPNguXXy1RMEs0lnUu33oTczkF/RZB8Hm7tpgiPUnm
P0cIMX5h81Uel/Gi/8U8ZaEtZq4rhiXAaxTO+F8e4BezDOaYEG+0B/TPm7GMlKCwxxwM7bTQUhBx
leaqi8pFGdilbHJAMcYg1jhA9WD157X7ivb6leFJuEREkDFLL0hfTFS+h9ifaTxGjGJM7GTIAS48
88+nvWUSjI4cG0dkkrbiCWdTx4d+8P9ACXJRxOM7CltLDXSTASceM3hyPIowB2NPz7L1Wce9IDxa
WMe++EQUGgxlCmQfJ8+IjB6zHvVoSgw+2I2I2IqZWW8u3HWzjtdmAljCJ/eWCsA+B5jierEaQqY+
9EMhVrRoDZBm+H+egobIv3ek7Urz97IHLSw7JyEp3ldBcDywclKR5E1Lb2sXlEtW1lilynoRiwRD
lRXd5FEbSTDXIjHTiKge5D9c8D/rP/HwQ1L7+BZg3iu/MsQhs5v1Zfrb4g9dZXZ79xrXzuKM3G7c
+teR+sv+oE6ZDYtIwWpSkyvRM6VxEbh/xZkMzOzoKuQO71UPOrxaALdWx0myIItg6mKBWVjjGSbe
Y8quGQ0bPPElsN+WRBC2pyX5DuhmFtdX5MLUno7nEq+DorPsP5ADTIGQsyxBlE2aIvMuR18YQOLm
FsWTk25wquT11p0jBgcbeEENee/dW269qiML/Ysbcw9rbk4RMTSYC40P8G+lISIyTqs8oDo4L4wW
OIbfBdRPWbgYhK2Py5mqQEtCpzBhpn9D5pwB6hIbKTV0537uXPqyCJfjlH9TJ9sSxeSIHZkzRFlg
TpnVNzTsA1ePb4djZaQLaxGiHfALYuVyVGbSb7zuIM5GjxWkZ6iZuEcMzx7xMqff/ciPedM30Te7
kEW64MLtNymFVLnI9mPHZVwuArSg1gtFasEt2z88SPBJ2Z19E3Qppa6Yo0gc60P8vIg1bt5iU7k4
aeWVEejBNHR2Kx4sr+x0o1bdVnMxiqE7MbzsCGfVNYJsbgzo0FYeF3WVzYULh8T2YmOEkXu4nByR
LBbKLni7msvSYrOvVxWAoKmOX+CC1Ad8AY+LJ2SLXF1maHkkwoaDOGwbMKtYDHJJ37ankNojHPrp
nypATixh+HN/MPGslD5+axUfMpZv71+Y9UaU7flKPJICdUTtnSKx4YRpqlIVuGmQmMsccuXHL9wY
6vmMO0CYCBYgIWKL4nYkkKdPLXe3EEjXxXwW+SU8qBK7l9wwYgdPjAM3IOyVE7HdQ/wgfDD2sF3b
VpFQu2jDJdVIFb+BfVlZmIvIxul3QyRA3RAhGQDAbegrvmab/o5itbl9pp1MU7UqMxbxwMvujerw
4KzLirF7G1fwB/ATihCXwchx5rMYATNhcl2Uw/20KHwN9aWEStuB3YuMwlW2c675HQJHCtbHgOMQ
DG/xqMqQhzMC7eD6vRzD6DipeVpOmvX7xccFRGOASbBL5HOp8rzSA3KaFA4HDWViCeAsEMIm27Rb
HAMB//4FFtzTKQzs8jHPpdkGsjZU7h9OTWE3LAzsE64HgDbmBtKUvSwHBAK2YVGWz5qF/heVMlea
Upr/h0HF1OGbOXtNmukAZ3swGp9uvdWpVQd4yr22U3pwFG5bgMy10V9opPLkoWPH/ppE7t97z9RX
+PMoWxrRTRnvRJ7bDFT6GueOHrptJ6H9fWCEi4G/cbWOsZ0gov6/wgbBgJItt7Dvp8rR1bL6gwT7
y8+BB8CqZ9rUwwIFUrARi4MCdmoom47ZemXTi94uVhLDgAb9hARD4X2mX9/FBZBultYgeM8fF95h
twLm1eRpxkYkg3/nr5/p30NpAr2HGAEf47nLCZ0XvWvi8osxv9B9imRK0ZWbNuB6PnKIcE2TleUq
7UBqHZJxeOKEUbKiQK8fe9TKIUuVhc+7vaWz1ZxsUmFeAC3d2JzVr1PyXdn1q2YGrBsTn1o7RDla
yeGakrUHsTjUQGSVVoQkoygahthkkD1Bgtf4l+l+WWxt5xwbpZMONh8Qf0z3y2r54n2g4pX2seAL
yRWnGaRUKON2G9LopDsYakYf0UELH8n4EVOCjCe+2AysMCplyPJMUfXU/Duuby6R5v4F2qm9RJH+
5gc08Ua9O0RwtL85j+ejCx3WUvrYnO5fWUt1ATV2Hgimyazr0/zVRx5Gef1kKVi4XcU6kYeeQUOZ
09Bd+aGPnEkU+kxFeAFzvqerrUI/eguUh3tn+T+AcvjLw+VdFp/DXmFyJ+PVoCssIFfU3HHOWlxZ
Avc0vBc0AQ7xHNYnHyaksH7MZuX/lJ54vr8Hjzqheca30tKdfpbJm36Ya7vF3OJmHka4NryuECxc
kcuynvZOXg8LW653dBQGJutWn1wxIXibtWCBFsv79BSVg9dTsNwUPc8MXn/6b/uZx9BxEwV4X4OV
99WnVrnOdoa7a5bc1jRriGu+52mnRH9HnlUQ1btm4oGvbY7VTLFJLmUbpISDwEtWxOHyjNQIcxDi
QzSdiSFcjrapoQj2hmGZIOIATouc+5x5h/eUy+tcULFATR8wImy+D2mrZ+jJV/9rXwRghQ3x9ncQ
xNjPP36wg8RxUwUg9prq8p0ekfJyf3GkiY3/vWCEby/5zMVnb5EmZxhYiYN57qp9fSlQrKrKxi3M
/r/rwQg1J7sbWLuwtziHnTlx2COOG6ArzhEEoX59y0rm5Bxipl477TcActFNzt8qRdLdRWU05eKh
VWo6ND2E3dMQLixshQvma9sYBhmZgy+nGCQq+rzobjmHlrALZOW2BSqJuPU9xrSXmYTvWez9OolZ
OO7HKLurCgMCVxVR0GxGIYWOuWQMJzJzheAhyb2ULxAdVqXH6pwVP6Y/qpd4SVhOxs9iSlfwlTyB
DvU30XM1AeE0T5a+4WjOsnZpiq8K8UNlb/yg5Xjv56BnfPcRUGU4Z+tiTF6CxltnemcaXQmxgYJE
/MeTFV//uMppO5l09eUdafq9hwlA88onSdNBbZpQ4DxYIEkHhKmQ3lU/A3DN46qDZBE6t/MAdIUD
It+cGC/SedaJmBjrO/pGmDspBuVxrPzk0IN8PLg9QJHOTwJefaW1Vo27kLb4dToDOhSGDrNWFOsd
3WwHHnI/uPYXUTggLGGutlOMVSlGN/w0x4M0M+bwtEGytQdT0XJPnb06ApVCZ9DIIspcyEtDJVgK
kxodR5IicJc6I5YU7QHP3HKpRK3t8wktpeTDwLDXeuKSYvkiR5nBflTTH/7b6J0BAr/QBnbtj5hf
nTidd1D2eVxd+991g9QdYClmrjQCr7XGjUqvME0MpSPLHGC/TGb9Y8q3UgUn+b9o+oLtcgG+MfmO
90W6+PoKAA024CkCJZIEVAe217s9m62w5gdutyTAPImWC5YqIe1Cxg3Uv95Ux6YgZ8Y0PrQvlWDt
gF+z5x8TLUPeEld8SJDZxNjUc3ZtkRBkn+oh0XtQVdYAzQXEj5ohTDUwZYCTIqVaHVBwF+xw1sfb
mkI+yNrWjW2BXhy3z3DAQwWy1W4t6DMyipJ6xKSrayQmGjiYBQjitHNKodLYZCLNCYbbOk70b0Sw
c5IUcuxPmkhjDUoWnYZOgmOLwnIhsZh0Xn1rQ+V4WURZGIihdsquMceuFeiFYvHpFbmWG1ZzqbKw
U5Kro5iETiiV6PsR7u6UtCQP1CVvPdDAAMmJjthB7rvCO+2T5WGufFSC4tk2vOzR6OeVVMutZmwx
KFWm+0YTqfsYdW2kS2ce11iN920cH1gtjiXKx2zgJPWaPAZEKz3NhFEfUcWUAsHNsBVQiZneppq9
JOTe4ymXMm4AlljgYyyCZXZrD3VUl1DicBQKY/DZGNIef8TBaqo13z+CmFGPCxYDJqANA5s06RUs
LDB1iXO8URBerc9/yhX0ER6G4K/dnx0Fe7D4nswONdLF6+bTkEnWCsAcgEgpUBdMG0rA4gIGyB1r
HrEehhG2N7QcXNsQgXexvADq770ENK25mvIlX8bsSLa68AQeg+/x2foj3Wud8GmEsven4Gv8XZLW
udar8Y6tjOnQbB3Nnx80aZ39/EqGABbaSuYA5vXTpiPglvvabWjuP1li3C+owgjpzcRVrHWt9BVe
gqxWbMou1UWvVLcKFufGAXbIpKYPiW9HqUOqdDqAerHIGHCaog8uyl1aa89Uhhvf8pQQ4uw9TZ3O
OJyeZloByraWd3Vvr2myJyPS7oES3NIxM9o7GOnfN0tWyeAZkRhnSHsHJ5f2YiApDeSlIRxU0DhM
istXHi0vqB3He8+fwxg6r1t3ay6gZP2nX43Ubwipr0alL5lmqyu/NJRP1u37whiJR61nai3SdwfJ
cNOtCLJ6ROZu5Q/n0+ZjtpCeVZrEfPZjMp4cD0aj1coS3eRwSbdEiFpFOXSVsq3sizAAnKd85tzY
KuixysP5cDsJpGoso5OXV/REvfj74LYto1qbwn6eSG+5+4xNbFqCH7toV3sRoRrH/Z78AfYiAK6q
u46nI8nI5K9jy8z8zyp8h+UIZ3UdJ3D13kEdQFH438JjxLq/EOit78VDhzQ0R5vrFxnRaieBLbol
c+kcp0F1Wg/ajEKZMFEqh3+2vBMixcNB7DZBJl5HhtdDt2ScmTK41CMIeETelBYNyp/CdDCf+jSg
/Qr7Qw4e56ZeBWJ+n8pcQKz72bJANFzSORIoFX+0lJzSNjBzhXhkfqBaPZhSnZJAcddMjT9htGg5
I9KjMYdWzlJCT03qXO0N6D+iJUG9d8yfGY+hnKHm12AdCKC0zd302gyaIQz3cY5OBgXBm4jLeWuP
dwJJ7CwpzCot/euny5D6rFFYvRnd05LZ1KmP6tI1SgbBJBCaUYHUeXP31/FaIIOZws9e/zB4Csd0
ZeVgJweaRZYOopJQZn7m/MwOa+IGnS/mk1SUaZkfBzAHWaVD//1AsyMLUSl0Ej6123d4rej3W4eP
AmTXYpknkTpWr3aaWpZTOLwGHekh8UCB+IqvwIGu85ZnsyuamXUEY/Q7IEuhFohe7xblquQ7eEzm
cz+aetT+ZiSjcFVBijQqY614IMjsdaAOr8j8S3EsJtGkvJO5v2T6bjrHIUiEMadGqiC1sZv+N5G2
mA10LZIUHeomlU88k8Ypz0UFC5qY2/9kWydL0A25ChWQy8TB+HMRigDLo1ckRY74w9WCxngyGCSx
uP5AGYFITsGuI27STFlkBQC/wksAGia3XeQL17paMiJhJGxYUrSCDVIvzXQYpUpG48mg3UxZsg+R
JYbMH4GSiDZwXAU67AXF8WMGLcKMxX62zPu4ABszuoUGZhoTkhRNarl1QtGp6s4nk9V0YFvHp2Yb
/rAX4xJgjbpnIzfoLsxLCsXCFbIseqWsV5BfqSZOeVYLsDfsm5ERceyt55qpX9MkFsEgFjFiOErE
w0PeTpvvzyXtdDXHBK7cVPuwnQa8b6RyweRkU0SJ4dRMHCADObgeCB48I4f9buF6rvyMuK+w7IJM
FTXM3Eg9BbhGDYjSiENPqDXumvkHfYnyF/Ek1z/uczyChF5Gi7dpWyB8IXGWkdIykFOTA7QHxjss
bgL3vv38o9VJp+P3/EkSaDmh7iszG2m2A1LsrFQQGBg0xULhi4JgQmkvW3tlxB28gtFzJK1VmUPR
07tWxeO4rKDugOmdn8PPrz9dJ0rkR6CBptqwd60pFJLCAENKmOexoMVJmwDTYKf++ZNrcDUCSBSr
LaQTNCaGyiduyobKEfqngyDImoEqLI544HN2OtETgKLH32Dlrj39lyR4/kFbo3ub3y6iClafRtEe
WNd6o+g/xWEREDf13K7aKsd3gZ9mt01kTVJ9+mltmp1i4zueyyhwP56d2f3+ZZmdCUcUpxrjlWjB
EnICu8RzatxeVCzyM9h3FIGKbzgsIXXfo+TdgXmwDSbY6vbm4gjg900iW/VMRJJox6b/E4QUwLBV
WsR/57e50XyGGiU/9BpajboYhAz8XSw2FAt+gy/UtVpxXCVR3UPdZ1xp5ITiQY1bCOvPSyn8uESG
zmm8dUXo7AVF0kvTX+ALd4MsO2qIymzca065BFgk3yYTTsUjC/I43gm7VsDHVYwkmdz40AX+A+Ne
Rcl2Wk6CtaFIitgqdWNNMBEananUMcv+iIM2cYVEhKhgoW+4mKzceIIX9Doj1rnNyE26XAmm4xLY
EJ5G3Dzk3WSM07IpRyAgOyvqftUuw5u2N4kHlNO1KBil/TH/Am5j0A7WGKY4PmvTqeeJCnazlm+3
uG56Kg+X3Fm6z/6Z4wRxOM9a4hsynTism+1VqD+6pYXr60fh97NLdjR65DW3wAy+LyIQrJ++qnF3
DXjaZY+1d+Kn/uD1qDC3kWYO7VqNEa1Qn3EzOZ9KrcMtAjQOPMIPdkqkz1PbHTPh0REqGFt5uUCu
sAgKAJea8zp5oB3S1Yu7r7QRDCTPb3MxJd03gnmPvgoGFfVRZ86rDxQhpwn0HxTqllQyqtq4bJGu
6ihTeYxgiWdBs1CRBUozC79oB0w6LM3+gkP2oxpFfmG1PRwxPhM8pTbeqQMiS5OCLLIPIULIlOXU
lqjI4H/3uXUnGJs8yMuKFkXRXkdLdv3aRMNlB9VCwu/3pCHf+JqLe5FNsAmsT9NN/6yp09D7FJuN
AYCsC5EoJQSQt/cBs4quudYoQjE+DdMpUrrNCK+Yai/c4hOzDrn9AA2Uy/9G5AlNPHdcM7PtyJMc
4moIaWpEiq4Q/WGcTQeTtEbTYrI+o3cB2Zw9o9niyarxZAxgpVhc/etO/edl8CgJvu+EX8oWiwSS
bJ8r2+0q5FiyAoPfMR0qXVRhJjVNGyJ0PTheW4TmJGPuBEiogk9nDXFJgujjkSyGRzjgBVeVYrL0
wXt/Cjnm6rACpzf3QxYdT0VG9jzpszwNfT3s5B/gisT891cJgyJGXTCPR4pYnX0lO+eT6KeG3Sx+
A2RtyMpKpQLp68EE/PR37iygvmOtKX+3+DO0vDwH10wSQiHT4PIka9Jqg3xcmrEb/QNJAyGKOjCo
2yw8maSdFjT7g6gG+vCEA1A/EjfJDjd/9sdOmkLKLs9cJNLb563coHJZETolD6M1yol3EBGldcvJ
rwE+yRXLcZji9a08frnTAoJstOhru3ze9lajU7geKEDyExZ4varO8UAUcumdX2mhu0j4XNySAfLE
c1O0Yeb+czm4/Q78chKk/BtLimoyC1+qnSm4oOzbAYv3OJHe5hQOrpTUs1DkEQaK6FUuCj0EQOFG
92Yx1CaYgrN8HqEvUNuNiwpglaCbVm20qBcVtrFCQHQlTWyQv4+lHGeoy6tjFyikWY75mwRYKJ+H
bpioVmzPVy/DZXiVR6rhTOUXV6x5qHFXyJ5yYx0BidRB1heF0Qk/0gaaLV2UNsKS19NQDmrnBJ+D
ua7IaWRKdMX6NOx5n127n1S9/Vk6A8maGAKiOv8WHZo7rworpqeo/jsjDl1Eel/f0vke/XGw8u6g
mlh47wOcToNilZPjkgj5htXnlH3jcsK0ljv3PEDSmixA4G9cbqFYpNUWW8zbaPXq2MShFKe7ihIG
lzqJWC2JMsan3EBSGjUrOMT4PG8knHKOIXkyLtE++ck9YPxsesN17IoSfKUjEBprmdhzkalSCoMm
rUClNBi6ClQqSnQx90v0UESWWic6NQrYowQxnv6vEj8mO2bvmpyxyWnMo4ijMkfV2pGZr/FdnNTl
6TCivW6X3uqnTwahUwS7tt+oNDm6ChNXzbFQfO8srW0xN+buyroJPOKLOjGbOVC5CEXgbCz27aRB
k5grDOR/QG4fiVWFkpOvWD8NPypxojb+2VOOlEr7FKakPbxqatQxN12kOQM9CrL1rLQNqWnGGbfY
crS/14BpgpFlXEZCjbMzHqluwG9QB7nHoQ3qOeWNt+C+kb5d8TD1dtQG82oqegRMdUTI+wbc/NXG
GtiTUkbWuG1D5gy7EF+3whg6UZLaIBu7I3qBH/JFMeK8H8yPfuFFH5Q4yYWtAr4x+D6Qmu8/2M2L
/WPQZP7js9v7HE2h0+CaEzvkQlzOGP+tJECUE/JJBv2lurvmmxMWcWLbgNSKALD7Dv4TpHcu0sY4
xQ2iZcS66Nl+Au+Jay9NgfWbmZUejZI5LUl2DZ8pyLFS48OSu8iphrGm4GfCSeI8Kwh0AG65bHLP
0Ia66qvlPTCSV5780PdZVe+X8i9qwK2MgD6yeEXO0+ggMJh1I1Dx05nWxeWUwiFEY/wBfcKlreKy
g7MqT0v3Beyqv1oJEj4BmwmFYm50X/2WsO3CxcS9QPM6G608KfqJ2GOBHAKpf55j55qaZvHpghRU
sI00O2uaydtfnYACqYtZa9A0f50LxfTHgZ1cOrAp28JlhLf7voG1ioguaG+m/tLQNtqrpkXpmYm/
RZbwx1rxE/A5ScIYHYC4459JxMKpoX+Pw77gAvueo47OQdlF8AUJ5UiyJkGzHhpyXvaLdwFLzb6H
vLp79mfgx/umf3p5mBL7kshTN0ZTKaLBEITllOihd13NN+bCMnmar4UzxUHXNddqMSA+BL3svGr3
9jpwa4uFNd4P2yy7Qqkur2l9Ma6J8dv0Hfpdc5UN8o/veM5ngqIYRyntjROBTg2jjDGpjRwg6Frp
2TPeysqui3ORjA1qXIaBAtaaMxduaJycJkn3/kTnu3y60ogpYeKw2fWVFMqJUjqUppxPmksyosCx
eqIWP1kuwNvKBcmdbF/eej8E95oO95TjKmtwLxKMygM9IxBDnr4zww7Qp2sch6XuryuvU4QSM6jx
koLcyB5IjjnCmf91enfb4Q8uRxEmpAWdVIU6RoAvbkSQMbPo2OJr4nCgNHL9P5mzvImKBVo8/MB4
DUILR9UhmCoKAN7Ix4EphGbDeQgRUFq3EkTWP8b9zqAyUG57rpOWL+D1q2UEbBsi2hlxTrcM+Jwq
t8sQtfHfrj9goMBpEWEvZFIuEt09QSkWhy2K4L2Yfq8Wsi/1Mm4TZBcIYAOqi56YedOKOAMFGARp
wtdmbcmWsGDeoYurMM6a82bWmDcBBvaUsgqYhrHj5EhWV3iIXUXKaGYyFSmgGwCESTD3CqKC3YWm
ipRp1OXFiUzGt2+Lr9lgv0B5dOF6CqSAVN7Cw1fI6tvrsMsNgmDWsRdBh8cD5x9aeo+iKnKnPZyw
UxmUaqlymHP6h8SAdmYsSqbw0tG4EWQFBGvybV9CXbRbJPSp9pNCxQmOORWfOAL72tWwSJpJWRg4
CaPR1DfpAvixMCvUnqamRxtLaFI92qcm5B5J/QCMLgxKOPpJlEEqJSk/yFMTn742THv/glzRL5fg
ALZb1zRnm/d3oS0ba3U90XfltPstH9bIY5nd+xrKCV4OYNeSsIqBcnvINW59yNk4cJrrRbh2SZ4u
MI+SB0NFCM5LVYPHqrZzTKcmDvdebzERxVbn5z2XnCReSq2dk0ed9mqAUaJcFO4TcTfuEIMUo4Yv
e04ZXD3ggCcqoMx54JwiZkb5/Pmwti3SFgQzdfxvY0PHYE2fKk7ohVGM7ILIqXY5UG7ILXVz3isF
5sSqXr6h1tfxioMBQeet7QySVWeNu6wrJD7cqtgRP75x2HM/IFl0CJvOQd6a59CTwLH87VRGrdeZ
XqmsTB/OnQqBmijF/Bi5iGl2Isek51Hs6KiTjMvBvvJSZNY8vy3c/TpUxiB1U5YdrNW/hNg/FVhF
OvdGwgoUWUG0bQcivpLcG5nSC+LGwonvP9nzd1gLoDh40ySE7E93GjVi5wXoD0MNffCIkzi0fh3b
jBJgG1aZtEJTmm9AjwHmo1N/ByFBscK+KGpNvspk9C9WTcSFjQrR1hIdBE8LeEyTNZooLKXbzXeH
5QFiD3B6ShZiY4NGVb4mnSpw7YMN+kAaR8E2SHjziimnC8GvcfG7XK9qdKe2YC+V8UiwWxSp1iq5
fCUdsu+/dZrbv6OZCXcJesPZeDdWw2+TUlhXmhU02Hu544n6HnvOxmxK1ijMjOiuy4K6XUiOHLw3
WC3bJ+gyh35WbeHjlRwhnHkxV1Bv7zngbUaN+GDtBnFeC6dymh/TnFTLhhb5Af46F21U337xZG4j
aBzYocfcVqHGJCUgZIl6Bt7mGf4LvPd6P7FTwhuSa7xXOnEzwvdVDAfLsiTI48glKsX9N+OuwyRc
mJo0L0tSjhJ2itYaLn9s2u1n4pN2u5R1SAk0pd8tXtm0jeRdAWyzx7QD/M5Hg1tAK4JZo+2nq+B1
3jRgsQcI3zRPHYdrVq+djAjpBsyZ3oPzTeBeLQl3Kpatm3RBlVNGgbipo5da3QUc/Z9LijaI6Cxn
BMBjWvVCE2jloGLhOqA5xlkjc8OCwJw0nkY/NonH1sjwFMAMBFCmafRVJIN1xC6O+jaBiBlXpBcI
LbBYm93GTO9wRmIYZvzB15caNrfWSLuSb2CPcoEIa3CUgQcgPogu0UirApV6QhwL9WlFcuc78+Ox
bBSJkvwqfdMZX1TXtULTSBCJG5iT1ZkeBZrj2grgDSu3Vaqx/+9hw6SBkjNx+LQiCWh/X1dY+Xvr
oPq5ZW6mmBvyAo+/swvKmVQvRDA8opeiWKg9dPlfLRranaGfm/3xZSXA7ays+EsLMNz5tUqsueS7
6Z0k8GxoEkDBCeyeLbtKaxPsa0+GK6tcyoMUKpm7W0kgixeasxCR4zX1Wfr84+x4Nn5ADpxDoxGS
HOBoijcrVbUP+tkqEsSXJRMmcIK82rKM1fCC1QyScbUimOL5x+jb35SQdrRxNRLc64Nc8/AW1oWc
GBsw7oPrqUXI1l8kfZIKNcUkTDhO6+LGzmpmnzS1O5K11iplhlRzYLYiJ0YA7/dE9PXWQ5Dy6AIt
QubSyhowLuKeFvV6/zmBrt88IAWuSCU8RiQIY4ZfavYutDvnzXuFgMkiW+uOviM3QXMcI/fpOTP6
b/HBBvGibZ8gX8Nf6Y+cAd+zEg5BwClfWn3H+OIa3Imy3Trw7HR5o9AKa43ss0hu1JkkbFsH7Kpj
T2SRXd0Tm8EvAdtmCBginPm4g9QHIn9cDRdBLiJPKUZ4Umvx06H3/v6N0S0Lt0aJYeD7kYqDupjc
eb6MGABuClj8TanqO9mCF/kjxbmPtaA4Iq1OqecLHNPW2fMlyAdJChB1EhFSKErrLpjfF+dqhr0P
srVFsMnMlJK3jYVYuHE9JZsbLsdfCxVw6SSgSFAdKknRuheAtFWd45PHMJxiieJSKCc1ftytJxFI
qNixqVVNV5ovbdEhMXw7IY73cZF//mpO+SEyewjeTdV0O2NhCwVshn/OG84J2iUKIQffYtVXPHua
edf37l6cig/EwFcOPESvuSw964KtjZ0Di8agmW3I0tzSn6RAvIomWvy2bYxNZJulHZwnrFISwy+7
CzshC1SQhaltMkepg0akNtMz97xR8+eOcyVxeaa/FpZaObEtlyoNDPA1PFjYZFkjGoZsMue+Jg4f
R67Yho9SuWWsyzsbTbxwFPpd0xt3CtrwXiOLIjSMoQPRCsT4BSYlt9D4P6PQIY/9x7g0FPPjmf1U
I6b5eHJN5T63HRw4Kp6J5NYgSRcSaq7rah/A1XNsZcizTqAWosi4vYuOruEAQ0Z87ZQkRU3pSWTK
hRt47B5JzZ1YKaw0YZ6ySxijj1mZNSgeqPw6259gjnGy8t4LCJTej0H27KJmO7AYe4YWeqk4JRE0
2KfkfLFhMjO4GT9npXVVUmH56VTMPQP5uuq/rQiurTU/HUOg6OulRY9KmqXbuH2iv+gfWi3sCeRG
FnCbvFOMWNXsz5C0VFFoPD445fHz0LtDjibVE047akG9vYN4LrbX996y2NxKRD3YNw/RcJtZJFCW
OzXfuLFnAAOmYNL9GJnfEP76ODRWeNUnZUlAPzF9tFlkC2Q7GLYknzjLKCB+Lm1glbE7fR0sMW+v
3hpja6jn0jxVL+bxfP3DTDbVBKxMYn4ppoeNU2lfFNP7S/HwZDHDPx1N9KLhllqY3uU9NfteRV5F
sjcry9AOUKckK0q1L9ZUHSFVHYKBSVdPRK2Kl9n/rgsPIqpC03wwpsRhTk+j+iSufs9CyQFFLz4r
lwoOKM1chvMdohICnz7gXR+EnsLGbmpi9ZSbpMHT3DaKnJilMRNovZQ/D/lBipgJRibGOl/GgVHs
ybORwv9NrTc9Q13rrj2WLAJLP17FHLSiUM6VeStFYy9nC2IkC9cd7K18UG0xnpml9FTgVVHubKfh
0wg6e4ohKxLIPBBmqAbrRNqZes5sEN/lrmP5F0szv38voxV+OS89VhK3OBsBmvDxTHglWBapcT/q
MIkwX8GRblnk/Dv7yPtg6wLqcezzznXFqdUiuHfYNSWjutmedZbuo+oHqtDC/v+7pd/ohZle07kI
ge68xB/+R+SbMo5dpgn5P+8nIfPl37QYGcKPv9LEqcAyM+mh1re3xIKgMw39vAMDSDs4cAIXQUlc
2cbvypVi0wRB4ynUWOE9In/6aCPOt6Kk5mqAA6FkLjv8091SUYqmsIiNYM3O0zhtMZRF1WBFC8QS
MssncUH3EUg2kp1vYe8UAuUfTEh5j2Ya/AaIt5NOp1Cakd1UuiLfL+JjE1DGifDVahoLsPK03T3r
7OMQbPgAc73YVoUJ+YPHq6IRo6Wiq3p//ePZhKAO4i8keS3u1t7bNIh/AE3DTzMZ3IRV2tChvYd/
+30fItMARS9dm+pLDFeowHnPjJOpaiapIsaYFFPAmy7KZaue5cyzrVaBEDC1bXM9z2KI71mixjUs
VjX/9P5I93o6AMgQ0bqGo8z6QZQ88KIE5jhWdn3fwsgrdUQBpHZlz55QYxqLhZozUoFRjczb+/tV
Dxs5y37jJheCiiTNfzVaY6s43PS8PhgyiSN2BzjkoVjSys8YJng2KWxDZEEau9x/CF4foHoLnyQZ
UVWoQCiRWdTsYFTwjucPn5yyFertoQTLat3BYNK9TKkyFmZqb+ZWLgrOQopIDdXkq8xJrJyDvOOH
yJU1k5W/7BmYjjhRHRjKudSyDFr0BqLDtqVNPeOVfKqgCMxOAPcpJIITwFsU0+zYw+hxt0co5TC0
S/2kHsmW4b1aUxwFF82AMvH4sc2+W/T56xF7cf6ppZOOQHpSrB6Mgo4RANbE9DwXWS577bU4jmXT
Jx2zg+jsLGcr+hZv/7ctoZODjl1VJJx9E4TX8GZu/NoAWrQXBqSBD5AwW7yhOT2Bd0rMC7mCW0oc
Ar/UP7+3CN8Y5HgcCMKCW4fLNCp3pVbIzt5I4SnTVr7jf7eJbbWeg5HeZpzbluECY3kiHdcIprn7
fRnzqRYK2M5hhZtLdIO7zwsRjr5Tt020xiKULf3z9fT7a2dyS2uO8BJP2UwaqvXiMX7UoLsbQfoh
YoThfU9iiVfQSVIB1Mt0OYDKS+7Ntw0ZqzagH5Ve61UtL+wRXDNheSQOo+W6QsLeHfiziQqUdzh+
6pX2yyEfR3mYlOd6l8CI1Y7x1lWmiSEPzBitgsA7O6+BUrti6mFYPbil3tqaEX2vPp1O+HKcbUtq
ru05IL1yOSVreUnfFp0S0QTAxYr73bKhn9NtyuaaAHRedFrbSEgneSrRa4nc1UOuGI3WRh53txqa
pbHGOHlAa0O5pj0BuKL02r1bVoTshqzA1CHAgK61EJnmSikTk0RgbcGYBTaWkBI3cftZ36OZr5Ek
HllO5N88OqG5bgMoKvS6Er2HoAU9cHHA40mg1ZMjJ7tSAxX9eKuv4sssgDQj5KOwOHm8Ys4W5DpL
9V/mri/c6a8XE+VTHqqVZ9CpuIICkjaMvg+BFIPdk/oEGXa1QQ4/PzD+LmJrxr9hSHTXNpeoHc4E
yPzJmw05AT1HnZMi9FZMiEdfUKeNdcX9yL5CEsT7sXH7wVGHrsXfc3TI1hlh4Xv6+6mDvO4YFR08
m0fq+eL2fYSa8AR/ioYHmJPQ4546NL4SdUXnShhGaZ5+GyWoU9BHBPJ15ocQiPNFBbROG3E9hMaH
HR+Gu09kiXCeE5piYF1sXXvtZqLw9sk1w2wA3/4Avp5XPeyIYZTuFnqgl9lG/uoQZnbqJiJyQ9av
7IL/v7Omhj3sqrNrKdC6VTb3ETStyij/ELf/bt1PyuU6cPvvRrXKGaJFxNEWL7ngayK2Ni9UGXyC
93Pj6jVzDkwkrkzz0t4XgsHkqugnjfP7Itu07P/WVZwd2zx8FLNxpoUTnx2qoqTXSMnsszPevh3B
Mr8/7YAax6SKjHMUQOl8IqHcMrqvjwCcsv3IAbM3rQ64llapCTz0WTDrpdisbAfS+jjXcg0+f1d9
GjvSBd9CZ4uNLGPS4BndeqcUDRTq5w8rElg1j/F3VnraOk8tOu9wjsnVbUzpSRG0v1dQtgHNDDpw
V87d3PYzKL5qOlOFvkQ1vBstChyDKKkDH106yZVmVNwnnWGltc0ryB9D1QQNLawVZnL4/43YqMgf
hnlNCeQXCuKwA6hZziCLmJIRLgMchFymeDnRy8BNx68NnOFdlT7Blm+5MZTcj1Tv2TzIBcZ6CIoF
enCiY6tYV3dbYyYSchgu2qvEcZl1b9WjQxZvdIxwl7ZPtvPlrJ8nInjjTOnRTXaJ1KQ1LXMqpxQ0
Tft9wkN6WqJhuWdNu24T8r8epKDxBWSZ2b1DN1jQIpUr/YgsbYIm27GpZLKBWIGAGOVAOWTfB2oA
vukMaTXugFQlUcuvyf1hti67gR2fd2kf67nmDAfiNlsMPECVnXgLvm2cUzy5BmZ0ozctSpEfDDVe
gwbMK7EPRrBlCCxLiy5LZdV0pnlPAEyC0/BYDehwIB1YLafhd8mc2CqKNTgSuUrDW2urm8b8IzAq
SSLAzFyhX20PbQUKzJxisj9ZLIPd5ltodadUre8pd/imZdn19a3NOdsJlMypXuZ38xWvYBTbuIVK
9GuAig6fgCrkH4xSIIMfqk5TaWJwaDFmQFsMugTNlxx4rfQIbXQvv466jA7X6qGqzH4/qVGPVmgs
Nx4RhrXjy8y1FPIv+r0Fzc7bygE/YvfGkWGZlbF2Vh8ej4WsumDn9I+4t8dIQVhoSWAQxZZBG42E
eC6gMrDdDnLSBW6P9VOORutYOta0hxYBIcPg9YfqIDjMXReG4t6iEMK9J/1qutHX+T973IUJocCz
tcTBarYNHbGHMqjL8Cb7RrvyZuYTBiXVlwk/dCRfg2+DyzbExmR3CyRrQpXoQousVMWXDhQnC3Uw
paPh/mYS08X9eFer9kkjLI92kCW9DyOL+3Z/iJX0Uod0n9eiO49K3Sd+FXxBqiTZpm3By7470D1g
2C3GzbYwINm4u1pXPifqfuR/1U7BnE0MU23Mi4PHaqQqRhPcsKOL+oiJY67EX6X9DTm4tj72Ac3h
gqkL48M59SH1l7q6G3okX2c4WemBkpMyviCHfv1VEqjrkOR2vuIQp4Tyd9FDMzqD0a7xFTg56uA9
xYsVVU+hQ/iBD5+hH3a5x9XUMxbD9jrXzl+CCtoUE9SZ8OpYjmOfdxiAxug3XioQnFkrk7OSxO9B
CodXxuGfDYvNbCnebK37Vt0sM300nfyBUKTos/zAdGJNyo/C/aqY+6DGwG+VIy3RAfRTW9RQ+xmA
Or9To2KOjJSiTsOqVWFYE+oE8/0kvopfl6eoUu4unnVS4CpPL4d+2pGamz1Xbq0bPDSA0LQS/frq
mZN4rlAWM+68zV+14UZwRlzqrFSaP6/43SkI5H3VsoNy3Wg1YzBAE5yj+YRPWYaooJBBrWrMIyZu
juqFobNJCsdIuB8ZRlfTQplgw0BwKkKwhpwBiIcbMAs5d/UFyT8XQz0rxTKpb6ib7OnxftZYFjeb
uFOoRCXMNWAbGFFo3tuFB5C4XfOWR9XhYOUTyJCBCtp5LweUgOVKuaHfG1pBBgEIAoukaJnpd8/9
95aAKbugC3FJhVv56Y62n7p/xhnVz23wZ/VpZHE6FGj6HQ68thNpD6H4qbfACWrxcxqATFs6W0ej
W2q9Tj8DHb1q+uII+PwRbyrFVFh8ZfTqJHHtDRPV+Hbo50fIK67cb43cgxHIs6JB2E14GttiV3OW
0uVTMllP0jZ3mlSLs3Ozq1mJ95Vx8i6DhgVatT032aCoiIBFsgSi51Uy/uRYpX+czMOSkmVpMJdX
x9bsqSQlv6LY0kGzYugDTELOC7IiK/t+tBJqslhfh16ylwQxg7CfQcSHTtwiAc52mlp9LhfyWcTK
OukTWXkINXc/7rT6BQYm+2XOul8n4ehXdWAO0t4+41lriwByolQ7K3b8lmir6zpwawjnwcxx2aT+
IU07rc464t+Xf1Svn8+fNLcE/bUfGgrCRrTYpYtomXPnVhJA6w/GS5WzamZ3YFyLFmEh7H614itI
xj2FkOwBvPVt22TUdVsjw9a2b+sIvh+P0uIhV5gErAZFU8Fwp8WeS2CjmbhBNrfCCDocxJV1FfvC
Jk1KyX2trJ836mjWMSIXBdu9qu86NODgpCoTL9JQBDpFLBLwUmxfBLpfZJvCyXKuX/6zXRumvA2N
nkaR1GRCVlEtkMQNepLxdcjyHjEDRJ2b9x1nh5ABAuNqsVOm4ZAfHxBljoDhFK6tT3cA22To/KTP
rNzjDSsYPv3s2Y5Gbj7EF2M8ajwQEA3xtRlgdRAt2vGf/Ki73B4Bp31AvJ9GUoo+pBjuDpw1McAd
AK9Kl3+mZ1sWJ6t3s66GSnEzGlAGKRLZI4dqnYDXLhpgOlCFCfy+qvpJdmBnR8RcJvsOLLFgUHrP
St3HOTfE7HtzwTcYoXXMZy4NTkcPZq9cv54Wv2kB8no7kRcFrX69qRulL71wTSKgF3W8yBXUYESv
Tw7iYB0L6nK3oLxhBWc3mHaZTGmIVyt/ZHZz7NmweaEgj2w4r6rSO5ANx0KV60AK88Gm0JQ8OHW1
+1r5RFjxYEYGibZ1aMoMGqbdgFEtfFsHcDejVhgyufDxB695LjWje12jH+ZB2rckutBxdgVBe4Ql
NPGeejhdki8JZz2u9IcnLxspVFHSbNqN74JuoYJofWayV0Y4KDmTS+gOQ0QzhXsVdsZnmOJSwM10
0liyEqYpg1j2EUhv6rJjMZ06MzGkHsj5EqTGHQ2xcuJ2xYcwSwsa9ea5Vwr9HLENur6OyQGVqGoX
8HCTq8ut+smH9xf6wxU7N1LoMtew+TiKoPe/UiiDnPOsQPRhYtoz3LGCPt2u7J1vJwC/dn9FFnGo
lhoKXdRhJrMvarWfDco2yGMI7KO7mly7cwF5V3VceMoxvmqWZYSQHFsqsEnpQXEMnKxQBlwsIYf4
iqSFP3H3B2jisBW8TY43vO2txLKMGrIxMTXX2bbnG7PH071yhIDSnx/Ix/WrcgZ5t3e5valHU8vG
KGLgfKaTgFxUJmU9wP1+qFobnVjeNcmv+tu/foGt9Y8ib4gICZBiJNuRwr0oMTCZDJl3st9sJvH7
ztFlPKwuaKQSF9DRRsNmwfG8nxzeASK3QvWzoTGbkcCv90MIMIu/iHbt0vub171tseFVpuoE4LS/
8yuG+EsKYHH2ZoGVZ6zh02jLx36E7CVZx11nCVveFAIcBdwSxcGJg6KXuX5z0bCxBY8UnCPtwhpZ
i8I3EWceYjHMyGJ0sIbqWR5j5BuDH6FEd5QSz5OJJoWkACmlHti/2Jx9z2uhJka+xXCT6fP+dxtY
ZdpNYOaox55o1znYkLe9PDrtnVsZpgYQcwRjPOv+MS0G2cY185J7kT1qBM2wR9kZdPEVGUF+01eJ
Ds7PO8c5uU0f1xBDvrRXDoTS8O0bofQp61uqNCN/UUCnVwCh7mEwY7Q/6B0BAxcANHyw/9CIiFq0
CbhlsZ57HqONXDXVT9gnpZLqrsFUl5AlNGI1HEgdq2NcJvS+CZ3XvUNnCITHAP/XeleDNO92cZ24
NflyQsOjsgyJ+owVJEK7JJH7wvLhInSsK66SaK3k/kpL+Nofj5XhgoCwjax8sR5hEXJy7JKhlC6A
9ObpvpcRNJl5pL8BG+jphDRyh9icgNhcR4/5IlZhV6w8GO9eigWlAnlqWR4ipDio+/VcLXRGdcue
MVwjE2zQMMltU0gIeG/v6v1Dsy34zGZNDqowuz5UIleoGG2CINw/oMDy0ZwsLmG0eu9IYnJ06Y3F
o/ebJXjvNGZNYwts7dnR7QgQrznRNLlGgj6actW08Ol25C3ykBIn75R3uCVDKqqfbpO8DQNJsK9C
yEOQ3dhj6lUo6vSZGSHLCenHaBk6QuQMUtNcE4WXZieatpyqkIThl3KvsDK0FO6U+nHT/MKC2x1G
pHHq0Bg0lAHt+mykXnfHpNmC4TGNteUJ3kr4JhJEVD+ZfF6Q8nHkcHIMXsu1bMrYi4pEL+9a4n1t
CSs18zvd1KsqScQB+wQhMbfnwCwDMe1Kz7whmKhZDKD6CaLRJM/PKECOix2pEIq0M/rbkLhb34SN
YNUe8Zu1v7FElx1JPTnuDFkBOgx7P4w+oklAp817+Wtjd3Fav0J5lS1AoCaFuQ6eUE4Wwh9v2v0T
KFSQ6cwbLjTJz4rfac1i8yUsV6WFcF2Hvl4xaSwfkks1fwkiPYmvMvC2E4VI0l2rw43X/r/HweMj
wZgoLF6kDm9lOTUR36koUVpsYLyiwXnKaZRWVBRLzC1lXqTCG5XyxuTRzWz1WlZKmCeStCKMs8HG
nE7NPkp+P3WbFNN3iOB5Rje5yJVjlwBh8kZuR0lXoBS6rxJa2lSmUm9GIadZ2IKlZEwA8EqsUcow
oVfwLWepdjoC8o6ZoSAUdgwBCpQ6vhMdFazlggwhXPYRQwRYizfRm0jaqkr5WxFQwe9bGI9hxuNa
4/GyE5kwugVSnH9InvSx6SmCAppehAfeICz3jRAoUYfOErPTXs+6x9cTYpURnmFaBzLhUtYamUZi
0kgh3AGruFCdWjZ2Q5icrXrbey1BiMEUqZzMtukRY3aMKZtHaz50u0LOzE8hYHJomPZ5R0maNe0/
MgAvIGQKXdo6nfDEc9yj5UMDW2aVMQW/wHlJ9NNNTgYN6c7F3fhoe3kMR17V7QAePENvniMa0Aa5
VigU+4yf67/3oZ0WMQivAETk86JYs+AexH/8kwtLHoUuKBEJdPhBXRj7t5JZQqrhHVaQLcZbTuqD
GCfqjGJgpHPSt/TjlwdPpq3h9/QkvRPfUjSaDkN4ls7xQnkszkuBY4onFMJMTDaWEMc3ziADP1aX
rDreqm8fqPrIuORt5qxb/2wzW6T2NrJ4qDxyGT+bqUobficUspZQ1GC+SJ5Y5EzllTR8M1PKV0Gu
9glbjtstj9yNAEExqyK6QvtkzBE2Iu6rkIvypCU6QruDfGyFIYgw690/lguyN+YIsgaywEd5GY7X
Q7W1ETuJFPg0VRJVAVtaB745EaaxnpCE5KMDe82dI1WF8sx83XQFNZD/vVyJkxA4hg5w33/O2ctu
k/llcwRqKj/d1LLf0WwsbC79QCXLM/NBf8FGKzrwf7m01NVMfAkOSN2Qvk+IZxR0hOC3dTSEp/eo
zAo9mVEcgMYYn/0r5IhL3pwEY5aZrFFN824BWYM3TyFOwzHFrwC11KgP8azwaLLfKQgDoCBLa/Kx
vabUtj/jrqQiijrpD/B4Hl6IE3gONgLEhKXRhRO5/xuEytyLlWjR9j5R0GlImqrs8ntzVQDnZpBo
5lO9jAwwEkiFE5gBY+z6iP70r7RR12j5hQW7LGIaD/5R89PzdngBt7KiT43PVjkG5l6Pe7enGmqY
yZxT8mIbywB05Wnw9RvZo25OoX0kLAoIapAz8fHJkBmzAsOEynZI0HcSiD0EMZrEjXYjEJEIeW0Z
YddZ8+VpdFD4fDF93zU6Lfmfc7r3BEtnHC9mk49hx9R1LfzaopVTOV7BheC4uGGv+ODq/sLkD5sm
74sLO1OE90cVPjNjsW64cnMs9utlWCrvj2DO0F1kJBVDniJcNCrWreAbFYVuVDtGWDwEa6V3Ds5M
Kv4DhBeWlzAaczjP8KSTvzHXhuNX02OajhWcxykh5ZVfJo4JIBilbcgMPniBYJLcHjpI/xtPIyEP
nziDKnsb1/A21rELAloAwleu3XucGBcBKB+MTk7f5WT0DCSXSlrRF9uFK12/kSBk++3KfUetJHyQ
C6UBeVjiduG7v9a9Aj6wQN7DlqUvTE52vvKEwG7Do9IFd9aYpOJ0zyjYFM2C2t8IfrLFKHfkAorD
HjK9b+ZsCWe7Ft8C7NUzyqudmWQNwLQD9JHsFGQ75KJGcnZszJgwI2wRnuLFO7Z+L3msVP1Eg57q
AN3I39SqTCreZET0iRICElZerUbTLQ0pIOk8vZeJiKSWFMMuHZE79kDEdBusFKpMaDjUzpyWDlBa
cFVa5PzpF0TF8h1ouAxd66/4PvGwsjY3CA496voL3MXm58YRACVw02kljUCck6U40ixGIgFhp3d8
ia1DalEvOPWvkImIPdA9WKZyrG7e/+Ii1ZC9LVP+dLnx+CJ95Qngy/MVrw3JXhy4lavP5u90/SQl
6d19XIAlSNZSAyuHziEc6hgQfgyn9ye+ApGj/OUYkZJkFUTf6x/IlIk0JQvmgrAUdnJjN+2kikHx
w0QxZXHMoSpP4QbOLLRrtqzgHqsm4WkPdpDCksESKmvtdRXM44RPShOquDLbu2W086H3/x4OgCcR
k7f3KH5LVSwPmHqOZvy1lM6oae8tbHZ/X9kIFlDuViw3T806U2Tw3/S/yyb2h7kkq9/n+agvvBhF
yM8vHvzw3oWV+fzYqX+rJ2SL2A8TfRbGoWf4EFPqitMruN/mj81YlY4t37iBnISp5q13JfCaV685
mFSF3G1F8fRz2Qd2XrfrgXs3HcGDVy9jyIskxo4Jl000kjKPafRrZU1mXchDkCxzk1jHKRg2rM2O
l5ajVAnp/M1D7pyJAr1iRWU0mCp87FTaYkyYxzCK9gVj6KTeyjux5EmmSzueKGhES2hPQtCM+OC2
7KaxZpDxgMc458gZOyCLiba4KNwPD3TTxjfm93q32q7SDTLmoF3k46qZgEMKGE2+JwElrMqefz+O
RLG/4dc2Gw8Nz+HaJHq7suI3MpScgHXbgy6FiSQEWkykKG9XMKaG+Bvus5yNDL4Huo01WEf3tDfr
NAObFXLYSg0GVsmy5p06gaI01GHBGmnJBySn+jw6qMAcEl+Qx8r/JvLyx/DEWJCS2JmEECghAjUN
xqzAN3SzA9NOXC6FqQWIwzfGtluj1cgDTF91ziBmwa21m9bpktyGXO9vDDPhb3iiUHKEktmiEJy2
S7M7OjEo2ivVO6NYfoc6TwBZud9yqsDG+k/Fo4RFPF5ZW9cIUJFFI0AuF7rv7n4p1pAGvokx5Jgu
08i5C1Cc+yIkbmt92MkotDyCJnsURugU2/c724tLuHJ4SH/KQaNSyUEk6IyfgMpTOn+Ayr0mXLyf
+S0G0f7aroZMmgyM1qF0JLoA1RONuKJuIwX0uMhg+VKb95YlA+7yVDsM27fOmKZJGEKqEFbbnjEu
V/Zwoaha7oEoWBiE+VbSI0+uL2ENYf4snnaoclT4S3RQenNFj2i/Qqi4JV2a0Nq02/SZxNl3+Nx+
QdJGDuXplc5OBnr7Sq3XgyXh1KhPFXdAIPr9wDf4xg4Zd2f+qnxwHKTFo2otzdEIv9LM5ad104Zt
ECokYDbAw0/BeYXnDrX0FVwgwoR/JOAjI9wkEUq8/UQuUEPjPM7LFI38x8bVOvnHqCt2iAmcMMrd
WsHvIIWd4IxfzWOAAErApzImEUmaMF/fWyCk5v72wYavctRGJr7t3rfkdK2G4wtufahT3Cl8H4UP
zEbMFzUI9pHAy3eXlK5e8sIkiQXddGhp8dJfDOTMK7ww9aQvE4SsfUy+1ruYPWu1x3k22LFNJj1C
1DQghBvWi4t/YZabPOU1kY9MzkZsS9pfHYkpp+xSrQ87hgO19ePqiFZS3dAPhw9PMFG2Q6Gq2sEn
gZUENbJQpAKYozo8AHkMgsZkhuGGai7Uv3dc4vAFY2OX2ZREKK7bFVMW48zWu7t9Oo3TPrwK7GiE
BdwNKwds4ry91Sj4Vn4rynwKs2qzqYJf+CYVLmk3USweej+WfK3yc9Bij9edJFNDFdfetpT2Z3VR
Wes6IOjrjDw5fXKQ95j0sOp4/Bx5iNccHicfFjYFRuZvkDks302+HlKyx0lhWhzf0vH1MVCJS9DK
5868PmanR9mp7Ta9iKDY6NeV+VzGGB8RCCpRIyAqgJk8LLrIXsFT7CaXgv6zfCqwrKWl/VWbQWrd
KRa/9Fyxk4BXRIyjeUd4Jg2j1QUKH1L4gMICw9ZxHLbrfeLOu8kkaLq3FzgE4S0mkGslzpqvO+bs
Y8geIrUEscyWe7JExJn/D3HLCZkljKnihwizV3SqhW7P+nPq8BCBMCNc0ksSUjiMXu67G3eem5G/
E+CssRK/fVi51aTheKgKg53NxJpZh1ISp2DyYoiwIupjxVyS63uaUdsrePKTb8a8DZtjtx5OsNBL
gauNUESCsm57Fi2US6DynNWPg8jPWRASrXldqvX4aCzKgyBFDdCtecRJ3yGt8yQrhqfd7lyUow5B
/CeI4wd1Y8zSEg068Oq9JT65OwJnsT9wBAMeI3ag7qU56EMUkNVoX0QTgvUZJth/YahrpNdwrJdf
M2QJZVRaMLJfKkyvpPcJix7QgUvGqm8IRFDkDbGDzEgjLip0W8++3ltLi1ndtOBQwgxp6ktoMmWg
AiBLp7yBJTnNtTAkz8/82V8dAqhnGwQlTQQJkWWocL1lu7NqpT99OSnE71IeEo+wBEnnx4L+C94g
fwV89bA0LRiwaTAVdUK53wC09CWZVMkBO0CoVm4by7CGFrjV7K1tvj6pE29kZ8VRLvxIwO3zod6x
LLeZWP8QTrZ4XJLUXsx1c4o+Tifvj6c26KYGaMiqr3W3pwJT2cT9gJ8/dtDHdF3afBVDj3GimpE+
EgNk6LVx2LHrKhskIAYLbFIOyg2ACK3CVTW4MmRn9j3DVZ6Bg5xYpT2Q1HoZ6hwt2BsW3FJkzAff
jsDy3HXucWp5nRp3FAM69av4dF55NIf02RdkfnuiObf/j97nH4HzyWlBvozGD6RRCdaV+Fz39Z+w
0a53QcRcc0N2SElEHXCI5rHjuW3zadlG1An/W2egNNtrKwAw4jyAje+ENAqGu5DBcv1n9mQbM4w2
CL/33OeyfGySx0CNqDQAIAGAHElLkB7+OVYTYUmiyKQCyzo1TUNp+Lz9Z7M4CQyVURxe3O2NfPDx
I+fTXSJNSEIhIZbdG5rEXPw3tkfQsr0A/k2kjh1ZW7+OBQCcV+XWRuvabdagbkLXhLlK3APKMxl5
jpqaFa+TmcTf3i9I4rGDof9lRBkcEUG8ffw8qyUQmK7fFqo3W0ONrW/43IsIGR+uvkVmk+ZVFA0y
1ArIKxXhLZxw5o0X+QauiTbqm8KOOwRbUq9joFyX4yBMYfTMG4vsA4BfvVTPd0kG0MlN4bLB6qkM
ZXkpbJbUuMlytyM9jeYwp5x8V/otNpTxDR4xghaYt96qpUlKlEGvfSa0WKfK1f4T6oHxSRSfmKbK
+Z/g6STOH1hmmOSHv+HmNJc+mdb7I+16c/M1hIoi4JMaTmOu99b1TK8y9waYXZS62Y093DFzTQHl
EDWsR2gJWAsIQwFf96l5jJSabCVsCVShwP3uz8FoQMLfxMoFD5ZFi41jJ48hPJQ7jdCAWfoU4rFK
NCitKA4uE7L3Yr5CJmaSja8Vl7+K4orjnRmIsnwrdrxa3o2PQzWdOPscpq46nAXz5LAJFoWT/h1M
dkhJ4SLv9LQdBjebrWiTyQelmszUrq8AaD5rS+BvvHGHPcbJlmekJXwBqJynZgIPsaMh1RlCP/52
i25MAPfpA5Poz3G8w7BAWIjtpMNKhuQ6MYoaVHPN1/f5rO4mBJnSVuRSZRq+hSX5dyMmKbRNEei5
OGui1AZIl5BYCv4OM657DCkeAAIfY2qKZPRPcTOQ52zazOz+Oi25SksIaWM+R0iJaV8EsPdQUIKO
YAFgYsnw+zhtwtsIKvgD3K7HaeMUZPv/vM4oGHSLYgTVrNUXI9BYZdk7Em07vlc65yXkffV+PQig
Qq02Rg8OJeQmRVZSm71XHMThjUnlBRkB6ffWJXGYlb7fHNRs40HEaEz5sL5JgGJbgc/mG8VXgRc7
CUioIJc9kjQ1CM/c/JKPkMW1I+/Gyz5Hfnb6+WRLIfGf65N+9xRozbA7gUpcNv4okZbi7+n5tC3h
He/cvdyW7zu6g7bYNI8sW1X7PvygbtMPVgLHlEOXo1Sq1DBsywQK+lielDdb3i2K6YOZQfz9RjNm
aVFwh0x+lH7ck0XXBiNIbRAUEKnb10fSnt6i1Rh+a5sZtODdq3tf3jpLLY43PLUjLMuW1C4iPMw+
HBoIBkAEajXe6gxDxW9MAdP6a+4LK3W9BT4ZCBOCHYlrB14a7rfuqQHK3vvw4yFczQ4WB55kldK5
xV2RFbjnc9hiEQFwR55y6M/X8jia+JVyTugohYfdbBRLzq2+L4ltpHVF9uW36Jzni69zEBZf1URd
+N3hQRA0ijZ+ZyNVornLBEK67+cBVmm5WetaXiJR7E8RCSCauAKqSDMHrisTL8Ln8pQ4pDqFutG+
L68LszxTlnFW13OrN30IIrx8xFcqueVs7Rl4R6T7QmkyhyofW95j528b3uoA2aiIfDpiftyscy9K
fktdscqQwPdwMIa5aldF3BvjVYQlO7XpjxP75Uaa/BPwbtCyTXmL31AgSvvnWX1xdXvr8qL1cScS
22K1KC/laSt1bKImovsYDGAkm/47dN1NM+87XdEQfO91A9r/cbGm//zpjNZJfRrslZ1x6pLDltTk
XYpPOFRNjIu+oSWOD3uRJddNK++9LppaXZF+AD0Tj35453Ul7d/WhVwPil45sZZAtetWNHIfz9qL
smkqV6paTbox0k2YT7N9Wwpo3TtPrAutiLovb3sPPj3hzs8unm4NNZlWd7K+uifaD6KnMOHB2sDg
+0kV7EaI3i2O9m23o3AZW7fDpyV594mhzXY9bMrApmEAcoSjYBvnFFiph0m/uAGMuHbKfNOjFK/D
RyUeynkbA21Q3/GgSsn9QmJwGlob0pM9XYgEmxzTdQSGyiuN3H4W12GwFB/HHSH0kI37jN8y24cG
RJpYw/yns7yupCaYX52IpsqwFpZFAsG+3BQWCo273uTSPkQf9zzwB3r+pQjADcMvfIMfMWh6OqQC
CVehQnLrLtQNjicQM8pBS5eM+We+6b5ouSj/hPl04grvYZ8Wlt+A9jOj7OuvGfkWQRn06DNalRgH
heetqRke5bJcFaZ9UFNok615Le2XU4z1FQmwXv4IXb/vMNmiDZhOAfDn1rjQRNDsEUysDu2kZyDL
83iwR6jKxWsIwI7TMxJCW1HDa6iJ7o3hSb2qN1VBNyQMTcFKslKwcecl2qhFTHXut64/AdRnu2+D
Ro6yVQjMH82DKjYENVCbfnOnBkUA+JITjpImsLZHsVV4Rm3dPB1ZhogaqUAUtAufHpGpGRHt/k+X
cNCWUQrD3gUcAqkZZyMNF6GHBqr2CwWpn5jHjt7KYV1hapHJbXLjgWI1/j2u/gM6PFc2zWRovpAq
HQ1Sz6rRHTVvY1srquLQl3IIjkhj6wpKWNh8igZIliB3t4ogmHhFxLNdW5Vq/RoiG/Bo4sh+9YnM
24YfyleiRvFPCUFEFqh+qDZ1pgSeB0ZQmGNfFKHrFXnn/V0raSJ2dC3OT1c8ac5wwaUQp9OjfJ7x
Awp6eYCQCKm9wrUD/KpqfhCiS9uOuxiZK37IMLoBHZYRhgbJKBogNKzlaqL05pnsQLwaopx9Nj8U
TfVTlLQ113fjd8ztnHYaHwFbpH6nJERkYaNqbPqYWRqW/n2E1Y3bpcjkkqoIgvcDXPjR6X3dKiS0
iecj9wvq8XeznV0d8l++maXCfl6PsLpTZJC52h2n0T6aQvt9IwBS1KMPqBCJ1NO7oFLLpcnaLbaP
5xS3dC4quXLmVr4qlD9Y4l772ufK5x2/qRbZVuwS5ZUUBS+3dHDLzyJMVRqhty9EsnENVRNV/PEO
SdQFEjl2dw4Zd+EpXBCETIedsaNGjZOtdWMCSzvILli1SgeIYXRIViqvkcSZyWG/0xuocJM2PpmN
AgQ5HrcF0J2FPm/j59qiU2s7z08U55otoVwdLz5IPyrLipKbHVRTeawQJGJjB3wzf1+1yoJ1/NNC
Nz7Ucc49C0s0r3UleeBNJ5ZwxTTlyuT0tDdQF/Zb/TZu63+aMXgCZi1jm4qkapo9YdfvmvCD606c
9O3akdlhqMvcpixV/7S0cp4PTUFPHbkcFdXfaFG5Tq8gCXE1RwFVcuYaSbd2MW9A+Q3TguyH0W7X
fW8NM9pKgNrgW997wPpOrRIbG0NK06tldk4lTCIocgomPkqehbgNGJKyyqdeQkDMHJdbp2b3qpOt
HxQMJiW0+ORYXabjm4pcSaB6d3wYOx76sOL99Wky2+mQDSeoGFyMUL+xSSr67Z2sQBgMdRVVZnL1
WWXjWn9Pvo5EcoAIAahrxWL0qCkOD3sJECfRWW52W1D4MkfHC0/9IcjFHfoSIIUP50ZDPPFNvFzc
BnNVZwSaIv/COYLeWkbeLJigV0yw7gif9k6a6rADydBrkzqfa9ZA2DzEIqIhmX0hIjKD7Vys5hfk
rHuphFM+/fMSAxsoTqBzPG84Dpk5xWNlOSZkzPy/5nGhPrgAX4XOacLvBubcM/vEIgzpFVcRaNBE
W5jIsCVr0E/ka3ZXRlXQm2keqlDc8JCEuaWikh2ty0uYec+FlCo/OsOSIvsYTGmZrWucyElGBjLw
xRmEYdP4Hyu2ZXNJi27PrZ2LMr6drCR2T6zuDo3Qx/rlbEyJMXizVtKIfaJX2uFIvMhC69dKeFnx
KwSKu+OLT4SN14y5xQ8l6hHx5aNf2FcZV0+ggxJkbNgaDPtMzMQk57K1VgVHmYTSJeawCjg2LnyR
IX5B+6YGfQrFi/b/apNAx//F/JKDbNws/TkJX3g5rYb60DXb+rPR0+4+1EcMF9/bLnIXB4XdRgmh
WyNuC+ZkghW2lsJIP9EBjSVfz8Z3uyJeQj771rK5/eQONSvaz8R/Qqo49RuPv0EvRg8MM/COHNb7
19DXds4vgcWmBzd3bROH+OZ/VKac9pTb7o9WW4WMUO0iLiXdytJOJoyhfRasqYDVfMEcXpzEC42v
98uDFaf44nYOg/4/s5ojOa1XeHaCmR+xRHsjIFSAwmOBjGCI8X0z9tvpy1Yh7tdFOIeU4vQTL5Ww
M/E7JgqxBwRYlZ6n6p5PFOTYvKP0bIS/6oprEwWk3q+Ko7kUYmZ3T64Aod0HpgoWiKTkOIvGgILR
vMxTskKGH/W9dDa7XMqY1iBDbAtwrHc4Z9rtKOboRvJaAiUTM8cBYOWk6OZEy/ekU6xGTpY0KDDf
x+1LoR/hwKMKI6OlH/1QaYPpRs5YX0dVhsYughvX+sEiGe0w3tsqP28rfNNUlpKqhQZOBD7QJdgY
lXW1qM/I8bLD/obhHl15vQQv51tEjtIM3cSTxd02WSVHCVzznqVzGHm7f9GdNygaw4Qc+TqHXrMT
4ywe2A7yzSwJU9BsJEyuzTtXU4+T3BpREIoVis6eeGArhuoTB9lJcn3neKD6NLrbLGMYxS7XsLC/
Y1pQyu0pEvmV+KiTB+KAr9d/+92rKPhBEcFK/FlqviKDWgSqUZ2mIWgaUgh481TNlSY1ipgrMBj5
Bi6VdTGwxmcfm2YKV/axaDO7IyqBoetiEEtus1pgjykvWwnAdVKLE6VpY/aNmrA7qErsBW3TJJis
rTjGl6gh2ZGilsWxD59AIu+D+g/YuJM/yBWvNhs9Ceu4XJL+NyLMl/Y8UpkWpvgDZz1ofy9y8ffp
O0TsZMCFCnf1FfsQYaxVajuGXjbwwMvfnNJOKMOf86Nu2wbn6F/5VKEke5Prhh6K4jb+tJAv3khf
jBmxmqlnSnGwEAD/m0XgJNxu6SIeX7iuPrdaOZ6h/d5sfVvNHR4wx3STOsXc3hGSI0lKLvI0gOtg
9N8TrS2dZo+2+UOCC+qv6WFyWfmvAsgGVFG7WLrWnJx9fXOcokVGMsgfividELl5ty6sqyPXAHvK
OoINYVYEe2rOKMRDUs4FnlewQiWtwBQG8lYyQqkAPk8EoPvmeNuxqkEyZbMgL6WKcOP0BKLikInw
oOh/UZ9ICa5BDQL4bfeaCedbHCqlfU4oh6REmUIW1w8u+aVqkaF4UsQaU/BZUdIM/7v3LUaPn7XZ
FUgX6POxF3eZNIXzzW6FLYsaFISnfsnP3IGR1wSQEKtfv26jjijJfWkM4cGTCH4hDlbvWJr2b+xm
1uItfyFRqnYC11qXjRCUf99H3CKRF7C7zI+kRM+XdQE2dfXQDtcIkNDkxaPFvurx4GNNbSUyY/55
7bEa+FiMiRqDvVSIG1CJEaHWLf0chHVLcftF0qOplsBKd+9pcZQncTc6EFT1KOBkl5b9WmoUChvg
gC2HbwoHq8cRXuef81Z2jUxh19bg8rWIL8QJ4isvR66Pc3PTdchHvRm//7kuUZ5FtkBd5qyL8CkY
WFfCOxsq3WRhKLAzqKEH0UNNUXV9EU9CCvmoEsNcF7AByK9B5eFnia4r9lBDSTPSqi1WFVxJEMV4
BC2cSc702wkC9fmKhn5Zg+ayLwKh3FgNyeVWjWR1INytNZ+oWDxQnkHipGmXhoaARi7Ym4gNALxM
ehc+XlV64bBPrk2NMwEL6Z00jiFffPltaxud61E+E2sDizzPdLz1HaK1M1Hq/3C0V6YQ8DjzYFSa
mYhdEXL+dNzzU/l++BNEY88wy5pF61I73gS4o7pbg/Ze8FHhKDWBZ9e9+AAV9MbgiIv4jXxr/J7C
XCMt3XyKNHmsAIEhlc5aC8XVC4qfQ75hcfgu7BiNUKwnjvMvq+n1YknY+oqI3iy8GslCP1J6eh42
aJYI+4G3T3sIKFVcDNEsz/jLZGIO1ZTiuq4vItwYe+40tGSBX5aN+hSrEZ0hdOeRnFCmWZof/sIH
lmPP7VvI/FqR8D5zypwKt5W5L6GES0jM8wG1+Y1uN6ivPpvZJ4O7eRnSYpOQi3hfKX4qxSgmgODM
hwBbW5xsWhhgS/ZheJJXUGNRSwyM3rX+/KpsQ3WNHWluHJ72H3RGKqW6dbnQG8gg7h7gVwDZs0DR
/14+xqbvESYwWMOiku+1yCTBTs1CSff904w8ebaBkLGyFVv9RbgI9I0VdWH/IGiO9fI2LHNe1yb0
+Pj/juAT98GC8/+GLVp0qwaopTD89sBnqYlJwDTQJncNGpK1Ywl7Mj3gX+OkmXo62fnFY3OtlIdZ
BlZyP46JVq/ip+RYyXcudwFGtTHiFlpb157lcWkwwo2axFMFGGIic4WD572wnlTrQuUQSWSMDOiG
o2yGUgy//PuWL4SeCnaH3JuyUDaOMTDTxWmzeFEBPMLbYU4vxCXvBnQyyzRvg5ACU5RzW5Zb3ZWL
568JJnptDljNyd1bMni1PQmbqwfuUpVR4hglJ6nc12TbJE1m0ROvOU2QGvE7K07hIWxwMojmXhxR
MfBe8b4f+8K69e86zmGyscSEaHeId5M3mj/tFOel0A/gAsl6HQIBcKnkGOruwOfZjfMDIt8sewgp
aP+XtWR42/xhx/c6++ZCvqVFXdC5YljvAU+vEGN7LCj+rw4KIHz/qEULQNE+0LgNS5MVbtaL/D+l
YWyFS4IRC2YBtnLBYIIK89M/Bdyw93Q9POgbt7h4IwLhaGe3Hl6hPNa0ANvWYiPDp+NP34JtMr+E
hSGF2Bh9NZK14tlmGfE9TOuTdIPfa/wu9qN179mly0KeUlic8KwO81dvG19QTLMzGzdsxbCNVZ3x
33kZfpF2M89YhUxu5Amc1ZEGbitNyscfVVAPw6DFOa/W1zEK2CpnsnBtRM7hU98J21kuzFPjSVt+
oPSa0GU1otk+iKlUX8D13Eols2Q23WHB0ax5yQFPKnaZwJBXAORQsIz0ojCQc6Z2GUOjqG2U3BVO
VDOQfqq27eWXHLLWKFD61gvILQt2TNA35seXunKBy9f9VoOIP4GosmA+7gF7DIZ3IY5EaSh2yIi+
ZNr6QsoOxWbbAz9+gaEHxJOyeYPVvhRrn2ZZ818J+0nwCwjmFXrXD/X0FTg2EcK7F8ag9R2AYxDk
YYr+PEK9Mq6gG1S9OQzoeYS/VZP860QvmuI7stwNjPVblwTCt9n+G1lQrKetltJUyrpvDGGd6k+q
wN8aMc9cQOjLGUxU7vkMOSPSyqRw+FQo2pjovG+UDxpjpv/B3rENlOimLq0oCQjUGpoLemGdPlS8
/1tY3ZM3lwu2S+wY6WhFN+Cj06wSxr+KRFN3dpUKU+KKrS7W9Teyb5YIyp+1YfU4PYy4pGKDexab
+wxaiGtxFXHExKDnTErpt3WlSelyZL1zGn7r/IuHkjbtcegKLbtxTvB0cS7PqvIb3jKskfrRXHqd
Ggqz3J4ogeecD+4AyLasfeR5/tqBGWotsn1eb2wPYsO2jLdFtG86toSWtoR5OoAL+DSr8CSFRRpk
YExTSeyv6ZDld/CY5MQ7O0QSoj5U5WD5UhutFaP6ul+5UrnOqd6N/TyCQSw3f3rntleMD+SQTOmr
dTkIsH3zfhCAGBPy5uw4VWYlet0OQJe4Zo88Yx9SCVFjymtRwR2K/i39rMhKDc8myldQcTqFJp2G
1I/CKEOk41T2uhifsw+CJY9OTMRIzsmqjbU6l2Vfir3jmf0SO8GXdiy+wjkg+36vkKK8RlPRJAGs
5gDnFowPpujQbsSthT0RdNT/njU10EUh1fVOSckYXUuXwHdOyiQDk6h221p2Ci0aLK8bcLac36m5
dUV6NHchfCD4ubhHsUB+feYFloC3YQm/ZMkWCKFflN0VkeuhKbksc3WvNAGMIqFY1s3RKGA2BsMh
7+8YUIU2+aIcdXuGdMXL7+6tFpKOBcJpvovKFImUiwSnz2DdA+h2ugjiRq+GYKeYqYez5fwnf5rK
JTBATnysS6vzvbhR59YkeFSos1SmSxM1K9HLR1SkG5lgqSudsjcAlzgev0Q+lxvXPwKNfuuDqFIz
h5Ixo5GMMQFk3bJIwaqJ9dvqZ4vpKVoQasISATU8o5n/WWnDbZR06eTku79tDtgqQW6N7iEda3Nx
e8ZntXY2ZdyrRDWB3jovXlCp6aG8p8TN5PT2WZL8F0j15lEcraXtZkbaKZ0cCgaT/z1gFKSzm/tL
/HsuAOlkxoK0xnHG3UoMpvWkzCY2Yr3pt/u57kAxWEZWGCD2m1dARXaOpDzmX4Nc0LzwfAYL+bGG
FDidtpNZDeKAnUviK9/9qGoK1l7c8eDqdraW1ofKKuV7u2KJjTlw/l6M0s3Jtiivv7JSRKwcIeAN
x7DTpzrl5PdAj+zH1Z155mEIjq1arJU8QKzS5bHsAQR7GT88evcbv8o97R7F+2z6nQI0k+2YeLBn
Ftirm6B75S+rcach3T6Hap2gNIMVd2f8sQffdATcHp3sQOEe2mXeYakmO+HQRYHxLbC0TVojD9X4
isv2VfCwO7XVOGkJ/WmhuH9mV/PHNwZkaRG62AFJAVbDXYk2KStV6gb+p01WmQcRJ/WvcN1H1Usv
dsuvem3+V9JGHxk34ucwy5rtjWqWrHCO0+kNctWv7s1ArNvWqgSjjsQAuYpBskb2AtlIVMzZ0Cef
518a3hdCilAJ5bxsLJM0EIE28HVTX3QYMyxEPk3QxW+9xcWDOR6Oeh2Qmkm1ul5SroT8Go7UlpYL
oCEfY5dmmUbxVVO/bMHeYFr/Vl4JKLVKXYO5efoLVDPqGkt94gPHljPIf6/JRaFpKi14Lyx98j0p
cWzqGQKGrFiHe9xsxyES48CD/jZdepxu1vMi3+VIWNCfIXvlV9qcZBSoKAo/1Jq1slaT4i/MrAWp
yD9ZWfpYSgI1lICj8A/KOv9f9T8uxHAMcf0qFS2ic5wHcPIDdR+gLbAKNAhfpH5irxvCp/81BcYd
rgpru+Q3baW62OiqUU9s6Er7zHo2xM4e0i2TocKjJnWfV/zsstv2E0STgpj7/US991ml56KA0jUK
X08Q/DHRcWa3yo2Nsxqc0TJtr8uOk2uFnm4H42w1lBKbQS8bq2fUpGbFg7zll/dBgUya5wtSzjd8
1fsVPW3XEcg9Y1ZMqMOSrA4nMvT0DUTYaLimnR6BMyF/Wg7ZqWmEy14itaS07B61gcuUnKn7Zpfd
aP5VES6ZbiY5xkHRo6Fgd9sNBJUTo2Rrg/qj+BwuqGj/r+iUnOunSMg4Ws9lY2lePX54N6n7S7xe
GwkDQ6pqHBjYQ+dEGOdBOliLYQ9bHgsWONcC3BCxET/SDKUwI2ZarV/1WyeSla8cJFzkRU/fsSz+
QCT/mqslafZ3Z/lJBClJ5WGqxeQnH7SwqVhM2LT5M39R+yvM259J/vTerWCHRP0VN/rqsHQRTcOz
e8LkjHqJh3QjDbQ4SIFs92RtiJQm+7JEutfeFkKNL50BZM0+rfU6xAMMfv/usLZ4G0vf1Nfjg8iw
1+7DVp9MX1zTn3F6fbKtvNnDb2AQY+r759GaGD2Fs87p1vIuDB6glMQwGuNcKlovWKS8hD/rjUci
fLxcJPseGgyoFFX/x1LLEF1DPDwheodSZophPkc92S2K7Hvnt+BuVf7kbWgJ8Zsetg9RtzbtTpE9
Lyr21kf8unZKdxIX28+qYHPKhU+ijmIrX1QCVHTxk3c2yC7pcEXlqUDRjQuB2rVhwkSdpSkvWOo4
FAglNPTXZpK3fDPkagQift8NmFmrNarOPtXF6Ai8WvxAWr245OrdrvTjCPt+XjpFmSEGbm9/+rfG
b+N5g+iFUJLr/jM3AsPXQoTonjC44i3UkCgbFWXZ9zQHfZEpGNE2tnZzsRSaN6RDrpI/ZQHdR+re
/S/gZrM3PFX/CljkLF2ExV9v2HPtHCinLWjqaxhm2hf43QK6IO4TpLAozKjnm+QqV7O7gPW0+75P
zgZPb8gByHCofqqz3VIhd4tWTp5j6HdJm28DvxWGPhnWjqGawjFCOBHAlHqzHlHUDbPt5A5Lksbq
55ytaavyMlUoiOn7fAnVhT573H5kad4tsXy9Ch1tf917/dlKuw8rtOv0AAxT1vfKPYspZoyPYeOm
imCQao21JKeqMC4A/yxoaOjGKjiDgvFyilWb9PuBqUAmSDVPxjLk51okROshvYHAgshL4ZpO2RO8
Kqfg+7O5N8jjatTKRSuWuW39NKZKIWtYJEJFUqyCJXbqhSrCyikeWytPz9i7vQZG0iRM/9PgxSxa
Ed+JOIMPZvJcV2uCgbhAzvQOfWSVqpovJmXVewgG9nSurTUdTScZw1RzljbdvWSdg6O4wR4/2oyC
CNV0ktKo6JZkeCFlaxLCfIJgCYYrGzmmuPxWzFme6g6d+14TkJ0DYK4yc5nKk+bZll+6xcgYqDU2
59mZHtrjF0SbDttxb8YjuI/q4mmGo/OeNlz0uGiP6tPFGUR/95E6eMXbU+K/KdNXaDdGYbUop7C+
zPZjOoLPpNNKNY5qu9DERCcFTL+loEIuS8Ut4p2PyUE6pcsnaioFDhR2Zma92fZ4v3twt+D339B7
l/IbNh01+Vu+iE/nmu/WS0mXLeVxz25y+fQIcnlRVnive8k4yOoSR1/Njhb87lizrTuInSjE69ST
ZtmTmgXFOZaVKrWyzgzB83CzJKk6fF/dDO4B6ZoCWXo+xJ8yqUHHNmixgKMZE0zSZ4j4gUttdwWh
FnsSGfrSh21a4/LD4KXrEUeV+9IapQ+Kol/DkovndsXgxDtIR5KFhxzQ3+3zgtXpNyYXiqAGhAzF
xDltOvWcCFHyODrbGGyJbiKBlGTQjQZfehBEYA/wfxweiPxk09ttrc1Dr8jc2kGT0nlD9p26esVQ
TZSLyYFBloAg9WqPmGu7cAJaDSXDSj0ReKTxeBO7t+up+zxkCm0TUHkQaum+olo3OC8A2ttVXEx1
5lsbcWHam4UiACdthuQWfx6Q2GEBbD6qDuxYM0ZKHTKcfaVZpWS+9wqsWeKAbqrke5FXgOI3wqCW
OlQEzLkxfqeWjVdLlMnHcQLLTBzUzhEDIqPyOfemtYirHQz6WKugMCU9gSuQBak+5OPNmn1hd+xG
CwMoUHiVhoVOmdZnkw4HNZp1xDZxAjTPk6LBBBODMWd/+knyhE5jCHQZx945qECnmizSbYij6kI5
Jd5mj+PxMMfUmmdjgFHba3IWJ7vw4POzVkopExfVp88K9yb0089EKxmtVuFzwj7gDbqHWb/jb2Uq
2txVrQXO01NIfpMnfLqqAanGSVFIeAy25JxChxMyoZYldVS3UrgWlC3VQSf5/4jgF1/pkvkhz6m/
2nlvzUrZNsYj1XrIKmv+OiRFTDihwPhwO3Si1PzlsaMSzn/qb6+4rlraWnX/4Uy0U9DvYwJ5PRxK
pair5SgbNoL4oX1g0YBh3/mqF5vc3NOATulpaPrxdOQnkT7IuOgrUavkwqUnmEKNCufJ0wqxxM0r
EqVziqeWGuYebsv2xivXEpw88OjFUaNE02SXuI9wV0Oto4LzzwDM2fr+XKTaXQsf4257zns3JM3j
WVUnfF4PkhAc1onX7nuPJ8XQyVKf/X61CldbqjtVEefoEyz95ZT8u9cG0CLUrq0jjLqvTHwAQpHx
GYwn4LaRzAqJY4XoYSxIc2cOM4VLdOtERg3JG3U184YP6nMtQS9t7ikDEyGX6wOeRFqA1o2II8VH
Hkc+dAcva1UmVtHZEzWEG4I1IDHjST1/v+nGNPVWhfAAi83cd/hbr4e7m9x9nFLM9Nn0paP3eg6g
5HMmoLi8XM6fQXJlaDYC79hXqsxNQaYMRFF6Wg/RV7s1P003KpicZW1Ue5caGAj5Xxp3VR6aaHel
nCjCxEjXwZTe5c1xuAuDSUV/iHx61UOG7PdzUAnCWcgIWxKdXgHiTh1mfobOoGbaE2/nqF7/6uCO
sEPE8A1fVt3VJSSUyt2ED+NNMKE55g1K/+8whZ1bXzB2f/sr3p2NOvUvmHzclhiXvdsluK/cWAfq
Abdpem020wVKOG1rkE3gtYJTyPdMf+NAI0ayBKJpL0iPx95cSgA78Sp/Slab7E2OOEW2/Nt5Shw8
SZ1SKPHm2vYQ8AmF3lF11ge8bqBjfz3x1UiRoN4aeqTb2hgLy4XaJgNSEqCn/JFqQrhEXDyn5Gmv
eEDWWWXy7y9xFB7Ing4Vr00RSMQ9KFCfAOhBv54GfSMsjnfK90xsv3nxBGUW/Q62yVDb3xURUh5V
4JNQA6Go5GTFSfche7wF6I19s9ta54SkM+Z5kRKdQJUq1mhbP5eUGNgSnKk73IFT/KEgDG6DrKgv
eUHQrL/39b+fDb//uaPjwSi2s/p14ki+O/4hsaf/aAA/1kc4ZBaHam6hnnKNW7+MAYYqEgvBGpjJ
9L445LlyKQw/xwhDQVLijyTHndc9/n/OZrAXi+8dO7CrIlOW+5FkaVNsZFsiMKHEfAD7eMU5Jh9V
WNhVorWVkdYR5cWkpjw6X+YpKi71vSBqDIQNVYV5UvobGBh0XwoWtuVIM+bgdXItgDxioLF+RlEU
ijWaAZO7Fv5VUElQDWuQt36GlcdACP2GihzUs9nYxovo018vnqr+9Zu3f1tSa8HLStg1ZecaKN3h
xVpRCvbhKqkXTOku2v1G98041MCxg/dzbm95+OaXffZFDu6CeL2kWOZ/OS/nzIIho3We7FMx8310
OtEIizwIYjERRSjIH8PO3L6DV1JGIlpcOG04DyrNRSnErgpUvtLUaUppJ+MWYSTu7oegzv5MQCDt
HjA4+8Ei9l6VTBEE12jcOl0PYpE3kcB6CuBMWSWJFvgoZjoK0WzHDW3/kX/87uxFjuSoVLRiho0V
X62HE0wnNqgi1aZxDULhrb96Ebry6wcqMlRqhboPSXRIwLuoecGkf04hR2YgSqKutxZ3jRWMIae4
aEkqY+9Rr/mGlF0qtPWPj7eNCfNdd+yUhGfKErtWKIjG6cIyyAcebf+ytQfHw2ERr5jYH9GOYiw/
PMpDlIAb6h0eDVDzAi09U3rSKoMfn5Yj7JjDNbci5F1gIVMh+2TrWHr0ACUF+0l2Knel8YfVNuwm
8j5w89Us34CiMKL1fYiLOY5XE2SBsZ3ejGUOeOAYXsf9LoW0qNZGZrq9qKNRoJkW+M9PrDiojLyZ
48lLXKadaefhiUQW0JgNUGfte+hp3FARNCM64Z/hAujU35kKc4NgAONW/2qyGEcucncxSqfb/Up5
ZKBcoeblmJsoW9/dGVcT8XGq3WMREAnEaRtqZn9N8JY8qhogRThwZK4eKbqrXI00q2duMc+fzPKZ
isQ1Xq1YD49jCWVaMU9tGqi/FJY8YVcpU0Np4rsTV3LD9CyL9vs2D7RB8BVa6UTjimcX0hveFySE
6gGlMCmkrG5re4t45wQFezwz9CMXyltv8Khk58aqEe398DH08n/duSxiSZG+KqGp1EjE4/x6ITLB
INcrn9j4e+6SeWVPFt5gfycdEEMjEGtf2Eg/gFtIYgzl8cJcD8t5FZeKjGwrxbs+Rcb3021YlgLC
NIyr/zqDm72i2Ag3yN7ukZeGvR/1OPVDB0/YENPXF59MX3AMI97Ao2yO8cXJRWExM3VfK7P7JrfA
6Xzp1z2MW99OwbmnCy4Bq59p2EtwqDW8Fd2kC74LlrnMdmzRyrnP3QUod6lXO73m+D3WtPJ7o7Gm
w5Fn7ZFCTeZQqXilRxGKT2mYE1EgecZX2Mdd0q3sVdDZTMBnkKZqPd5FxTu+ssKnDX97Kj+Y2FLu
T6cNqHzhms8XEjSrKqJBdP2SZ1ETNXe9j3KpYmgqVASjUvh5f9mbdntOLsueCwvTlGPSmfxw1rSC
VAAfcdRj6Dn3+oyRe5g8trt6XgYDL08C7OqmjRF38KeOQOcHcWemESLe5BuddxjgSGxrptLPgMOF
bvZubfB5UaEmdduktyXOxkbUbrLglXvAuE9w8FjW38HH4Wi89o4m0HYwJaP600oeoJxb69QbnwgN
FEj2n5blNvAySyN7q4f+my1hxo7VIXJuL6zKY0CDJJLvdOMBnqmoF/c+d0Z7hOpM4acwTalpWQks
14hXS4fsJqFuYHTMRpvyqnFQg5WDMOSQDRO17W5ca5IeSppsb3GnKaafWIFawQPN2NfBJX9buIJX
5aoMH7XPd4KENUveeyZknXAXwr5/7GSsY25d/Js9UOkGEm7CtNHiFQBUk9ZZsUOjNR3Dfu1zNYaE
UeDbKWyOcK4bXcV8FF3UYcOtbgq8oS5p3t9Wtv3X7CAvIauGkFcdjIDcmqCXLGwXxUauGtD/jYkY
UODTRbwuCkkhca6Da3yPx3Gg0VkHD9BgQcjw0dgVSAL/oZHmM6JWtHl4uWoiP3EbNk/39YA5KbHK
eC/rb0qCwOmN4Y7x4K1ZCq+LfJDAhd590tQ1UIIFVb7b8QDLpsSx6zHNp31ZR/ym0Z8BXMNcvrG6
EP/sKjIsYC+YJSzhbUfOx676cYKWLYKaSIOoRhDO45oPJs7yl0yp8NfWOYJuvBe7IgVlxBmFzWeJ
dnhUK+3/sUbcfNyY7XHeiKomsXGHke18P+PwgUab/WBoVNE02is5xC1iOjkf7u0L15F5M7KQRJes
5dcTQ9i61wYiDZ/f8jUeY/X6Bl5q8h1QwVyELoHdGfus1HAPPPkjoAd2Hq8mj8eV6Xx/ugnjg07y
XMS/JnLvjJtQzM2CdwOX5ajqawqQuh0Rq4vuInC84kQzZAT/kWGi5wy+qA6XEpvbAyIqyPqwcXns
7ntuaufoAqZsrccXfjou+gmhGqTCaEiAK7+tiWofKGyV5FxQt78v+liGf781KOzkYeyXkv84tqFs
23Mou6Mk3to2MDXU8uuLyiLeYY9VJjJuWOXP33nHBon4Y5I3X0CPeB/CAjZxIq3O+AcnJlGKHGQ4
nuPVWVuC7xLEmy6JrBy4ag0LtcpOquosc5AIsEA9AJ+Kr0KIAxUsidhN9jCfATfDxzWpY09eSvE/
gdgni2zvj9dvgBNHrD3M1jqXqgyy4qpt0xGzUvf0IRlFMa/3Gcp5eI1KLtoVuztrqJys3dVqHTgs
k73viI0GcLvxPIQK4fwsg2QJhVv6YC9gV9mwq2BD+CYUq3NL2FKgVS/S0V+pfjz32LR92TjQPcl3
xwnwiJOPrWl+75B0zBu5c5uqD+/0QXck5wgtHYljCJXyTCXycN2/a9V+71UF3eYZO+RI+BasQl4t
fVEVnvCbLKg2Uz25towGFTd9jMclcBYGb+vR1JNcPWaMwfjw/KpHvo+hcUeSDSAsZzG1LEzZV8KD
pVlAX2wC3LiDo6MuIRTKOj2m8dv2496JJpEl2NYnFkFmC9nL9TuNN5F+bDOWo3Li/L28OCzJ4GQ6
X/O5ET/PDbzDWtWoo2noKujiVEqz3+FQ2el/Fdz3YbYL32Z0bQj4g0D9ukZp92kSwdzd7mQ39+un
TQrlKnuXLzJPNnFwiXgzBr8X5dIOavVTAGQvIDLrU9YdEaD32OTGvYqbFyp/tdPF3pSY3MZapEW6
myfYU7JUgZ/nuJoYIOpUS5Pv6u/CttNV1fjt3B4Xr9Cry8cvds7N4/FkQo6I9ltnqBrcejn4iCSE
C/mUtysMksmjStma0dJiAP8vN83ZGffnax0PjkmS5zfaae9EszVn2kX7rF98Hy/DMcSFvxiYuBUB
74zA1zRxRVEwJrZbB77CAgi71rAqe3rRE4Pt2/WBDGxYJxzIVjALchMrbetyfNjcvqw2Z3RoSzJs
o7cgCLN5DX3150j8BPB8FcAaNGoniqetz3TNiQTqaIaew0J03uCJkYGtPqMMKK4/HS+EVUPvQgjn
QuSTJs0hLVCeJXX9w9nuiCx0N+Cf0qeVPrdmI/OwFRp9I0Rf7hSl32UKlFl8mH2rZA3y4qA5Nq9i
X3cQVpNDQxEPgOKOCP9Hvy9snmon69N24niOcNiqcAU2z9zL7NEYevyRrBzit3cDpAd4afGZSAwt
tHYT7LlJTfKCTduVvsnRrHhwD2i+8Pr2n+jIgEWeNDBeDxIolP8wiWIkcRsFsW0ggOwfJ+/eIyRa
yaJ27OjpGb33irdNCybB4EnjQ2aWNNwcw0kruk2F8sveILkOrhRBNlI0Sh20s/t0nrVIczHdTM6r
g1GjpLcXHSxdgBT3ShGyD7cuadwJ1wwG+sX4Yrcy84h2qgLCILP04lF12axMdn2NnCg6fFqFNdND
ybXU21N8W7M8wXr+ykGqca2Te3hhIdsnrQK50wpZxRSYwxsJhUfaeqaOSzlhUMp/+UKyNHjP2sn9
RSibzOjhfaSn1FFXgeIuccj5Unr3HnAkdjN/7G5A6e6oeV85E4Q4V/O7M8ISnexXsfsUENIlL+PO
51v0rXW//v9a4HQgwBY+cWkNDDM7L7QpkkethVpp+ykMpM70JmTHrD/hv3MunCb5Kz8LTLfys/b4
PU24PN1GAxiBboxuy7HXpSftXhW7w6MNTFaT4awmCtYCo1iVdcGRsYAbGxSk9Jhkk0z8KIdJcBt3
xtDcPVJkQac+3Prsv9Knk5fkO9WdYei4H9yJawMdm1PEaIpVrYCNSXU4jVvfoG1CJSnEHqM91uYb
D5VByvBp1WP+I6CinsxWP1MhlA1KIry7VzlrQlnbJHA3oNpAuyLgmWW40t2Oe31C9Fryj9A+BpoP
9zPim19LJcorW+1TvSgVoF6FGuOcK9o4m/1L04jr8dTWXjfr7NowYnKaFyKAO6TJcv0iiyA36T2H
6PekBGysaJ8YPiW/SI/Cf78ScZUieniLD4hPq+0znvGkv76t7A7RYu5z1WTSZNFOqLHD+RQKEiMY
DBIjXwzv7H719M52+1qqhJYpeGCz4F89nz2XdBwmZSLhmGV4EN2JlIWSjygw37Y0oJRDcRf2g2ZP
F87bhs3ZsIJBDoum74/6oE5CVD0eT+yAVHoAPWyn0gwEy88CDWrVLY04mdoXTF2elojKql3tHuyS
Aap3Hk9//142obCqcRSCJobRcvLjQ9XprG8NhGJ8tM8uq/dQCqkYUSRFMkKYsHYlt8ocmTCu8kx7
/RIc+I4N801L2udYYJpQAnNef3O2nKfudcxsjq3kaCSgvZLbOQLYl2DmwrrsdFayzMvpTIeZPrsM
9klztF0BRvmPRqhYOAb6v7bEqxCoxMneOpeNJE7WlXNpLOGBpC2rT1QZYMy1EHu2vIbC16mehefK
2wzIVkR3vySSUWJkrjMHfAzYyzPIlkC4LOsoSBtg17Ex6vfTewOsWqvDhz76+bVXjYV1StiIEPXA
IxicEcoSv/9JnesHbZMEwfU1bxt2dQvKCe+qw0wyrAM3Yf4nSemAzU1UWXz+czI5ttjly7y1P+O0
+roZGWigf3eu6oyKOaPnezufmDlZwRqbxNycw9Zm4fyz539zZXLrFkinTDTW8pkAQHj1MkYzEygk
BeqsYKHaJoPWZjxJP1gzKCVkVLk9Y542H/vLDe4QGGcJ/C088UwY3Fmc3cUSEHAsS/R9NmLsyREX
MyDPtK6z9I0pTaxbRRmhdW21h0bFrmsKjCnnZffIRU/3kYK89PIc0SDEgNzknI+rjpz62fwSGFzx
tuWT3d/W/hRvoHL6V8szC1PwSoe9LiF937B1ZWILjvCQVq4NC/bRld4g1zioZ4jausUBc/ysyPeI
thdeu8k4l6w8opRAByy5OoTdNVkFbDqiIXMRugHNRLDmaltQfmcbPBz77E27Qd8KKnz0gonV5gcT
rPNlh2Uk5zqANhr9m98ysh1mc0M0ucO7YhPcUNavB+d7TcgolkjQ+buGqx9PZxOZtxsRkHJKgtkc
GIcZ/3bNmSCP00PmNnkSA6/2wlLwBtuNEbUH9RZdJ3CnTSUQ8G4MWOZj8PVsKcOopWsjqZYEOgX4
5Mj2jJ86zah6w/4uk0FbClxMfRUjF67E/GGBMSmNbkmfkHRYpbUjggn76AkitVhdAwWHdRI/yj9L
0eIsM3HNoTGD1EQIVTO/X6qE+w8folqKm1c8khoMizrnxQP9k4dWufKvQOYvfZyRJqT1UPlOHf4J
4G3fADIVlTSn8OgZ4enX390ydchQC7tF5NFN+HrS129KEX5b05N48SeeikuChROZ5sv7Oboa5XEv
SDC7I8iFRzr/8wUYsZh8T2MUtGwlPdjc8xZ6VN+YRCzlx29TqlBemzxh3UX3SPysyyhsIf7kBpdx
CxBxvQ8AM9FHerPJDezwvBXuI68Fmktk/hWfgt51fxg+OKV9Z60/uKZ07Ka4s7MNcymOzOhmyNYj
+FkRrcZkwFoWtlIqk7oklJVNk8Oshbykq2etZj3Db7mpHUd8dUKVgXw1AOWDTsrvh/cUjGtyXqIo
GWZjImlmWLVzV4037w1rwAdm4IeKdSiZffuwh8FdoCs3XnmfSlg0B+drngrgiVv8U+ldnBcyoQWm
XAOFJHq6+UJMdhZcjBFt0MLy5NKR93a/doG3ShTu1sIz3TTtwtg92UKYv+QoW+ATpBZ8rphe1CY9
3xkwUi3BxbvMPIXgMclbUKToTb9uZRO+X1GDVf+7uvbuKs+I25fDDHvv/HfTjBrOHbiSRhUgTsXh
w4Z95ubCxhsH6KG8wByNfWzao/r25nzd1yON6kKNxT8mbe3KgV2LjTtBt6rVFvx4TrZAyN9oqI2q
Q9tR4vJtKST3MvMQTz7feSo3sD+ieggxsiIQX+0UMXMyn4xhmwHdCVsnXOxtx+hZxqqeMEjqdtqx
kMkSAkQGKqVlUeeIvowzgMrHEuqJjIWb4nM7yLs2w4niFi6T5LJf2pArydPID06foIFtKi7V/9Hk
Z351chQWIKcdmxbp/yk7rShIVUOLTa23nTeuNSoBgyxctbZPoLM21E2/HDxJ66+epk/W6WDmSSBX
z+o6PI6Wae589qDsE0mTcbNYU8pN9BbZkLohVpj7fqnidzd/kaTLosdbxjAkulALfBJ87T+3xj6G
MvGpjuyoK0FXL2rQymVy6i4xLFuIBhXgY5lZ+5DumNkl96KRzkjUw2StVeFXQEyoJc+XqMn3hYZm
1qisj0IKJa7+81PUB0ddHe0IBfc8IQHjqv09zEVVgrXFiO2icIda/PkHnjWsH/UMcKkGsFde+VCU
/N3CFTFEzgeh+otCZieSGXyuf+yglbHgS2sM7ywgFlkcOkkZMytMB6MJtSA0nN1X9mWY4AXFMgE/
Wvesz7dTk4v2Vpmx7cFVNraHHwg21hKtvJKzbl2SdjDAeaFhGLnKY1lBhA21PAkN2zdI14aBquDK
mxOuD0gjyUKRYXBm0de3bZYkvvGue18sSbLjhm+pXjyay77+AH29jPAEZaU6LGi9w2LWd1ip+f+6
9Rpt4CW3sKZOmKsVRyuX73imnH0KLEXttAiRT2Ak0PwKLeklj/G7s9savyPN9hpmwEb+7pkXBvfk
PO1tgkFhJ6LcD7v+4y/itb0bDT/U9t16olgeGJ8bbGJXukZlKqeZV05xiZgwkq87bl5mTfCNv9dI
GsQ2z0Rpb9arTNqeUChVIGBuYu3OXjLI4hMjNyOfGKHcauaIHhMkWOMYLYiQQtjIJwA186yiE+6m
PWBiGYrpeQgjNxkEEKyfJVMeYefi3AE7v7HItxi3uJSbMRAth6A+FtbpTmKq+ldyb5hfpoDIXSgl
eX18eObjMi6NM06DKWYE84w0dfsVYwFZLdLSo9Avbvk53e1OZkUVTMbgtVHM1cdlQy2yvdde27Ma
lNcs5GjLxL3C44ikeG5iZlxL7W7Ji3WSkVMHGZpuX7k7BbavZrgttm5CcBzGxJM+D67M1k7Rv7st
tVxy2e76i4UpskQcNaL2R7e4sO1cjMkDyK+dtg17VAMt8iIqFACkuiDOyOjSp2Mijf1v+Tl0izBx
dyR5S3dNaNLFVU1Wxj9bLW2GZST5q/Igba3PybUToy2Xw84xNpppx+fQ/7Mi2nd0WE/Lu+Zjtsql
c8L+iNEIHOaJlNRYit0jVbBMU6tqXRnf7IFDLYAm/7yCe5EwgIHoIFKfYBZICEXHyUenJ16XGSv6
AKhl6oiyKlNI0H71E/294iJdL0b3fAM47nEHZEZvXtv5Xi2SSEtQw6Vc9LBQvYR5A8gZZaAX3Stt
W7oKHWjHsF3XzfTX7JvD694gW9rXIgubZKLeYuiYVtXwH9KOTAMo2UsAKYPwKj7GVdNWpb36ATNX
3klOTvqwqjgZKM87Lr4U0t9FM3y/5QvfD3PlOUrB9qmGYIldECE7NYR48iJ4+cB3DS7BylYqbHZg
7U+xaFo0aRDQf1++tlfRWSQEu0FGdFszHr6GAn+GjvsZ5wZcbTNwy9FGISDIHi/xzLSZyUHgcO7Y
pPW2AFgk5FA/i3CRMnkcL53SrRUi3QGUUcV7uCGj+/cnd/d9xY7pmxuwMC9oLiEpkXhWahhJPQQ8
URw04+c5vSfsTFpcCKE608Jcnwlh8DU115twGL+fFRGpQAbfKzBGdYRqtWdS9SqOtIkrKM3s7aWK
wuOX4qaGxiE2QoyugckPdtRDo66+QUvkm/TQ7QCzwqXqjPy6qY1pCpyuQtmnxnBka6kSgyae/blH
QgqGzVScIQGNivp9R60CCshY0fl9K+VWsca/rlsU/cHFB+ZSSu8WM/pvV/yg0TtF2htfG1MdrRzv
hCpaxy1lVy/9h03r9qLteQZ6COSBtTr+FAd7nGkjqBBNCGApu5ibMvqu/niwkaECvQCJaKTsGIZT
3j6CQOcWQko6l0RXx8xxyl7yf/Vh4uBvrTJtOyqC0iU9H+EbVfWpUYUktlK7KvA0QnK4regLeLWw
m27irP+MLgP7yLrv3/YEhM9dqMzeVsbhgSdDqeW+b6birKZ+IC7Z9YRJS5+Xnb6DPAcp9y7wa8cL
Juq/IE+hW1DkImTwvvOB8+XIAFYWMq+LehfaxfafgjcZ28tgVhVwb6StJvK4ORb29wvJ2TcVnviN
yqTHLfI2NDYemMEEFrlZ7fd2PVI5+QfrKsK6VdJxi1VaHObecW3IMBjtkUdHUrVuuSoD6qBZBndD
IVo/JEA/fiBb4gNc/lqHiMrYqHOGmeaNl+2q1m23iAMPg5s27VRDTQZ5sCfxSVYMr0z58tBOFPte
BXeStxkFuR/y2+gxOIytwWW2oYNNmxV90n4lKNWN063ZPBh2DlqRTEdUFiAa3WmBPLG1wup4P5Vj
ts80uEA9d8oKMoTVhCAkLASdOGIGJg5r3zCsI8BMmdpEgU5BRaBRFW4BTwsB1+64h9S5ubVo6MyU
QPGtt1WNWE6UgL13CzFL5fpdijixAJnS5G+ymuBuhXSPwNJq84iWuYx7HKbm0KfGbOwfM3AZeLq8
FhySd10b72z/79QIzrCAw02XjlwMPWOEUhMkV32eD+DE9DR5y+d8g8OiOKZray5ujUd/oQSIbk3N
xHkrvo/RDKF3nO1uuAW5KMPsjLBGFli3i/TMHIvxbSbV6Yy7cvzBl5StHK8FrehKMKxgUkf6Zl0Y
ApaRkd41a4QrNaTs8XuHopjO5fWojXGBtaZQ16WJCNE6VAgDLW4CH9jnpKghOIwkB6GJsEtxQJ1K
4eiUFcUwOROkeYPLXIB8WWksyMd8WBX0m2hpfBKeL5OFEBb4+5GWUzcO/jDCsZ/WaP/NVNjQV55K
iPllol+UFfo+WMsEY3cL4BLemMmxF+ZglE06fC5F4YJGK4dJ4oqCqYMFAVHV+4jwhSqIYcPWVVIB
VudzjDlzLrJqsNvct46MBgZWpiT/cP1X9Jai2U8/oRgaD4l7EAIb0yY1ieNljUC/o7jf5Fb0jsod
9qYxMCVqQUl/RIQj/Ljwp3AYo7tSeU9WzVhK80rUSgd8lyH5PDm7EDc/Hu7SjveDYEiw9ptnmoH1
gnIu4ZXuuJfpcm6rj/PAGrHzasWsVcICf376C+MlMpvyBh3NNV4ofm4emEMmqXpZdqenKH9kXTk5
X7lvnb2oLDjv6vdH1ZbktXuOme2JdfWpGqdMCxW3C1F8Ugo6N1eVcRmtwnY0xjAClVvw8T3TaXTF
5KATCbcz3XXQjHFMS/xPsIUdLwVSHdcoLadZz7eXK1ubWBq9ERpOCKxV8I64nN3DJaxdwjdmqST0
X3+pqKj9MFUFgP/zFKA2hf+gY6JI+a4MRvzc8JHcx1zCb5Ee7x3IBMO9SoUnk7K3U1lgR7ryJeuK
sopqFeZIp2hd2nxAfatyJPY/m1jPfYFnqgyInO0sv7BR3zQNSyYbNQXws2PZX2zUh8c8v8U8gIDG
silV3XLT7AQzfMx0EXda+qTN1IgGMUZt1yLyM5rGvtO0gnjlNnKd0qTg6YuknBHTF/TSDi5CoPeE
SjkBguSMVtMVTk/KESn15euqbb4QBVYYU4RgJaN6CY+zlW2NTPzynBj52avfe6uP0yZjgHSDcVab
FfVsNlEkpPCqRK4BvQMNaU0dhwPhIrVZeWu7irQqWQf0xZ56uBe+yIVLSUdVDAT/8LlQsh6Oixji
Eb0nQVbJCc5mT0N1MWy2c9e49h1lXjWXt/R5JNRXHESaNxJtSTL+tXwTMlBchWHjAOelFhsfVeV9
fAVa35PJHyIzPxXsaPLZCuXYnE2B9TIkXkmeXn89A3YB9OAc4WY07rFMiWF5ZBDjr8a5QTjETHS5
cy50keTGSWZU/U8J27YS7yrn3FWIAwLMDK2h4OPcC1K/tGfIXGxaAQhWXKIMh3ULdUC5xB5I3cYX
DuGoCRQYwvap8FL9RZJXKwlv3pi6nMu7NsE5sfp+d0Be7ijrIT9n915F8UGhT7WU3129drre+Fma
dhb0YSmdtDRZmXD08eVeylzjR5ktMEMY8K0Tq3zJEdHiIav7H+tLxgnu/dsDazb6N7aZH1h5eTcX
ssboPaT59+6ojEQyGBzjp6goWHiHdhpT34euyxHdUkeEwZQPj7pMC49WlzMdwkaV416FX8Sn3ET+
+VzaKt6nVsQEHhEOi8Rf96e4RSiME+x9LSXAyQlYB4yeYjapBBOSCXKynJ2hzgTNUZYqyHYcQnu+
Up3PK97A/9dn6pnQaHe7M6GdR3rFeto/9pRnHYGKyVMWOePbCh5NxBotv9zDCeOJC1m9os6ppZPo
cjfDESfz2cqhEpjfhaYtzdiinF4275hrq5N93u9XpqQqdCcZICdaFlctnLR/fF/Y37811wK/Dkhm
sbgjkuXccqIFTPsVZxJJzJz8wtb3eK8jB73Rc+JLiu17L+LpH6gJkoWR0WWz9JWL3z+y8dkT0MPM
H/lH8Qw6LCg0h0TkMdmRCQpJj3/eTDWMC1si6VXAj4OOE/PWFlxTdJI3arzDftM/ZdDLE2WD7wWf
cAyJbLn2y0JT81uJ+N0GYkXK/UoYY5o8HVRQ2GcjeEfK9gI6Ayfi6F7G0pBIloPfAHeW7sWIibAn
4BOhfK8VkX4tcxDNsLr2PQRNvgKrbtyK09RPKiXnt3rX5CEZzRae4JfnS+I4DbLofaopQFqjm60M
Deua8LjICPqTTLlhvtKWUH72DkTcJQ/xj4JoB/SlA/aCCwlXxl/j8xdcn35W4d758XPBMJD8cRyI
2/KPF8cwve/DwJirAaIfVTd4xT3Rxy6FwBGxPwlbY/9Xo3sc1Ggw1Ra198hCLT8kBiCpq8iENqF+
0ny8RLH/Squ9WhWQbotabnWvhCO/GGd+S0N9WRWFIjgPo+LEHuKs2jxpLZLp1p1c5iaZGJvAueRG
N245tSGqu7Xx5gz83sHABWbFuzDvqzb9u0yauS2rFPxNwfMBcaHIUD7BfHdNct7Awa7a9ZEeokIQ
j4XXLvUIa9tHxkzjcOrb/if1J6An/JKZkLzn4K9FQIijQ6Hk5a6I3wq8b62iNQPr8zHS3z6ZNJUZ
l9+BB2FjqLtOr5xRg90G2VjI21xD8yIqe6dJOTCQLGZngLxOGvOD4JnkHyl8YeLM7epg+FZmsGHe
Gar7gbIM4fIMEWv82G/TfAOD3L1nhpPePiWj55MWf3oKk4/CJYZDUqeQUdCEWUjgiZq6JlOdHh5X
l0Ppo4rj5bn2II8QdELlQq2kUefNFmQCYKvV1NdgKnLYFy6WIJcHdPk4MXsoVNcoot/mFIDPfAyo
EY7NIq0Wt79j5Lr5lohBGbf1TrQQdFjZKkL7GXi6jYeUZ66VQ4KEN2di7g70uJcpd7v50bmAgJ07
70YJfzKrgN5i5G3fqcMezPizEwUmq+okGadUoz7XCJ57uQEkcs4RYzh86PdwgxSOD+i/qquTMzGY
UKz7Q7YwVeFXy98AnPTh4OPO87Jk52JKxtENBYgS0jMRpWaNT1IQosdYfXWZwebusw8aWqWge7qy
tMLwcV6PEOVthgzipqIBq1KH801zoT81lOsigwFi8fvC/NMWASe8cP7anNAp/8noE2y1ui7/bhPa
9VnIdi73qoPvnqZwOmiRp//WLN+VFNZqDCBpi4SQLnbibnSz6L7JQ3iIkG7w150Wc+3UHHxwJdYw
aWjjWtA0xxS99SujnXP7fzmqTBu/znz6JSqQEp5J90NL0QYfIuojLs35JoMQ09SOMWf+VMHOvUi7
uevhricW596Ekm+eop8/lI+hW1QD/WS7WsXVmA6Edk++Ka7S/sJn/ByROfrel001TcpP9ZnOBy0P
TCgKrrvRWxXQXiiILtKKg095TmnnNgHmcFI6nBL8BxGgyyLk7xtDDlBZS3dO2Af/ibqbpAEvYxlJ
CwmfcZvnVd2glDno5huWiuoP67VBZDwwny7OGUa1pb1MTFPRm1cRmmytflOt16+bGtIo8zbnbX9b
PX+uZ2JaTrkX4+sg21J0YKvbUN/Bnfxgs+xKZ0lskj14NLWAyx1//G5HCycVebWFRekfySHLRiN3
7Eui0MY0kM1KqzJoCikyl69C8LV6p8/tBGGhIUfTRqEk55AhBuej8qfiTZloKekYm4eIKfJmS3bi
EvMOhFC4cenzWHM696J+UE35iIYacJzhsLFtcerZyEPhF4tS2tsMM3Zk610QJLnTYOd1ZXUiIXuq
6eLnxV5PGzYhW0rKKE4Mocovz4qS01zZC4451ouGG3Jqrfsd6/+wfgeVGSbeNonTjZw025xdMPYP
dkg0BWOzvU5r6O9QhIo95wYhKwHoZER71NWWr9wKllnoESN0bjAvY7KVEV9HV43nHKu90u/B0YHA
b9o8Qift7+Jwlp5mGDi6+DT9JGmHaZd/J1Vjxg71cW/o5lpoavewGrDxyT+/z9YlO8EQ+LLln/PG
c4i9NSXAwCjqj5jhuVAlVBZWwnKtCLXb2+xMnpCZeSel7iL873nPSMgJccsoMnhZzli0AfaMMzFZ
cCQ9abg+GKwhwzShppfJtm+lrieZ2dSHGFJeJatCmW663LqYLN7TwtKMc5vJ/T24zplvjIUVylEt
Bvv9hf521QyRt6TmnCm4kjQ5xHKstQdu7ycDVpPFqh9F6I2/b435VGXdk7za2Dr9ImrE+Js/pop2
GMUdg8lj0KLwwTWq1JnOalS89Ft5AhDBiiG5Hq1GLqCUlT7NHS2QC/dn9TJ+rG+0dmKmKYngZlZD
iOrL9ZCk8jhNS8lgh4RbBOLxYlkW1AD8PMIkVlTAEFZmaXEJx69+Wk6u8v9jmQYSXewis0eAsxoX
3GdWp+OX6kLo2QDdsEPeaG5vAV28kPmu06IgHzSooOK0UZOjXOj8AsiiqOM7Cmy87HxLW/KWobcg
HDXF9/yCKxD1vRmhSea6yoveUqufsoiy9HxQoGLaY0zAtxRLkQtlBo9sjcuXNRiCoCL3PTpD0lph
DtuPu2RtNuMUCqbVfFj6iQzt2xc4GMDlugmT0Y/1sKtQHS6f06f9wZVMD8BnNmic9qvsepIg34S/
g8HzptikJ8EJYe2dHgDTJVY3GxwCRw7gdPSmdASFi/RFN0jKlNEyhC80k1DdInZZ+xChEa7ub0pi
3c17QSGRmg/e3/b4ZzvtRW2jFir3MoKtQd11shlfWfX7l8n3gZLqs1pey+KrM6Sl3q84TsN7k9xh
3zuxiO/A/ntN01ktbM20OWZlItqqUDFGy3Zro2Vn0ZS7LfiXCoWh7pfBwnLy7xNXzyrINrrTOs4j
gMO0dDkHa1TADZ1Z5JXfpr94CpSSlihezDBPhRMmB3fHAr0yfouha8UPHnx2IzCv+reXwcukNz62
xY0s/VQFPIWUdGTk7Ct/iY4Kqi8kmQ9yJFv6n69824kyS2TTGriNroHWVtzvZ30ZS8pVNhRlegql
HlwIajeVM5+dHSReptlE5hw67SfXbXqFQuPhFN4ZZDxPHJp7cA/g/2sCRXcRFfw01hCmI5NCbzbq
XqN4ekaFD57QU66VeKQT0X/4qJrGY/Mrdqh2KNQZ/qc3TxEHPHwf2VbpXAd/ZIA3FxX6eY44SEzm
Yru7uLvwS3SRaNPfH8kKEFyfoMDBngqzLzUOy0aF6yWEqqMuyAME7uYiDmDne1zZGXHqnOSwlAr7
CTdWbKLBR8A94pASSnP3RtnA8ruE7MJZugqRLupBoVs6/RSCYo0PS9SeWp96CJjjJg/vusBmRMfA
DbQmSOOZ7O2QdwLsZddh2gYsfLMLtKECFQ8hFFnFMEEZ7NJRqCRCkemIJE3032mZH+1zCxd+rVnI
usFbMdsKbZWcqkfJ4JGDfRW0Y/jZJFhgkNO5i3EFDT66OHCNu4l8UXsH4HzrhMftCBct0XRlmxBs
NCZ5YDiCNWW21+G4eWhdYiA5r/Fc6YKFeiITzTKgGMelEdElbviediMZNELkVq6TRHq1Hj1ZJFVh
c2bpLYVmzUkkv8GAB4Ho6uY4wS2k0K+t/t/8uVR0O2/6Cxht4kyyuk6rSyDstcbG7d44DDO7aKjn
sJSAohNLVdkwDHczsnHgVlFV+ODtuGF6hmdBUqMHhCArNsUR621x5hkYwuJ1sXgfupWb6kbGrdPP
z96XYeeLoewq0cpRDRnzU6X1DoZETLQko3H/Jw0x2chpt1vTGHnACJvUBABddE9STYhhOk2Jue/8
u3X51LIhBf4RSRl+97Aua7EC/ksxk5xR+gt4TR/gV3dWlOeDWoHnwDfbKm9NvWYzxrhZPFWHLTUs
xAD5ih85ErI0FPBsmehsTiDhQGOJotXlf8hyFkFC2s6e7i/8UcsucB5ruVizpexikoCXoKJTFJb2
gw878QMLCD/+zDwLjuClI7RngAp5JTnQ2i+iH1lw6An6JncgzPrQr8ALl1zwu888w+vI/yIdxnpF
Eq0Am1xY/PAAwhR2WVddZPU3FNp4cpLaIZb1Ji6MVSDo59pIgUcgBlBp1WX7yonTnZtmo6ceEzws
cAUeTB76KjtZLtta3J587QuXadIkgO0SLHKPAIaQqvPPobUmp6dHJzCValuUxFDN/v8f5VWt867R
1anjBv1ooyOTqal22NKOP6yeJtCDnnyGigv2EwVIE1h95Ugci+w0YojvQuuFFUQDob3yDtjFB2JC
GDBSVu+IIGXrPUpNTyI0+LPHFsnyuzO7lZk4NV7mNShrI9YSt3EMx45wI8ZvfPZHPv7Z7rzOuKo0
4ZHiJyydgyEHqi9Q19B2xSoiajDRk8vDJud+tWN7XQ4xMllIUlAeV6Z+EBjMeTDGQq96DAfmQy/6
vb2sCO2lwihtQYsox0+WcpVytdCCh5HepLeFRmhAoXy3TqAVnUqrNb65qBhjGftVoKo+kr+38aRX
BBLfOUj2CS+R0RSQwtk/pmJaouFeAbcrtINFURaOBMCsnip3rt3YpNTppYAUyRYCVNohrAcPLJJQ
Ya94IMZpUpYTmMVs52LpUph5ErNnByP340potsUGlCrooqemdjq1iOxD+UHUdEYNN+V6rDJ2S37q
U/zZ3J2UFUYNwjxISQw4TlnatZvwefOiBZDx+Gb4GBzqNf4UOmM0YoMP8uww+Qu2fweB/OL09EmP
t6T4kNKydeqmU6S4P2um7HimfFLQC60PVCBZPwYnyZydOV5VPjAWWUIky7bxm0dKbcz5axHwKljU
+Xa4Kxs3UXtu4S7qDzvBgyWBegVVgSqRje+Q3ki1nZqmnZ8Ne0cRzZ8a5cjzySvCwCx/X6AqbgCn
p/0Ntp+LdPXQwnjWQ8QtupM5P0pHCEdY48hBOtJNRzJCeZ6hkOVOMw7jqRlbfvY2tLChtyFB+Ump
kIAlX/MKbaLSwABjNurW9yiotlhcCuPxHN3zgeum17T/zwLW8H5Ku9Zh2DowHmm4rLjUzNWD5Ucq
KN2OJsNkklyeYER1ROcM+27wqwpjPi+rPAgb52/JyVR5XGlW1D0YPPCZ0xIlv2K2YaSzgwmJJyVJ
uOOW9HAmAvcr5bnDh+H3/z7Rj5HuZtqu1ztuIlhHxvgdikZuQS3jxi5mlQ081HuI9FH2/2LdlTM+
jSUlTwVOgAd8bqWDLmlmyR55+QQTB4HieENWb08Wb119oVCX4rkLWcgtOSP3G4HPlb8CUEaBvi14
rTL5OVkalnYOHfAlewweP9b1FQj5ibRxeV4TfedANW9/Gr45TEOOJ7E/nvGkYjUuKWPOOFsWHZKY
igcSdNp0wj0Z58P5PNfAh4MtqDNTOSw+dqbsTBYrgND8g7yd84dLHzHmcFJS220Hd4lS0tQpsR4d
EZ1dSGslAw7389iuLNWFIXPqHyD9CMuf7sUr0QiOV/dpU5E5t/NFl43hjzZtxUemPVpOyzcUQsfl
u8khfTZS7t1W2HiJ7ULN/K54MLJuz5cP2Ko0CITwiUomdNaO21NwTFV8wfh22qj5vY/4xC8qu2ij
WyGQVrGGkREEOjwIx8blCpdS467SWXkAMTWcPv2muDMsPzN+W34ZwoVWgERPvmgzS4Hgb+Gt+5WV
c/+At2iiuc4/EPnbjISuvpB31F6uNcyVVhapwzNI4mkpYQK9RsuVRsYw4C9Ln3MVA9yTgpmft75t
rcYPdUv4FME2Gy4XJ4fjGoWoSiL36mpws08q+U/5qRVjUpamzLuO/dq++bo8pPsy1t797ixSU2P1
dkKCKknKt/O75OMSwDLlZhgy0ihBIlAjAYv9o1rhcqaxc4P+1RszewOALf9KSxHbA4TeO3gbH1oH
9r0zXKijqgeMz+2OT+kBUtLgY6KFIC0iFbSl8eVsMYauUl2z+uEqDTWlUuQdBoKGnXml62bcMtGZ
YwxZiDhlBYbNuD5dPl204yx/jxm8kq0AP7uTAk0Q9Gt2Kwa/97NSYmFbvj1kL7GyG46KL6O+c/He
U36H9BcqllXqKhuDON1MsVGNW3FSHOXWj70LXxtZwNm07kjuH89y3CV7ha7zXL1wChpwkOh/0jBZ
rkGAFaRlUg2nzBrn/U65SHvjlmW7DzWANvLU3b+Gf5HhD4DavgJxpOLbR5brnjjOlLzWHEhLvMua
NZMjxwu/mD/khxWOAepiYK4Z1ZLxlqZiijYCOxHSktvlpz282D7omGraNr5vqsN1A/ss9NTSkQNi
h/iHqNFKw6i9nC0yMH6e3yjOMye/U268qrp1rn6Prhvbmj+Duz1wMC5w0Kd1hs8lPLfzVUyrxuZ0
PYcR7G0Z0FsvUKRmHO8rUhtu8a7cSkH1d3/5JNMie/rhDjl/vCp7PSJ6c6vChxBAPSMKcG3RCUpn
FgkKeQJxNRQcyjj2LEEZ+FnJ3zTg+RK5OV6y+7DZ6Xh8PpzJO0vdcPSf/PIgcnFj2Y76k8eF9pb+
6/bO0e6dhGE7pry6nGA//79tr0j9yEbWlk99k2iOPu3NNo/vhtpf83RWPhgMJMv88H8y/nzej0NQ
6eC4VvF2nmgi2OuDRp4xdfFatSaKzul484bTdea06BjJBuHsU43FTost7eWfLR9XlqnogFE//QZ7
8URxFKppyJQuVaxS2Bd/cAV+0bCXelwv82FCBvdWSMoDJt0YF+3pqRF0zLSkU341rSvkdOmeYN/Z
CyqEJBb0vG/HScsQz37Ykq2RaQKSHZR6a3cxbkTd6ETpxFWlYy/ENSHjAoZ4lyU30EoSH1+Q8XEk
VzwHbXD6nDIJHZ5hLKHmUMM8WG29blL6P/FHG9A058JygtUXF7l4J5JAMGN+3uzPJZnbbbnCrWjC
25bU5Gxj5iGg5a+mePNcgSX4dpT2uCpAiAbA5Tv336XWzqqvvtPsow50mxXlerIry9DXjmGY8Miu
VRm8d4e/sXgM9s0d5FjlK/qqZhxuEVycSRgxe4ycuZcuID54HJouE3cQLLEE8F4SLhFVdsjGEQ0E
S5c7MoEeMOlpFP10Me48LJFc0R5xLc6IzyRGY8gt5SnCu+7vxO7+Kd4kp5VaSn5+yVWhRgyviI4b
560OEbaJIcEe2IVe9qEStLq6XrDZDtbu6ktugtNfQX3wn7YIoNrRdDlKKvMxlHH984Z8nz1ni1OH
+m09DJsdMl9Vu/a+wt+Odu4AAhYJdbg60U4WyFlazP/WrXXvcFQFLrXLXgEfk/EZqm+dkqPi0Rg/
Aw32cnDiwOzTqNF4SbrEuEwHMyE9eu0gMQu5T3gKYXeuOtwoHfR0GkhDTDFjR/1KQrFWaxxh8EkY
nDIpgC4dJ5qRm8SyK4bsgBbztkErkE1ZZrVN1ewqLZamDlC2ZdjB1v9A+0X3/du4xxGsqMzz/RV/
Ktwjx7AugCPheTPtTQxi3YfQ/p+pRoACNntGc3kOtrz0d+Xv///sIU83/Z3xREEFd6EH85uwRdRE
7nz2GZbzC4K6+mKi+1oKwanpsP26dXHB6pVbIEqAuB8KJP/5Snd8S1HDsCdeh8QKb0KOIwPfcd2l
EBKHgCpUpM/zyqHAJJY9fCKlM708YY6HdynKjx4dfyp93OVYvLPMCzpzVuZBGc2w06w2BZ5kRURu
a4lScoom38FrZ0ypQFK4LrrRBghr5ApLqcYchowjyUk+wQKpS7MtVPtOIgo5ssahjCX15Wp1kzFx
PoA+ZO/1KwQhqy/q73aCwh7cbow2sIUbycGcJZ0+G+A7PCW+bSyb+RobAdMzHbMjWz8RCSQsiVmI
0XXy8z7RiE8g3JFkVg4eiKfQqK4hqnpVLSRnoO+2661Rnns8CazEeZbshXNozCkBlcNGDMbOUYmH
+ZoZixWK9KLQEUrQ05NJWySqPkDDRgWBAJ1+cSnkvX/LjuHJTnLH97/3OD60kJWUEoiocmUCFxlW
+aObYKbQ4fv4nlstgA3suMT9my+YHRxJIf4WKXHl9w+aiXFB7orVXR2Btu1Mpmdi2QLoD3FfDHbo
0ZFC1rh+sK9bJCGn4Zngz8yAf1nlytsrH73NWLWGfSg3L89pNxSk7+AvUfW0E5LHH0sfqgZBBxHX
kZ5rFkoPIhZhSfSXomvjWVm65XIv/mYx9R/Ad9r22nHIMJftJRmiwFsc+vaN7GMjWwuJhVlO6rzR
eyP8W3lnD2OYMgvHr/E9unh5up9nC3oF8DeXxBxf3ySF7UUge1D4cslY/ktWRrW7JSQToOgsGgk+
9djWG/h2W7JA+QdMHpvC7lGY0sv5vhZebuL1USTym6vfytXe2Hmo6ye5wMTDhqSQ2L8zaNkapT4U
kfO0fNxU9ywxFPoVYW9cxeFUVKkHiVPlECm0s6xF2fwSGEmBrN+Ai8Y8bk43HV5FIy7G73ASwkHe
9d/rLZWMWOkZ4SXEJeAn11CPS/Q1urUT87z0BECzubczlpGU4aP4TIwGmBXCsIX6QJOaw6q+V9Ke
IGraf1Sy0J3JxN4zYAVyEjHrGnoup4uqUfWrBR0sZRV9VIHJDGdLXmnJZYHbi31l2CT8rqlQBwDo
yF/YaOabiNzYGIJSPRc9iXpwmf/okeACQLFl5iJ4kMst3kEJ/slIGzSy2uoo+xrhneAnsiyP6Awa
bsWAxojXWBgoAWJv31Nw859CzuV148CJKf7fLQ6rSdkMASbObbSCe3SQyr1yBdOyR7PAPZ404Kyj
6kDthiQSytSCOj0CkAjqSBBO0KGaea2bMLZZCphWu1UUsOgP5cR6RQKoJiKQQDFckJnMElDWHlqI
Xrsyp/7GBncHKhvmVU7BCOuWxQXVkIAN/zpLRTxh25sIjFoR3ntTdtO32yZIxgfTnk8uX8Kuo4uO
tdTN1F3MDrhnHgKxXv0NhU4U64o3QWFPl378uLLJ4Bk4vw8YNrI5DzikZGGO+Ta2Mm4vauAP1TkD
rQpa23V+uDLVA517rtmDVIjdv6wV7TenDj9hN9EvXVU+w7faIpnowGmVuAO6RpZvNa215PfeXLGh
9qVEeRUEMSlJbOlrCS4ASQ2eFykgJ0CAFg0wCOu/4vdIj1s6u1/+Y7dveINAQZxQtGV6UQDEBHv5
a9PiKMxg6uFFpfXshXa9TDn6f16Yfs/xcA6/UvkctUVx2FHvCj/0Apg8EauRhJqHhVnpQLogtaoA
9Ha9jEeg9EA/KmQDOmuJmTXOuW9nLZps7DR/JLM0uY2hb3bc/g65c7eVzvO5MwKs121sIXAyuWAV
E7Ep18mFHFDLBp/R+wYnpUCh96cGDmblmnL+Tjo7Vo3Sn3aN2rW6CywQ67glP+hP3flnJ2FKEhdv
xteC2JwVtPJnjDYs16LrhaYRP9Jh6Ow1OO+D3ltntOrDJCRsmNPqMeIsiWEMMejA6QkyA3Q9DG5m
hctJ09+VGFHSobIK6rh7TtA04Oi+VmvIcWhCwoVPDmfbjBV5iiY2+FFbo5/ty1uuCnS7pkBAimCp
7BQh88skIvtWbmOh5Kdu6RiJzuLB5AKQGvMB+3N7CIypLMppzpbXIqMwBpQIuORa7AhNao+tul4g
ImyTlK1c8a92/Ypq+LbkomCe7zSjOkcDbfF3BTRb3AB9xd7iNK+qZkxoQyK9bHiTu8/FdIj/5n0j
FhADIYdaJaszQNPumtmwQseCFR7wSLbCC7Zd0MR6fLRZvMQStW2tgDH5bOwuxyzn3UkrYO1gjYHy
IpoDRzqGtpAuqHdeyP151IavNPifrIO1pgY9HK8XGXo/XhBuANbPyQBWnQKWpf1OBCADyoEzacg7
pyfGRGrItaR2/B8hilmNHKjL4QDQnXCws6Z+3WP/l8GkRuB8FroQhmM3KBAe1SYfTsna4PIO4Ptn
ggaKIfs2kG/luivEC3YSANjEBMzvzgCFxW8xU6n29F7wxmejruecp48Lj9yXVX3ClfkValKbxnkL
+LCJzpCUjE/IUBdzAlxia1fVSSUgKNEKptFunm7eVdQCkjysk32tnM4tfwnw8SR4ou1zskf4+T+6
2IITd+P1MaM/IFy3GY674sUueoAjSxeHxPcTpBucnBefk60mB6LfDtG7+/xJhC631w5cEv/WCdcd
sx6r2ZXqG/IdiXfOk9orZpkWUV3qlaB1+dSYsheKgvW0KnoxkJg07SwJ/KBWdPUWwSrOWpLzXI5+
lzMh2TBLzndfFeXqI1NIM7g0rXjfsQbHiVKnTFUyiGpXo1rihpzlYpnDLeeqzNoY+1ePSueT3H88
5gEOv7pzbqmJF0LqISutI/kPljZaoYbjnzdmF/HI2fnxzS4JC0qmApQuezsUiTzJG6SjPXzBLumT
0qugGfdubUqBI6SGuWItVlDVs5asGpc2J2fuPMfpWJo/ytzScvm59P2OCQTvdiU2VORjLiTlQ7u5
18ZAeMrLxvJA3vxKc9w2vZPvIc9R9KTLBxgmV8EhHXxnC33wERnL8f3kehiIsv3EYm0cmi6pXBDB
7/8UeJuIjAhzTcnkSmsnOWiijgbpjAv9KF4+3s7ijqJPlt38h/R8P5HMhRlxo+8hh/WXK5rN0ie5
RatOAJuPrB7xJT+61ldaPGB2IYgdDz/Z1i5Tmwc82HpylyQHb77dzfqDj9p1LBOq7qHRgHwTEbra
Pz8z41cAGX253D0UD+ykxaayUnKRmBHPGYzQ4gobmvzqaYkKDqQTh+WiEWtAcabX6BL9a/ZVvFz1
MEXjS3F+12TuM0xjifMwxHvYUYU87DiXa97Swkeb0/HYRiWvJ+eIuyguSvPCCeByovgDLUwLD/SV
4fSWdvyHKs83Nc8hIpSHRnMC+mkdlFYvBmo2VW7+dkdnetRP21g8WRgDVFdmYdpbI2Nk8mUjTNQm
KLaAnZAIPfpoiTVbPivvPZ2OnaCJmCLIyoubSC0vgqupOzRyZUnbZ312MEJH4OmOiv01lmrvdqQJ
86aOOansC1VSANsiGvjnuOE+YTjmAsbgrfXF7Tdc4kL1Dpu6wogtcPjkrIM6V2JZVIe8d/EXqfQw
nHJPl+wdfaQacfTgNHh/XrVY7LTQrO/gsbuG+n1DEFdVGGNPmlfgdyU1yDg18gdmUVDmedJUV6+N
zlYlmIpLnXxpML6rtHYGRwlvRuagt6qUrRXegzvl0ubO4ACtWVFKuWGCYbk86O6vvL2AXmy7/Zu8
g56T9g6nVC7JQKOTiNeLTAmZdx14uGnoUvcJL1ANrM3TEWKniwN5UQLAJJ1Gg//kcZ9ULBDK0zuW
pm2PCcUT6zsztMUoLVfuViH5k5nPbJmiWQZE5zHxcFFTL8b4lj1o3i//tPdOUQXOtoxNZ2tl1enM
vBTw4dUAapB7Q3Wc/6p9dsbm58ZLXW+XcwGqjYER3yuXIgMEV9Yszjei6lq3d938d/07feVFPtOK
K6WY/K/9Pjq3ICD55RwyVrv7AvwxYUTQDhNNsxYhIMuoIi9iFgd009g2EFdxaEUbauQxgaeXLURY
IRR6jjouJNDWBt3hqRWFHtJRPwyifRcykK7dljdj1kMddpto7uwCcfcMIDsuiZvz+4BJ4IzgVYKW
Qt8olkYxkG2XhEoGy3pT4yZhtopJAageY+cTmLdlTSuvxlFeOfiPJCM0vpHa2gTLYAq7kPodkE3B
xNXthdt8QwfWb2+xFlNQe/h/sdYMYdU4Jn2Q1Y91Xc38CYhUz8JB0wJsQjIm141J38e71cPNOsP3
b82Wu6XvXwrb8g0PyY4hdXm/BgVsitotyZ0gRFi0wEfJK7w++jyljKeH73p3+YIW9ikPatvDx+oZ
72bTlVM2adFHABykzUxJPPxyxPyWh0GsVOSpaG+Dunkrb+nVNccofT3wkfgwxUPB0TUegrYPNs/E
ONuOMLvxgoIt0OPR/q0ovmJj1YC9wYaJYfokubVGk5djuiga8MZo79vnb7SJW6Xx1HPVF08IN+zT
S5AqWJ5gaZhafR2ybMqc2gxm9VG88WwhO+zmChVlH9LHLzkNBQ/wnRVPcBudp2MSJQ+xM0fRs0sd
kEw/Ubbt3eZbpcHqEUNV9Rti7frIBJvCDRozy0j2Ld2O3whVFYNkmDuPHRUPQ1Ig3V6Rb6NnV1pA
CBrn1/cB3AwKeNSfoRh4zTo5CjP+KUnr2DlFwoqiT+rupAM+FXDXpO2AEUQZCRHRpaZ3c53/c7Pj
E/OApuI2ZoAfXsub5NkrK0vBGEH1m3bjkqLTIFtSgycdH9AUwvgirpnbDKM1AqoYH5cM3mFxeT8f
pDWpxtld6NQmbLjNm2LxI9Bjri1GQCA8mRHugjW5jlAgGy0Oh7X84jrZhTEP5DS7oMgdjoSIBkV+
KtDxFPvcD/EH8Hq9NzWveakrlcC3CGb/gYIHYJoM9p5cxTSE4N09nRAHbGQyVWZtjrMNcpvIETnP
EknPJ/9pDerplJUc68biw/HaGBqMGbkPNOWc5/aCapROHxp2lLRim4TrnH77rBgwETalU4jlVKHO
n6ZaMeZZZVoqufZ7qlO1dteBFpPiiDT7cA5sOFA0yG5DXRBUnWJp/QhqFq1QY4MJ0KGXRecTbt2p
aXpXC1NlOEy4w1eM6jsDkhZXbauXQUw0G/vD+/UqM/ANuMgr0MoanF5cpu/99pJ3xVnspXL2JeuW
+4XWNsMbFk31/O5YvNd2MWHCPG5vn1vm71wPPvnWZ/+GWzG6j6NUyVELa4l6hJR9NeCjNNU7QtO2
DBqPYF7p5EHOn0S/F/jd6Q8IMFRCRMZXvduYaHIfP0Al9+FzQCvjGfATjhtkiNlYYJRFj5Fox5cs
8MQZrgaLcBkUnjmzdnYlovnwaQqJAGfhDD2LffTWEafHT9wO53j76A75eo/F+fDgLAkcUPUsC691
r64ZTuDQYk2rpshk56SzTgyGcuVraWCJ73HAvgbUEdTuR75zFr6zzvdPYFaOvNF6kdgukIxXpZgg
5ycb+9K2JU4THmWaAgkarCNk+W95PtJ58FIbGktFKIYVlrtK3W17hDJIuI1V/Di7KP5SNzFDldp6
ktBqlMnOXYxyF7IDmp+q6dlLyt/MjeWn+hdUmKu6dPYCAAtQL07j+HwJlAuvTAPTBki0VXu89TU3
QkmLUIttpB/xJS6FvRj3e5MB+nnqHQ373tJUyOFZdPVMJYvztHvRN0kc/f5Ppab8ur/xr00z24Cn
Vz3Gauj2h/rd6WjjFQ+1I/Cwhyv1N7L3CpescPxbBG+28ZlF9r4nPCRSCDkXGn2tb2L3ev/PMLaW
2pqQ17oMasEA9EmFvAhB16BLZXxXB0RVje4CksmY2b6akXo58g/FXxn9hUNq6cHLAfS4/IBDpPdL
xdM8YIxXFAZHIIKGeLPpWhJLcowgbivHveI4Y9xstXxQYcgde0B5SesF+sR0heDIPbqt7S92GzZA
5Lal29/NueD89OrcRL0uCcx3aW9h8e9quhKmR6c762vvdTEMdvGJP8kw9o9R4mFNjCguZs8ZStji
cS9Xvs/BoXju4JQOhqNCYRZMjOJaL2XbgWSDhFio9Y8tfBOVqkyrswh2oqE3WT8AcE9GekM64C/t
vTOpfRpcupP9GrVpFayqIpWfkpAjdZEtljFwCbm6dqN0ZMCSb6P+LY3F/WK/j8ucNprUwWI6u6HA
h5jQs6WXFJRs3dCHamWLVn0E/4zRsFZ6Vidr/2NyYhLXuiCnQXNtHKSsgs0G6eKGsL292xS3KVdv
O6CpUAF5rx/7RyuFZx5WEDI1YQInjbsEaAiaHCoW6XXpIq3r9xwgtmf/GP7bcs68fYSDgpTOrNP+
ZeF3nLQKgJRyfVmpvWlugcUjl9Pb3U+p5xirdH4sYdRXW+eK2nXLGwoPQj8GQEEVb48b7g8M0Db5
QHeqU+S177GdapmYT9uxTkJWVLjVCmAoOojZWY4Y9T0D4rEJb6NwAqeuHAUvCEzyR9zngrntg1t6
ETVXQpgnVF0kCBVMVuieFpMPAyIsm4/7SQ8bRcK4qr6ynZhk1uV4wF7gGU1U5D1qHYT+Ri5TWPaQ
JswZqqoEdIXQCJwJSNZ4SLnLXiy8nHhTj+cwiW6rYRzVtEqJ9y6kRrI2qVPByJesmLW56zo1I522
8kWT4iWC27m8cqLHX4JieSHeKWvj/FwKtwDPHWNo+y41c7a5SsJgpjaEMmN5eX8oDYhpcud+SFJK
iZ4rS0HjJR4nZY6fIhbidLm7ZkzsKBL/ZIz7nC8eS2gVz1Hq6fVKlw132YTyeZ7tv4VZ8MEbz2UI
6K6wvgI1KNh4i6vx+UPX12oDQm/71dWAVv+vRaBphqFNxwRbzG40eWz/o+gfUFr0SrMIPL7Qp/61
fIrsPxIvknhQMqLD4ue5rkQV6ttEtlDsjTjwRW0ze/dqE9eWPyWm7Dd3erH2VOPRYQeEhsPodhhx
1BPeJdLCE/vPHGYCjKcUfRE//SGxYZ7vlRTWFuiL9uRhBwv4xLCC98z3iHmk0swtKAVnJIa1GkYT
WzuCyUkS/mPVlQL4T5CE+XLXE5l1fqjYQTd63qcy6Lf5RGJ1pwinF/Hr2aH1NXBVNeHUYvEBpwRy
/9k9HNXzBS9VL63c+AGc079eEq14WCiCs3os1qCKB8jnzJfo1XCZe7Zvj1q7PlOOmL7Zk5EMdyzS
as33dQksD+AbbcyS8vLf1l2C3OUk3VfSgizRRacwY5SiQ51lKRNzqi2gutbbFtmc8uejzjAxFW0N
FZX7VNDaf3LYHaTJwIAVWLt+7eycwA23wxeWV/gWrpNuKm8+er/Q3HhxwjHWF3HuK9YOPe3pg1S4
M6tblxXcCLI2ZDupOn9Q0fOiWiJ4PHI2rgKddu4Bpn/ufJtsYyyPh6bHLnEXHrvj35wxUMkKdCAX
Gvp/HQUguG7+g0DzFl2Ro40An/ucA3HaBG9n0N4Tgu8Z9VTKtEBvMV8+7+SsLGfRd62dyxdC8iTq
fMAnQ7+EF5Ss/r9KBttPJZ03GKQRhkvJONzlxx/aG0OHrvFvg+qp2vYgt46Fm1vC1C68zUru/jIu
KyeN7FDtIyqW+cCXQO4jKVItkpTjnvD2wFk1Ml+l1U7/EIoDxrA2NkXbXCc9Xwru8+tY3n/JJXPr
+bjiKQXH+DJ396/Rg+z1Z0vKzdgXxtb9oC0uc8qzRywdskCzx2xZ2pIe9+UbWGd6lWqKUbmB9BOb
cakZ81oIkiiCWmK4Y/kCLVzw6CVyjpIG0BcF2lVaucc5yYkxaE9jPQycjCFLXLk0XF9uWLq9GBBR
30rC3v+rer+yS/LTEw79FFqvamuKZG1aY4yrrOW48nP/BiDPxFkfj2BZICMRZymwqrx4MLWYaSd0
4+YmF/RPuGAi4CYtpxBzVgcoI7Zd1KlprS/yZU2TJBropN6vaL2sXCPC1z5THtLPXU4ecUjlkWhc
a+Vcdl+4rBZO7ZGo/NzaZggpzBrP5rURIE2CdKNC7P/ayTs8aaxO+MteCLAPk3gkhRTIXhUCuYiU
nndsY7rHn3qVI82kDIwC2Nm55HhTKLU3tESHMjWMxPHSHrTpQvBnBewxewdchPe4kLRnjH2GcYLe
iEn8kHPlyyZLvZZG9qG2Quud+SigNbENuWawIURrK9OVNw6hg0scBrMe6aRcP9sLT3TwHUoYZfr5
JiZd/iZBbr5gyOMR0SuZGWMoJRWJEHjrVa3nq33iswuFa6HwcIHlLwvXcc09Pzgj2IXrLKOmPeUp
5xvaovymvKj1o+wR/KK2UMlRdLRtfw0ogEV7aQFfGmL/Q3Gf/GK2fOQndelF1qok3Og7YQadmrdv
STH2JUOhJ8nb4bF+QcyNAKqquHJJELcZtmlCUdmq+IZDBEUESFS1K8PcXnpLm+Y1ATRogyQEMY2a
a/KPEij2YOuJbkNsI8N80mL1ipeqCMvpNm7UDOLcSvtIXKg+lNVeHTaIg7Qm1Vpb2YzVVJsS25D3
e+/f2kpYHByI4mL7+LPHL7TXKRb4lDzMlsvb5i9FVX+c1ddFOSgAfHYW60R6l8P1Ur6PaQmNdBlu
djjHBIXMsxkSvd8slggrBGRB9A2ry4AS3bCJboSvmK6jGSwKWcaH+hMD4cYqZnC4N/5tvKxQipUe
UhFay7GL3NXK4Ps1E0ujEFOQxzpOuY96yIkneKGw13A7BJIf2wQ2g9ih7AP7CRY3mYdN69ZefPtG
ZzryZyzhOsza060WjFuSryZb+DuCr8AzG+Qug/Jfi7ZTJWrSWVEGnPEZVFkW4J95EWyNqxHTCbHA
2cccUMghfHuKQ+7EQmGXvAGmbbuuywdS8BosN3qK4rlYNO65CRhydpUJOv3lkmjElnjDI2s5Vv9u
4QCDYOmZ8K5hsjH8Ek8m3U+TZj3c6m4E457dOf3rnfyZBOfDztHYCPpkyHFB5yPcNOKsfRHJHatS
2LxSZNW2Hklfuxv/+lwkVwHEbPwZNlS+nUx+s5oTB62ZMtWJJNiQINYYfPuSUV+7pYj8wrZraLzE
ekqtowVEcTHEfEWR88ULdzGXEqaT+jqkDFZw/A3xw5Q0tFOsbqL+TiMZhmwDVsNHQI6DqLurWQrN
zdp+LdvLjVeEImg/CIxacF8xoprQV3vNOcsMX0EPKa4J84LcHUZdT8dzbWTiHoi9fHWeoodlCk+V
oz81d/AvL1BSzhPUWE2EVx/BAOa/e3oNrEFgdfK9pmlYmi35BjJjipEiDZFO0sOIUi742yPYrq81
fTqlDU6ii2Nq3pFAWU25A/yt8xyowzeeI5XST97AGmvq3S24HIi/0a+T6HU377CgMwzlL1+DtaJM
SQbf0l0eTIvnj8+iol04jkZF8KTi6o+Db9/G3taa4Mo2LyCSn+btdFI2RYcjZRuXwMoxVz08GuXI
dYsi8G/9QhBL//0xntG5DVu+VFNAUh30qnsuW/25Iul4UkuPV+bnZi9OLXoShORyH+a0g1BzbBR1
oYFFZFCJVoYptjKi9yokxpD3pt0SEgBryVsANhWKjkUTnFnXZrjqlIEK59TpY8uROPovyR6PBYvw
6KvO39fjqvmkjTvdTsMmV1JZQVuGlDrKSC++3zuDusZaD9ouLoEZFCwbwMmmRhG7e1oKfcekvp4+
6zJbm/t6ohD+/6Kdel8fZWJXSropgsBdjc5JkReDRAHv5y8+tN5qGF2hiwfCPGrjedE2ehY9u2hf
UnXkrFs6bg9PhkM1i2PaxQfFcnTehtv8EUQtKIR8n2dl8rhp1zpaiGgmjQzfl47p0nRx3fl70qV1
XLL/uWUi+Fjbfz8tfP9vHj6uZizKQFs8Xmi+ku8ZC65dXW4WEMMzmcudvpf2ki5Q+C12hO5iBaYG
ybnpk+vrSbhPvsJ09RLPRhkREH7wNUd94jq8TsqTQiG/JoBRYNQLceJqvMhUVXuPIrR4SHUMOr3K
2hItm+2hy9FY+vL2gZXaFh1O5ObQ/b8weHNtG2SJHYHYztuHMltoEbq1sHx6I9BRvnXG3dt2oXB5
cPh0cfy4TBJAVryoGj5iaiFlF5Sf9k0mvdOSwFqzFSmH/1tcF74o1BoSjSNabH5h6zpWLYH7yaHS
1obxNNwhM+y0pRR/FWJnSrpMQa0tAdk9FXFHi7WGCAnZ8s1UG76XnHuL1tdx5Krhjl/Xynfaix+8
04gt8gLsJ0f1igrwM7zAv04TqWeqvmcAk/XFLTXmIa9WLrGEGItvjL1Id4qi8n9YEpYWNTxoj6md
WWm9Eb9ZA/d6CdTab/IJUy7iAJ6bdzw86GYtjunfdbxx55oh0wd3BZA06IjjJogMhcdLM+LJ5swl
n/BJbJvScqE4/4gVgVkWRMqyxf7F7byzeQYCICxODouqoj8euoibc4waNVDDYgQY7g4901QD6XZ1
sbe67g7E9YqGPkONlc9vXSxV+CSHz2U3IopbSYw955GMj2IUr+qxSHE3icHH+xKC+PHhn8I1qCwx
3bkAH8ZgTwYpv+rOO98NLrWWsFkorfcU8TstnUpQqaQ2TUejZTeNs9xp7TJ9mqam/eOpHZHe1T/A
27TA/ZiJx2OXy4K9CecDByWCLn0OPRnLSgA0wNBEaUpYSCL6KXGy6d4tZOF5ibW4WON5t+bCRRZf
hDjT/cnzQpBPh2G5KChSfdt85zQUaVdqnd1V8Jm8dP7pTVEW4km1Cpqi2eDUnr5HzU/+UgmT20yK
hySy5hUN6bfQ6arkwiUUWWzjrUy8Po6QDstU6nw/hbY8bqkXysXHvWC4XUYJ+3nFq+GdGyHIJEaU
ERDXCbZo50Q8OGjH5Kk379fNrOoNR+YGsHIHG8/F5p2TxGdhN67+RJv8dOb1v4RwiSIbItFe2inK
+5SF/Cm9W4smPuU3n9HqnVvlRy4nTn8Hk6Nr+7eKqz05Mn3qBSxhLSe3ZoQQpeCQMxS/ZKMzkdxA
+l5yw2lGxshUoVXLYQ7xvROhzv9D3NpmW9z6w07BrB9KzNrSuD8ERcKbS6YwGN5rCtxhZaAlIVJf
LPN5qZtC4KpxPp2Vr/4SmBTAcWkQnSolozHsQWd6hUnBWl68JLzF8FP1iEv8Nwi2nZmG27viaUYR
fnbqF/LL36/5XvTTKq5uZjTizxgTR4ZSjAan0+PsCPSHk+YOVxAYzN1cQ3QU+5Ba28o/FqiiXIUb
Bqib2TWY8t/VhBy7WLcY6/sUoCPvB1r+wnQL8OKvvONhHI8dik4k2CE4FXjMp3wvNazZboIwe5Au
NzXygUtzvfJkVSzI5QMXzWirOa8uLbi45jsjI3rZvYM5X9mMFC8EAc3HpVk1xIt/QFARtSHHGSIa
LMbgDQ9t/4kD5D4ehms9g+Kt9iRPwxsWkZjqat/5VuntU0OPRzTP/EX7HKQkJeqGLquNBoVIAgPr
A3jOL7m5SgPb8A/y5O05Ue6izEQ4+becX3KGGoswztokJG9AdnDh9lY5nVPLxNZ1AUYY8E/mmJgi
5mKpyVA2f40NqPaPPnymzE+Cp0lKSqtJL7sZJMlre/2hVD8j62HHnFUMW48tg7CMI3/1krO/kLVp
dNpIRcvUDWgwRE0WpSiYjzlwKYDW7tF2dFgcXcQdx1beBEgIiWJ0FSvetURLUP42/jCbU/Pzx0dT
RT+uvOLmo9IEgHldEz4DZ7cij+bmcpl3/TRSQbAByrUJ0HaFFzYmElSioDkQ9kqx9MUhfnJWyOiS
w9WzRQYHbPjor9pu4yje3gWPAchdqTSpRWiH5+LptCURxZ7n8o1/PvL7Cq2GP0fjMCn+bEfVz612
sSIPQXllTUb1HRHNeGLAM8w42enIqHQ24aZwnaYV5qt0QMLosvfSnRvwzY4veZYEvFlBGhZilAKY
ap5ZpGVeUSxEVs6kzv3PIVmt2SuThZ/6Fi7Iq3Kju0krKu/mkHrG2UbaLWxlXnsfai/smirYuOky
aY8hf4P++ts34TskWhTV+7rXxh+xUkpEPdx0RhVZGil6MSCCIUhgZh+a4Zzxk66up9GpMHIZXPwj
VP53yjXGpzwrjWeq+cYlDtNfCNYE/NTmdq+J9+7nCj6xO5mXIznhRagUZBntHiMyySE6wt60GaII
QB9lvMVbFm64SZ+3x4RLl4Xjv304AQ4rgn89VEX1OG99gCvZ734MIHauzDwQ/7Cohz+u8AG5kvF8
/ojq4MyvAbRWttD267c++mOlr9F5a/8XZDfgD7m/EiOsiBhP4EgjLZULBGzUabE+iwAklIJTTz+8
sSY90Ma3PXmMyNui0iHcTN0Y1EOy69wP/sM+wt8xgddAnxjlo4ZieNRO46LkXScJQCF8jN0FhxZ7
JFhalvIaVRuBv8h+vELN18fExjUMONLGJOaJ39KlTP/elx6pTYiKDEUH/wXgl5xf6kBuCCk9ffrs
hIjPfbKzXCq+Ixo5MEgWse6HufmUDmyP+J/MbeZiw+LZ1kJwdz0zVdOClba0/2MNaLSD2bfOoJRL
oK1fBroED4pOtsis6UEvSbQpvw3HB+POvjNew4aNVQWmiir20kBFE9ks+uQYZ0A8jh2WsXUZNV+d
bguZsyPWuZb+zWAMRq4CP9vzbFJ+MVG8WbFQmTb6A9yKFE0xAz0hVyJsgW5NArp4LlcFVZDEHEzw
64Jt2w5buRkunhzyDaw94sJHPOE3nanFj9cl8jQEPb5v/baJYeXvFlAUdqd6t2iIt2W9uC26NsFV
AB2sMWccNDfZZZ4JRy5w9wkVVgXX3H3J+LmQu3FiaRq3ucp3OEMlgn4LJxVGxTqp8203Wldd6Mjj
Lss4CAEQhzl2+oKRZK+Kqum5ZwJEEvoPMv70d6/7IS34AKLiIwVW6RQHvyB9uz2W+OlCos2DGDLU
aPcJDcni2Wa4qxbaWuY5y2E3Eo8Li9ed1xR/RCuOs8dUjhaoe808jgba7ZEXcyzz8TKY8R94M03Y
NIDSBFV8QJyJ6Ygt/F/MjPeh+dWtV0M7xsZNTN6B3exJKUyncY8klfwrxg0jHdzMDVCXBsl5s4ZB
vnCYPrNxnr9o5e6IunvBsVtNokWsvaRYpcMUcH8dh4gV7ilgzG5m7VSR0DeWsejkuHiYKdAWzhit
Hd8MMtEhuh7T/QS580N3kjMB891Pdndi4XtogDCEjcUdDdeGBXDgYpTQmvoN99WcHDKROUQYKESR
aIGJqRWdmW6oRBUQmo0n1YDCYXhCkfxxBKkRb9/irMHIyOlEpW+0N3AARzEG62NF/PUBfiyKf+bv
xDH1ZELP7v+c4/HWfuLz+TulXEt4AwLdMfplaq7xxiNJ3GnOhYwAAOvB8kOuFkL2Zxprvz5XUD3E
GpiDQUbew0ZQZ0nRggL2BzeY9CPbdZtlOcpANXeJjD2rz0FjE83sSB14s7pejjHDyZPxo/EOkvDK
3lJcD1GcmDAbVupALTZQd3hH9Z+qpqWNWPuXZVHu/z90MmDbLPkxzBlNxVg0bFcuFzViCYoibLhw
PRio4APUndA96QPrDh78pTHOoFV4qWMNX7l5nLhhmoWdAvwXs8FMZSweVKVyTNjX4nqnTQu3f/0S
72ezK/nmniYD+rj11R/tUUvWF5jJgijtOX2wTkaxhDFtTvehRgvRFd2k8MWkT65aM+S4M4jU+I25
KQr1vMw7wZ90EN0uT4okDV7Fv0mOZI1a8retDizZGA2NbHBOMVXasHW/42AcS8Gm7k+fSJcPz9H4
67xJ/ZxbWqBWg3OzJCkCa53A8v44xTd56v6TAM9uN7+d8oWW+7c5tMrV0NG4LalIkLd3TFrVPoJs
Ym/xQTAA6qM8u5WH+55HoL5pr+YiE+9MFR2V7gWX89uwd5s1p7OZFrRAHP1sb9pDgF0DwXs9P9Af
Vh0Z3Srt/IcxaUxGN56LmbaMLws+lc4WRmZ8bfqoGkguhDAQjP4paOAIyWOsKZkFTEyeDJ0urOto
3vInN5BLDkQow1W1J0Du10utpCwsktfJNKtlK94QUL6QvrqKZwqG17X4RZFEt961vh/OfLppHUlI
R+W74jG4FvR7+S7V6XZ9weKyP5wyDdSJ1wj+RxHNnF2WEiJOaGXRoYKidzjmnpbmKITaBJSt9YF9
qE9iphE1N3+rtXmpGNCvt47faZe7V1Wuam6PUe4ovcZCvL2bY6+si5hlQ2vhMxnq8kHcBZHJMycE
coIXDyyua07p2b6WN9R9j+9GMRYgGIYUASsR1ka8ZkrbvYbKSF0BeuFR/qQAxOT5t2ELr1pYTkvS
fnGxf7i744CDwZxbNxu4XPJsg8JXDqShr+6BraIIVlYlP6ZB63BLVIY0xk/9/JVVXZE2z8SgDJUa
9gsYkl9vLlLfk8jpo7F9uE2AaEfMsAkkv3cVdrm006cnV40KDhHPPsRmQDgBh24JP/sWwRf7zITW
jxQWMzN+mw4UGhHZCdkXQKDaJoIDjv7WVsLHIWZKOU3VtCrDTSvr9fKx6wo5VrJKYvogGFno0CjD
rCfC3vJH2W5txuyiyW9qI5othHajLAF0NnaODkiJ5GylOVyXLyrxbi7D2fOiOZIwDRfFvVsR+2oj
8tbIitmcE5EmK5808iR+0sec2q7InkTVSkBQTmyim/vNSHSnEZVQnmKKbvtnIUgUoc/+uJ9eXqMj
7mXA0wLb7Tyw/OlDPFGD88HcrlxtQLhpmyZccF+8nhZrWLj2UfyhvnpMcxMekf93PYsjamMi0/LH
UO1TzlgPwUIs2n8MQMwK9vS5efCYvkkQY40lYbwv/p+oEWqD38uthRhIOAuEJgrLquTU0YPrVaRr
hXTXRVi1t0Qx4gh9BgwCC7FqS52lR+XGcUzwHtIq8gEjca/NR5mnUa6iEz5NdMSwcsWGyWk4IxM1
HG3oOgklmGRjVZxagz1dR52qCuqjL1fBsNBV81mGmI2S/2BkaOknRVgXu+gh2XxPEml53rHS9VJW
XLxSBb/O1p2vQrr1xoakeQTuqT1UOTtq3yGyhMZdXLoLXDg+SIbONhP7aBNP3jqahdE/BqVoNp+V
ZgrPI4V882JPrWP7e4KE5xHGdV8CTf0t2wc7/N1RSQ2ydP+fuF+r3Ks8nCe+ExLAgvo7YSCVPtqJ
Tspslfm7wA+OzvF5GoQmd/qsM7nP/eN7EpL/Ov95xEVSOX44zvcXniDRlhFoLMdz2us8EFVu9i72
GKZxBLXrb7pVK9Ju7UONKLg29irA3QtJ8lz4xdKK76llzszEGM5e4hKHXxnKwA+872DEy5jK7kNB
/TTHlr+zjCvknywRSh/viVq7zVD/8svJ61UdxeEpcjiByNMHNbiRL/KtmRVTOzd3LTqLM9OkIpWM
/j6hZIGfOSwNrTOTX0UMmqlZndx8VIt1oewBnKd7Hk3eBFcQNny7hYncDy8otA98vWbZaQWQw8+p
M/XfkdIkgK1HIbO4m9O2TMY1ZJISFEZTwOpupT/JRQxNzDPq+u0eZD1lhotpFRHbajp5czwPR2qn
lacilnMjG56gS6tYe09BgHGhlU7lu80B38eWNlY0weXaGLkrIVRgRkp3cbiVW9gxhTU+FHaeacqX
5sbUHaZjccIh+AkCJZK602qj4A3+LVDh7BZc7csg2yjAu1tg6DhZWy/0GMyW2nwKKAuFP+19QfYd
ac84eedBj4teqvYT1rLifhADHH6I2/RnPT5KnIgvSDJcx0WiCqkNnpGcMKWCInS/GuFXlVt9tkxC
QscVT3BE/coMFph73FQn9Bf32CUVpFD1tEw1baAVR/2BcseEckLyYPeRu9pE+mjiWwFn9mS32aU9
FVa8p2YU9tIpWN3a0bSz237rbBwWn7jQ1od0Dra9OY4VCwTbveLxzz+u6ZgkOU90yjelFZ7Xo+Ih
BMqnQ4kArS3Zh4WGIgL6m0Ag5Xze6g0yO8fLzaNl5Ac3vFLoyYViexPv+Sqg2aF3QNSSyirJcXFq
f+kYWNd8nntiQiwqadpTxsF3Rc1hD9M4Qlj9MnRCWX6qjhHLsBdvZpUdhOdxEcUA8w11oE17mrqf
Calzy4OMU+l8pbpqzVxmse1czzHyNohhDbnkP99nZ3uj8QUNs9TKJJ3CUeaEv4IJEQISMoS3nFXG
GCDnvAr7JCBvMI9OHMPYT+KM2vPIPWytJWedKhn5fG1o3OfnyyxQd9bp10LTvhSy1rpOaeLj3dYg
Wqo+CIqo+kXBesKbyPX01Jt6djTdGXJUJ0EciD/nehQ06RZBiBYEUy1mHDPzh/Pi9LbPAzzS8LJl
CeYaA7ZPXnSeivHOwk1WPXnlnr42Wj+iCXyTOeVr91c5eDvhm2sFJG/2yhg9F47h0pzxoddLDc4S
o0M8548LTlfeptkeNywtU8naJveOkVk5pEfU6ge+1I/fasBrSsEy229SXAXjZc+7QHsBtyPY924p
03d6DAoaJ2ztfL/fiuskrn6vBL9UYfLQwyf6cLG+sIDsLOxN/jPmCM1iSB3wYudDTMhIC9dr8lXz
WOwExFINLGTed6LlXtGRTfTSdkM/Iw469Q1OE5PpaUPmPyDt23GgKvCJ08PZ77JebJdGp49RNrK0
aZzug/TLuhq75WmqAYMhsx7otrfH+W7OWxi6H5Mmutq0+JT+wIqvIUJOqh5hUbV/z0f+vhlBZF5q
OZh+3OcIHXl0mVEbV3g+686i0FZbBmAE4tJ2CIQ7sKeCwC733DQdhpIR0/mb6QyuWZjjXp0suNOU
90cx3XEPtR1emxm7CVoq5teuq7qbwqLIXI5NzA9+WDNLFeCNcHB/MqqWOHAHW7Xstuv6GJ912Nxo
yOfMVJVHppWTzDXILKX1t/WLV0nhCysQA0c+DbypMKxAettfax+XgSaTtrJknDL2oVhifsWOPmG0
/siVDymd5bOhlds8vJ05/5z58L7NIJHsZ2vymyPgjEdAqkoZZC1lO0jTtlBwAuCFSGyn6IHdJDuz
7WnBUEgtAXCEnpQc/bx7hIf0nu9cKcZEocbfKHxxwo394YIcnGUlVpbDlQAZlo/lVHHnCw8zhwMd
ucWEqQx32qugCaeT/oFUJeo2t6ZSBamr2WgDgqlrIKWcA3Izd2WgRBqTW+U8pJbNf2NCV03Et5VS
CM7JAc5gcjQxIifARG6Sq+6qpLJkGT6obQ/YKHrytLDU2eqDFErbBzTsEVD13N0fIXSNz1NkgI3F
loQbH+G+f6TdkqT+yw/CamsnmNYxPoSPKs5wyP/M2PDIi3O0eBuoMTTv8K50sEOeRdUu8QXFTQI9
UQhSisX6eDzby//yc8SAY6+6U2SPW6zIxNDMVJgWkoFsTSt+YhzyiCpgz3szbXRCSxzwFkE7FC/J
Ii14+MwT7eBUPc8hvHcK1C+mQZNZyeiHSssRIC1A5esvvc2DAw7QodW16NvliUE5wSad4rtz1CbV
I1glqQybsiNKyIR5WgjyYy9mjE8hd/qoPalm98dbouk2yjoiqe100Fh8UprfcgxJnasWsmGxhQKb
EZ7giySINUfHK9XXROHMsaZUoOGieIUKhsBGc/qlcsZCWLLcC/ofU7pR2StSBfu4leqClpZpdwBL
DCWxN7GEkQWB/y2QEGgPbuEKngqFFRSjAgZN1lbVoW3OYmbhZDHFIL4Ymq6QWnX6ub1CF+hLTqOf
jyxg4bp+wtA+m7I+H9TJctP+FjrnVJruDYQAnZCqllm+EeJibxpijzdNmMKnhGTqrmbsOtIrClNC
uXgq7zjYUYtXOsSNG7UDFgFIWqv3OcS17TaN0h3Ca8wS3flJTNWVmju1E/34qIb3ZjBd5QIkslfO
BUFbar4Yg5P6FODT3b113KS8XELwO+VzwmqpVE6EmWXAX1yGM941ID3PNyFZ6X1+u27TObut4/P5
8+ksf8JIhQ1HL00Via8KJFo/QLqUNlsDVJKzr8KZXu9DMEgnWdhdCA/NI8xSy9eZcW8ywHIDLNeh
knT7Jf3poAeIZoUTWTT7ctPRzA9FeeQXtAGfwtHnXBOqunXUfKagk4HB9slEN2hG/1Pyk/YN1BTS
IUuZma7wIKzqCAxC+7nGZqNCSpOJ/6SNTyYZXytKNHV6ZzB7MXG7wa4cRYG6gAXBxyLrmqJjbHLh
auTecp0D9MH/Q9XsSZRnAUUDZgpNfpPu+qpjbvklTICEKjUgeMOWxmj86hMqibcap25ZKtV7qjDP
KuRVlUr5s44Y7uhbX5P64RV6FHlr2ae8hWQCJ0I+1VsuSost8wu8s1+bTMZ9NYQxixEuau2O2Hil
OCSTU/Dc5aI+j4bIIh+M823g+5SvMNc+DKMCsHTnX7z5OxD7d6J1/L6wTtHzuL2FJrpjYvyk+tko
rVtm1IjGAMAU66fdyHE8I9+jJdLRT/lYUc7GESv867kSx9z/5YnC4vpFLTES47SIa/A8J7aD4nqe
mxtNJu3JqiBbpZryhcwgLE4p4qxEVIkM80TzmsVZj0lLs17xn2479ulRS8HLHbUmmpQx9euV3nFB
l7aI8bwaT2lgwW6OtfuBLTBrYANErf8Y9ewgZAOtt1HPcNqn0VX9752OqL8ILAiUTqqGK3PCO0Wo
bxvb1qXUzPMK4AqJ8sWPsAsrIwXFhT9Ud/FkYiMGjZLrjz0c96j0z8tARTLLfxddBJNu/k/3yaW8
EC3IbqMxwvB3BsXjkIup4Cdnfrvth8crtu/lTuykVb9aGw9rAvy5YugJU/x3IW/MP9xksxMoymg2
obhWHPifePL4Nq4ToQBYuFY79/irmHyaz/XwCZWpqHgooJU/McgJT8GP/+83bEmXTeG1DGuCDWx+
5XKmDApUWTWZmJbd4WfxmO03hS3VWHjngfSxd1dNJw1XCye+gR5KhiaSeBXtaP5zN5a/KUrgi/JR
Xg5ko7LVSCCu9x/+qHVxqUtuFhOPVYFToArloPjSTHbxdcvk/TNEE/VpuHg2OUenDjytAyhzM1ju
2Qhy+LGvV19hHbPVsczJXBSR8haFkXgvrRYxi/OT9OUvaiwQ5F7/qZfH0FdyuS6yWDYrbZ/nAEqq
BtxW3x8uK+4HXZBNxgQ2CvcrcX/4vg8zDgRiOGmizySaGNCopnTzdYeDy+BsAHlAmtq+wVXvbXBt
bl/w5zpkE+oM2vBAmgSxBFRqY5M1LQWmp1i3lDinzzVoXzxZGz1/c2OHbAYVxcuxeF65+XYDUGtN
uuEeCqsUs54o66f2tSb9qF5fnTp2Z3QQof00hjbV9OGibPte3RRYHfYTEldZYV4E3Lb4fyMaxkP9
jBrU3tIkOcVnYVa6+isoaoUye7HspqFIIQpm6ivv6ctxPHHnmousNnOOAqUisT93nUEzLcdaVdrV
FbH+Jbse1LG7l5+koPs+bWVKQswkFqJXU3UuuVKUc+4GwZ2igeGRNe8iYGfS4skVyuMqQsA8pKWt
mo66KzEtZZnoSXs6aP4cwkWU+QTnC7JHHjWi8o9y52c4mygZIwWoba8bSKMkR/ITqCqG6csE75wO
cpMQkJOQfJE1W573ciFSOarfg8/9d6AIR0/c0j0fNn6V2wfCvOfSZSYqvgmr6/L2l3AANgSopFq0
6JkREtk+u2z3kBhyex0gzVhwLbr/zZAKEXnorfyTWC1e9GQh+YjV/kg48WBkCUA76QzyfeH8uqad
0ZRNTP3h4OC+i1kyduhPquKMmFU9wBolaeFAzorSPqsk3v717zQJf3AVZRtejOXiJ7pv6zmWtubf
0kPDEpgotitRsjLZaKrpHzgkPf7N5QEGLRRq7pZWrSpL9Qj8vDSOvc2CxC72JyXAcJG/wWo4fbL3
noQevEgptHX7AyncgTsM5tJXZ1T4jf0AINvLpTDUhLWXNl8Y8cm0Hoa/QYML4FNPuVhIwtWcK89K
zOh3MZEbBI9sx8q43mjaQ6xtuJAq7VdHGx86ZtpRE9VQktkn/qBJMw6obiKFouE//9kZY7rl+Khx
v3WDSXeneqAkXRUOahaDN0WDAN17UiFDeA+q7maRrOJukfCqTQ90Tne/Bj3SQTJAwN0JGz6VHKHj
e7x9tDMhaaZYUsBEeLSfeJgJ8x55ylRJE8jnhY2fU0TejIYeYM8IjKEqYFqK5B1CIUlRAP+1NDKx
u0lPDNX0YOpbMySAbSva46+MOrLhkdagRd0qf9tisR/YvB5OCjCITQTbymcsB89czgYe4H7JNvdx
xRv/7barV5orCsuKzhdDa0Kvq9dYQbq4MusmZPi+RxD+299/1RA0lQ0HaQ/eipJ6gkebgmQC5V2M
1D8PoeUnxy6xaU2nQY43ZNmvT4S91yoDKZ0DaiBPnr2iC2o2cJTKSduM06TKRGz9U5Oo1kj2giGS
jA5L4wWuLdtAHJ1JRkpQOsOm5BbYcVBIJOsaAopgdNKHEBBYOFVBS2sImHV047FXsC+EbkzSMEG7
p7htpVfdUtGaoKBTt9M0Ke8/4+qGoGQrHc61jMPP02o7ufOLyD06NZgaQYjJTs/Lei7KFGvLLrPQ
WEpAfS6nrgFyxQVMzwh3FLKtw2M5oDWTZcy4h3MmAjoY8aknEdE3s7KrfIwqufLShcVYUqHiCuUV
1NasCtPu5zekfKSP7pFNQYssmHpnqH05xi6CoCqZD+W3ELwGx0+BIHfxnDBpjn/+E9SCNi9spaAN
81zIPo4/+1xdYqVRkS02HApVlMxFeuYOFM8z8cqbIYNyaZklkgiqVDZP7ljSWzkI1HiefW9mg/jx
248aWvAYm4v6u9LUjAYhZ655WLD0w233oYalrCZ3wbmgdggrO/QTwPyaCX5g+Xu0AFZfsttxTN/1
O94JisLQiRHb7un2U1aLg7EGqfHS9ANGZG8/6yMOiVxcUiW3Ia2QCEVeSN8Q76iiqGiSjrJXNjE1
qzmbjTxOh8uf+D47V5s82Ptipcy2uNRd8i1C6uRl0xjjhM+YTCrC61UTXyto65uQJ/dxBGE7jxOk
4Dpa35+NLoUqexX2ULP9a/WTUcgUt2kq5ULeFWH6D6HNl8Afl018nQ+tasUGVJ91gO+nNWjh8nMM
3KVwSEqakcc4rkHMjY60BujhBtRxI403jo2MvJv+mI9qc6jYsaogIIxj339K+KoDAH9V+K0R9hR1
zA6TLjMEK1KVf+9HFdZSndPQL37JMf8LxZfb3funFCOf1kNUVZ6vUUGxLS5yRSP405rR1pCta8RN
STWBLvu6Cck87mZm4qPBbA9RQF2VRgVu5c1Dn6KyXzF7G51VxE2kZKVD3BroofpeYpA3bQu0ChXK
FF6eJ1QJH9NqFoNf+n1QrRWTSo67dAQHMSGHP49tnQxFF6VlGKNDp8IiX9n4FVZbRC8zffOOTDhV
t/R0IlVKDFWMz0xiTqsa4f+km4tccMhfm0I4OeBsHTrer/m/Brp/hSPzkqvdlel9HAZCq9nmmkK/
7azxXydaFUd5RiIzInvcKKjjB9ZDPtcapt3ODYs14Neln8IMYnWrqJu5Yt2eIpXfi0T9hMDkENu1
grnMg8KvW/EIzLshFQkNwKQvC5xbXGcgOmxmGFbqUgTmbGZZ7Cs+Rt9AbNHqaTVCKn9DLF6UL4xs
qpTfJhIphhbpQgGaJpuO73ebozRNuRla7UJViC9NeILVWf3lufkZJ7/ObCdlhLltTU1VXYIMQSRf
6F7VwzmT1byXaQhAwEAf2aUc15EI47xjUuclauPmKlsc+FELMvguoibhZjOcmTOhaIFWzo6UoTLc
Tt2bQUE/ku8yyUqbE44TV+A+TwQmJKv2bJQP7eghNb2quzJ5uBwPIp1m22lgnBXKmRR+GNrLNjnb
JcWAvh5ZmmwjufZDNCcqmYdlUGmN8JQTz1xhAD0owPHjPEK9b7HxKn7n1P+AWqEWAmmOJZwW2qi+
x6O7QCRpcfkI2hLEWEErlDlYRMCEihLWODohuB1+rsmWhM8P9BFeXhGw/BRYn8zyukpI1fQGvRW6
7w4j1OfEPOeKBGNqa8G+YjGUVKZ5+6LKWtuuarNYFbCu98sXugSdtIZLIwFX1R/Cf9l/wMqHjnm3
P87DwGvWMkaJUrOqzakQkYn1HXXJtD1qOFLLOBhp3Xz1SA+lrvV812g1hT9JHr7DqdXR9kJN1FJV
ceSbPRaS7vLloNhfmpTW/ArlwsIgaUNU69Y2pfJZ7UUWvKJKSGHYSlOgi9+rVZMLYDsQ8HqzRx38
4B+WQYk/fFNYcxrZqpftCWn9zIbNZXyUqiCFAQRJylO6u2hT57iGlERaKLknoZVMQcWET0i0I40r
PZ3i0EmgU/yRX6GN5qtkp565H9OapWk5wPVDtK+Fu/KFTLh4G5BdHi6rIHk3l4nXnRsC9nrCd8/K
es0MLZggpeUJ2riF7qJQvF26KAYcFMnmyFT4tJXiCUFNPHqjguAzILtpJF9VKyACobbRDPBT1+hO
1210xFynqjlWsFB4N5j3XOtl6ihXnmOdyU1L++hOoRrAe7FJHOpP27W2Px6hbR7i4Tw4QxApExEV
crobh+fYeZUGIVAMUBLnS5dBGxAB4HlF1D2zkvCk+Aw6hCkG7WOdWudoIrhEyzLvApNTP8HKwWMd
m9vYulZaorXXVjl/EjdHnAeGfdxg02dboBAdHMc7KUHkCQJDGKFKcPOFG2mNCpfMm0tjqLZs6BzC
Yvy+Z+lgh6rSHnp5pjgmJJSkA7yW6yImx5uMhuO0ptHZhNBj8q2yH6FKFTW44pDs6KK+O17ag2vG
hxGFbqKXLX1ASRoFdWJ/tKH+mbNLkwtlrMEk9EaBJQ770MveHuXNMVWmTi+KLlzLoyq973UGHoHk
Pv1GXF6vzHpgQ7bK72VaV7PuZxnw12g65BL0xSvYJl5KSNn9uivNvvfdSqinc5Z15KvUHTkW8v25
i6BPP+E0hRPcehnU316elhoWUPoMwEZKguVcXhCXW4b95SS1MMZxhNyde4dLCrmWo/mRSHfLuJ8h
uiygo9yxY4bmEwKqiMFUslxo0D6I3Ta6xTaIQrkpNIhpwsiyYS214nqZl3VSXN4mP9+C3BTnR9Gx
Qm4aMd4E3SYx/pHjDv6EpCV9kDbuPZqYJarGL06eIt8dpmap07UbHYI+u9s7YowJkf+fin+SYnDN
KeFanl3nhRROteag89oKFGjIuWaab3WPXYKqxE0mbIj24htZKD2NqLpah7WlROYo+0s/kpYisDMM
0Y+wBybY8Yg/JGX0uzaA95hMYfwUok5WPG8rnUCMI6PUqASvOwgNhSVNLpn5K4sahBrA6rVlgAv1
JvGaOiN7SuABVXVadYJZYlax3jpfxEElPKgFmu/GGJe5oTqhTnZGUbW9wwkidNjhOZQrt5AQETM2
nl+IPntu/PIAlHH+UL5/Ylhk0uDQAlynfBHrM9nmrKpEEia4BTwD+3p8sbnxXIoaGpDW5H3uRzLi
fkJDdFlN1Cr5gHLCnklTGyZigNGYCYXpwZSFLN6oFlr+FqEnh6mQEcfZ9Dn2btWqTEP/jUt8MYnZ
UKCJAzjh2r+c3AnB8bcqOJTLnxFrQ6xkMt8D86a3jB/JNXNX0bggNVh8eo4Hgh/pPJLKInytBVv+
pO0SkoGxNh3Z6fDBPDrzpGQ1nuSYgWtcD21j5fCD9RFH0yiqJwzYukwSYpdbw0lmiIsiXmrYV2QQ
K85Dh4FKB8LKGgyDXywxyFi35JlQp22So/gFgDAhsseMrqDfvdp5iwRROIKxncwLAlqLPuX6ON/q
bXkXt7s2a4NhUJPUq5nenWKkyfOHBUww2MEpId4jxzGNUzzLAC97xRHYyY/EB5xlPojXyI4q6UcI
1tuxn9xxIWndt8G6UWtvDg8NM1fK3I1ltRnSKfAW0UImKRtMd5ROg1I49IuF/a+U2MVPFKurFfV5
bULbixFTgt3wMUJ1pCNuKZaxMd5Q0DcsIk2208zWKXTqcUjDIJMIxfNBUv7OdUvifxUY/JEG0HAo
B3mUlCYV7e+lTV/5SvL7pPC/QMqc9eZo/hZiVPKcUFMI+kjjys8Gc3j0JQwdjdwa32+lZA6Ne52J
UGTtIq7Ci1H10QDSe9/CszZB+5OPTG5QHDT/wbOvM5IfUuT4Sg6gygG8khPj8YMnB6pilcFYxnnl
NxA8hAdVVaYANTRqCZQreifHBqVvkBox2Z3xyIJE3v+U0yFbV7y/d+2RoVvzANrC2+TlTvddb8eU
2P9HIdt9UazCsRdas7ARqRmYMBpP0t3XVmNLEet1MKQiQtsgjreLCtv3485kiDBV2RxTrsVhxE6S
vOKreec8QjU+UZhgI0JubeyDSKQ3nXQMFvgtxB18fJd1E+YjNHLsy+z+RZI+Uoa4ZbPbozFWF+HX
4GNun5AadTkudQCV44znhHchaXxT8roJtLf3JEMcYAJMbSh00vV+sTQHiooxJyO6jFyEOS3u8/AW
1WmMR8AVmYbbzamgQTpT8HgCmvK42ezxLAaqx8da22TGIHfwd4OerVVZ164fdr2xO0urEB9R2dWz
hwh5Tq9e00euUgObFIk8U4EfWatvNyGbWd3y1W5/fhZUSSOcWMF/da92iUd3df2BnGSCN8YYTIIE
G40aC5tlF4L3SIyvp01Q+fTxLLqAHqQ8Hx8zAzy0hCw+qOSsboqZXsLMEtavyWPN8F10pMoElHrL
lCG3lFCXbV/Q3wUVeEpB05vcOBI594Q5SUBV0UlaFyTmz6HBpdAUWNEnZpIqUQKlLoIEInyMCItK
NtT7h0OjV5RU/NdVBACEd0Js6TBCSnZZWjmKtCfquRDd7dC03zyhxuuG8WnFHqQMSZG3Gs9DAFq2
l7Hna73eONaC523ivvPmMSFpw30LVcOqoREf+SzEMXlTuv2PiB9EtHJE3QtuCKVKcPjgTcSwE6Oo
+oNZ8E+rnvY+CbwfifQHdVuPOFDMvKB4mp/0Vq9OBPIY5iejzCzXLlRhEwrzGUZdNbaJX9+BWrAr
+G72CtaPHIiUemu0sJ60CXpg+Ha+BPFHPP42OWv4STD3uSPzmUTXmFjayhSX28vjQj1LbQqzkwdp
8bxnwhSbOC9iDQWTWVHWyiHrdnSzroLQs4rT5MTN3XooGNt+/rndKlwPbpqJxYkvwrxiigrP6r+0
r3FgpCOpSyMlrIOuwkDUc3BMjfgHJVNBZm7er8ikj4/HHZo7FXy5diKCGZGZjFUe+QN3v/o54kN1
oMKVHaU0bu2ormnvZvi2ZLUDTap8Bt1n9B8XQLpNG8UKboU51fjtecZhErQR7uL3kiIKejtxsTxb
uNL4afnjkpZSk0nGOErmlgKgQfUBWXPlFMISl/t9g/aWKy4KMRyDtJJM4rIOMa0Docgv2eWPFjIP
5SVsmg+OYqpt94Gpil/3rIfYRS6riypg0xV8DJSS4DimJEd9j94/7ZCxmwrUEcWp6IFfA5VroFz2
5PWeMfjCNo7jBr+igr1yTQ58/ywSppEQ086TdNvoSzh1cNsOlPLRAjfCo0vMV/A1c7KZqUkpDe1j
Q9wABE+6yFUgvwYFJOQ7sJwvdCEgwnce9lsVqR/e2k6raCyvrZXueNIH2SiDR3Pf7UvWMsCznw6v
bdwvKSM3OfvfIPy6PgAWwoaGnhMs+TbohKKg+hEdUBnMCh08LAa6SiO9iFJNpEYpgj3LazqIrKoF
bXnAtLD8XyrYESA9uTyL2hnJ+VpPZIs87u5XB3i4uH4AtDSRuiT7Bic3RQjoJ2WrR8C1BMmvZIHV
as7W+b6jBn8vPO39UfNreZzPEIWD9usr2BdSEo4Y0gckejdnveB07NoPfzOvoL/D5LOmktBzQXeK
j2pqz5z0EYN4NMGFHNAhVeBaCB4Sioaj78GGUDiTcgDnMn5U6lGe4U3kwblv3TVu1ITXjcyTnLwW
xhKh1XdBrg5AdVaQMlNs7JeUUFsZLUVRrqtCZ/XtkEViRolyI2laX6xULgXmz5Ff8W39LMvDV4xq
hXsfqRPTYEvm9roJA+eKCvo260Iz7uTb0ea5OVufzsUISqqx/ZwfLPzCh0meEd36S9bixx9HKHcH
FGBChEqHtH81eZ3oEwe46Y3Hd3CDB2NcFPKISznFAmf7yWGKKjvP1eRQATI0V9HAOjcUeKtX2Mfv
KkNtX0jGZXeADTieAhgP5aHYGOvPUXalIkYyi55KpxbkE27I09DDM5FqV3hK+QC/rmjC6kzqls4P
CQ/y+ri5XX+FGCWPy2tBJJjgBHtBWFcdTv+pJCOVZ4gI5g4loqi/DOnsbMiOB52U7/mqJc/ZTcYX
YWImFFOv31JVeOvdL0uG8svXA7XwhyBKqTQo/3JesgKvBDbu2dE+KgIXgMKl/I5xnsdG+ciLYmHT
L7l7NYtUuww13meKfwJyiaiABagbwOPZmqwjAiZgArTSU3vJOgUtxtdsLynXatqA+FQzW+3vYxfi
5fV2nGxrHSkQhh8GEJnD8akW8xGsZi5jVnqLswSmiIX3MLe76vOK2lRrkP1Lp2U96cysT4Rjeuaz
cormJGeJdCkyPv2rR2faLdux9vhojPPTmJbJdwBIWTEcdDLOJEiuKDATVbqqoEi90eNLk8V9D4ju
GQWM3UI7r+bGzsubFyOJb6evWod+hnG4RcX+xWORiqS1neE7WRN9hQLo7Na2hUWqvniGMgm0yGoM
zt1R0+Neg1ZRtvS04CiOIAUYc5v5xAy5g0n5a4AcpjHs5c7eISD+zUDEUyBJjLXE+wiFfHv46exz
FMonRlL5qrWGPntD6XBHo00IcC87ipf9ss2ShoiAScAIauViJscz8igqiLR3lFuAUpYsP5mAXH4C
BJTkzWHAdS0dWvN0SvcKVQ+r7EaXZWN5oSBiXQuQQiEz8NR9L9v9qLoCegft8VSeigGQjYyA7eUy
Q4Gts++IKu8o8DM/w5kKf78gprgcBKpkOOTMSvY4WMGk47LHr/1OmKUPH0kgsQ/An2PcEe2QyMe1
N5HQVMxxWrI5+22isOv3evGT9MMRQZqe756CFJd/IYvkH2JlWon9+Ezk9s3SD2DeP4jA4Ur7P/ub
zmbzvfkLmzVt2oVwUaZwGxWJlm9NrckO8CgdZnJnb4FFPQGDN9acgj9zwUIa8Dbawjfw7r3FpHfE
klAX6BKncMS2KAP8jgfNeXlXoeX090Smxgy6UBOo1Hc/yXWB7De3v2M1yO57lA++mnvqmufsqldn
zFGTCc4JdX79b5gZLW8oaCxLYS1AgPpKJJGIVVuGuYE6JC7Vp4XSMnyGe76GZ/8RSDwNL6P5EiBd
USEr+ZZt1Skm+LGihs+eICFbHF3sGPxwjtivJrSTfgwc0KiJvK5jBd9XUZgJbcElmRYjF4O9VKS7
DqyJ04yYj0h8lQnQbXCwk1t371QoIDf+1oL04ZV7yolKoGWLNmC/AVMCyKukt/3KWzTTo/FrmJzb
+IzFLimbue/WoWt444geN2lq7OV9jySu8fYF5T3QY0DYeuBZxB9L0y/6sQXKckJEfzoBRxBtePxv
MslWgAAAnFe7GtcCys2l4kf2ZiJ3/aruspzJ2LxfK8pBuw6lCNdTZPqFcFngNh33OnOc1BOFKaSR
mSjxFeY3N9Us3CnZxw5UPBaGc1Qasy+wFnZUWm5gSUIfGLc3wMHZDGW1q+OsRP89AbtglcHKvWp4
90YNs3dDF5w1DSPpz8XtyqGVAAhRwk4eQBrBgJci0C2HbgaRt7RXi9GO1K1Ad/BInKEmTJsgqpmI
y4RnC0Oi4LprQlwfKBaMEq7i65Ao9wEAaZ+UlnJF1xk7+tG6QJ1tIBKUJi9Z3od+1bQ0uwJw5DM0
fea+xcFUg9lqiMUttDxNOopZO/bJYsh5F5iRVdxMD7EGGGEmejAQhd7k0U8sMrreNf1KYSkIO8LV
qWbS3GlhP1CKh/cv+drJX/TifEyhpUYAGqjTV2hXC2KrzOD0GuawsJxbAFoSf4rO+F86m6RfTMhl
Y9cWuOEnAfuqCx7zZZ5eshRsU0HXQqIcbXLSHJGETWM6e3ByyrAxc0wOce3aQ8AA7TixpQOqenbI
uTrYmxq9YLPl/XUa//KA9Yt3vfyuCTJEuOlSWsq3J9UvcPBbhjTFIznHKQhHHCXuMu9vABWyIyoa
to84M2apZQN7E8N9RVAwFwWy4rqPYPbE31SBWi6761HbT8RP4LVFORjasRdlnRFkEAPFGVc6iWof
LOYo25t+H6aK6Ovqv034Mr/52W2XQJ0wIuMqxsfy4oo0T/SpSymfdqGEB9zi2u4ZBO6V8EwOslZm
2AT7v1oA/t+ilq1SZWHpbF66iU85DL93HhHYR1DtdAOqpLd3VMGincpiP2JddxdTLhuNQdotqgmC
Z+pBj/9IL10p78b8J51v1b+JBfREmqG51BqT/zpSal61YWafWLjN6sYoTHJPh7vZx4Q0LWWgHhvc
py3F2tYFKz/PvFWc+w32BTILxOYz/ryA1hBEZJVvDumEdQr7kLTxZPM0oNT0iGi3AODY/r66e8d1
bV5ZIumu8aKjn7Lv6KiWw+kQZ+e8J+vrDmS9vI0UXzm1j+VNXTEt4AvIQXUH16Q3W1Sab1CvUvs8
ji9S1fCLbz++p0RdxrdGxWBdaAM/n2zAQ5ut1aM2p79oaIdcrCnnIS0lcgR8CVOZkoBJT3f5jxtF
H6jw4FQ8IJsHYSguWOWooHEbAQ1UyNiToohy+PJPOGpR0kofY13EJ1hOC+9H9B64YXMlfswbsGsi
PHbPbJgazvaAzFjgAP3rNv9mDsqJyF/t9dZKbRmce+F3wNJDu0jypjZdz+UKnuHnLEoLfRPm7o27
zDlTXs9mFUJD/8TV6obbwOBwTMWkcTmIyPWorH7FGXfrkXCjOcploFvWhBHVNGkC9dEPrWEahRhX
iMKOgQe8/AWOhPu0v2Gkj/6aU3AzRVfi3/7Qqu2ncwjXtkq3Tg18nn4tEdTkIQ3vJEUWBDvaWoYU
tvHEen1rtLRD4X5rcj4D3Z4D0RowUSOEN4Ot/ccEJekCjvd6L/fT/I3bAUWlZm01qfxmMrsgLdX+
ZFX+KmxcmPeBw+LgHfRomNzVJUtaF15d1WyQVjUCVkZ4ayUHL0dqX/FpoDx0m4IbSro2bkIZ6Fap
MLgRj1kown28b0QlEatprCkfM+AwSmxkLSLUDnQT8JcArODNtfEW2ocAG09HWWdDTe+nVeFldHJY
Ug6VnRMJjokxE4x3p6Wc37aW8tEKnRcET9TdoHo4E8m0aQ+lI20aMjvG7nWA1mk7NxGw1bD1qVPM
S8MWxmibYRMqP3cYRhIvKeOzO5xtRhKWZyQ3oBm6Ym14YOhquJDOlLU9OooChKlxI0VodvJF9jIA
Gimo1RC4l8BkQjt1bOhsvbGdGO1TZpNSF5Y6FnpTufxPPE+ZO29o6bjAhv9GAlvy40PnCI0H+11q
bgS1ZNlYqYstEgnu/4o1yfrYumauLQCU87uu+/SbkwZX33e9IHWLkDOGyB4rR9YsuAr9FkgjZ3P/
MtrLtGlPOWcY8hw1o4GJ0qHCVuBO2I3zvghcZZ2kUj6CKLLkLEb1zE1pd6OyBSbmPyLWu7jN6egu
9VIGDFt0Z2kZtl+EjEQDF51ehbOta5UMLpsB+sC4ebWvHVLmHO2eCvDK2o8iSrvpBTvCW9KoKkPb
Xg/yjoeZCksR0YswZoVgz4kY4zbhnPTTpCGAZFh6suIlVWqj4rB2+L/Dh1p9Z6rECi8CVj414QBT
auzab16N0PvHrHSRCcg1oHjUUPFhsTHfzF5TxbVHKsYWn4yAD2q4K0DOC2uiRqJ+pRmEzH4S4gfl
ZJu5UbHVhabILB+WgmjmESWgdl875FP9cefUe+1+wWfVOsyN0tgjrAov00Q28pNKttGY3NUfRYGc
DuTZRHBGK8Ur7MnosiQ7Sd5HSJjBtTbKXHU/sr6eFmjqvEIAkkqZJuvD/FfvBHv1IMXCeZm4raaC
JCi7mWZeTi2cL4cAiTx+lXxHK32MMNdHOOvqms/q9V78fCzQxQzcK3mk1UJV827KcwSVbDKh3F5s
NmEF+abU9fCnjKpGlwvqNJ9PBpLR26v88LKtYb+gGmxwvEz3m+B7w0L4C1AborfR7VVjH7+BdXa6
s64q3WF/o/j1WMFJET2J02bzNxYkdRb4QggsHtB4MpBGlNzZMCSiPiAHIHwWQk/TxP7OK+WOqxTw
jnUOkdZaG6C/6FvB9c+U80l2CsimkFlCDMri46vlDyRMeNqGKmusD5oQMdLxgO4d09LIECfL8nUr
WXXhDcQDQXnZpDhR0E5kCFe+MLYH5/wlYZ3g9uLNPHr7eDZnhdC8bcYhFEDMXc0uMsXFOFqXlFWI
GqQ4bELy98D5Zgm8A0I0Y9mQkzc1AMO6g2queMltdTcf/FYiuH5iLpSgWIsGGCDAHcfPLiT1mrWK
n5pfZD9eomhIf9Qu1B3DAqgS0nXRWJZEbk3HWDurje7VocVjtdaj0gOh0HLTTOy/PoIcHMhXdqdV
/JRPWR3zAL57wlxVArnIk+IKtvJSCcHQRd4EJnLEOY5KAdUbMDBKHT0UiXMg1yibq1UKIDplwQ8J
0LLnc2VowsIFy6t73T8+KGKL2wS2grqhhByUhBgplA7emsFQcqKQ3hPvnj/HbVQXBfJNyDkd0hA8
RsgRk9XlUcogJLH1rMpLY8/IBANdT38OM2bfutv7OtV0RE69SxJd92RDTSs2uU74e3yEhpK+5NzW
BsVQDP3U7feQcIzEStaNj8Ng/MY9dA68HSfoBx15eqc44zgEv68EkP10Y8VUTPxlE6oXX1TihxT4
DTXfiXoZcEBngj+ExRd2pC1RoSFge5JWvhxWuh/uSgZH0yenA8zCldHX7CJM/3WxcMx4URJIrKNC
Z4LRcN1rJ0RNpAQTqVLuV8ZyNbYi3TCk5mlIFfmOeNzppekuXh5/iLewPoKA/2TjbHkcDFN6COzt
uyFItCNfOZ1Dxwg8cBFYedPgnTFQaCvVtaO1AM/ljNz0xjDzT/B6UI5+PrIJQAy61f0c38pONf/m
JewX8rfo8ZymmeJV2oo0Db7mPEPGSOMp5dlfm/F8ZztSRocwuvGmCMiSDsHUyK2+UFhaqAuMPq2/
UnSLPBLu7ZeZ2u+2QhED+Xv6p6QdYfSwKoZho7i8qVuSjMAvyw2JK3XvZQCnHvaN+hyzM/ftKOA2
VVVBgQmPiNL0uswpKZa2xjCkLgWmxLSk/WSN0zZmA9TQpYFTEtn3yVanXVDNLX2HShfU+hYQyXSE
CDtHIrmPGZp/c7cnIZ/aj6/47S0KxUotaylZ470ErxAahwmE+0Lvz2ddOO3rsEpWZwEM2aUCXOSo
OB0LHeWlvzHhTApRR0XvAaXDdNIky5jdjscESiSoI6d7c/06UzXQLCY0EyqkSYXMoXpjdEWfWcw1
yms/+ullLa4T6GikmjdJYXlSH4Z4ZnG/xh3i64GWxXxZUOHHAH/gkWWaHy+FnrgLBVp5qVvlmrNB
3TXOmW3nuX8SaqUPU75wfBzDqocPgtn8IwjcI+mNk1R5K2rWhgWBoYSIYfXHHq4TvsvlDP1J4/SH
9n+GEkuFBeaKf/0nxh69pX3oXlnGptwS7TCVSdCzb7bZZ/1h9DWJKTH4RNIHjVpQZftJxwnScynb
82CujktXt3kMNY1/uP+rNqg/tpeGcWN10m6EOusVbfG2GSByK/6xLwY8Un5trVxus8QG+RHmnCBZ
UAmUGTMXslysd6ONkMlHU5LXYA8t+qGdDplNuU1ZBae2dspg6HhF8+iRE2WFcNYAoMDGhMp5fXiY
lUbenSSeW3Wy+XIBy4+L/ijO9XcWUhzjrUTw3zKoYwX/6VB0B6T8w0pPza5vCwKceVfuqI7qLdnZ
WzxT48oH5mPHPGP8FIEYdOfF5O1IMuKNNi4bmewc31MUxRYQTZMaIEyVFkfxW0oBMvjbEgcAE0lH
Nepas7u85Smx1TcYXZD9MAXDEYg8In8nCJd3c2zQfDqq1ivhCBPSSITpv1gZsWXnLjWIpj/Wif9o
EM5bz8xYqE3bp7V7W8mINkgYCS11Fz8yf/j8IT2Eoh8hKKWOPZbUyVm4rkz5Zs7l3Igoq648Z/mM
hVtTpQ4b/pjZIf8qpzy1JtqySwJnrCip0/4F/yz8oXOemzQe2iSB98RV+tIUcYNXFoTJ9MEKmCd1
w0jn9T+eEM84s+W0aQfmt3Qf9lQmfkExtpfDdBbU7QoJfAf1LbX/xEaDEt9BlRWxqkZt91TGcbGv
DtHwC2OoVf8VE2/3M8F2WmonQp0nHOYAHz8/uIsy8bB6YHYoRjPuj/O47JRET2IFEBB74XUVGbpK
1CYzeg3skM11RCfN58amLy4dYIH8lbGRMDoZFTY06rruy8sGeSlNQ4xvIWTNBkS34ccK5K+nb022
JYk53KzJ+M+M3lmhLo2ZX0KOY2uMHm8ndHmYmhbVOZIFyH67tdYxWxxv97QbG7iSJfZC/xbF9tZr
II+d0e4IkeC+we9I4SLiJ17Ra1I1rfLwnDTIXKklSyvBlOPlrOVIQHwYezh9pAM4DqFB31qz3I44
tbQawb/dETY6Bvx75glfjKoGN2aCKmAZK+ODRVeizwNWvyqGjjKIaVSPnn2+WYzCpD8FykQ2EsSZ
3fnABI7xPfsNrFhfFZiF7hKCSOR2TMYUvzYVyEkGTXmlpxom18Q5EnXOY455wJc7ijXnCPCPYL9A
jYm+pTWtfkSicRt1fnCSlA4DTBzt2y6wPy4qe1QggXLQ2rtd970fwcYyI3+OWD7YEIzWVmSDS3ah
jW0lR0edh9IMEE1WXhPzvXcotV3OTpgKYahiWtCADFxmFxBIiNNEYEguwk/kksFbpmuSPgUF9B3d
XcWSua93AJ/ViDtFF2rCQ76ye77QNbKLdxsKZi6+eldDkHqkjmSsimw6sRM8iR+CjcWPP2o5Uddf
xPB2Wvoty8rVfPpGupNi0URBUI27Ss+y7DrmPBAv+TRo7KRg2+HV6iAMdpH9JFtIvyQZAmXU8HCL
0clmSsiB0C4OgshDe64aXUqQ70KhOVNN1KSQ9b1vCJyVRkuurR5PB2GM+7IY0BBT+iDqyjx6SD9e
tEtsoZg0aenlODu7s3MEzsBVQEcBbNlN1XGjpkpqK+U5Lm/2INZ7nA+Upjt1rSbG5YAnGDKrgF9H
nNPn7fDp+0RgmY9aCG0DZ9WUNxtAAO7ojKccnnkJujrBIvbQHAmiMvPF9IGSJirPEdyRtpeIDpH2
kdP6+XOhl9nSeryga8c/PkOHFUm2vIQtAbNrK3RFTwCIYR4Pw6w8vI6Mbp1bteZbqDx7XUcQ0dY1
0f58asKL0UZ7xk5Dc//vXLyXLL/bDdBtB60l+RG8DnBOqvR/ySVGuHPoR8k412PR9SUpWw30IXvv
acF1juyDJmnOYWT2aw79brgACLwtXhy1RSbM3R9VN1dDLwLksnbHG7RyCDYH9cd0P2Z1ZyVIvAOw
/MXBH9+DG2U3XVT5aMrDrDrGlknQpRSJXw0xenmkR2vTLBpaqvA38M6Nbl4xymBdgwjVwYHw0Axp
fG8N8sHRe/LpqwhZDfbXgnJGOvg2KwpELkDPHkBiFem4n/SDI2NN+zSs977vR7O205kcnbtYzVix
VbmFaBxPWQFc978WQUH8Y0tJGSCU0dsWKKf7r/CEsupkHOJH5qG+DGVbHx6Ky79hhwVaFqnzC+jx
dApsLDRfwpIRm6CphfShudHfGSBhc4S+82vNmBfWmVauzKMBGqm3OLcdDdgAmlNOJaiFjJbUmGM8
7mJ8E2IiVQY8PC7HvhaWSNniiogsglJ5Et44Y3nIAFExhmM+SLNBou3YZes2WtY5OKZlHPK50wXG
zW6S5SDfxOEm+lGpEVPOXetBX+vXqM3PlfKsa5oR6URShGAT+LCM2Hi70FKiiPEl9CFE+B5wjDlC
h8IC757kJooiyQVmL6NUun5uzvId5qrn1og4GVil0sZd/8Yqq6KZyOvw63dSF7uzSaTNfJXu0Pe5
mbQ2KdDQCMLt3H9cSSlNdpW/YXDTqJUOQCZLc3PCuPeZ2sv9mWkRGyXNncwgAlVUeGHNVgoV3cWB
1bD6tFjPQOSC2YBkJ2hI5u03EcSjV/sQqrq8aHqIOhMJvT2sLKmoidmdSOaAG6thFhP8l5NjouLl
gIEJk0p3I9EK3wcLJfsytjdk9TFo3mI4Thf3f5hfEkObeoyoK3WoU1SnqhPEnUIUuhypAc/A3uTJ
5gycI5qTFMgLdg8M+GPZIeoSIG/HoktpIdgZR04FQeY65ackBz0VepGHVJlqMsf87ktyg7IIbmZT
8YOPLL80NmgDOlYLT0FYXQN2Rpc6A0razWIeW35vHJ2j8or0Ph0h4qljB4540j56333pUTh5kAaO
DIU1WCxjckpe2AF4DoTZx9QXBb5L1EBAWNQQRKUsDu6TnCVdfYxHTMlC7Tvp2w8rKqm7K7NXezpH
oVejwqDqa6pLpMfU7ulGmE+1TzzXnCYiTpxYabABn6a4IUBvns4FYgc4IfhASBzjVp2U/Xp0+T+v
826eiBR2D5rBB3LFrqlziQ50esFDhxn9BYJA6Racb9LbUzHERbIYZj8QQavK0fVHr9uWJpQnhkIJ
gfpWJ0MZtEXgHFfZD9zJAq6kq69oHTd0d8PSZaOJcMyL+zhraL+55FQa13s3GrG9spezsF6UQJsB
e3EBA1KU/E2cc6IXAnKWxJDOShPakeGLIwqbmqK/YoWZhM2na92LjQrV2qJ+VZ2jlMcDWgfcSehZ
1wgVl2/YKaSPztc/1doHnIgEg0EwEC0iydWYrZGf3/kjSZsWAqT/JFekt0hJYhnFEfMHn5gEjwTt
LwaX5QhGyMYMTqyJWDMvdNA/KCXkUi7c9IDhLv/v4QEmRfsilxb/92+u0ETx9ehwDAW1r5dPiTLl
PqNbim/oBkxhWhR6EmjXPkI6gnH+0Get642UcwJxElE2PIaOlkJz4g4f65Re4rpq+06GQLvFWYGs
Jo6I1sIeo/dABjuzQT6bYWl6RWeIHIWRZ15Jloimf3CL3kfvHP8kS7ge9UPB2/aXE1+DBiQJjE7D
vnlNnEvTpZ/ovZATufFomf8FGubNymbFVxGWEGv9hNQLA9WEA1o7b7Gpr1p14ubdq4ODI7z/TvFc
qU8mJnHSXH/n2ZKfkZNdS8voCrUMWpN4+1lgfgqCPALA9jRKiof8VqsC6j2m4C1PcaN8VV4aO4Ha
LCKmtnXXpVPR7MFK5B7pVK6/rhvE4P57RBGxIR4+mQNe9rSKKl2bLDC/jGohO0FMFC0/6NpLBd1G
DBFB6FzK50jBF6b8aQTVlWxZ+iYv9CmSXnjQIcqp1e+RcCRnXnaZ0mSCnkcM6ub+Xx/ajaAalrGS
BwL3u40g66TLf+U5OTckN2G5JMTFglPy1emt4wcGMkwDWFYTafQO4d1TYybM7lJvGOd7RCEJxlXs
Oc0w2BXtLKO1QLSlqm2PMlZvPHLe+1PDCX7V8n8/LdVo7GwHMwa7pCYCbqT+MZ+rOU0WTnM8iiiY
7SAtigRM9VBMmTlDxFKjf7RPhcQrjD73JRO7PrKmY7QjscDqgJtnX24Tj8BRasI2YlWSn1s7JxQ6
uBAeOq7mRyIeUPdZ//FnsN5SjkiHssab4LlgY9Zu0z+sJ3u2t+nC1oCz2ae0IkbtBGtpYAnEQ395
Nf4AkUcuf1IUpbQhME2ywrurPCfOhucessG6dFT0wygE3Gtir7E493+tOE/hkf8pAau3/b3bwfpU
Az7eTiMbNioRM4YJp6JMq/l42We/nZ5JBcU+qcMnGUEj7JmPtt5bmYGCcmyAahnR6s0OxAunUshr
qH43lpUDCi4DYU/+OeR+oCbupGeKFm6ej7oeSrgLhSvzPS/blNozJzXbe7tfTSt0yCsePr3aHRQP
0hksU1rkGPxWfsN8+Kc3gBOUsAqocW4jLRhqFtJEipuU6Fi/CrANndY3KEtHq/QCPLicxgCp+/8P
RSfLvA7ay/k2WoUQZkhroc9oaRWSt8EqQx7vPXESI6/0+jx3cQb5nyjBUq7ou1XwLalCMiUqbaOq
0MQEgMdVgOpGB8sDGmAgXLBy0YGrBG3nsdO5QGKDQxH+kMSq7xJI+XKAL3yR4bufFNo05jRQsDpY
MKicES25m+a0sp3vLtBBybMPyQSIQkQ5GOnaGgYld9BOSNx8JtMqGXjtmXMjH48kewG3iay9f2na
rIt91SdcVfMkhzv+9rw3wXQKC0t5/FIEhVjfoeNCT9KH8kmlubLeGu5hjGBeF0GgTEZtBAEYQbXq
MqKd8utG7mlJFtYABydXdhZ4dmpnTK29NMSj+StChdJFNpGMAbI/fDU3GfK++DF6zqDv+rzZBsTP
tpI9D6ERsWAQzqJLKAvgsrvxWa0mlXxcD1dcf+WuylwbEcvJMZdnDZpzJh3bGYV3oqJ6YGHXyWa0
iAKngQ72BrQmKa7bfVwwJae9Hk2iWPvWBThwvvQcUuJduMVpPH/8duQ2QCW6Q1a4Mp0hNaFyVmR3
Q6e85EXyRQHk+xwIVeb6txFoGFNPfokVvBtGPRBviNSxgYxc/J8zW33nJorndvMBZSlytzO9OpGS
smUDoAanteygwHJghMzhLJlQr8TW/31iRV8XBq0nY2mYGDehYFT0nbr+8lfTgWuEwWqUnaUALtGf
SJMQORkEgDJco3rI/hFXLV5EHd+3fX4RG2/Sir3vtCBisFaoh+ReMjxhpyRV06aW36Dwkek40ERY
sQjFzPHR5keotnVZSxuJKXSh56gsi/qkHRewwIlvDMGIJ16uQkS4qjEDjH+99jXPU+AR59tJSbSE
w3I5gIeO+cRLghGxJpOoGsV8mRCGZCU01+3hj9UeXobWNK3BPPYDGoyDxvndl7thTcYQ+p892LpY
zJ3QqhUg0igYPobnUIbKuiUl7EKJmQZgdEezI1g4F7oMEhYlMMnsChurWnhqq4y/iHfnNQQf2MMk
XqAZTBeIBw917n/BEoE+ehLYwopS8Wqgf4xqGS+1g/3aaj+uFnuUFEUuoeak0M+5rjYTr00CQ9S6
QlNXxiQTxZy9PzpeglRPwjsphiKAXMsx85HbNem/rdDjDoK7K3DL1n+VUz7k0FBcspIdvW69W6np
CaJDr1pYnxKXB/yUEUgsbJd8zIvUxq54fEnSPAByCGx2+iW0G5KwgLJ2vHj0oSEpsTHedLK2st+l
LqmMooaAyULywuaZVlWCKzyPItOd38KGDHxEFjmF1yZfVJP6dN5DQs5PY4GxkE92vyUNgRWAeAjD
4nmrUKd+hpF8ZHoqL4Y010mZXovDt+Sqr+oDVlHwZF3mce3OJfedHkEBe/8dNRAUjcMyYjdp6hln
jKKvfhSwsRofBvbpfI13swNedqLxAdrbr9es0PnSJvK4iCQ85AxQvg0B8u/tsAfD1/MSCp4L6QZS
uG9xt7+iwTVXWwzVcagYc8y21KFV4nx8tF6sYdnuoGF2/pufB0qnjKSUFp222FO8mhGMucdbT5HA
CjjtMgmwf07IuQxxHrZNyS2kdBA1xpWyJtB55lUOuyMm2KMltgYETwni2etVAD32sODykc8u1msD
DgEiylFXjtvlheQHVDcvuQJ5a6d07Gm1o5MLSbYzmpntdKkXPNCoE58WAwSWSgmLMe+Q8Z26EEGw
VctfmhuLwTN6WtZiL2yOD3EIydGgI8WWXVUBTZEBnT6F4yTW108JgSWL9CkSTpYsGZ4zor5P3jDV
i45yZ+KL6iv/ZzUrHiDGNVy03yQuwaSAMJB5CsQNX1jpiJw6XIuewU7IPjcMKA7nrMLhfKk0WGQF
MHKGK6CRcUGtQhYkiVVTfiGGNqOa8ktIzf0Bf9c3sgPCry4MSPON3Y/a7xsa0PIGmSAbujZdqn34
8sL3Hm+lkSzb7Av948d15EZviK4uaS+Gk9N47WyvIW5DQoYfLKaNIz5Snj7wlQVKagWbBalhp1i8
N+LdptSOSKLkVoDDidrH43l5/DebCcqzV0OOCUQA2k96kuM+5N75n2h54Kc4+1lFhey0/1G5wmnL
kF0E2Ge9Nge8i2OQlyZVKM+S3wBxKUrI1Xs+HRQx+V+XTkKtcExl9upNpqNH1rqWmqjN4IyAPidm
9UyZXM/1SuO97IzQc2Hdom3ky3Hm5mw3FKeSK5VUT2VW8t0Lv8mKlW/lLzuEp8FbXKYIgtbgUWhX
nTNZeha2TATjoeVEGyMeqlzzKd62NAnuHV3ApfVemqtE5K0Yx6wW4koV+r4mAOWABwr5BqWtXyO6
MoTkhcZ0v7LNxJcxh+Cy8F1e4nIha0AMkYXbinLujMQbLsGg8WhpZZGw+vVeE+EYtIXRd7HRCoBP
0qVdKk109Ot1/fDC/Aw4Nvxv4Z+hAiQZhbh58ywyil1grbX6Px7Z2pRdR7xbqEd+oOjknrRTLkhn
WGdAdwkGzSMVas6ZTq1LZldbBba/luLDGv+14Sxl+Hbv0SMPejbfJ9T+KH+aFoWxXU7aUl7GpqWu
j1ffIu6NXcqa6GRFvtN2DCwzAw4Tg8tKwud8OJaA2B1mLSXr10uzpTAdaTiJnIPHemW2KjRcNxwi
d+rwl19/SuOpHiwztp/rpOd4LTv5hHUywELuVyvOWYrDJxpGZ2YyXmN27WbUbzbOe025TUZuk5Yt
WPUXzPzLNnvD8h3i2DC4qE65yq7d1dCcCV44+ePYaD770/4W5xmeWkA+3XTvrZSRK3I1q8/gqEc3
Y2KrVZbW4FNG0A9bb5cTzVktrirMQP1NV4LfwuzCDXUFTpk+0SgkvtJn1Vggt7D6hP+mSYXY7djG
KJSTZlbuXaJJUfKRtIBW+DbLC8Ly2UhpWLOZnrdGimDtByXPXpdnTGbS4pHCWIZNs5t9zf6TmEJ1
MIIYNojLFEBEL2N6FFZUiQ+abX/3Hsjd7tEfLcVVaGvwEcZ/56/dibZM7h9+Gc5p/0YPD+UmrfzF
6rBczQhME5iPQnLuyzTBHRcIW1D/U4H0o/yWZHQLftLr34Bgr18Nld4H1pa7bh1Jd37BMISnLjrG
JdiuLKKGZK8TACshEqFW6f3MQ8dDutj8blSwFbgYTtJezqml5vJD+Hw47/YZN0GWP8qRQLDyl9K/
MKfL2ggiz65efMzqgD970KUyeYq1vFGEi8uRDrrEABn6jnX8IOEk34JrlZA9fd/CtgmulmVU9ooF
YrT3+ZZp22rfDGOdD+IEj8wHaeQJLdLBxR8nepEjNWt2qCUNppFBezS55pxZ3CM/DGmT4rp6ynbS
RyxPJ6WzFtVr6iX5OWXTr3rLaAhQCDYnFEjamI8A/xKj0dNVhysemnFZhmBgCrtI8OK2YO4Bo7Ec
s5IX57VYBCqwi44V1JDTPqXXHwFzURdk5BQ3KaeVf+oBKhcSsSPr6k5XNTMDfB+68UORFHyIYI//
VFQNeJddinypRHf5uG5iVqfElYwf5PQVZ+8SQD6La5zti+obR0MxI6Ct/rImHVrJFEWmVAhAOza3
iw4wrDJjW8NcK1VY8E9D1ZNR8SZ4WBRAAifAlqW+sCkS4vrQIWDzWP7I4HGOatcc99/FQZBIzBdT
6pWkGdDs0FSzsz0sNIJFn8tHfO/BVnUoQerRBbzKpfRODaOXOLZVAigdlmLlAqM882vrvrAycgvh
D0IAE12nQNtYAuZWLumIVEbp5j4RoFHW29bJz4KyjOtXJ+RHAoO9Keu+YGnt2imoxFtnckpTOp/b
a67ivQF+VIzmBfQXN9HjJvqxzREnMsnCHauWRQ9DYjU9MAG58rRCj9fdw9vlfTBpHCV5iP86ZOq7
NF+jrhzlw8VbR0YUXDH42sWpNdYFQZo8t75BemOatHkO7NVnSFqLpz0WH+Ivj0fW4GDU+aviqpV6
YWdVL9VKCKOjP1OT+fwVN3vNLyyfNk3NPgXbS6QiGOCtmX3XP8+4cUm3eOrYGvh/kmVqcwGIY4SA
OQXRa6CL4/vq3Odi+nOa3sOWhYQW61Em8KIppINFS0yciEbNFA1WR+WtEn+POSWNaUCb6vZ3Kr6Y
RMhM/R6K6SFNgeql0YTtN48ZMiJuizIOxDX65xCGMxxKQklPG3YNNJf4KJ5iyjxvYyrDyt4sd+o3
V26pTPb+55c8aY5pfQv/Eu+WnU6yJ/QRvQzpqi1exMVcqJW4+nfu2bgSxmiHTbiYWSPSdWosSJ4w
UKZ+SfHnUCXK689R5pdV1u6gSiYkM5KNvrT1mSfmRzL9MLZRUf7EIsBRdc2iyXcHu4Y8cnl5YCB5
NZ1lOMrEHnJRMiu5WNOSuVEKR6RMJVHFhwfwKl5gHm3VZfdj3Cvmu/gRW6JwoudU53aISoebNN5F
UZQveVNWLZc7GYLBvnqTPOsdBuJqNPu15et21wfHYn37cJaNz5J+ZWSA4Dx1RRaqg8aEj1ZTLMzt
zyU9S2TSayOrc1km/eV7+85yBRUgVykmZbGNusBuRRxCViu/yHXr9JEWNvwcXI0fr/a8rhwJDQxK
4gh66uReHSi6Rubo+JHQ6aYfIWpH79eU4DBacMxk3rzI3CLSWjzWmRBy1ypx2CywlPkELA2MdHC0
UHTk4IdpxxW5tO9d9fVCFA/JGjEJbrjvTg/tUMrR0PGW8BZ3RkpV5SecJDxKKHQ2ucricwqHAjU+
BU6o84cgHo9TCrp4JE+s9PQLOvmaqwr0TRT75NkOAGtmSQ/DuJ3d1Nyg1/OwlZI+hcGWO8qTSjwd
21j83dtpsd5FyIQ8q7uFVbC0h3zXe2H02KQU1DrEUfZC5Uu+RG5xDIsDneOGoqZ6XxbnJ+K81xW4
2D9O/dIuUL8RbWxklo6liuzBGtHajIMrAMKK7h6s7SpohnNaLSRoXLazSIk6snnGC9ZARzSNkHg/
I6aC5d3hTNtvVdqMx7EpEsTsq8TcvmtdINuC4fFGq+ZpNurr69OKgWDRx36B4F/g0+FyNgmkcGFD
iF6glOXzX3oGuGwO0GTglMFLICCH8XEibH+4tEdxEQjxLvksXFAgRFNqoUlLI93egxPORdi3hzw/
E+7BeVB1xVTrDSawFcS4u8iI/OjxWFd6XQ+iONw0kvCu6ZCnxd59rz3pb9bDbDTLC8hzqvblzp++
tACXgKzz+h/xg4Dt6qU2fS3WOmNBjAdg4wOh/3foNHE9hCz/3CHlwgFyZimDsND46zASQQmdnZ+4
cN5pRKjhQ7fJBiCWNAwhGwn+ZJ4u4hAFbVHuHoYzFKAZmQMp25YANmwiCbfXf9AeI/i0CmB3rGJa
oJJuHwGSWe24fO0y8RTs93XoQdcgBZsyjAlVVc/Gaqc2QIb4C1KEDGPnq6nAw5bKf0ZVBoQyXOuo
NdiU6FyOQYTSuxNpvM9DEaGiADi1gOjSPAyc39/c9vzIGUs6M/JgPs0jXF7ORMdJPa81wfJ1mFHU
xQkGPx1I4ElGl3kcP3qu5Vd6NaYiQlMV78uwIcNsQbl0sbhY8c29yARwP+ebAj/ymZ4O/2dmRz/J
ejLHZXuflAxQp8BGI85wEGsG2ETfoywO7PAAgeilKnzowCdU7RatkoanhQfBSb9i97gD0WfSgPAP
LlflR833JiZNidebWxZiFv23hSEp4zAqpsQxdP1t25amWhCYj6lI0xSK8380qmf5/h/sxgfQnv34
xoj6Z+J3w9WrFebsZRIeB+Ha3pEdrR23NHM45a5UQfzsjhNS6UCrmj3OHG9j8OEpqYNof+DGW8RK
yi9LyL10mPXcGVhzetpxjE6IwkSqkTdbKnSN8SEbzXzb5KoGzrTZg234JC/K1kYM5CD4Osof7ZVn
1WzxcZhuyg0Hq7hNttKOKAj/ZijtHzpY0Vl04vaSmIRfEUnEhiszdH2mbzzWLo2LYr3h7ZhrmLwd
u6BJTdTeK3i4/vk34MGZq5/Kh2CIo9EAxDe99Y1ii9MoPl37nptKeZ58m1cfk04DcWsBF0esoBJy
tAN1gAMBylFioQ4A8yzl4CW/ADrN3kcKMqRxfHZW7otS6y1WHPHKAzftu5itfB71azCqUkSxtxEo
Sdrgm/zoKQhTJhUxpGoB3x/GC4rRu1dBdt0yG6Zi9OeTO6d4esuKEjnqOpG9N9pzTQPG1DnWbk93
cne1C1Nl3Pz+5fUvQ3Y744neag3LGjS4GcKf+PHmMT67M8zRqVpoNn8O/aPMlL0vELEpC8/+M4dX
o37peNqvNXIwq23WjeZrgMfR0+DUfxwz4hVb9N2LnFgLhfKwzBULzQgMJ6YDsoSiEzsonbXkEMDo
dhqBT2mPb8LujQME2YfdRi0qL6cxHSvsElL9keeBnioQtRvj/+zk476rOuwL2iu3N+OruxsIGSw1
BnGX1CVZFsRrJAFPyMmdojVELa7YHWqW/B0uHCrylU9pBiBg92ma9Ph5dankxrqYuPCz7Or+srph
1p2fdjz/H9BU/X4m9BrByFAw6ikSh92un3dlO2cWmVi27ZMdbVg+2H817XlecSyJtkyHoLITtZ5a
ZlDTmmEB3LurvxZL29yEbj7T2Rt5jq1HYPrk3dohz/R/gEB1hpuXGPtS9SIEJCC16UOwFtCy+uTE
kS3SEmgvl/31HCwLNV1wnbLiUaQ1sZLopVhiMnwWvQFbR/+W82L/SxNGOi5q7XGRTwsVZjkvVxAc
1UWJ+qYfIUnDYBEcQYJ1uuuj4AEInGpz0Lme0ZRRmIB3vA5akXEIRbpsMEPQYcUP1Tq1K+OAusYg
4PpnOd87VluajiNwCgKDFwka1LiROM+AijUadU5tUwmdb6fOadwA3KeLwkNMHNKyinkwSnnnRQzO
vHK0Svab8STuTIuNMlCbTH6kEFC57wg9bVfNw5w4rAHVslLHIlpWM8JusJoTMalq0V81+/+mnABv
NzGlPkca90na9sRMUPDRmGAjfbf6Ac+EL8Lz0hWJqv2x1MlLi2pQft4tOZolkMTvzfLzmuftMwO7
aN/hzx3S6va9XlO1B3gfI6ZyjS7whEU8z4c0rVB6a5u1pVnBPqECnNK3NywQu20f+y6wlQFBdnhW
tuZ3ptCePyTLCCcdlsiSwnOvgBiziDE7Uegc5+VnbNadViKHAOJhWtWxGGtVxMEVm71pmxEp2l1U
+aQYKTZyqlOPyPm9hFn92aiEzoef3WUhAfIxG9HmFhLKiaCpmSzmrocIwwclvPHebc4Y/sac1AWV
JfZ+D1tR5/pXHaK8J3OATBTReVGkY4FjgD3ZRluAazIWXDAXHb+M2pOgyLj+MpdPGd+OP/ZlN2cF
xV4KnKumxY3tQmM8fwR2q72naLJbtLTYC9QWq8apJoJ5yVzgf+p50WXEAElPOkMXnc5i/ucTGBba
eMc7JxhsTS6sjBVSsSz1QkaZBKx3Iwy+MoX5Wfb0K5mgfoe+VIe8jXQEb++o/wIEm+X1Kr1rUmC6
5wMp663CBGg+Ff4g8dJQfcwx32SwMlqCzGLY1vRJ91txpMkxXP8pcDiRq2TxDMj40Q9MZ0kP9Gxu
lC7Vw1jmO9fmBnhQ+nteS5gIWWj5ChJsR0vshnJq1Ue3/ZMrTAqusBoL2LBKWrvLT63qnO+0LwE5
erg4EUVuqj4K//lcsiDJiy42knsHQgngdqcrooDvwoqqPGaov/S7rSNqMK8tgJWoypnvpUWsSSqm
r+Mcwec7ssny0sMbtzh6NX4gK01zXbVboI+GNaD9DagS4Z/w5cV5AOSqCtASHbGYnQQoq701k79b
Ju9CBd04POmTvaYRADR5n6qJiWcqQkEXCIiaf/MQsmHhQ8W3QC+IV48aNi5aOTutjhz9zAyRcPDY
ODpBu0/ULoOdaATNtJLHqRVlf0baFXqOB5jLfAGeJR70OT5+SDeK3EREKaq1zaIad3IhdVWwIkEF
0pQIrbh1YSslaYhx17ehu+P5PVxqJ0sZtF4gPnxct0jWdwbYLQL179IyxUKlFowzzcdjdaABOoOs
gIMdePi5rIQM7u1x8kgdXbxUSfF0dYLfBYGV2HJLoGsyndSvfMIQVLOBWQKTtUu5/98DBszL+jJA
GRlvALVtqtAj2Eck/2K3z71nn7EUM/ZHLK2BeZ1AL7a5gHMvO+Oyvww0EeLyjvPssToP8uEKBG/9
9IzdWb6l1EAMvzkGkLrY22cFWuJd1u40keGdRhGJ4rhk6aTust8IK5JtYsRHuG7Lp8Ixmh5HPUNz
n2O1emrKTOnb9FPmbgpOrayLshIv2qkM4L8PmhXBl/w3Mu2EmORvAAiUcw+sxKlfElRTq+f3CIuh
WxvlfjUGmpTaYadKVXR7p8W66gcJlEnWO31VwMVLaXJ+X0mxuXPOFU2p/AMzyf6lWcZv2B34M5hZ
aA2aIJ/jrYHVNdalBxHbXbYUIUuFW/NwkkK1HsiCkUTQwrnLV0wveN0g2nvbAKeCh+szDSOSKX/J
W+V9iIOhBlAv/MpoAWlW/RqcpFpI/YvklB7leu+vYzIWvQqbzu30L6+pJ+G+Wdu+P4NwzMfyxLM2
AHJlrHKkFCeoqYOlEZtPXKhO5ZiBzU4qfaSzT19VCtITHePm+5KskZduOjTrgZsdEQ1JShg/Ko5K
pVBUa6Em6dlZ2vmrEKDt3nv6PWkq9l/gOmSZQ8ht35Xi6iIP/+d1o6cFf1wrFdol8x41W9h4S9zv
Btrh3SU1h/jJ0JLl29swHKpfTRu9HThcIEdLB2QBJg+7Vx8jtCrCV4alYFjMOYU98Tw804UG3puQ
WR/ZwlGMU+5QHHnE6JEtnluwcnYij4aw8dB0rS7/LiaJ47nppZb7R2qsucVxAqwBakidiFkfHem3
iSS1e7bN1LISYwsvcG5ZoRuSLhfqNu3h25MhNfYwaATbzj0kfuV/Nj5FIEX5EgVHsfGItR8HHt8v
Kh62QqVUWFD3hAzAg32Fb0RplANnvrIN0/BDkFimckjFApxFkny1L16ai0HTPIpa03347FJQBUUi
m5PdKtw4rKvlt3Pp8g8lmcrw4XnxbaEu+cszBkA5yGQ3rpH3rXM3A1TN5ZJkOMOfJTIaT1ZtU55/
TvbXz4uJaBlWnwJ72PVPh+rSJn022RpvXuMU6wBeaMkZTjI16vFGkToW0GmE0y4OjZDIP9IZ6qw8
kt1rzBqRfe4CrzgPiiNMDKKAcaC8pr5DGzSS+dieEeRYpATG0QaLib/Q5R7F9jkrejJO4q6kHBMf
bgtj0xwPEIfimLXcv3PYoNg3UwFPXTy3NjHqtIk/tWViPLt7jI8+df2zhULvmG4gvkoswjGAEVY9
5e/n9bORnZ+jPVYB2gAGHBXAf3oEzzS2cnc8f8dmRwEG9Ca5175VWtIgvirxBhFm5LgJcKYDjpGh
+ncj8jyrWa6BK+VuHfL9phD94uR5qpxfhaIuF01obSDiwOxp7osGomk37Dp7FeElYMOh1qDlUGxq
eJmVF34e50lkW+8FDU9Dsam9bzSaF9C/fEW/8vHAZkuXZMlcpxGWwd7iCmDb4Lk4Mb0SHB0rtiH/
sc08opekjyyn0qKQLFVl5ct9Y5of2bhNFPPyLkNRRkYpf4vK+yp9Cm1yQsrscBR4HfNfjjGqxIZ5
ALW7so/RjdXE2W0BFQF2oKOefDdYQceKi0aO6vOhR42x3NlZ2H0IY6iJ+jMIxLTvoOjPnORPdf4r
GcNbcfQtgT315i5xy6wl4qGDZue8kUL6pIZ18DCD1mbC5dP4gY5WRqkq28AODQCTRKTjDIEtb4/9
2DvxkeXoxVPsmAXwXurIjSqV2XvOCxEiI2gknYZizOCqv7K6SCLR2QgV8r/jx4yOL74K7r6NqbS9
L+HcgRwJ/faIQ5mgrWCmONoAG7DBPLeOIleL1trU97FlVRemFFfXxX0KA/FgOl5Qe+QNuqBiYlyf
wg3XXUdDfHZLC8z+g2XFbmdxet+4CbmZEwR5mt/VvBW32W28VdWf4u3CtY2/QyOABJ8NOKS92Tv0
159CpIPyO2PHD3DgXU1jbhNvq45Aa1BvS7VEWc2knJ2cxne34iOyeEWM8s17/KmKdN76po7Jy7wx
xuhsienQJ8EqPo0tsJihzAL+CqnqjY0nLKIJx/t6hECctLI/aerDLXkuDKhiEC3e32hPHtyxkCTE
T8ILZR8vDkZwosh9OzZoxlEbdhLBCmJQMQG9KSdJnrfKnH/QfcnmMo9lOeYS+nJnx50pGDP14vCP
BrMPT0uzB3WkCGpPGNbRFruQcFoDpKIgJArbw732CIJoUw43CYQ/cioSb6esp+cE6UtoedW/2rEY
mp+U5yhyB/MM7ZUHmp2/noCvMLyAwOev5dtmfEZoJZMiEXM2TcHIrknlkFOrnGZ99lcx90iHaocK
CUyINauNGAuT8p05SJXvFfKLaP9tn/naqUrjQTgXESqBqPjjgLEJ8ZbSWossU6lyyrP5eAJhKkHS
FSPhNy6UM9nlvc2YTGome8PfA9xuYhDglcxOsPXdNGiJ1pSR/tlI4NoC6sMyk2n2b4YpHeTk8iU8
D6lLc50HiV/G7iKbYAJwhfQ+eLFUUzXVPxqM7HS++/qsJBAGlhbx3pT6gZXJX8AOdqt1BcukyN6h
xRS/XxJA9Fxad5Nv4J9VVlpTqar2KTfoG1/Ls3UXFEqslHCYKO8v8EGcFd4TpfG1jGarGaMSFelx
N5FXMOG6LOzi8LeNg2KnxQCRZIk4Nt1DB/3s/CAJDdadPJOBedHsgJ/MiVaZqI2ePMV00jWRVNAi
5Pls3P0HCLwg/Doaj5HbQxEDm0A0B1DFamdNvn9aA2mhmrjLnywTPuFeqRkOn8ZGtuR4Rhc0oJaH
Q0LfXnbWiYYE/BuX0FCl70zD/3/Iu2NPCxCsICi7qtxl+0a2KdEQ8Lxgr8BLlfA7bAXqc3gTKOnh
m0pY//RA7px0v+nELThHhk8LCY2WjK/heYdwvojR430KIFlCzwAjoEu3e6CN9/RMeCTvybgUXOL6
7ZV0Ih+M8kCcotWOJbMl+8FYoGmhGSjaJwh00Qzn7FYsLGVE0M/WfAWVB/xvqWhXAnlgOfMpmmBv
U2qrMEv4ytQ9oJ9NFPNortdVRUJGCTIF5Q/4SOBDPcdpid5lEeYvwXxPeOniefM9XG5dOsXLmg7+
0G31CwIc0mdWqZohkcCbc9xXj5FGjn80fFRfU9yoClk8JPaYw9K/t4eSd7aLgT1fuLMoinLEQR0a
vlDzTGR2XqDn3jXjqvyVOZvOYgx68AIiuuccu6EEUBNc9L+W0hYdh0DPeOq/4qD/iyEPpWQtGLPc
spbIU5mpT5RufZh6FMnWt5UZb9EN7NYou4YLrdQz0+vlKZmzkuGz2yguanO632xvXGYs8px9emnL
Eq+GezaSNVIsA8lxi72a+dRIMpQTgpIpfz/c+SSthursljGDaIxZwrqcQJ7GSPUk92yUVpVEeUhj
aOnjFQPq9rAv1cQCvVDkNI+x9kuak9YLkWZ2OAZR+jOgvBjyUKcODyo3PFsbdospof2EhXBhfWw8
XyOMTExnGRmfbn6Gvc+8V9IUgqmES3v7IWqEzIu0S604SQpfsmqZ1XFm1m2mbxzW1tNdWHWT9+ag
c77z6QMZ085hF50TYDfH5qHq35W8gU3/syY/JtF6D/PhtI4saVl3Of+YIXUr75EXR7HWCJgqh11K
ZAXS74ixUATKX3KNGY1flOJDaO01G+9CmisQ8/WgtY1+yBDDJPg6oSXTLm2lSaj6vcFChjcubNvd
t1bNBAgs7Sxqvygy2z9pyH9yHSCZGS8r4VrzIR6TMN3tNhikOgm6Pageev0TDvs3f0YWryryBqXL
WUeZnJo2h3ZhqUl+M0i9JmT1CWGZPFQj2xfNNhTmztkGDg89EB5x7Z+QQXdtoK4+CJ8RZRUgW5N9
dy/9fFZ5G2w/hrsZUlcR4wxKfL+0o6QNZ3hdRp1q3Hn0+shJZVA6ZWOzApIfQD+54jXXJutdtlJR
3I8lOCCWNI/TZCaJtympwopQW+oj/HeG9Ol0+8oBElppgkv5FYDNH7pbjjiGWSy9hxMGhhqqn5wS
z0JrjJko13kwEG4hT88VVZu/yHCJKekBn4rJjG68lhpdzzTEHg+hjJbkzCtQdXOy1ymGiPOGmBvT
KfIS+nSOpJVxKl+nxOAEz0dPTpRq+HXZZLlKUYKiTxidOp8vLbfuHeaFi/NE8KwxhjeyDuKRxQ39
dgQejpUJbe7ljEYd60l+86G3zKfm1Xz1uL+0EEWfMRlO0DUYVj09S16W4EHPF67LGGRy1WQrBzXn
6oho8s9zb7h2w9HAC9bzvr/oQxm88G+DvyJTPeDvPK/XAsWp2IVto4yl4KWU0Wu0f63WRft9C2ZI
4mApDjWqZsgudSCTID5GVvU4Mxu68Kt7Ud0zIg/1H29c4cBB9fa3lnlPoHRm/LFr2Sn/TCtcT7To
Pis0qPFKPKDOiZ+Oo4ACqcjcEM2PZ9NaYeH0SNVSRsb54DuZSO3xx2LkBF+e6/WcKhU5ZC26KV/r
c3Ah1dIwwnIgkvhaA3dlLqJ9KHZbti8axJqcBP1coDstDkfGLu6g2d4ultw8toDyF8/xxjFi3G03
EWCblj8WQ+o7JRGHCtPIgiHHD5mtgh2zVQmhlzuzO577NjFfCJjs8hpm6wsp8QWtT7rcdBwHYU4E
kCHmkSXqq7iqTtWqc4zNGlf6qNB6eRT6cOBTUH9KLkaxWfSrk227wc/y3TwScfm6OfZCGIf/VOOi
dy040HzP59BZlgoiIBMGmETL14+sKYBNfD2k1+cNREb8QopF66rD+fncSwon1fSCXH3aEEjF5FbR
aaIyfdF46/fak+7dbZcLyiFForM7d36BnhpBYRFMa/MQP9YbXyFhp6MyE61oPXtR1NV2Zq484oaG
aEK3/5yXJxFhGzHxF5YbYdQlOhMbHqBv8Utk9x+rqLH/AoF6PccWBDK/i/bdwUGqrmfvNaHCbdsO
UQWrUaBViTOHCg7sAgAMR/Wco7RpMHma7f8jmcyanbE9pCmd41QFNNvxM6qkMNBjKFxHmMyil1H6
ScAHXwUKnM/u0hH5jmr5cxz655zLl7Z/KOX2TxAaTDoXfK4b9DBHyKU4tFcMCTQzedqNFxQBmoQ0
DxQkvtoOaK+E2pvYvOjKR4cZdtXmTD/VDPWU2kq4ZqlMvsWGK9DXMQ0B4uLLzxHKkUaKOggukAet
5/AS7yfHduoM4eOdpok5DIJm4FB/27PjvsTj71uxoGEac0k8IQLRFpZyJkuk6aWnrH4tzt6mbGeR
75zkV1uS4mOwPVHst7jUMa4Ep9cF6fS+gdpJ/L+1GpVWRUDrGrw1sG152N5/IwblM/l8e0hh/Ffh
xJGx3aOC0OL0dNIBfUO5Fda/qSrOoCwhkL9LEbTI8sQzXz+wAyQ4D/EjosSwX/2RNAO5KMXZTojv
AnRuzBBNLH2VkWzNbxNYK4DK/vfai13A3ytTFLw3/9t4Z7Vo0DB4uoRzT2yDvAIyBfj0vM8ZqNj6
mqc3LFW+hZtsu9KaW7PsuOkj7QDA7IiTckLXZmclAqxl0USdwbcx3HD3tTeiDZZrHVojxnvrLtwN
/5PKLuUuQ7j4fPvcUztq6ck+NKMkxkBGRrBzfe92RPHOMPz+8ggUtCoCwbP3B9vTrCvO/VvzQZQ3
yrrqCTNL1duG836qkB9lRTiaLr/0w2pLVFhD/Z+SAzi3+vSer1ga2g/JwbuP0JjStuNRAITINYgH
KiLA7Q+56jR0BP2uXwdASdArXE19s23vFHsdIxBlFNRkjfMNjY5O+LPaojeIaAGBr9wzeaRtcwPM
FF3jsjbxNObYs41gG54aFR24Tq/nEdv/pBzx8T5jAoF+b7LpF63paQjwqbc/UP6YmNWE4SkQRONy
kUWouvtTjCPmJ0BfzofRBGMOYMpLNcNhLTaretHTR/jqSI7WNxYkM0uRajDaRek4OzgdSh1MafaM
NDQARWtq86n1HQXkP/LReNTG8EgRSFaqA4icdmqX3aL0Le0Anf6ax3/52oumo8wWbbWpH80KUMzM
iumSAPpeWen4WANb12/d3XbNIQ+w9W2rIsKpIU+AsDWjPUzNyyiF+1iHtk7B7T+jWkF+MbtMjtCy
dSyOXW9cvi/m9GgvdERU0rwXcdEx7YCjWifr/BoTbQiojlnasQUgsZC0RwMJEDdnYPuvYij2OP80
zv75/jZpIH+fxoDXtovSYgsLcgYy9udW8z7uHC47YQzBvecgvv8kjR990pxT+vutMYX7MWNyCTTD
T3CudN0P5S/MEW4yYMGk1o4g4IfLkpx2dNKLD1JKRJkYR9SAUf+w3KIAEiGMenDqLPKb53tfw1MR
RdUDftis2CjLBoddfi9VDibuU3TLWKrWJzwQ7bQ5PHNwM4ZmOQtZ+d7uGYjqx02S3LaSGpyd2Cku
8vkwldGpafpP3cRzXJY7FbaYtcGcaCAgB3JM2CbtrOgiX4uaxaxt11F6aafH8B9R0fJGmrxrDjff
0vWOXoqm3G6F7YfWrUIc9xE4gLqsbR3mB0CrMaDn4jAKxaBycUecF8teX8VFhg4SVK89arnqakEB
XLSnt17Wqy7/pisqT6ymLL4G2lZx007nagUjAAsJyoZ77GR0o8zjUHytPxGj2ZvjkUhjl0y5wpxq
IzRefFn3ULI1BdkY4qeeU6JRDLOs5Y/tAQkzZ3xek9W+REs/im/bP1pf4RpYnhFg5c0kpng0CNQC
f16zZk/XHeYfFfGUtexBfh+ow8e63Pfk0465JDpId1JxZWUZzXn8/eUzL+Xxwk8YukklSlibLcLu
nB4+TzYMGItOy0lKKiNdgOEbJOQ8ndk1XFJ1sAwxuU6SlUGoxw6Wqxadj2c4Ki1R0Xg81nAyhvX6
GwerPrADyslsiWL6nri+acY32Mn4PyP/KUt/Hit7TVHqbmQU8N+pa6ajas9VxCYfyM8gpBjGBm2l
UEbFH2zVsor4BUY+N0sjlb6eVFdlz9SUS7YuZCq+F2a28nfaVsrwAW/Oj390/qQv6lO0KfYJZc8V
K24vgIa6b7lORHo0dZiTHKRuqsUPAeZ9iEXuTk8NeXlpybKRaapTV2NBrLTa7VAwkBj0VbAgJbf7
LaeA/j40me4krIkgGra/CA6qH0XU/OFqtCIycHdkE3gWpJchLxvJqYaMYhglT9AHv8Rh42e+Xv97
VHo3FnrufcdsMPbxcQnaHrq+w5Qg+yYfqc8LMv8e6vngr4lVwyMVr1w9dqE//4GXJlWSSnTvmxft
msDkN+7I3PjZZoCWWruQi46tkpOac0IVWAd1pfr0niTIp7CfZsY1nSz//mYeS4vR8XPukvYUWKtX
2M5UhqNMgmpRfHhv4psU/EEmkQjutIINRAqWmH2ZibrlByDfXqDReIkX061Tz1HtAxpYyYhTYgls
LTMe/3tRpwdLNe+q60aFGb54a2OaraZY59h3ij8RVV2Y9Mgk8/7DPfsIRQdSGZuIpHsxdYleOY/q
Wp7OG1kN0doQLT1xfLpE7gnzNgGPJooMx+5ezAKQoRid+PQaQ8cHAI7i2mTEBWBtlsNAeattH560
TG5w2cs+4B/VJT6BsKBVni/hIDGRkjvCe1uJN/sp+GOfG5tIQork2jNRrKREbjGIvFh7txNjl9Hl
jihG+00PGsnzuIxBI8O+zgm2dxoAU3avWbeqdWf7FBeYqiEmJgkzst+Fv5Rn1CejKjPJf1DKPWht
xdh9au6X9pIuoacWDTjiH03BkHM2iIh0s82s1vf8CHn3LZjWSOr83pumJkjMBjQP9AacM7Avy6Jd
HFkUP9PFT2Mi+jAwVeiG/mtdieuhcgaAJ20mWBybBLcu/I86ccY4Reh0i9M68lua5WSNy/twK+8b
12njr24q8wE+dnhzUEYoGGi8wXkzZDH6pn1zAb1AACTLC/OJ426ELNpHdZffuzwmteTsMw9m3KZD
JZnn0K3ZiQVlvwD92NOP9MU9rGKCwQlYZvtQd4Gn8k4oOEV2GbvEZxWva0vmhje/3TCuOvxTytcC
DiVWivVGlDDllJCtBQ4ZfxnOM3dJFiE8t4EYfbgdtwNnfazetyWKEPIdqDrWO2F6q+rIq2zohkMC
FVIdBz6460KbfrjHiub+r5O+5aXm1SyGkrGu1fLL1B7jGSe7aawejdSGgf0m6cQZy56aEx1ydUIn
67W0GoRh09SuY7sephjmbBuuzOQnI283Qqnwv6zDzHW4r/wVwgwRDJZUsHKFg8/mYXvmBEVIAVZw
er+HNx8MjhLFs++vrfB3w/J3zin5IKj1HSgabgFU0lBBCFXJKAwhAjh0FxNgV2E0bxwORBnQlJCe
NzdAFIznbkDQzkRpc4jQVL8HcdAsJqUW0wR1scwa/HMBbZLR/a17DdgZGcu/ytlwDYCgWpvXmtPF
QbbdDlUo088kG2XrxM+4kEDCVT0nWgTwCXDxAnAFj0bO5eGP0Y5o+4uC/bNSWu/vTbjfs+xmewGI
1BxUM8Gn4cYdt+k5y02mSRwirXiBSLmOrUusprBjV+Y8Iw9iiU17wzneBHmdVU6RPLjGykP11KsH
Mbkw26n1q8+jNs4mCVksysjdAk7sOS3DV1JCjdAf4SEa3YoiR4ZpDoFDVjvkjIMEdGgCyOZtaH91
I32bidV7Ymzi1WZW+I1z92rbsUxVXPxZ7IV4patdR4pLByDO7d1f3kovY/hp47w6OaQ434l8ZjYK
k/I6R+DIPEMgrX1zV1cWWZVMvWbGRdQrkO7rw+xSjZkHumkR664F37zZbXB2DIavgaiJvtg371QQ
yL9JksV2An5EfNTEmNyAYnJt7EUs2TiXZugMP822WdyXuu79ub/IYnxgzj4b8nWhEoq+ZAQXO4lS
T9CViyC/lyvGcesvrmISosOXMihi4cwECduI6BoAGL2TcjTcOI4NPGa1syUibjjNtNN321fZefaQ
WOhB5VsWIWDbJHZhTIbC9+Oq/pFZ1qrYS3AVS7MFS3nrnh+x1CAcfkt6dQ1IcVsjRHcP7JgcqENP
QR9MCAoWFECD3LWTXLhtUtzqWBcrl8ikbLtv20roEDOhtK3jVErHifiUBE/jFBotLvuuD3SPwTL9
iE0ugpbRjN9SeiaAOHlVmKKYfMUX0z0tZTfGFEv/VwqqEcs4+giHXLP5FGahxSI/5mlNEqwSmANK
d9eFXVP0OGzvNh6QVMCWO1COolfJ56/QIexguG/9MsAAokhTEwAkEzZvDAxSa+XnbTgMNc0LXkZY
oy4NYp1SI6DXjW+s6ao5xOL98IsUeEn7slAyGIQenB88+czt249o8yPJAmZh6/n+aLCBel8Y9p5E
Gy2nvptrZ1k/SWIKCJTWdteANSMyOtsvb3taIQfAgYDIoLIR5+x3zylp5y0nGDSriROqlZeoEMcy
6ZKEIXw6kq0qpOdxplo2YKifSjYslyWMLFdzU9TbX0jbIOhg2sVvEMidH2JZSiiyZtlDs85JZDn7
HfZ/ym8B2skDC3X8WCV4IHYYp9zuCbO+ZbfyeWiH2wiZHaze/CgLuclvWHNh0iVnqDtMejXUz8P5
ECBbbcU/i4E9FXuAn7sqe/bAKLjAa09bF9ST1crs0MZPQTFRWKNu6SKg8y1NZOrydhvQwtfEGngS
Ih1g/PHyUhsMAaYWG/8hatWuCnPNBnBG1YRkFIKeboPxvji+Q4saI1TH+szl8l91o9SUGrC3PQJI
DKy89sMPzTmkcpNWv6B5iRzQuBosx55eHVb5D0TE7uQHvRpPDYVVGoEdepdoi9wU/WWzaE9Evyx9
OHWxNs3QKG3Lel27Psk56eAkEkYAbZ7JXlwCXRTq3Uah6YB3EOa4aGmQ4IfGG8cT037KUM5u8w5e
+wcfPyJl4uz0qSXBFdeqTESfWYmlT4F7pa7WNftLb+qNy8TabD0hu+HGPm7fm55P0jxYnG+9yY/g
7ZQ3PZQY9rwTEs4MjxpUbMMOgtZ8jv169tlZPHwGee9FrqEjErdRMEB48cdEqipw05HYTIW5OfIw
svIoSDtY4vYiuLHCrCbFvQBl6FO6y6t6VEuEOyhY767IaoCMi1a+MDRZn5gQ+cGFus/lqiJH9pTQ
iwQVr9iQ+uycWvm6FRHAhjnk0mQQ1kaylj5aqnNDOzN+P55XJn6Kos8AtzXRLB0fE8wsvc5mEteB
dN6ykLK9MicJX9sUQIfHoQ5ftmV/dKRhlZov+zF3aPdB5ygLROarPabhVFr/cykhPL0NwoW7+34k
WBdAeqcUmAnrsOgqEvycs9+K3kkNFGBozI71Es+cmFB9kt+LZ12DVXtNe5D24c4uNJ3I+3dMQZME
X5LbzSPYKM9M3lSpNqf/FAC+qJFp+hZRBOjfMQfi4awFRPeqey8UTnHbIZqx92/G26D2R26LRMIC
pmXex/3/mKcJAd0cfPAjH7OxV+ERxV5uHHD9J9bR9xGESn5G4ZZV/kxN1GWu2xQs4fwzavTxjLer
e4BDpp655f+5JDNqo82uc4R4h2f8893M/kkXTtsWwi2L8eD/q4JMeyDYlUaauuF/ktOi0y2p3+vZ
+lI0arqNf7rxz1Rx6W0RTa6Xu9XzSh5RxwfzVq+ARHKl4sIn6Cved6UPPa545A/4MPHCfJ13pIGH
5vA0cXZPk+uhh5/Fz9y0MyoHeNVA85IUWHFzfGwg7aIuwl/aU+ICYvhYTsSKq5ZZK2QN8TwA5xPm
A2Fv+0vZGC98R5NyFl8WdNb9k5w3/q2G2k6MAHWhh+P6njtKLy3GgJ2osOxWu3zKfrOUkH3ySfvF
jgkFE4nCFjVX5M5oYCIR81QFa8c/YvWm6g==
`protect end_protected
