`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hZClrjQL2xcvpkOw5/Rk0YfU4cLpkzqVyCWW+vyfGfIwRXry56MPNeJiKWSo2kvUzFNpnQa+st5p
3la0itKKWw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cJPY46dnrBJ9tXvtxt0uojXUpj8Xad3TGOGCLvqfcn4WvGhwrOJZFUe/HwihZ6YPBs7rBkt5Uhyh
Xkm+k6ryH9Zyr/Cf0z3ghL5tiNSKvqVnr07tvQetVbBj1mTMYyrz9PaJbZ2GSQ3ef7FulEtNjb5d
Ef3ip+c6Tj3HkCyyiY8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TFQ0extCZz/E4dn7YXorUbY21QuuDSbveq26pUf3opJgYPyzCKX0OQxTJaKwiG/DkXlSQ4470vtG
F64mjUEEXYREg0yfX2fIKjT3/pF8aLzpCfQ1udOc8Cqg/Nloo+JsSd2tPEDJWk2su97x6eFnk78x
PW3TR2MiO42VBivqermCpO29mieSZnNoskYUOHLuzvhIR/J/cMXMmiRcjbEh7EJOVeq/jItPudpb
5A7hITRte89rFpkFg/VWLnuc5MEctO7uT/RZTQKLJOglWXp7f+uSlAE8dDm9YI/IS/OO6o9HzTnl
ZjoPWmmJNO5eEka7WEI14Wnl+k/UI8CLPr7knw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vcA6tVBzywmJsvOGZta29NRAU5c4+e//Nq67cIVRUCEbQtu/TBzGuVvmTJqBcU2b72sDpgdn6TWW
HdNlgPm1q0gl2L3X27zzFiw+iTqSprZuK9pz0e0O+7oFIGbnzvM76Betk1rhRGfCV3NKsrQsUZ4u
rDVDPXN7BJIa08/V/boRGCX5871PZGtOEHw8dBNIr2CfDxytdwsQYl6TPm+s32UscdK1DyJij6yT
56KtqClpqYfV67ZmyPtdLKDbmf+XaEr/i5QPah1raC09d1fb7MNxnT1kH7oV8klk6QbDqAwl7To9
5v+jCauuNWvCyX1my3fzbWm8CuK5jAU2vXrvKQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X0GXe4413l+ZBbytkXE7IOL3xzGFtpeplzzSs/s0NIrsuzQG59hJqM3d6liI4/SHNkEwiUHF5fcA
qPHT1aga/AfSC2fylyJNGOz0sQfh2IYqtvq5E9GT0jShxRibVeFndZ+Y3JIt0LKOKaJRH6y2b8xy
6wfF/6pZIu/XRu0+C7TwIViyLBIOEVkhGghVsgslnz5RcdCiMXcPgHGucu1btmub7Xd0v11aqvjw
nRQYV1gduDrGtNJFU50Dx44Rm8IdndMJI86N8vZpVgUQ/OMe8SMOXjkeT2h3y/ijSSOtaOGLwc4J
4FjK+n1vUWs8aoq0C7jQl8iaVQ0ALnmzBmX20w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
em7m0sQoFdMSKYlp8fNnnGHtha7+YDLScVsLXUfGGlxdfLt8ouCJKEWVOgI2bd9p+aNlNqsE2wgE
0TfwWzF8YzQRyG5k4D71zPHOQYn/Jz0UmLVWoRmjot05b2PQFE7C+HkI08wo5c05ZZCxl6GDqV5l
4gtb5/kTvmII6wfHYVw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jnQk15tdONqg9/ukBwbkokOqw7S046x6VLYIf5awLeVUFwP97gQPSyGyxab08piQmf8PTrUAKX72
uf2gl+T9YzH+MSUDS3lz9X2ZIxf9dJ952dR2W7jJmggGx1ffSB14bOmNaMusHDQuFAc7oIVIlV0N
BQamQACENzbxrEWdKe45iLSoK6YHZ3irufuSJGd0q0JgQk5V5ZCDAo3EeTV45HBV6fY/7cH8XdgX
13Oz8nv27TkWrLmJhkJ7DFi9uNOrMz165v4vI6iRZqSkOSjRpL7Kc10mXKFv7RY+K1N27WQyNX0l
GYRoGLAwwvJfLg9SAlAh9XgCAb9ZxD1SGt9wJw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103440)
`protect data_block
5zPymDwtcV7Zb1kCs0qBiGgd4EFt7k1mmYVKyRo4u1RkTgVSVDDoQzPhuO+aVoF967wVpAbCx3mZ
alnPElmXywX+wNmzIny9tBfL8R1Qi5KzfjxwP2vedwE/5sfSnlhGUf9OiA2OYZWuQtxquY6+iQ3G
qHNX/iPFYtsJt5HuLxzLfxsp1mJrqcMAYllUVTLU7KA1+3oSyr2LcqCc1v8J7KJBVPtGZ47o/wYL
F5n2GI27hk8pkhMeUGeneujsCH/5Drg5A+vusC2QR1pDO8c6Mo0J0Nmfcs4rklTGjJ4hYMxk/t4M
18MLRmXrK60eTyRaJCZlP+7NCjKq3w0HHEqHBkwkLCoNFBFleCSot5bdidWGmOMQAIY0hQ3VUDNJ
oH++878GFbGPq55ZYwerYI2Ovck+BfFtCs/vt1Iuck81y1T6rzrJqq+/+zk8VfzNNOOCGDxjT/Gr
ywpGKP7Fxk69wyQSXiuiNOyxJfEETAUH7h4m9SxUIDcOsug68tx8D7vUn9PpMuao9L+w1qkl4gkK
xtgzF6yrAQLPB7GpzoTCV5ErKo7HPaEHOtxulJsIDJi25EL7cdOxclE60s+vcuy58XYtSIPIsnR6
xFlP+x9U0Yr47iN2ztzNez1Kt+jcIKyTrE3tSzTtw1RW30TUC9Wf+tYZ2JHrA4IUHBUEY2iF+b5z
yHoIo9lxkCLz429kRb0PZ+FciKs2KiukkwDEUcu/XwNcRXFVogxUI+QHtkj9yjmUJ5dSMnD5WR24
Xni9RtUFSTROSeI4zs3pAQa5hrj2mUgUFC7AdvgoAnFe2rRH2Ld4WvEvP8ghilrAmPUI770rqdTI
gguiBF04ijCw2qLdPJaO+fWRdfe1YT1GiIB6pQG9M6ELd7FUejQlBr/nsqPqvYNHsXvTJnSbMamZ
bliHtoZF9qaS/oUAYkZFPqgTJWMKSLV32p0DSRNbdTPSJG3Mi37YlHXKIpaiIjZJJIZsV7S7VmmI
mUqjFAObJzDSNonBeguFrieRPDswVg+Ak5aAeq5HfLp7ZXxgOjHkEdbQz3cCzCybKERmZsVtkiOy
kRGuFMZkrlMGl6aDko0PH065DnyjFOD2qB7tLOX0mkTa8kcDy5grZWhzZVtFl8BnevRvw5+YZ9Ys
jpSlFoa+1/RsiWizq89unSKcIBRkCKJrl058uOtnbDewlGJMrwoSDDYjFXVJXhfZ42NpidCdBv/u
uS9BEjHVg4NXtoJfiFIAHtGaEyKhnRz6Zk51OW6Ypzj3efbzh3RNVVDOSJpN7RetNQa8P+IP3NEu
U8/7uY/5r5CraWKrYR+BFI3KGLdTKvZ9Fr4ZWSa4Q+Qdb3EsQdBojAyqijoUxni5PSD+28eVPzlC
g/BdKj1W8trw+c3JaHnp+pM+kjJDxnuEr/Dm2SOc8cittK0/9We0BlAgZ7xCfs29ynkv6JSCzhHz
Ng6NWPAWgXIeKO2R9jO2itGDtzR4sjTOiSIabkfLRMXdblostEhaoRamQvvtx+ehd5JQ8oGGcaDQ
pSkTc1x2h/9fW/f+oeYe/RcS7/Ezh7goDaFK0A7PEbdXFMAk+uKMGqjYTT+RLiFVMpIe9SwCtBr1
sbDJjD06my6gGq/mcrnNbdxsHo1TN9LlscSA4wMdT/ZcAhWNfCBcIqVWITuXoqEmohfBgsKMttZE
UhW1OUdskxflCVgWSBEK2rEtGo55lQh5yHiSigHVqkSTU8o+oMZI2Ulge1f2JKKs0y+nn9rYLHzL
U3dXFpZIbgwv0vd8JD84YHWZMs0ZIQKNs6DOoRgZe8Udi7KnfokFfrW+CtZ0zPNekcrOMpWT220W
A4Ss3a/9v+U8CGTQbYrc7iiCzZkAkeI3Tj/EdE6CjFsahOl4GThhOK5IeaZVwP/ASmDFf/sa+tfL
kIZxCAw7bSzb3c2Y0e4x1JYI1tcn2e9BafR0Z2T9OS/qRRmO+D8cTcbXBiPMaEAQugkpz+daBznT
12VvIxNQtVvI/6fuNB5xD9+iSS3aO9ONdv5UtF7NJn9qtLNuRGvHJSSU/bFfw0EY5GxaDIewRl3R
YlaAIP2g/T0Y8ZvWwejegEgoPQ75vjDKvrbGf6Csw1pwrHl5Qm2ej+EDOyIU6r/JfoUwTWm/eNsz
xd9t194ADxCK91nzJlEjWx9L7uEE63YNVCotHcDNf+9A0fx8aZ67FvGg2ofSJ1mWfiVYUPvy5q9/
DmhBre8MEjVoSGOI2p+cAKaRofB5kmCVV4c/YAafsCCIe8lHfAWWUUe/T00a5pXGbc/8JxkcEBSY
P5L1a3SqfDH9Ih42HZRXdVl4irnlAcmv0cIlYwLFPCqMAnQ3oPWYygGnSgP/GO5n8I+5WB/i3wRd
jmiUeQAh1o2hiSPAa2RjI95XpJk1MjqPtasf4nJa4uIh45JymxGrRxcZv5CflrDsge5b+WxpphsE
UJ0Q3JHMAEEYntOoo3lrQy/2Jj5LNk/GKmBDEuKPcWsBpm1AKryyL0WVZktItJrs0cB+4zkqcovT
sjXoaTUj1Axufw5+8sRlxuRGbit7kbG//MQTGx9T0hR0xLmK52DjC9jJVnJUB7V4e5KzzlpojWER
fl9QYd6mkzaJ/jqm/P4rDUP7k0YQZo5Dp+seW9MoOZQZQzlU/piji3AeiQvjXI9c4NepcMebsgEp
IQ6xmnpZxyCB23h7TT6hMwLAxiGEGP9ukHSuU1NuUOA9cYUybhxs8ZRjihRD/W61QVS97dxEyXUO
VYqWZvW1ql5b9ATJnvSHXOxIYmB0jUx528RvQ+/1W6QJWmh2Whd9Tum5jfhxrbEMUNTBYU5XFnpd
s4oEcRsX65I7e6q1N/B7Jx63nQq3RGqvygimhXCwTG2VhzpU6+qpDGBv4dwO+O6MRTLTPTsPW0at
fbj5DZxzgwDNbX/5Hm6NpUb1IQ+d54CzLjWBP9S0gsU7Cq3E2smjCU9hR2QwpJRSYuYM9iEm1ghw
7fyciL/gjPX3VRbGjcxqOPrZc//fSzqZyyYrIvwOErjvZzkScoB+MfjIBmGBqz2dkdmW6xfw4JxK
tbml2P3Lu5SwvdiG59640e4y5tL5bNcLHSpmtW8FIXM2dv0YAfBbPvHO43AnFVZEi87+fXHWpwfT
7bBeJIIZYWS9cDt7Q9KQlUohtm2E+FvCgGW42ifKi6tt0hrTmpz3jGG+fNWwur6JRPQ8c/1RVBV5
uUOplNdZ91zHNfLZje/i2TJN7VIPrIgMeHGwPXzmUsbOit0eOGBm8desYTamG6n6PVkJOD8KpGgy
jPUIXy/43PyCXw0hI2WRctaEbgQ+eX66bUJzAeg5q3OZNEc/ha1pNYLsFN7eaS76wUfMhd2PqJH/
sPiHARPwk6l6dh+GI/BWJ+mxg0ANEOlL0gQb3s8gmF6Qkm7QS3KhwWxVy7Cfh7HmGwLG6BkF5tV3
vO7rLoRIInEW6xuUDYCwlQRclcs9iSkc5sKSj5qzKZQo0R7CNvYG9XHnIf8e61c821XtTVnFdb6F
mAHKSnwH1yCj4vb75431KUf7/u2f4M2GEKw2BN3Az3BGp+g8W35Aur5Gc1pxwK7VbPIDgxt2iUh/
lRwyqOZtXgPlao8uXMNUmkvH8F5o5GMoTLNqTLGuTr5/jgoTm8MxhD8qXPOHkCaNktmueASmJ/Z+
D+wEZ42DD0aiVOwoFWvBX44P9rF8nWFtqszObXOpNoEWEmde/GXP4wHgrjLTEXrmruKEKCpC763V
ATSfLKdDou1jn/HpKvWKZLTLqI2Je1Mqs31uTvPCDGd0ud2MVfwaU5WNP7F12PadJgPx4yXOc3IL
mWC/ixfgye299hTrBJ3CgS5xp8wtkRIZcekiAS9nUUwhGJGpeaFrduvl0txsXgb40tnaT8n9hcmb
rmNrVtPGvuKiw7k5cHaQ4MdfZ4yzDBZIvmoiS5GQxTYVhgrKVr8psu7cDFJAhefzDwQua4H/0Urk
eis+mXTtbxYpAC9TA2LPJd8nat1D5fmdvW3UytMPNUnJQU2zxLaHEW4pHLHjm8bLTBhq7rQG2z9E
GgeAx7zR28yTFBZWmhtrcArU6BbpVvGYcYYPt0dMvz0UdtakM92l/PJB9YyQHmA4YPUp+HoPWNFV
qC4kYb7SRfesXZx5ZzwxBzC/aHkTX1LSNEd+F0gapu7sLFjIAhl0nIt0unYnfE53sZhC4FyTUJSP
c9xNExxmxpgefmJBWKcvaies8FqzHponnPaERjcPtJLcroYuRpjXS0MNTYA2rt8Vm/r1UFXepJya
m7s7ExbS92qXADNdIgn6SPsN4AIyggPFD5g123uGdM3BUWOuyxTfad81rosllyxc3ONUfXBHYfzT
/kT0xilJmDwremy4XAUp2fHFOi8BPDva3YfkX04MoN7cKF3a1R3PrGz1Pa+SRraLLfGEUj+qbkg1
uV1DasJFrnmqESZgJjnsdl/RFFqA92P/1OlJ6f/vO3LJo8MetJuKgASntVjyXZVCIm8Y5dzLl/j0
lCezc/1XhSYvscOYckzqTlZvnxx6L3i7Jtxfy47f7vCQlaT1ZeRftpV+Qgou0MeyeyAYLW7y4ThO
fmXSUYLnr40AX/4Zq7sWVe3IbYQezG+FEfVy7aikF3e0k6pUAp9KdF+Vg2bDvKtR58ukl6xbUBlH
OkTvnrFOlFb3mV4vG4A1HJy9wFxwXQPnN/bYsaY5hjYfzQtFSM3Gxe3VzhQ2mTIlxiaSwDYWG7dS
TExYwmuUNMWmzTrjUfjTvqKbW5VjyowOt4ELgYvYXjVSVQlsTr/BswKTFun0EcGSwA7XO9z+Z3vl
mTpHd9KA7XAt+cYroMfqJ2naQujQuRldNYEeSN9ZZ+0oUpQuWXubGhD53acZWfP9OY7/rVyiNpvA
augPILGprcx6rBcBnVYzLzGEwhMpjEUcPoz78hzdU5EpubWiKNafTxg7A/hQO5PDNN8gWvYgAIgM
c83lonT/FykRGwygMf9aLlVGapr6aZxRJcrYzSUum7iw0+mXeFKZ06sxWmAXDBoTSmAh9Fpj+1ds
aCvEuhAeHTUJPYSoV3zsLNTQNrZ1Toirejj9kNldVdGyXhlcw7ypF/h+BnkVnseaCS6ChYMmIhAw
7eW3NZnau7zWWsZ+J48fNLXm1F+KyOYx8Sx7xDrPnk0Ravu0X1KALzo0Qci9f0jXN0wO3YDDBX4S
gyYS+NicKdcc/OitlwoWNBNe6VUrR3K8iEsE5ayOGkn7/qLYRpde3J7EVOBEv8raQe4trFWB2NJM
ryY2dHK0giqID/m2OcbieKPtiHpwPNQ2ViujaFTSRUfUwAtzsUxmosn60D0/tqpY1M+056yh7awM
/x4cBC24qvyT/+bJU/OzxHUR9nxbZZK4XuGp5Yd5BxOWum1MqaNqVZbiS75WhpdBVdcx9wvny4ag
SJEN4shJTdFtcU3zOAiIMWpA3F/PZZDM7KGNKBeb6c6Xbgr3MF8JOq61tP7lB/+nLjAc7HC5EHJj
XYn9tJncqwAvsmDV4OO0kCdujE0Q/Y59r9nKDnh8pvBmOHotP65WN+D/+8qe7JpF46T7xjXzEE9J
nwT7HrskKqAgM79INUn7unaDg8xmZ9l0XmInJDTyoKVGakSv+I5kRG/4lh6n8HSwjMLn09tzujOT
Nz+7Z+Yzc2m3er9KAy7NCpZPGJosxZsvYF9PdbcG90kK4J3DgOHZtm2/elZ/MxRBXYbaVTXPd06u
Us/HD/Fd1Yrl6katy51oKnslXTP0UINxGl89BfPJXg8EcshVpIMyRDbpaNEveW/Fd110uwpeO4VP
I2ceiKa19/mK1aHIG3hLh9HgnOjP8iCfF810R+CTIutY783J49LLpwgPuabyzIPMbTAbxIbqrkMV
5Lwzx3e0xmTktt5kfy/VglmjSwfJ0N0drUvqQQTomk1fmNE/ztlXW9DzUpKKQG6y4u/kQe2qFYAL
c9aXfX47lY5hCgiNfb3VOHf8npOBbPzhpbE61kB8hVh27t8QZsCx/cYNDEz3SnrC3mv/W81y/ezC
ZxHJ5PFqWk5ssEKwAj62RzD2jKYGQodjox29GqwOUCPpgan6JgcyQ25WlCtkBsiwYTalKH3QfNks
AtWKUXlhcOtCJ8HJJIkTSFa1in0mPZfT2mp2mJsvp7Z+zzEVCHrVmVptlMPUUe0hehG/ttYUS6Md
1CLlVMLUNtMpBjuDR1+9PWsi6WqTnbVwrgEFmL/LsCP29msLiA/vFmbafAeWoE/sCpCDrdOLLluo
qbYTS8prJqiLWuFxwI95A3dKfK7neqA39fRNOotwDarmRuRD6WAtmGfL97j3G+dOtLZb4V7dpwlF
9ZgVvYes+pvwVwVnlEXkirgpJQTluwz24CgweRqYjtcQy00/lIP8WesZ7arIfHD5G1UkF980TsU4
Qwmng9yb+7cZBBbPoeQity9DrBj1aZgtflPq5EvNKPNXWGVBo0zKw5gcxpdADTRI9X+ehDM4xfIl
Q7h17P/qFvgwk8PTmaxxIf2JTvvujEENFxx94siGI/eAimCkBaGnKtNNUOg8RUUSq1Bnyc+ZDPyZ
B7Zxg/dpU/k2horpdlgnY+pP4i0OPswUb9ZGOCyj2xfJN+mQn/EzvwqXmISkriBtKV9BVvy6AlSK
Rtt2pICfFaNAofRffDQIlqYjeexHJ62/DLFABptKu4ovZvfbijlzEODC9jVi4Ol8N86GgsOfuS7t
aiEmgf9Hxfc7FQvJY+aeFpjnRjGDkqCY3xcpv/IEQwgVUKD8DMrsMNYI1/eUwqooTush5YjGsXfN
uqulrpRIrll13byI0rNg58s4tFgkPxPm46PlMIobGs3G9slJcXBxc+13mSiZ6kOL6b2i2eRwpB+1
vTUy1MwUShnwW3lur9PJPYpSvztrjTizHXTXcDOkpWalX1R4JckTQ+826c6EjxQKPp3nIkb9mxzo
Iv+egWlIEV+1qvRZH6NnC+RFEaD0xTd+esVWvzjXTdUVS3/J+X/A2tabb7YTcILH0wLy66qeiMx4
V2dAMCThLC1T/Xrr6plOteRQbr5UavsmzsI/5HTNHWmyFIOTqLSElSqJeRfO7KAR3t1Wpa8VcQFo
hmZRpLqyyMXW4M6PSqlbBJIm/JE2FIhgMSG2RmsA+iSsYDIn2t4DHCdEqRonZJTKexrTwypAkiYg
/3BO+KVeySEIvwiKJ3lGpE1Y9Yjo9WVD8nLj5E67KsJ18H/twm7yAP+AblhEf2G+p+5IUQV635Tv
R9HSFWs6kcsZieG51OgW/R3HpBu+gNoX5NkWzQU6jTxgwl8OLTYInp5aJ9jnW/haUXCOjgY056Oa
cjLNvHh/FaQ1QBKvUu4rckGQEeEjJakxdFIFEmPvH4snVX+gF0JgSCP6ZY+8LU3V2egCjy9xOEM+
exdv7j4IDvkmZwvLNsOk/2Hx5MBgU5sBvmgJcxkvwXVFRy0u+tFymo7auF2HSBNQqaSx+XzPFFmU
xVuDLWVc77ya3r1NwHW5UqUQtwd/xp5FYjVPHZiY6+VA3sQ+m72W57qXhs4ZtA5RvcpyFnttvX+e
K1nnhKdQ34r1n6RSOqs0lz0kryN6lYTmdZAs/kP2p16i0R3yRPMvpGs8e/90OqGY//yJp7YVvkVo
CTp53nxFFmBByfGbi8Gw159wthmVpEhvJjr5FZWLVbR4iXapDGPkj/rQbdJVFPJ69m7fPUn8gYcW
b7qgS/Ig3fsxNd8kKqC17rkCMsboF5w5gV/P3n+oCeoi0VnPj/0O74e9Pm1XNV30P7Utxbp87a0R
a1gwEnlDW3gtxlcffoZFF2ILPsJXp+HJNzQGjhFC/8ywsniVumBfKideCktRrFFmkll1lWP2xrzN
YyxSnQaX9B2nq747Bl36tV9zGsmsmpMb33iUzdQegpJQqRr++BGUfcnFAFx285wnyjyN/1nDmYz6
MtcLvsgHRBgw4/tLUOyL/GylSe3P9/Yy8r36+W05+PnYr4SuvSRpFVCrWlgatvqQi2ch4bOY7thF
e5Kks44xG5DIVF0OzwniuRmBItRiyk20aWdL2Md7vN9C6dAfbkAVM7DfZY+ztatqljspJuDDuYE7
yxcE+ecWgUOIQjOjPh9w6W6DbdO1vj49O/c17GYAKuU9B+91sL9JxZeOcltJhUW9vt8rUSfAACDf
sy4pMPZefj+zX858cVVuV1Uz4icpdVV40f6/pwzi+Uzx50dIIuPOQvq6ngjgfURYfGPN+Hg0Q4EA
4LsZNmQSgNI3gxrjEqi4AWyzMvuAJjzWgp7pEsdwPkFj2GbELKKZvUdPsgiVlp2lOJc//iml+U0Y
4bNPiaEBmi7Qy2HVycbthq1T+4TgvHy1S7FVr6BM6F3b0uCf7aDn8KDSJ8ZpgbYzcPOPfPww+2oG
F3RbmBD+sZR2dK3DyellHT5vWl54S4U9ws9R8kwmKxs4Gn85EXfOT0xxaDe5O64347yKq+rJyG+m
/SaxLW35TRSWzVxQp64DFF6EeryQEv79wFIaFXT2zlw2i8d+HrxOwfu9zmLLrFZhy3y1hbmm/0Aj
1xFipoB091zR6ITXicIVSo+dHMILqNkDeJiVTGmUMtMxHwJhDw1y52Ygmuu/g2zEYnZR2luOmFTX
O4BoaJ71nJJPoAmVEDbKDNUlItnsWct0l5eXesEwvGD1vU4jWva7COgs9labNRK1+zcP0T26JLe3
tYC9gU3C75IYxhk8CJO7va0/w1NHEpBstgcJGtOTgQtDHH9krX00c4oKd1RWTXABVW9LS+0xNjAb
EHzBmTkQR7FzVcsUzDOvFW/70niCUDJ/kjYCxlvVTI3dtoft2PitLc5UKdLPe4kP+3EgzAaFcduN
txacCr4SZyERakoZEnCOFPdw7KAIP7zB8N2DfLeNqh2ti2Ecjr43IPGcyG6Ubbyzg3TKgWsxkG7j
angZ3YNq5IftSC/PtxtZ2i8U2aJFS2JMFp2sGV4kreGcDsggz9JpzD4PSPFua6JI4OEtyLgXAzct
fMC82tDSPe/wlhHjQ1NvFx7QzQkxnQsEqXLjS3Er0fWhoXhNicdgB3Mqf8Go/ggnZp7X9LUbra4f
igxVd8O2hOfibOZgB2dMJjC5Kwg3kbgeDMoscv5ePcUi9Z6fmEou4GG3VR8938nGYxtN+Swg6T4p
7OCQpvHZcr+j7NrXFiwBDdXxIjGz0Ni3Sojx+UC7rkeacxDAobJwZOPtFJsA1MPvtfQwPvF+TnNU
/8XJP4klMTXz4joew+8xmhm9ibfCRtLG1EFTmBzPf84RmBn5A7leV+pkRPHnm0nuT10sjvmbKql/
gGXNkb5X1wuW8gPM3pvNw8d9POTqrn7TzazFSfFrBj8qvRrRUjNF+p1FFil87pwZ+v5Zo3f4Kdjd
75J+a5901YPJ0yIz7n2Rq0XuudKqP3ITwsO5llq5Rwl6hqcd2Kf0K6FcDS5k9jJaqNSzlHWzE3Mn
XinPGzTTUPk/Nwk9zq8OSJREq2Q6WaGC+PA9RUCw5N10BYauWVXA1aCUyxa8wRmPIyWuUWv2vEl/
xjOH3roqFUeDjHksXnkDc85KrQHr6EVLamNt5DgH6vrpJ9DrwvYh1Yxt8quKt7jharHwIa6Y5gpd
h2LcH0fUCxgtwqJ6B/exzEwbZ/ZUaNqDohCm5d2OuA/b6bOzEmlVLDHi9wK9XJFlyGgoushuCMmx
x6/mDhmq9p7sTujN+vHYbmvg47QNayAWEDLeusVgGVOrSWZWhA+5GSnI3gZ4Xa6UjXwe+runCds3
O1cJlClMxtEYg3TVokeg0YRF5ZC++n6nEuoEi7qlcYU8ys2RGKT47kqkA4cw80+eW6sEXqVrxVAF
9VcQVePk1QJas1lU5rQWL/aGbu6RGieBx8a4tW4JbNppG3Qe429/jmx1bBHhuaZqAV/+CoMOUygq
kylD3cvLrNbBhqhKI88XD1V7dyKkcFkUAcgCvdlbAAklGMcOkcY1lNBoOf0wM7eULc4zRUT+rK2b
Bfd+/lIJgDd5CeqQ9BvrgBBS0dxV+mKNPsOvgv0ybLsl9tG4vfv3ZxzbgRHPLpgeAggeynRTeN5z
f7U1UcqhUTfmHEJqKhAOj5pXttV3eu6aBs6ZNuluiCoMTbSEy9ynuUWiHFHieli1qhwBWVuLueLs
IzR1lxnIoBplY7uMIMvn3Lge+5XfzFDr1SOQ3+7ImGYNR8pDLuK+KS1Uae5szi/KSmU41gve/KsN
TcT0YKakZrvjafGiC9kMHU9vV0Vv756Wrxqw+yesS5BO7CZNd4CJHD0GZvvQeQIc4RC6lj+I3Wwc
u8Jh+5qqIA0TxXOqk3Jx4JmsXFcHDlPIv/twv8f9Kmg1XgFw+Mz58J5PkohdTd+CR/ZtvZdDYUXA
ntnE4Dcrqwv61joO+LRrgt5jGxO3SFXV+6bI52boF+Cii/xtCPsNJcbcfhyL1EY9sfpjDB9fuc32
xS2ey/T1VeR3h83uBMiVTwrDXw7h+xh1ljkNkneudJyiZVjMY4xj4iShKHU6F1kfD7LDXH4+jLsY
4jRiik3kJxGj8p6AXyDQNLZUUXKJIH6H0otHYjZo1dFPim7HOixt/B7itIBVgR3yZ32ZrbwGbiNA
lHuQs+zHkfmMOauBwVXd3Myz3pepx2l0nRNH4Bst44a6Yfa3SVWulxeiOOGMPbvkit2MHqzX+clw
8otH0AaTpQS/8j6EI8nbqgMlPnqLQK2CfBE8ivfcTrvxnhShL4YKZjAVC6GmWlUJVgsqGXlCvc79
eQjQ2Ab7pcsG4lKMWNtfbCQeqqB05VDhKEV5Uoxl2v9U0Wm7a5spaWByotoVYhPLSCjMGXPEY68i
yqkwncugoCsUQKVff6MWYBKcO9olAS6sL3fbI4ZhLc57PiEI/bImUuE0i0s12uqh1169qsERVswW
SPmw3Ea+rdnDFOm1UVnpquqHhmUOgWY793Qc5GXaE74504ioZavSRosUealUm/41s1vLlJR1+I/w
8NloXRBdn9utPCVKTAZmQEAGjTe8UF3aVxZ+WksuDE6NgfoPXtNVIeNDdmfkjkXxgsADIX3XbL74
NKvpXFpXRwD3jZET3YIbClhzNiNkjT91bOQdISqaE6gS+JVBxuMjaITHYctrx4oyFL89V2grq093
eWw3bFlHu+EeeLYDlgQbKQC/I/0P+ZhbBuV+uHz0JT2b23AoerFgAPa+32qRdFHd/qCaacZQSYgM
u70ImlNZshjyyX8cqt3tYNhT4/igBurQyJ1q5EYuOaUkFfNptDuOVD2yDINKYlpaFetqzMVI92by
PsFd0cixhxH+yrZAJSnJ0y6LH0VmzyS99DyqqlAcyzwzod2IyotH2swpDrA47U1HEOrSbWw38w52
A7cZjlM/2Y3FgNWG4aymZuvWHb6Ync+SpgeKfUlTwZmCcjMU51s7n7zjKLQNANAzM8I8TfiTYMjr
COWdKa+sauCVF1Q5XItJdadCtgF1XioKtSe/allUHsgexGacD2OI0SwGhNtUQS2O9SwGW6yKcqtR
rMRgq0ycCgIhMHkzKaTlQOuj0ofivvvkL5uEe66AmwctlijUVzc0tfRtk/BcVXcOldYtKNxx/21l
AvRq8LRMaCU00H5mRbSl8grA7Jb32IWXH5eXw/Sc2sCBpNasDuM5O3NrrjdxVG7nyS//3chWgDwf
F97OODlqB16zIqU0zfQ+WHicnArWFJxO7x4Aj6Y/7Y3Yg8KShj+vMzBZcDQvE6GZwVbyPCp/GMC9
voqyYjo0sAW1EQoYTcYMfk6wGOUz6FEBtjxkRMmqzHkoB1j0q/YvF+27cAF4FwTfCLMLbVGFvaAK
nVByRVFIQgZ4IznRI8Z7A5Wdcd7yYniaMJtjebx5BA/FrB0Qfr0ivaT/eNcfR356PVV8xcuJL+sK
GILTu6AC51unQUTbWmdb3s2kqeqV9qcBJwEj6/c8ny4reO1e0Y2e42QXr7zC+Iw0h1XRdEERUFGU
gmmk3TiH2N65PPjNMmWJrXLWRkJUeaT4soJJtr9ij8sj0l1RpvHwSCwJpqxTcDqWaKFBm5a1GxXH
HpomyfozMy2yp5cdO3Rd8wjdXjm7hh6gVishMfne4WtgPaHAR0q0x7leewCp6hJiiU1hVJ+xpABq
xC/uxjVGdRqf199ph8eda2NFTiToPAF2gFuZ0jxl6l+e6ffY9BKnU1lt+R8/VlwkQoTq3qAZLPl9
3INc1c5sNdnFFE0wq0bLNaw9l1WWHwT9lXhhmOFXluCOF51kOhmwtk6AFw9R2ZM3OSbf1SKrabWn
WtJ55AU6h9acOvId8/1lXZ/HIhSQaely3fVj1GCrZfEn5Il35tXQch5DITVDBHr0GxSOUjajJjfR
u4gYUbtvP2Tdmuln74RrjC2V9q1MQ74pddiFnv+pAkOHBKg1nVTB8yYe3H0gwTriRi3Z2OlGLbBM
Gl58++AHPwPARz/g+ZcFmMgf5gktW+gVPdfee69i/dl/AsTdYznRmXFA+XJu/AQvVBGnB+Fctdjp
XBnOJhSo3hPqHfMYazIEe816sXh608ThOgvVPmCR7J1HH5xMMqW3Pb0t6sdsr6bR/H7llgwCR7Jd
SQ2ujmrPoEXwt1YMxmH3EZ9hhj3Su4YndZZEW0T06nlV1ELH9gvvLpV6fZpR0xoUwGbYyYM4m6cf
+JJHUPnntMpaC014c++Cn5N7Eqdrn7MDSpFgdJIi3u27TJEvZORlXNYGfBFFEzMRFZZaiSxTu20F
Da6xhwENtUQidOhHchCTdvDZBUdP0W5ryo+iBkRj6bi8DVJpj729k8oSWvsg7k+uWDelPfNgmIsr
yr35z4JrP1dSVuc9oaK7Ugiyyzi/TbiudFGXUcDK5vM+yVbBXgaGjFDHIty4Zqpk8I59g0x0iUJy
EU1KNg6wd3M0ZpbtBuXwGeXTBaQrwShfWT92Wj4HMSBw2CQ6M66x/gbHTJPmk4+0TLjbpxXG9hTF
VM0aa4hpAuKcnuMEYxfk9dhPzGBS0ORu46ALdz1ySFnppSstL9Ts/KVILqEMi9tr6LoBFucXxuIm
sRSql0NS73HkqNf5DiX81XOE+pd6BLN2JJ8MjxVrVmx9Ar4Iwz06mUcgxRsNI+JgNvEIX2gyFQcg
isGXKxycCPDk06tgRFQf1dNLcFzrlZzRxCewfhJDKTuCis0e4h5ZJSPsHpwXCZzne8tPeQ+vD3S8
5l+/PPAg0QbUIsdFbtEEoJKMr4X4qyCvo1gzYdQrgeqOMURKN6LfWGgcpzo9S+QbQUVLnVmwMq4L
4xdD2BxznSCU6+9rrhhAtNvBAYzxhAFxO64jSNg7tKugkV+cRrDp37dYid09RJso56n8OXu2eTtQ
O7RZ4b55OJuUmv0V56pY6HXHtLwCy/syJ7YOd+mCBFagmutbz1pDL864TpyP04txqz7exjecQg5G
5bCN3eu85JgN6r8nUggLRKhZJuSgVm8s9DhM7qc1FNI/V/9UBio2Lx0cUGw5/8dyaPB4iD/Tw5MB
UaXlH6EPpZyT4hl8MVXg2552PJsTW1Z1wBa3FpFVEAuVVBDouFWVn39jwgmyA8MPg70ftQTlVSvK
Wm8ww/Bhj3c/gzBqSjPefeKB1jis6nYNX4t2W1yKaDJdcDW8tq5z627/eICww/L8DbzNhQj05VMu
gaSoYqTZREXP0lEX2ShtqpPTI3CRVFCg6mzyuz8dfVqUdBejQN6g/kYMaD8gpxPB/RvPkGi1908L
lzGErAjr7s7F4u9YQdyqcAxI6U3mLra8Z4Nl2FIrGt2j5MVJGsN90VzTv5QQm7AT780hp/Cv9cPO
w0qziHU9KY9M8MM525mxZ/s/kRkuDuv9mUingvECY1+y8J9USmgWs21Dq+q84gxTPxvN0vnLRVuS
vdrHhzg9sLaAhGE2Jy1RIDxASqCS1tOVVV1kDmZ5SqWwboNznS/migbXfoSVRE6lSRu/YRFSv0ao
xu9P6C9c9YZfOaGOu34FBZAXb9dPysa0Rj8dk267Foa4TgJ3BQ+aQqD0HeOg0zTWjoCr/PfZnAFd
DaP5mXcKu7uzu+fW0eBc5eq7Cb9nwDlekIq3+B0zv9i6IHSAELZuZta0HNDPvHCmsyL+iVTCAdVq
NENGGJQKd7JW4WpMTZziYcLEocLb4DNYEWbas+2DiA2O0yTraqichTL+9OtZoecpzQAgRLvcdVPE
S6ImHyyp5JVQ2IPFsnjj4108ct+VimqdTV6Wl0z+XlgvcP6mC0gQs3GiEhE9pXfKcMyxRR/xKs/E
gw8wgMVANNltaaWdA5NKQNXXFshKA+0RDP+L7ZaHH5YWuOxM2tWLdlXq0SYBN8iz16c9uUol86dT
G4Pe1f89gR1X/+fnYe1J0V+Z7rLWx9qolSGkSMX+2PsqH/ZgRwAWhog0Xzy/RRx+M3kMIM1wQ2gF
KJj/GaLmgvEjgFm+v3LVnkIS2JiH3ylmZgz+EuTgoING3SPQZcjlNuT8eyXWAAKhEv6U05DH0tYy
0LZhOLf65eLZTXjsRkruX8We4tjvcArz+Ota4lITc3fBHfTXOX6EgNurQFdeRevdGkXsuSC29DZE
BaMDMJMrudByIdTlNbn7gBSglcyN1y+oni+t3GXjvcI4+Vk7LCinjEb/Fo7S8+PxNJWpbw4QU8bm
ESaZGDARP6sHpv8akGMJ1n9oJKAMrEyDHssdf6t6Z0rqE5Ukw4/E8g3QskOZCPhxKsn7eg4q9yNI
wheJVSx2ZVDAvn6LaCOgDgulRZ7Y6LNVHIQAtz0GQeW4kDxW1d72xbsATbOUwYCMcZ9WPZMQDepv
bYnwSTh5JYrNjHo6R9en7hUJfPiWMhvMGHF3koooT68IcioGuXU3qnnymMs50bji3li+olZf/MY1
rc9UogpMzIzqr5b28JYRvkQPfW3iD5puBgpgqf8IwgNg55jdwK/SJ75SNiEdjPnI9AFHu5QkHSFG
7gwTD6MLBAw7y8gv9qOPIlxNzIxXdNqDJ/F76B39TWFbAKzyRHoa497FJ5Z9oU0w5J7MjBAyUCY3
GRyMjayeuOH7wdpqLAwc6cu2nB1wARfleonnSZrfa3yNUmDHQR7nRbV68p4Tc0EW73f0/EILFKxj
63COogNrJeMCRV1SmY0YsokDr9urGs9IOSNCoAVWeeea/ASHtAfKvevB1XRPOb17Nq3pgtRWMfOz
/FhOxUVMNDFo/hymLdzGcXf5sBBJGnGtvuy2NfA9dskt/KTxJ69Ld8goxO0fRCA/0+J4NEa5hNY5
RE5btv1SYipMCNVPqyCr8Rl03LNxEwqEJRfodBLYkg5TL4LOyINgcmdGgeXwt/PvOYgCwtPcvvqH
duSHUp+7NoNg4cP18TkHWdU+KTToXKEzXgpWmOiZx9QH1btOGem+/bcLl2hBIttBiQdiG9uE5F6u
UqjTuOZtNeKVm51/ctcxFM82EQCitrLttCYHWNK2RNY4h2zVO6k3XHkB1+yDE4Vd3fEmVEy0fYTe
Wq9Sb5DQLN8B5Vl1TDL4BB0AjcF5sxqCctnYxHufpmmAjiRQ0mvjw3d3S8BHmNtwdPhbCL0jKF7M
RaxHLsiG7++9S5FSE2gJEc8y9yxNR8z3kbDgkrsMfgREg4j3KL9wY45IeVquGACNN4Tr0u1FP6eK
2CgHwECxKOI9aH/5xLf1IqUXMT1lZBiKsUfLqrlQTtpKpCCkFREeRNJ+ye3M2wDMU2D1D9nRylWs
6HBGuIluh3TpMf1LsJecPVGKIaCVrmGA4X46ZO7/8iEVfACnPWAAbcH7eK8aE2mQV3XpBsUrJdJE
rkQj7BGS63kAg+OeOywmFUlCNnkUe4dD1c9b5ggXG/he0pLsT1pyUHW4kkHwHYxc2tweNJgdtyBt
V3I+XZhrfTfG0YXOrXWkkNUd5l5T7FX+F0ElvI5MvHWDJZWfOdzgVc8Sk+okr4ac4Q3A8XNdW/Lh
hp8BkFMtADHlqZbrM28Cz36yw3vE5U06wUY2TZcFccrWEnoNu8D0n4RbtijXTjJoLMmPabJzpv4q
NO8pKsIcn1aKbtEfIKR6U2U2tSQCeRtiAtxk1YGva9MWvT1DSh4LqQwVCXAH3XMiJEWyHMhxyYJU
OR+Q3gyamxvQ3cs+5aSi5GZ+aAzZIUtbOOwLw1/Zubu13VFBRVPNUA/GkiOSEPlvpcm9mmKd0i2G
IrwJa607nbjqJRy20P7TiFTbngsaPGvfVMccma3YaiDg4O3GOG9IQQwYofoKaI5fhVUFXVwN2UTO
/SOqxPjWT1zgZakXkQYD/VDeeEYAvGg2uLAqpKqAsuVz0j49VcJTyIPIzzuRC9zNRV0m+2Ah6uJx
/YtmB46HWOzx9/WrDoFB/9E2lInydetGtbsgefZlYJDj0oMXHa4UuKANmv/xK+UNSn3diUMIdfOy
iU4gznNERVrhJfa9NjfQaZpvTJISJNwMPy06E0dx6k39zMoL/lVLeuVmcs4uAVQtjJ/0wiKQa9Aq
XZO2jW6Z9u2JHGutucZxmUl95t5jY5X+k8AfOP89jacQfPnWnBCOaEsvrjX5nWCXenoqga7Nhqpo
w0LXirJlV0Ar6yOO+J7GJQbxHReJgr2EZyyVL3tais28jEj3scNbZjD0i4xaMb9yeQB0WAv05CVd
WKd4VJcrealGMcP77/mgu8VAh8GDVTFNfwa6wR55g/gfPciGT0PBEmJ0Ta3m5b9WIm8EjMPYwaA0
u8eVTYFYS7v5knJHX4K8XhawRzaiDwf52XRN2cAjO+WYD87poLsPBFPrio5CW9hbIeFVQ/5oyuv6
G49d5DEDXnpMEQbzbgYHTM9st/Ae3mFA+M5XML9tKoyEhjv88ioKZ/90C9psd546AOtnEAapjGdk
OUMOwvUvVAv+FL/FiJlfybuM/elQQtUnfcFKgiVTr53EZJWelYT3YfbIGo6eSUNs7JnQIVgU56Hr
/vsCqbA6rEJzNXdN1Xc74zOjuNRKY8NSjNoN6WL2QXuZtNfsg50GhSe+KdXuGz+yQvWOhaLHU9pQ
GZxOYi1wGlNuW8q4rI21ib1eoRt6mKIIiN+wYBscwPBFdMiE/KrrNkmjdAQ8pGt+dA4MHBEg2yL6
Bu+474ohbE9gwZb0opxi4LUZCUZE5VSn7F6g03RI3dTKZVtq7azG2JBSWk4B7YrU9ucoia6xelNk
rf6S2iK8WJljSoUCFoFScbQmr2lj29+vVbV/TktwzeCybrJrjDrJhYhdO7ew9V/L4iPeIS/JGPi4
oY2kyCkdtnLK6AKw4oWQrgA5pdITvbpeNbOWQ0TbCULi+iEBqJhvwwFIw9mRHd+wCviMuWdNS3VA
UMZ1gjwLw9+cSZttvwZ2XrXsLnbmTYgWk038GpTVja/Kfq9aiPQMSf+O7Cf6E3sj5/Mgyr7vsJG3
ePbsI8cD4ADGqI3K0HT8oTIaE78ImdH9Svi2JsvAVKoKEUP4NtDmENKF4eZezZ+1MInMVhZ9P6Pz
i24DHM8/gYw7DNoKpfYknge7PRq7itKmNfbT47iQNuG55+Gb7f8tFcuZYS8Z4tcCqhwCwtBgwpZG
2zMkF92jQW6lzTj7IvytYZHmdr4x0ylJNpEVfEPgwks1TgZfOYSdhk7d+HPn74W8pT7gA85s7dlm
R5ZvpFEY6QNkd7pP3BVHBDLsTXGvh83q8BMLYKAcfMUzTMQDMtzPdztg1jv0Dz8t65K/eUhfCN50
3udLiPWI2if44REjG2YhQoN6WpQeWqUSLM94F+bhLo/ZjUDSzGJc6+SoYr/iPbnoJLOl/Z7s/MqP
K48dTtpvTmn7ZY2AIXIPT8W9D6Mp4pZCbvznGj542zv8a5Xq0d8BiNWVHJIldLj/AUt7fSrtQWo2
YXIJhkCBvLkKvxt+HtVYMWs85IETUttkmPF+F931/d3hcIg3jkZEWhjgOrZSa+h0LDF/lJzLrrKt
uRA7Hf3E7q+5d2hcloGd0eurkvFFZ75IIku+PuR9pAycwR5toQ5KqQi5vGUaJE1ZVd9s0+84CUPF
ZrIlqJjc9dA416Jk6hpBc9a4AQirxlot2jCyZ28fWsimnYEqzBap9sM4kuwBkwvtBdYfYHHvmL5d
u9voYt49djez7OknIv7mrrtFK3N4qGBJaH3+lS+nIlksnesnWYxbv0Et3/4qTNs9opI1BV4I4YJP
KnGrSeDuWZV5AS5WrJBDbbI4YWU1kVbvlhAC+5kI8dgqzxfdM336LvpJqaxoGayoapAgeBXWkrk3
xlNLnx5+c9uQsGJAtht6BXhWeCIpQjNutGOtt3c5hIec0AnyTbQtcmQINYWh7u9r53W1Hn316H1f
pr4tCL1goaFEhLTw64DtInTIHfMUQRL3bqW+T3QRuaCJ914vrXAXxBMU/L4teKAVjnWe1SotNK/V
kkHUWlPl8adHLV8F+7wrTOxHV8soS/rU67AtrdVHaMcq4Q5I/gAV2uNYoZHsPflCTQKeejefHx0B
aXiX0HB8BNToj8Xgqp5PrnFgCFtxPSFAxvPfKy+R8adyTfFw1/yMssuVvBVNsQ62/FhA6ubmaARp
rKKHhw0yFd/umSyx64bjGoRacbvhDJyN9cBMPtQC1AX1/fzbNwlbPIAUz/x1GvmpM4+P/LCu2RSP
94MKiUQVLBQidycP4Ajv7kqz/js1/VJgH/KbIrl2m+wBOjURruJLDRjyfGM95kWQjrHGBxquFqNQ
SALlDUDEmboZUkPR+PUCjl9wspchDhzBABiLx/buB6NNiaT+apMxrDHtsHpUFgNebBXkDlf76Ehr
cUQ8xdZEYkfWzMyoHs+d0ZNgtMmCZbo3IoQuhIv7NEkzkU10wPIuwgQv976NrZO5tARXFfiZa5kR
cX4LAEDCukYrHUsOoOrShUwCv7XP6kfcW/Jl8CUY/H6XaYJfqQXEwr3YTVpSrAZFdmi7Td76hq1P
qxanWg7lUnjtm0RKiyyqxTweb9HM4Wsl8c7fNs+mCSKAID7efUNWyx7mdDuMW4qyPI2B9O9ezdfb
WmVUwfYLG+iYSFVK98juKlCNkey+vbjlzsE2d0xN+zGXCX8hZLFrkNHCaOrDkEby7z5ntHSu2XRK
klC1s1FHWKeYloz64px5t8fVO4cb7Cg7qqJZIN40fhIDAW0LWlNLr+4zqLjwJ3sCl/8nUMCE1wU2
Xl3UZiHWV2mni12q1YVSCoyiseYMqoW3vPo8pI/nLfGql/mpI6m1IyGVah5ragLNqpoCJXyyqrz2
0NRRfpKGodc46w59hsyWvone5NJPIVNXNgIZl8xegh01hyFIDW87diWi8LrJa4+Y7F7TTcG6natS
u743rQ0S1kbk3UvDBkufQjiCxS3RfmgvvJBy7O1NcVRZpw4jxcNCgqzlQz1jykKDHzx0qJNjsO0M
/NbxsF1mb/Yh6B1mO3lHl1JZRBewH/uyS+TPqTLjuzCVkWirLkbXdOj8TAM3IYNb3xz/MFHyRfZA
KmqlG4nEHCac7PWPLnpwf9xkEK1bwghoMtcQBj41xyOIu6elA6cHKI6j827nnhNx+HtSNRWDwpF3
uP2SNszwKtcmZZRePMuU2mVdlO7D4Diiq2XWjRgMkeEvyytnLfJRiiGOpwU5sjLcuqcURDztEa2c
ogWRQ/p8v4upv1ySBmpWwXB0ubNfe81+PIDIQK98JcjDDly6gC5Xm71Y12L5+NCuvEmvfYBsAIcQ
CbsVrxI7V89p8tVg9JCxoeebLv6nWMrhbVzlfC5tGiy3UQ25jUPRDhMQeMRaIoz8a1WrLIx4etlS
JoHDb3yBTTtYJBbRI3x10WhYY35JmHt0CpuexbCQ9yRGT9vaJ9ecNKgnmtTNqHnFisWlKWvzAVfU
IhM2/MOCeRyPcL485XmqLQ0ocI6CEMfy+9y514F7S1YJAnoyC4rt6mtZWE5WWFBPrkUiF3roRLeq
fdEGG/T/vkudkRHiqwixpmTqGeJnbGnf1N056X649CytEfi2byct0+6yq26GtSuhFaHnBLJIVLAx
JOhx0Nbpulh08Mc+/DW8hxFSmgCeoFl/Rvsl7KfDUNHiNcQu+lV2ezh2dNrO8Tta66x/toTZjtTu
XTv1XwbkzOtQLUfi76iFEF2vB9d6w/rOUyuW9Y/Fv7APoDcDfqoVA88N0P1gl589Tc4AW7bnq58n
qu+Cf5IN+tPlgrr/LjFIIp9hU9GMiDMWOLcPYQlHHDHcAvry1vvr95u+jxYz0uZMeO5Jm94GK2fh
l4/2MuCvm/DdN+8XYMVvR32bZskPBftTrfMdyNl7op/5U5ex4PwvXvwToH7oXIrx/Eyi7NYU/+of
u6Eaomj7ZMAoC6FRHHyzsDTGqXy/UhLnHB9izHEMgarIepINtqCLFnqTCaGA8EwieXma2tWDhJil
4ACEWuE5du1tKFU0gEbLxjAK8jEBRTS9Xu42vbSlmuWhH0Es6Ax2rDTKctAHp60OCnnuk/CcmtVa
MCeJGoOnOji4gS0a0UvQAdhehLs/euJwrItkualz1i2ruZO4+1VTURF//gkuyd+UdPpyHXLb/yod
SPspyLedUCB7FdwLpUbB71p/msWxTgydD+gSXNZJTvao/xI5rA5VNhbybQZap34YdPpB2M7APZvk
0ssavr7SpZv3v4zZ1eZ1hGGe9JWXxX883teOIAyDoVauBeBEBVuxPrpyQczUJfRjU3KiumYavcp6
ZkeT2pBMrLzwB22rsPtcpStkkD5l+NhjZQAzJhopDIQqb9A6CnwyL3OHsi/7UPC8MSXEYCI7w7VU
A3Fno1SQ+v4zdTbLXj+0ea0rnVObYzM6yaar9HER54vk4nvbhHF2W7xcw92sbuxfZjBJbC4bHvSi
1uvYC91VwbSd2fgEFUa1XPjWEyfyY0gBzn/txJM4ZjvCHSOOtSLYovXFuTOL/lpXtNoIVRMWEVNN
9eq0feoLrGX4QGGhiujWvhWsauMgwl3I5EZLm1yo7ZSdf2pfRSPC80zvUSleCjAx/ptXaINHQyvw
y2kL6aew1gAaYFN7NgjzEzXN+hr2m2m6iYjLbcgM21XPbcJr98Oo1QIMly79laqAu/Axba5oW+nI
cJS8csJblx7FP+ENaUs7NELsAnuxr3EvdSv5nFcph280AD7+h1yEd58nggP01ayN4lzyVYY2BYoE
Xmcbx5aH9HDYTAZqHmRwRQ8FGUFZRgvV6wM1afi0webNdYwaadulgbNik6JZ7ECq3WiTJ/jkXddn
QDJANlXkZG/gOC60jeePEkN2SN46EajGA6n5wHUK1LWNJkoim3oxDC/K8ZSaFa6ERaxLB/TpuLwl
zTSohmpJXewc9pSrQeNy5RSr9ZtxQP6cSwelsPnnds9GGv2AxFUwE5P8DSCfKS1wjfusJbO0Wpg2
6x1ckskCbnK6vSCYjg2mpZWwAv/0G7D3BmJCYf5tx33fi6mNwu2KkJmr6gqtLWw3+5CSQiqGxfKL
/QmOjJF0wu5MF6+OXX7Jvs58cTvTSzY1aBAsC/4zmwgpUxKFNzMmVbH4uNsugrhTjkLGiBw+PzAX
JYvKzY+/YHk0/QGT4sDwbCnVJh2ml6190hvQYG282IEwracEOZm0c1Y+hMsu7lIydpTLNuqhwUeU
szdeB6a9MZbz9qLmEeovvIzXW3qDlasEOJwMWXZAtneXGX9QZ8D2a03J0hPEqVSbRi0f90WO/+zB
hlXQNe+3/m5if7tWSKR0bXjhjazwjdAl3NfoKKELnu1PW7vfJpRW9Og4mNHzQhwiJRaqJPQrWla5
HlLHdvU5MXe6FSc5EhRMutvs8aHnY+LX9D7X29cQFGh33W+/2ZEZcn5kqRZq/i4iudlMp3bc8A+E
Bp3V73D8Yb0ez4Faj487vdauM70/QLFOUpuvpn1qESgsmGUbe0CDGbTVvcdoAok33chGT1GS51Ra
lQphZ+xxGVx3/Lujhgv2eSWiXMRGe4K15tnmFFSa2QNv7Kf1Iu6v+XYhPGxY7EV3pXm2tT+U3x0f
hukRm8j5uD+b0Dv/c2rkuZ5q3lnywTMlb3CY8QW9JZk813k+69Bg3zAc/wVePuBxCVouX/nx3mat
wO6ui5+vnwsYRW6Fas+rAuRSM1kEqyIBMojtc077yfH1OclUymja4CCF2MR0XCClW/jZJomzIeOi
udZDxBHih5NQpK8uxLB2p7XyUf9a2mpgNIcqzncF9NkU6HkkAHPNqnqSco+5ZN9gVqgZmgIEzfvs
Rci6YwQXHAPseZpSnk0elUvODz4sIXKRFjn1RgpvJTlhm3/4+93t3J0MHHrKhqpRX7RsyGHkrUVT
CloFYuFImKlBYskupcaIzXJn/IneKyOGNvBOnCn7R/8ZxN2pFQE4Z48vkZ1MR6++HyNbE+qerFwQ
/0Pc4KSkz+WA0Mcz9lvnnLnUS1n+5FJS+Js5GnC2F/cMUithstrTgf6olPUCfgo9Em2Z9+OWQEu+
vd037a9PVDizpF/swzF1tEG3oINTD7kXyu9+GGctz9pSAJ0EhEXgR1px4VcCpvnnSKGcNkmp34YB
xzjfMfugzer/lV/y+3Plawa5YPkYUwM8WSk3qc3QjkmVz/UHzmGM54sUYc31/D7oqeNnmCna+n82
YXVRlpfpxEO6HELOmAPxqkZ75oTDZmKDGHfWPB/R3igzFlV+rnOG37kbJ3A/iVsH8LUpdpPtAWTB
5Oa4AL+n4RBx3PMtctMziGm8xXsehrHUfzAYHEJhxQVqMVrn6MUeLCe/N/eGYfdOsqbG8wdYofF6
brcvcXN71KkU8tDB2VMCy3BR2kq91PV5sgwwNdtZ1nilSHrfsEQ1NpmPujdJVvqWPAgL7+CVMrOg
ojkEIdC8jImM5txekwk9mHWpUaJXRSQ8QICg3JGK85cf68Jjc2KR2LKAQr9iNhQcnSmn/iG1Yowy
L/lQ3WM3O5Il2DV5MeynM32rUN5Cq0VSnu9rem8dCB98L3Jb6FdKZt88zQt04hnNINbhmWWteoJC
oy7Mr3/aIRJV0ZzJACCsrZY6yb2TSvZ5PqCSmJ9xE0q8HRdQhT4gl7isbBS0BxbFK/XBHUBVyj7R
6/JZjvt48pdZZvEIVatzXj3AEnj0afic1G0u+Q+WcDSti+SGP32BUJWeLQi4fSf3qE7i/N+TISgz
gplGKYwsq4Q5VydfLbDjDQWbvNoK8P/kuS9KQKGdkr4bV8JIqDDsfsBg1clUV0qG7FfZYQ2BIuxB
f1xTNE9t+TW6GsV11MDyRXxkwv6IZB37ZP9JTPX+vsITXMuSj5dDlSMXOsdX1v4bvkkQ/iLLlhyT
Q2fD5dTcnAZ85glJm6684sfrLJTGPPu8bJbjXUxD1dVkAOcs7UeUD4M51FB+wyr8xOgAuC1vV51y
XcDwgZZhAvDQXpRercJ+6QZv4OVp809/8rRgzLqZ/X2G80sjlZandOZtSPR0IhPfSa9yuJ7oMXg0
gcw05pAxg6F0qLLARV7kSm/8TOfhxuOOuNop7iQ1sd0EfmsR4vL19Mhrd+kiWXiawk1HhNrfo+Ba
3W4TGJQQh8E8sHXskTrqhExmf9RPiJ9+88rMVqzHLEJSw4UMpvgX8KsV1fUfntiX2NuoIt4TBR7B
Z3JnlcMGv28Udn7cdNv0r3UMgTY/TuajhzQdfIPdIyCC8r66rnGg5NxaVfJdfui/JqfdKebNkl7t
z7C7oGT2HFLXmDXT2FRwq6U8nVhauSR6fUrTTcIhiUBlxHUsD7QbKjyMNV/N5sZSNS5fO7nx/Pz5
MB0MWWysbfnAzoLC+AEt7B8AQ9ua5LPDk3Hp4PXGo5wepsg5c0SbeoPBiKKI8II7hoh8zU2try31
Wv3hEidmc0yz6cEd9E48Os53LNYGcahrNQAYncexUP2Jfk5vrTFCKUzynOE3aKtLxTv6Op7C7TvY
N3DgvRKpoVvpadY5mUTXSO5l/hqMhRI7KizhVi6LyDTnGxwJxT111az5a/A3RttA5dfabTeb9Tw1
re1wOv1smP72Z0zN2d/Dwlk44XmiNQwKPA9HrlC/BOkWoYDnibcJRbaKCvuICroaclTUVcEGG3GA
uX4nvCogvUYQ+aMJhOTzAimOeqJem1TRMPuCBt6+dypXmvK6pIEiCHLiM41rOi5QqjUjGxZMi2Iw
HuI0iuyKrKRwFoOKZbjIYUaKb5NknRiC4dA2CACBdqech7LrqeB9KmPyjCV+fL4TmHndQK19UIhP
+7+DUCRqBseQUsZ/AXTermFjrl+AethtiZJRb98wiZ7Qc+jDp497xqZe+eXUNxFlVZG3qduhHVke
h7LkomHkUGvSJbn7r4EucHYcibsNVDic9st+FdYJ4vsx4aQJJyEldv5EZf25iIjf/e4b/MLFXZgc
VU+/bAkYPWtuMjDsoEg3cwFb8wCqVe3Lx8BcDsrtx9Gz7Iv1zZvYWFoEz9830Va58SR/jpNRjPwo
2664CJIWxKclet4jC6E7x+4SylA4sUfsgQJhAmT+A9CTIxHC8CZZe9g3ped9g64w4xE7zg98X5iV
XmnXjL1PP2HLNkGxYzgiMoMbU3Nh0SaX2Iqu5CC6exomFW/ZACSP1IfCnTBizPN920nG2KiZnohx
HWEU7CgOWRuFMC2rVwZ3rXTKSRiuSEBe7E5d2H4Ib586HN3At5u/Wm7iz3Ph+9ITq+NHs//rcpTx
L7q0xwDj99Ej9spk7VwBQHuDbYxhqatvO5qNHMMQd9OTWdMnrx7XukzDlrdUgixAxeKUqwNFaHEQ
PM0aSZNn6xzV1Yw2swBm662xnYzcCYt/FAHh0ekh8JSXXXAcmVyTJuLGjhqkF+7o995NnS/kFuQ5
MKcUyLCg4IERAf26Ahqzz+niC/MAQh0Ap4c8Po6mIrZz2a8thydjxYes3zk4tAFkCBuceKqG1i1h
Csft5cHqLQMiK2z9Vkz9w/x1IkYc+Y+P8CwzkzstsFvg0NHJFqg9JOts9ZRTFKLFr64jinT6k+C2
Qt12LxdhixvTrd4STx51FKyB6DHWESykCF1kVkBgRfJWjlraCOP+5xHqu7VCJ7Wq/uuCVUebbpzi
QIyGQZ9GpmFq1xkjuu7wQB/T+PrFKYlvMjpvEkRyQNSdLJrGQebGxgxn0AsoTXAalU2LQj+DpaO4
UdGZtqHhfFyfEwaBHEMbSpvAyn5+lL7iA6TcDx+JF/1r9DWoxKg8LuNtnRrVadpKUMJa73t8+9/O
QG4rIBH3rZVSZ30t8zz/LJl0ht+wA27/qTjr7CyRYPS34U0Npy8hbOnt9tEirla4E4KwGP1MjfA5
EEPWybU4De7R3PiOXL0SJKfM3jCijK4+cK1vKQn81o0kCwJivNP30z2sBAoZBuFn9EQjKTtc5ndw
EC5Snc6btRguTrI3ijSPUnxEE6WGC8DICB5PTngN14WZP0Yx7NaoE+TpczkT31+94/pDl57suMSI
p2kOTr0tDdkGfiRpkIGkMejKr0ms89JQNGdx6t6AtJ6Kon6tDAQ/TkLjvckQOvnRDby9f6IZQAKj
zfF+8KD5W9/UAvmb4TINzsXU7lHYshP8wGe9gKSAWzU4bgcYl1AoyYGluN41tIfc79IPPF2n5M4k
m5uK5kgGxdGpi7W01kFxKNVjkOLqaI3HtZa30uJUBMfIYk1EZ9GoYH7dt5KTuKdqpgn8pFu7T2wH
SEznVQFRap6BgRCOAMWbC61nBi4NJuGRVl4cyEmzFzVfR/Usx1CfuKiDrw+tGw2GqYGdGvPZNuc5
5Cbe/1sL7QCDyaXiwq+/dRZSJprfkvBfqkMzUVJcNoWPXA5D9598kSowdlyS1VeLpXL70usLEkYY
C1zSs/7ibRgj0xg0Qo4q2ldr0OHfu7c+uhuEZ/lQb1wfHPXRQHTrkNkdsbGdGnczoB1rDNLa4id+
xwSKBXd2sJEwiYDAt0Uux0WWENxI6f5jXWEKKSQBiHn4crM8i8pTTf1EuQ0uCHSNeWRLvPPonlSX
eJjNto3qozDA/EsHJ9GX/VrB5ZOUPoTQP/oceyom6ntH6CPzof6dwnutUIpJ4HWo/6qsfUY77w4g
sHemkbxo0SW68ARcgOeDDBXan6MKgPkQfvyAHrQ8DZIPrqMfJRXvKXo1yTlVe7nsjlvWOkvj6zRN
ZyXSxkWNf1t5CisYke562d0qHk/i2HJhUruvkD/9kwcvA6PQSuvQEt7l0sDcnFYCG9GbCOTGLrkA
Dw+fWTgoo+m47TRu09BAtn8mlTLw4/jJn922EOy5wfrtFOJHmt+q1x0PU3W2PAarz7XYSNKC2cng
tq4eZtvWvLCmVLjIr32VVzuxDJxQGo1fo38Uzos6IbCAnhec5SQ+sF5+61A6nH25tW6zJY2x44r/
5VEWRX47fqAk2urihZ4JItBvthOcCPA6PE5NshGa7XH48jCt9u5sXndxCO/KIaGqP8yZnHG9XEUZ
jMg6hdb08aMFLf0FbcbyuiCWh9ZWFaxjNyPHpKysoGuGD061R4Fc5XvGdOWif6my1l4iBgYAq2Pk
bRHZ3WpOr2tcrKjr6Az8G7FjechKlV3eNf4/IgMkognKzCJAwjn2WZkJW8cVQm5cyw6WBwbxN+wl
ahBcU8fBbEUcN55Aw6AvxD8JfkCIxuKd6r/t0IktNeDqiD0MbYmbpQDHSuWKCSVczcOICxt1HMQE
DSUm+OHXwbo+GgD50sR3mFJM34fJA7qY4QF1hUxLwVZhH94QABDt3DC1MvXscyhGgxtxaTnJ2nM/
y+I/3L1M+iPE/vbH53uJI99Tojh0U1SBGSSIlfM5Ty4Mr9RNtXCbpGHhKirWBynGTVoYXylZF0Ut
mdtiOfBzO/HDJlLPJZF7H1g7kXJ8cIuCX1+/qB0XSTFKHhHassso71Ba0eDb6VYHlccyC1X23cXQ
bWuvugkf7cSqj549+NG7WcLlhgOsg37vvrN1fdQpSlOsXePCKKXyUOnNnyYabqnJzyTq895KpnBz
ztzmpiZL/ARogG6I8p3ih4FW7TBl676jRfMxoNzP3FF96kGdxZlJnyx8QBklVghYWWzFEz3WoSsv
pHlq9KwdbuzKdD+N3OoxnQC8JpHkgMNpOlgf2kcFpwlxZ6BeNY4eYuDrWZ9UROwPEcPXeJXtuLXV
fXrF+JuT9Pix+OetyfqtrdiStwFngcUa0lcDrzBaG/udj1tcvJucTyWq8WOd3zuchs1oDlkVrgHX
KNAE1gdINWsc4ZmF4EkdPxa5+vyrpVqATa94hvP9pNIeuoE3Qwwo/3VbKdwPxS1zLdhaugku/pwQ
xMhrOmv6nHMqr/i7v2ODwk4fPLvWzDPPkGlGuIgYuGSrU1njwTwB95vHaC0d+EK9KqApx0WU6Kx5
o+ZEMa879bgabuKtdmfUQFXw4V73CyOm1/P4FW35E+tfc6BzttzsLU6+jtZhoETVn+Pid6d23mvT
ZrCkG61e7xfVTKLGf0TK6fZF9zg8ZFCcO2178IuR4NRVlJ8ryAa1uXBBGS6qEjpr34U6qQ/cCrDC
8CzLW6iiPggMyQXpr/O/4lmzSFc7bFwHzp+srtQsWRDDZ2Nyp0RMH8W2YpBa4uWWQtBV8swHEkIj
h3yHcL5DreU3Nlfd53X2IVuFxLs1rzeq4biAKFZPO07fXyM/M+Mc2T8cAnXY5hP4tlzkfsous581
PB8Cu+F3H9Z8xrz7OFd+YYptj+9QtG/QRYgLlmnFOLyXAh4QZvSNIE9dgBaqtFePR8ZSTP4cRCeC
AmNfsKwHdo6WddMDAsK0SxQZROGFZSOIIqbEXM1J5O6BQmzDWbtFa3IyU41PLcA3tHG4h+vKwcAQ
S919ugj2AS7nJEtdAAa3hporBV1d0KjC/GhJdbx5hmhAZQoSH37w8HljjabD8ZMvefN4xEbVgQkL
Bu/2HlftNrhAC/jC4jl3+dwKvZfJIkbko7KxpO/17l7/rohu+ZgaAjrM4GvtR9ObU8h9pCINtZs9
M4JDuSlzA5oZJXhlAfXADUnfO0y2SfwOrKV7nTWzRT7Ip+KWDK+yeM032/FPB8ntGlyBU7lvtPFS
WLcqcbARh9qDQ3YRPhQwmMgUe67jWuoAwOh5DXH1CJCwXkCQSMzd+kSLbjCC8Oke6KrHZH5IBelj
hugqi5aqfKOlrt69Tyi1c36ZiO7iQOBbJkcNUOjvSmxeO6YNyDRqkmiNN5KTERlwZAvv8+MUQcTe
R8UXEhOth9npIhWz740pdEfGLqADHjMmoR+3FktfJ3FTC3lkd3uvsphLLLQuy4YffiTBTgu9zCrH
rPBVmRMAgvXWYtSBUG/zmNPvBhjNtWyZJljfdwIF6YXxoTyb2dbGVt6gDl5mnEN/tEJti80ruQbd
klpycYkGWFr6QlMRP5BRic9qb8gdSLQmIeGfUGnlF3L6B2UzZDJWfevNP39Am+Uv8E67HI+alsb5
asUAX1YdQL31NF7U4vQisCRv1HeDnAuq2NdmbWveNKFsYnEL8Ka1lpmjk0TBHFo/QQDNAQe2lhPR
SlWysMmLhiqVkZWjNh7zr+Js9r3dq4qIv3h2O79kXKlOe967rXgt/tynDJsMCUcDww5dxCc1Tobv
uSVmq5+a1WYXLY0R+AFwj1Ri8fcjx/r087QWXD3fByGpO75jVNS8HqH8N3aBCVtwjWOrBxVKiK88
DiRl+aOpx4IMgvE9E4ul8qCekdeukMMoCOFCmjn0sjFm+U0iSXD5xzvd28okVvw0dNBtHZqImI4h
6ipzrKJM2oebZMZaL57527I5vST/XA/Th36s8w5WYYgnaRZTnjWeHgHqbgLm2N0hDJieeBVE6SW7
UyMuIOjTdNW9Yc3DyzKRHA4fDPSeEOFMbarkfTQtPzsdO93oY2cWS2YIWc1zlccyWDXxnSFod/2t
2rDKFZXiud40hWMiDQD3f6uQ4v0glDdZX21NX0gP9bdnjnJcHpB79pUSWSJ52qq2MjX/PGVQIN0w
sLV++PUeK/wJ+CTvUVdfZeOQ2VuSvLwT9Ai7wMUON+S3i4NT2gz2sNGB7HOxMDULL9QmD9yGqWrx
Qr/XobaMyyPXjJQVj4/trVnp7h70L9NqRFysn5Cpe1iOo2NMuaqYnDRW53j5ikXbmN07z70zgefl
cujd3S7tSRdgCi1DMHNV0aAh31TIujtkfVeljhayWadbfli3Ux8q9gFLc6q2hVZo4g/bno7x8X/u
JVpbEKO+Y8qG1tQiNuqmhFvuUy6TUIzXnZglu9mknClSSkR/FTanuGWiEBRPHH9yiT3n84lLj145
efxoiQjEyfkXD+t1v3B79cJgx3Ye+jgPQXpIdGvvvliIUmBYbnU29j55ETSjOY7VS6xHgZArgq+8
zp4OA/JE1GGH5oFBiav1I4rP7zCxJFW2qOEObxmxRV+MA7sM5/n05mUj+p40yq38UYOpDNCi4YYw
/nvxnaqoph0ZpYi1hjrM6fLDYjIACox+7T8mUwGv6tW39IZ9rHXnXEUk1RiSzQYuRPfQ2bJiDrzu
kfCcJ+aqaRTVbtGWS6WN47EhEq9qjIto/a/fXIh+e/3kyFUr2d2ogWD9Xq6MKsusJ+xipIGZ5Jnj
Ha++3c2hKxVHndwid/dnXYNjc//qRyxOBqNxUp7EkN5F2jRn98j/YqdAU4QoQBRRoJYvyq/KwtuH
i0gLpJ+GBtptjQrGF1cqVGqj3F8ZhTpNtgxCaHXZCObLsjQMaxBOgJnY8bm8cpr6BKLJwSucfO4e
MI3VKbzSdonuwMliw4iC3lAfH4rnBa1sTQW9Iu2U5TNMfpQK1KwgvNP4Vp7kapCkl/CLUoXzQlJl
T2oyFMpdcdELdhb7HynRXiwW2QfxggAOiny9MuCzaKTONTaP3aurO3L1Y02SQ2U1CPR0+ty8acqh
2NyuJOg/nJ1Qn7iN9n9AeovZJz4PZ0bmN3YfT7vIZ+ceWT/DB0WuJPdpXVfwJPMjqmYhck52DjLw
6N98N76OwnJCEtJU3xUwF6dzLeVBU9hAVGqy4fNVdEihOMYJFp0/t1K+uhnPFtz0MxZwEWe3nI12
p8eufsQuoWuLs8Fi+uDAWfTokI+iz7wEokn4oEKwQ7uPDaxJtYSzYJfkVhDwhUbOg/G/jeBRUGNV
ILYNmeAjOnjXvs+jruEV+Tp6hstBzMmyEHxhDFGCNG6vAhtNfectOJj7uk7aSBWznNGapHq9RxrL
1CE1x0mUH+k262+PI0qUaznBB+jV6Pf+g5vMZrCBr/cf6OvmKDSRdOANscEP/RpvTx494pEBunyM
IpyQQSUj2xhg3GXri7juocQeXUdD6b5qtHlbWmNUKNe4s5loYifN+IQ3KF80wsBZZ39qqzJ3n/ns
UyT3lLSaGhUTkP9G0XUIh/vgHGYoRCI1FAWgogKZkMbT5XDxWm2wT/v4NM/TBHCMnw/RUhcuuayN
HPpjE49vDsfCnxKxIQ0JGrnLnNYu+X3iCub7viNWWy9Jkdw3jl8tbqOsHZ6+nkvKhnLrWCMOaBhx
IlctOm44U4IFVReangBHf72FrLmMRkP4j3tevmnuLbzugsHtzHdTeWKN98dGrI1r5TO1WxXI1Lw1
5GrHmwz4Z6+3nChLBZ4UR34wKckXNb5S2RKURgMujF8HBPk46w909S1/Xe0y0un7kUjGgVo+RHb4
/i7qYqr0v+Lu92LFSa/rO1AkYjp+BqQzyqJfI4SKlvr4DyVpvL5a+E75rfKkj8Z+/2Z4N+59qivW
DPkH8G7Q8Xn+0ZmfDGsrhWcCEbRdgaPosD669Lhk65+IBlfEaI4MX/JYrlcCrv1lrcjgG98LWrbW
9C7X664Hdr/FFFw4Ut5w0sTSrMn22b7OYjYGDLbLCEl8CgKP8dlihM3ADNGXl7SfE39okaIQ4Vcd
ecxyLOID+FM5BfR0man3wabt13cUMh5Bv+bxW7U+h1RmE7s0OVJY3LOoGy+V/WFDeZTJwofkLcFu
YwjZ0xHWOkwHmnOlFSAgkRLBO5kqD0/KfG1Oh5PR9IJuDf0P2VuT5SqZJM92qWGJnByT3YKFbzYj
48pJpI3KOOHUOOb+eg0wS2nQnO2ecleElfy/bcJJrJn5r/vPnHSbroFyvpIIKlr7TvTN63rkCNyS
7s5qct0wKpP70ch78Ebz/CTxGkxBxp44I3RFOaqp7B+4WTj/l8pZc0yp/NWf/+qQ1mvpXu4Wmd7e
szHNzWEMjy47DLaIviIdrdZikfoe9QtdJJ4IpTVziM5CbKi48RIR2ORxQJmRXDtlL38jEHo/ASVY
tmsy1Ma/gB0UAlreFWKIBFaqeoi39IiNMWJ++MAdXpUqO5R+iTaRmwIIjtgs55QnL6n1cwrOrrRP
NDyqbFswCHkkdcsXuFYjqYnqw/IstEjfH4S8GavX+CWDSpG8vdze9iql8wXTdq4yhmSHnn3gYZoV
ZFG4ML9OIBTWJm52cRWM+8TnFqsPFPoMMd7LiOKrZu4hPc3vidEmUAU6Q7FpR7vBIcmJT79VAcoU
KwffF7yN7JQo8unSciPaqwfHsLp5eLNRliSpf2yiktMwC4x9uTDrlEfWjCsu7irjO865zO3WiVXM
oQAIFTCOUSrf2+v9VyZsgElhMXiFFpyjxaFQf0adqrxhURXEEVSTro9HvqKDzTEcx13/6EHSlJq4
ReeNTJzGyEEDgFIxnhFVBTYgcmO+VI1WqQ4F5Ua5eXToV2yLvU+znnXsGyZnFeS0cAVY8GRFOz8V
25MbyQdPqiZPPUiJah1/cUD56oBlT1SFvoQgK3tWZehrp6UugQeolSvctHOYy4p5rT/YBoW6Q3QF
oVOGvsloDaGMgjJ7LIgQkyIJ5vDhFZdlHDrpQRv1EP6m4HIGF2j+FWXB1r46X6+l7XrPOrqrPr5d
RqJOyK/99/BZ3U+4Nw5hWw1UWTkHKg2xuBABCiw9dz7S3L091jSPEQreXWIQCH2iGoUgQ1jii5/o
YtnXxSCkktVZztebCKnah7KLeOO3uF9b9t5RTd68lDW+eE60QUbu6jbYHDdOtQOP92SjMU06iUWF
UhOjq7Mlr/485otn1nTdzOvlh1ObBoevrPoOoQQd0zU1jzR7JVVfkr0OV+q++yefg3nz3kpJfrpx
ok4FYjkaSNaBlUZfMJKJtud20npcYx4+ulPglzw+ydT8hFTLNaeTO8XVv7l25yVKILkMTI7bGSOf
iVetH+kkgW5/g7WFs8ENwkuAwi15/Qzb2R6dZ+cRYJAkWbjWaOcZIEw3R6DeG7C1srzWqPB+Is14
g+Z/VXSoySp5Hd3rZENYi632yBg3tB0U+ixCM8cT1bBSSOKfB9Cmy6BwLi2LdAIG1E7c6kQzD2J5
Cjkj6ivvs4CKd5f4i3GuTLo1i9ZBCbGngQrQiqHu6c3hJuTEF4+MdTBUYBOdMk7ZhnJUuaT1lVtm
iVyypKtHEGGNmLw2A/092X7oeq4gW/YI2Bx/3oHnd+qS3tzdcR+sqQ9mnKwc8AvIe6Bb0OKGNHy3
Nqdkk2Pu6JwS1KZicZnlvdTpUE0ECJCJyekHIHxWW4IUgHoSbU6jCta4K66iIOpxwplIaCHkHzGS
0uOEdqwDbi3Ax8Qs+Ax4amgBMiMR1eyBwJtoQ1cbFSyag2S6ywouiEyZZyNIZfGYSwH6eIRGWZvr
afGwXbyUKfLmPv99QbeXrfSsWskL83pye3/wQgchq1BRMDEQ719mpBOMSQI0VAjUvbD+L3knrdrH
i+CH1Q4X3RwracgL7bfWzrkwqcowbhEL1a9DeMi0KeiJ/zvyYAQyyoVXnljevJ4Yi0Wccz184Ako
HqUw/E68jhYqb+3TKEFc76ltF2GV3MQcxSVpmJGa1B1j4jVHRdJo54NcZQVe0iXK2kgoc9UnjL53
PMVMCz2/le8GeeIfO3lfMxDcMF6RH3tLy5WUpLzFMBRVcAPyaT0It2NsIhQ9fm5AFZqNC3q+5JHA
nHvQQfLJ6QXHgsX6mGzNNWI64IkyIHBQI2ecZqz8SwdwCRPnuqegCkx3nLx8fTY/ApicX6jVc0Zn
345/oXMoLWLrnla1y74dAimE1O9d2A7UM1NyfVroPcI/5cS7nKdelHluXH3Gv5R/4PuQchyy83fn
BTkqVVX7DuvuF0SpnmR5iboCDMBGLNnOnmII3xYn189kJ5L14/EdAYjyQ5CdFyWNEofygxxQyMN8
GBwtQkS54MBbPq9eLP4FiPXDnMLFsvXmqyoLdFZA8JY4B3CE5pAtezDoZc9ccVYNbII7zeIqePdi
k7ntNqhm8UoEaruOAXQtS2VWWnPveXRnHCRK9XM1u8Fo888qTpeg21b5nxT/IWEbIImmjufu9C0M
3DD7wqdSYiuPu2eagpeXM5XNMphA90rus10ZY8/zs364gxC1r6ZByLOJ6VPBVvdVfUq0UPKjkeDX
SArqCK+KF48Sy8KnYmxv+hd9lXA/lEu1s/1SSzs50IMxSgrKB+mZ1xla0zcFsZL6lPZ+Uf28UJyW
X+ElpViIqpojRoiR/C50zkbGrH5JyNw6S2FEdMLXiwrxzrVz6Yj+W+hYt0dODbA7/W7P1XxAfTQE
ragWLQSs/qZt1wraned23E7W75wHI/GtA7yWiRDuxLE2nXe82ZQb4Dj1TspfN3obZkEJb2uDlJzV
MmERzTQOdX7QTNSfev3SVZRq5BHQVLJE7SeaG1KwTx48tVZlIpfPdmELRYXgWsw5v6qbDingZV4D
H360FS3Tbyh6RooQJl8LNpk70gV+o+3Gs9liz2aRQ47qz0FAuHt+6peokserKKJUrCAarhjQ61Lh
t27fEXN5FZTV7zU3V9j5iVJI4Mg+jn5SOlfUnwyRf3Uto3HzKym92SnHATZNKUAiVhl5SNjnkZfn
FbK7oNLNNBzcaOnSAD/w1BDMzIzeQkQGDR8le8svaPYddEmIe+asB58pk9Fu7WcflLmWFQevvQvt
obFAb+EA3q2QMwUfPmoEayR4G/rMVKJGxUJiy946JuCIl0DwVx1MzXzEtzvchrS8Z2EWi5tqUBUw
p5Ge2zYT7Hgbda50Sz8CTSHx1iIOZAjfXw+ostOzowrymc+h6ucfzqer7Z8ASuckPPpIk7nSmMW5
PTSD6YHARcaz2sAc6Q0WaoqcYn4y9MZtXJ4bltZBJ3ufrpxAIiPAFTcVfj3pf5jn9y1jvd5DhhED
RvZ+NcVghx7n6BLh171TLD4Mes3rbXuIMPKH8u4Ddope9MjChjPLByNgZ+1GGAgf8UtSEOaYbfRI
XFvr1yDn6q1UnQbTz0jc6K9rOY3bqGEMPHrsfit20LJa8Dta3A+/6Ut6AFTgliXesFS/U9uxtBfy
5j8ZMxulw3YL9KjwZVv0ELgzG/37zWbCOvjsnvAidDTvQraO2ZS3JGBQ3SoanVjLKOkGyQi0fl40
CsgPM5DeTXalFsw5TtLrYM0I5gC3MTGEzLcSsMk5U0F1Lfvp99Tex/dE3onkdsBJp7c4bpKgD6IU
fxoE+aDJEMpuMFshYwUOmDBtk8mzRoZc8TxdSEj7apIVgDfapKCSYGzrnRZ8ObAW1PJCw8z1wPUA
quJwj0ZQ5NEyy+vHsEj3F+HSQy1iXMY58GnUMI3IX/4dC/91ECiVf9HNrnFr1GOZJR417ALJpoAv
vev/od8BcIs2B5cImnzDPlw8MB4bsmaoLozzFxKaeSJ+OkWiEDKgXctn5d9RTTE3o96E7X5qegvD
pRZlcXMI9nbpLtW85co8R0EGUcX7rIFNpA7mvjA5sybjQGXK1Ojhx5CKrxh53jurviSQeXNNVfBu
er2JFeNPbi04zsyyWdRLcc66WdPaZg0GDyQopaf+00nw3Py+xaTR89mMVkO9o+1sHLQxWclHmmIu
I5NqtTPaxLIuth+eL0v6nUB7oXR6kJ3NKuBAZbHCXPOHYB+G/CrhviQZM7h7ud3K+EpCn/DXdMvt
BufbzNI8ZF6KxvXc/uwL34KIcicOFhUYDp8ehyAQrcO7C8I+68jAJN6cHk2DbycsMw4IdrQqmVv5
yXUNSOqBE74Y1ykSKFR82ijUQ/eg0RLJcupKRv6KCicJP2mVnSwWDgyESTwXJ199owjJiLFb32KG
SicQpi/Vk0/dnV9W28zTMrA+kfdSv8ubJz39Wjmgeh8FZ8rMRbR4KSl/2m6ScImQaOvu2nz6/htv
R2qwOv0KlbtkMjL/ne2i0p8aPNFBimqtG8YTgnbcziAFnog2M8S1z5gZMFeClQs5sYhlEjSlt+04
aAM+GfDajhqIl3y4biXnUFAnpCS1ZPjwtG5QOwd9D67gG4pu1jM9/NnIcPWTcU1D70pkm0VGuGpO
P4W/MFWHOKeRq18uBiHJ3euUbDn0gBWT6P2WYImfJJ4KkfYTTtJUh6PnBCmhSD64nGDFxcMK+4Wb
21wDbDj7L/8JO2P8vZfrfLA8p2u5VmcuXlmGG0Fues+1x17ZoMXFxcXunLnG/h82UQ93P+WE+Ggn
jHSTtVEb4wbyeirAw1i1I3YlIppSbWUtdUo/9kr+Jn3IEiFuOiD9ejG0jIs4dc8+wWDQXTsiOqpo
EAnJg5ok7rnG9t9nl8m31k+HukpJJqR8N5tO3oEkyCjBNhDHs+k5PAicBbo845RNXkys4jG2NCjR
kLwfkLOWPAytP2s9SsYL/+t676h/4tf2gDiOzz16FCZNMxFaCtZt8pLswGXe7Co6iCSnN866xiIy
F0CD97QfkLBeUFMrdTTikt/CtiqUMKp5e80ZVVqufnbGCHtSMNTM1i/ft8kjFNw5C+xjJuk7urxk
SId1bbB1ACjDKA/8cdnrq2sD5NlgYTwaFvMTgi1cBCTtiA3oGPQH6eX1AqWdiX5jYfO6lvWL7WSu
64qVHDDh7BmZcATpOD1xR+yemXPZQcUaBeOeX/BbKLbuon3lB1H8TyEvOh84DdzLhzBZS8UvAxfT
WImaKKsNoDqWIaz3JthL4kVwX7YKLJ75BCeyvpx6iZG8F26zCNIv2Ry7t0XCmXUyL3+1NYbE+Zv8
IcUFbN1OffsHIn9z5iDfOupT3QJjS7xXWSEH1bbHuD16unRiVnrcoIS1YVh6S+VXAOlkUoS0IhZ/
eEoVW4Qkcl42QOzO4g0QIwbbsFQeq9OxEYrDDOVUdJwqGGdQ+feYiJFKEbIcDtcQUsvVyigmoFqg
7Ch2kvn26PYPRmcifdgtI9jn/JLwCWGon1lk4bqjBi+rIQp930SlmTO5upzXeZmxBKyVA+GgV43Q
xkJecwgm2mfoOWVhHYKavUnX54hFEukdj73OV1/Od1wSakuUfiZlNYmJqlaUnnLvE3BvBESoYBGv
UVevKTV0ReKZcS50DuIXbCaoquz22HZjo08L/8M5H0IDG7QNqU2NNVzbj8EUHqqLAFCM7pFwcWDb
NKPgAYiC/V30TUyZL/6i6t+B0nIw+vmyWMI9YwwWK/+5zrgVz8saGwGt5gsjSZol/LfSl7Z7uoUf
WGmxk8H9jCD6Umto7hHoldpC7jtx26gLKgk+ypvxNrEI3hGbFcpgi/QI4+evUAGacCSfGcC5qVqJ
3EbpgsUxyMo7vLXAY8SlsDS8jUoCo+19vBJU9WoFFprYkjpUa4aQMRvEePuJP/J2A2xQtwOCM0iZ
LDiUGarI0op9ATzTqEworn4vmSPakaJ5kt5VsHMZCmEcNUAwu4ZENtYsstJaY6q5MmbSbK0betUJ
wsG/5zNO84kRutcBoLxhpZS3wIiZ9bC+PJYb+GinXA/ysGHM7slhuflL8leCVY5lkU+Vj+KLdfxZ
fF5pSQ1dR+Ty8po4AHJoYiix7K/4BCU8j7OZrEOzxKQo3e6E4HrELeHnc+FdMpxYBl8u6fMaAzar
2lkVSpxM0Gv3Gts47mE0Uw/PdXg/xstHcROsiA3ts4b4mmcxBofFpQv9g0ZEJ82HvcjuuR45RoJp
f0Yz/Uu3tsBWPaVjen64SqmTOAZFVyBXpWG+4sfO2m0YZj2Dca3NieQ2ZAMyadA8OnvXCSefC1F3
5TdRXSio6x9YpDPbpnl5KJeTr+AgeUNsiolWtg9rjV9Q/PH0BxnJJDQv5rpJHgCPSaSC0EqShA+r
ZWJJHOgtejA0FZu1bBiRQqX8NUegFhtGgmuziLZtJHgz4aRZQE8VgLfhDP7OI8dz2t1JL8okUz6t
ogChcMnDvi0QkBrTUiL34yNlhth0xOkZoLwYX9HaO/SxTSItUr29MR7e9W6BWaXQuWORd7p85J4S
VAhUeihzs16sHaSys7D0z2aH750SCIb1EJ/vAOaFlUR5ciynl+X4eJMu75ApXnxnYn/vbOCjPguW
sdPQTCQGO3iX2HvGFjoYg/6euqqIXG9kE+nSI/nezy5QRA5cyABERgUlyguyC2I/4x4JiuWsPS7k
9+Kcd61ehsuzUAEHCwn8U/T72yTU6s9ljv8hKX2OkG8lS3s68xVh1EaPw9fbKIQIfqow/m3MBVoi
2G1v7veY2L5SQxzgq1noh0tOXlTOeSfT+3bqWTnQnz5zf6CgHmwD5BQNq4nFoT/Z9YNEQ7vOFhJl
ci9lDUH+NP6OmAyA3jmxNu5bL4uj3oU+KTsjuOJF7t77M2qJoTZLsaBs0N3oz0HITVu3BAJHqP8e
ih56xTCJNsdBX6nIcG/P65umfr7tD6TjU1vvuICQA/N8IxmDNxp6RX+lkYlJjTH/VoiA6FIUUFBJ
3lEphMjOYwINs9Za2EpeBaNB3bMf7aZce+uxoiNp5rU54RTlv1SN0E5hOgshbw02xvXrnjpaiXWJ
3T4j+WlUFFhWKuPz57k0ZxX9iB8w4AeEADcGUHWCadyIxIPBcGsTn/aiBRm16nDTnLJZyxeD5YiD
Q9MAeZQkciEINuxsQ58Dfh447NL8SsixsXOVubSWXTqySlZIiUTNkgvded/Z4665LJMnFJsBl2tu
6x6nR9UrhqWUhAPOXqNv+pLyZZhHipSCK03s8glzzT8ScAZdUXPrEIUO/bTd+HsCd5jshF5fwemI
LKARDChBB8hxVRM3ZYypcJn/DgwRKfTbT8K0GkRsrtBW3/9s8VEQtsEnX2YNdDL8dpqC6PLGBCbj
1nHgb4NRxeR8uVvxCmR9gs9XqIuQlym4ISxT/Tepk6sisUyjTNc2Sik8ncxDHTUFmNZp9OPJ4M7t
aaKuUFOXU46W2R3e+yhazDcMr630KPCsgUFVIGPZOyBAv91escma27Hv6pE1b/6UrgmIdL61oscw
yGKPhS/h8yG5IorPro7YPADDfdaVUJ82+AudiTXUe7sJfyKiIhSlR1c3m7W5YFyArbuBA6LC6quj
uqyLqnatPxCLOZbhfTsa11xOO925BWgBfBckRkqJOmciFHaeO3X+jexa8RFRBuLJIMoVLxUtx4Qk
NN3LgGKPOrly47R8L0MESO0TnRUEu5SFKhKwQqF6wUyC1HX+tI3cGPUR6t6k3IHvIzn/1AAvshYY
zpYTjjHez0iSt13PJ3iuwZXuc3AwMv6g9xQhDV1ltxTCdvxV5x+WiKXQ0PYEg1PLd40D0pd2ISs5
vjybraQ9halB7HtMOndMi3JyRB7nLsMSY2cu/FeNgq3iruqIpS+VcjZZSPpKy01BTuQW2MGCUZCh
kDsPHoV8Ilk1jjXcFsFkllnzhhW7vuDC4FVHO5kD69YAa81tlFJwHQXuK10JG8qXmoWw21zxNzz1
3tNUl/vQomBpYgl7V5Ggfq9IeM2YG0RNz7SmuEnRpZqxcktCbyKHL9narTq+dLoeoZlCVtOSbmNr
tlx5KuuUrKqoXzyTVTQW1zgYtIxTT7ZFeQFLURx3QGFoYXhvqvwTgelWqB25iqIvkDCZ7T6W97cx
8NIVbkKUrG9tePe3TQbwP+BA6CzIcB5lj9pAMVivo+XnucJuxWlLPFlkpY1Hb9ZWL5/RawB0MvBB
Dv+zEOG62tmXQ/MJSln8Lu9qh3iQdpnYXaEMxuzkd36tfGnQgg6QCWjxhdJ6OWReTamQFPGARahA
BxxePJ+csxLBySbEa1nC+S9X+AUrwPWafvOgB+ANt14HW72PtSj6nQDvcIdlYW5+p3f9aSMVcj5i
z903jFkhu2knrTT00jGxEGk22i/gKPNwcTsUMoxZreYyNVpr9QOEeg3rcrK+qVvbjnFdmV/duCqy
pgyaUPEjJZ7NmJgtTzdMKqSuk8xlHriIMRXA3VIdKVg/qLaGiSpnpDulLBkmwEo1PrLvrpMOZI4m
zvANwFqcwi822t++B8EVRGy/7PibPIe2NCdy7l9x/4PV8I/X2w9VR1v2Uo97/45LtOPeKz24ksI7
+/4AgZCye5Frvkt7ms69s7dg8U3qiU1bTecbbu5JKoa3xUpC0eQY29eVAZnUAMa7CISlQDMwinaF
rtHJwsVR1i4fjK6AgGOxDIDC0UGAApTdLcWAP0amq0ojDS2qFJ/aKegc4i/+jw+L3aHSE6dQR8/D
jqFpvMwtNYzaohDYpT6RvNgYo+qd3t1fy+/o9Hu7Y6pyC1sQfr2+9eS+OrxqfP2cNv94lFAnSfsm
cTdbVUDL/Z4ZoELl3QpxPt9tkud77rmkbNxTdBNpujU11QXfX8Af3OrNVzVQJGwL6LFBsfVKoSgH
aiOG5PWlVTG7YNHrLBjSGt9YRZ1CT8fTu+YuQ/4RqJz75JNitM37/G/66Q0vZ4j5Hoc0TGB8Gvgf
ZoJ/AU6dmUnSrLWAQfUdoJm+bSgwnCiFeUyydATNazDA/0wAtlqGVjHdQ2dl7UbXvqj/ay9L81pJ
vEKqE1VBduYHLOUF1XSNWiJAdZ7N3/RFvrEHLuCD/vdxI8mKJ+2zWw26rjjVPwZo6EofFkhtQp6s
Owy3Yl6o+Q5JNjkKVZw0rJB6+HgZQ3xlYavI2nccLjozju0gL3WnXDpFXILWURpKtwP4D2WVG3Nh
wsHmjn2VT508Fv1nzAHHJvXo9fmX1iqEFALwDRW2PKI5CFSaUjjkLYlif/4zsb7RNrW/6n9JezuP
C8InjSwhGV35k9XaupSW55InaQqDW7YIEkihH+ZF4lAqXFlMu+fxVktdZ5TDsUuYeDVvpTDRFpXD
kGJuwIV2SDdjdPb5mqVcFXB0htfWI8GaH5Y5z03abVzSV3+9uyMGEh8tc2EXOwGDUhV/KcyIc5bl
N+xAZfqb2MUhIrOa4mrdzAdNWBRPOROv/6piwbFgiCnz6SPECh+CqrDGTsqtoM9WKs/iGRlFgIQL
4gH0K07EQwBw+wDl9oY1hwTQdqCh5iM/5/FcKI8eepY1UmqVOnoGSg6mlRx2xvl20Sb0mzVfdNtj
c4xQAo1p7gGudYy8mj3BYzlxoJs6sJrYPDN1fuijfH4VMY22wQoiBDUzrNjzz1hNYKiyumkd70jb
WofF8hOCwne/scl3yn/2jirn0sy6dHY+x5Efke9rxKpbsDVdisXcYTELf4NlgAuMyIruBQr4nNMm
I39VlYnLt7Ch7aZ0zngkfLeq+LjyDzuIJhvH2HOHPVKovjdGfKVr1WETvTt1osz2sN2YLp16oM/0
0lRjdDoP0BBRZwExG+2LAOnpRShGVu3kJq3niha9cOGzyhYca+OgcIlGYGnGiMI9hls6sZ/h00hi
KbVzpgQ1/KyvGq0VJQcAy9CPzruThpkrbr6LcJFvEq0fMyayXT+7HaGLfJdnF67EbrgllORG2dYT
cWTSIo1wn31GwXNKhwEouuwIG1ttrTlMOX9zol9LOSX9E58efHskbcHcWdQ0a2uVVobkDmmI9nYn
zrMu0p/U7vx8PPWwh1CccQaiZ19fKdlcnsx8X7z5Ox+87UkrgNv3XMYt2PXWl6TbgdpwJ72wj0Eo
vkBEgxR/NbjpMzswVBo7F5W8x0QbwbLcbeU1wNX9FDlOJNJgXQLDV9bDXcYr9duMlTho1Lsy+Qt/
QRuiCrWmBs2GnNeX9FIMz9ysC1EK1IU/ObXtjCh8CnI0cOv/xVR05ku6fhG8imfKSpEDryDFyV66
RFN/bQOvGnTM8bSY3MeTbXcoE2qONmsrqEPCE2YY3sdK8eSRMdPAKjTemIkd9TMo+EyvZ1YTEd6B
6CYg6mffCDM/wcwNsB8/jFG44t+uIT+Vf9hDJxVr7xyWj3KQ9EpPGDFktS4ZNgHh97wXMVyroQqF
hk/eQe7gv1p3AO66+XuLI5x6Cksnuq7/mUM6QInzjUKNqpNUTma/3JGWryXY7xJbomHY/Hd9fB1F
S8pJCzOPEUWdQCckjvrqhw9FDgtjyxpAqddrJ3ZLWedo/QK1uI0AiBO5dmDM/TwbPQEtFZR0mver
dwZk/gslIlhWVs4vSvbdYi363Rbx/qmZS6SfG0cylzddu1ZljhQSlsjchcrHCXYBSC9DNmvvgnqi
eA6lQE5Ur2WbHhKKEGLqAIqJ08Ia576RufiWqdjtVjfw22AxuhuWYnLFGDXlbCNFiy9ogxBxDDhe
gtkmGws7uoBTUKCZsJUqWVptOK5N1DIYryGlml2PjhkK6BP+v8L3RwOqamJWPZ/nUjHE4WP9/YxC
rrb6V3a2oleqxlyXyRuzjU+w1yFLyavWzhFRHnxDgbuVkXmjhcYG0SxhvSBFBM5XDPjoa7GIVL1v
bzHHqi5mV7lxADDlhqvdWX3G7zaAze792w87hxgRLo0fizyNj/TmZNVk/zTTxxK2+wqDFoSjdtBn
bbitlurA3qekEB9koe3X1+nWMoN1g2nWkjxHihYUVPNwj0Os3z94sdb3gYW5CKdAdLYpjmvCrzOS
cRIVWdq3hchRo3UQ0xcGpTh3jRm3Wyk0/1TcBAkafxox+/0bCcGSBWJSzcYuN6G6oyyKubzg6UY1
aMOAIgCAwu0Dnzj181TKzdWu/lGs2mVpYYrWQI5txtgfdfT1ZcKKZimsYK+iDiPLZQxSaw+6qb5o
dzg7eGPO5BoWPONIfdnFg3VAh6a92+47xb10bnp6kc9VjCbeTwg6B/4QgKjP2L9fcuq/UDLhd6Xo
nQsrWUPgSrpWvhpUy6QyjlcPzErvvIw5gmlkHuZvBUPUDA0Wp1zFeUih+9RTgpF+SyA7PIg4X84w
8IyuqMH4f9AJRrRfpSJE4PdoQMTkc9eS5OBLZZZbiBhHi12DGhju+AcEianMqiTtfcEscqaUlTFH
QSYi0wWlOIkMsiGty8NyadC9gma7vvPBkqRHSaIOeeL+iIo/2XNvaxERygwOyO4NPcYjht0yVDDX
J0Gc1KBaY7hbvxpleBuaAQDGCRZ393lN5uabhWxGGGGuFo7FYTNzylo2PUbjNpa3e2HQxGpDVFfG
Fc9EMbVFWYhbCcF/Un9U2JAz0s+Z5Prc/72nRwQj2LVUbsxTMlGtUGP1wv8RSfv9tWEN3NlxRMQ/
plG4cWRz0s6b9va+Oilrl6TerzGZAsnsZuYBE16mQ60vybqAvk2i1e/3VXLzI5/wcuR4nQqYnaMn
SFQ1vTu9x3zssozN3D6OiQzkQJiStDk85h+iI7hKNtw1wVkpUkhcyFgq5MIfNS8zaGVw5Fci8Mvp
ZoBwt5itoJKDbm+Itj7iXRpZmT1Rbw35VjyDq/sJf7F3WGmPfqrlAXnQmKhxuX14SvuH/XOkk+yd
svN82E6QhZxYDJYV4JcrD9kyirz9/voOL/VK/u/hr7G9teLAuw02Ge73I8dPnl7kRupd9SAJV9vu
c34Y2ITXmIMH5+FII/6HYPWpxMY/2Npw5Bz0jodZpgIWgrpswr3JQhoPqm+jNLknyxTU2O/52cWe
xjp7yIj2ljpCevpLIugO7zdUHqxMYNiGtA3nn+WYR7nHFYRUG5ujDT1k1BvfMPDUBT9AlB/rI2ZJ
gKSxvMq//1RhZD5Ry8eyWNd5yPZ6dJU3XeeMyOEsV6PEYZtd7cm51vJBiQdQLi5q0WaJh/KmEMdf
d8KO39cqRGWQMUpYN7V7ebfHR21boAipb3TjyS9v063naVVsiWDbldrF5goiUAyrEw3NBgIoRCIv
etNKy8lJA0zhCx2rze2NPn14BzZe5lZSm9kfqfYtQSpfFPKhkdtnyhDHX94e/4tHpEiJYRHfLswS
unEvl5ohrEdzLezQ9qrvge5MkS1oLKPMKfJgJzrMzmjqsuUgMN8BxHDgNykk1NkaKNh3eJWZkMw6
xrgggAVJLtvWOFGhpZdZd2BZtpxv4ojofyuJQZudS7uncS2RS4CnDqtbcEtiJl0fInymA2btVOQl
qTF9AemyN+4H+Eg+WacFklzIlbZxrO/67gWJYjOLnBf82jTggYhVDtIW72Shc3OjG5wpQwsomn8G
Y8921YKNY9dNDTQdCeGQZXS6QEessEDJ4R95/e25LLKz6WVvi0j/Y/6uiZe4ySy5gsMTrH4P84PC
qogGITGEtLw9yMJ0cVtoRdCJfAmeae/brCF8b2rloY/TA1BKVw5DT+DZw4DbugyMknJLonjRflAY
p34A/M26EeSwwCDeALv5hmyFmQddddat8omwxnFb6ZJxrhs22AkLfQ+PaQNQY3i7nuUnFdm/AJQ0
oEP5tM7rk62dRFvEwSc+PnFEFBKxmuK8rQphOfpfWNo+KOfFEXTn3H1xnl5/27t2zaHkKh3/SNtK
BHEPPghNqI16/pQ08PqAc1VgmievvDk7Y7BS4ayxH2iNxsZUnEKysz4gbRSfZcAZzFQ7p4pLC364
w5ZGgm8YSTvqo795LhrX+155OrW/XzPhi712U5uEOzhZu+R9wD+Jzvt8wi9MNyVCUNdAdvGtCbST
XesfHvWHDOF+pKa2v3doWu2WDGYXP2fV+nd8uhWfRq00TnwQs89MxOgYOZq4j49BCNaxsW/JV5xN
GWTO+A6YUmuTP2NNzEPsCuyX9r9n649kayeWGRfPgnp+pDp4zPfNCpgFSENvSBbURa6c+FTLM5+I
7b6RRzXa/a5i5Bn0cz0DRLDJsIKpVyX1pbipAD0Hs1PZYiEy1t/gQbceClwbmjzBoram2WyufXAT
qTLn5I5ZGAiRqSJULZR6YT26Rsx81nyNPK5vfiY28Nv/FNpq9/m3N/NqVzPiNqULxIgTcV/JM8P9
T2g4/hUkjcREPiwSQQ/ifRPEGtsT23SSbjhkeypAi9GuuALsxOCrL23tVFEmmTSPERP5Wvo4yS64
ypx/WvBM3MKinQf7VB8xqfxgOt6G6CKpZjTEb/0gU9e48rMyk4NDR+OcJtYy5q/qzOJWzKrMxPN4
BBxJuftObz5+3SisBgL30IthUplVxRiTyDGU0MQueepDfvw5Wv73hP0pjGEGgH+e3yjOypz4+2Ss
FE141qd6i0tqh9Dzqq1qpAABvdcbYBgFxAPxms8NX8XbznHL2eQONsSmGERJfAOp9r085KlGaMaB
XwOk3B0iapvsHwNA/EN5/DXLtPrsk6itn7UxUxsyToRB8X01aVGn1uAi3NiAdT3bEeDma7+BINCd
7PCN3qN6JQfzqLo7Q7ccLN0Za4SMG46/XE0/P4BhZcXOa5FJZT4FH3ysUiNdZK9eCqhI2SaAf3nP
hoc3jVh/Qpd+m5JTKulyhPrQz83NAiBNjsOuiLn/7+M2Y+HXhXtuS1ct0OiBSIfQadgl4xh0XH7l
7O0QuiOb/ACr2i97EgPlU4X1XajrWqaODcx+bUo56bUkoEGCokvLoO5CriJnMfD1JpY7ThL6I24Q
c9mtWPK6E1VkPgjQ9kghLYJ4C0qLaKChvBVwfJFyyM40QoxTIfe4hT+qOJ67pRL0/KSY0SNylHdG
XOnq/ycwp89C6XckbSnLXn0FLbviYjJN2OkLwvjMEeiKSNFHqCdwWqdziJ7JhDQ0kfyxzoc9dZY+
hiIDIRml4IsjHaoWUJAkIuN+q+U5WDBn5SchQutYqDCknKvQlns0bLn02Ya04XNovCvH1KkmCD41
0a4lz89fB0YyMg2QwNigwFPjh1SCS4qAfayMDojSTUFxnl2aXYQ7Ew5/a5QCLyYFg4/BVJvFke+k
aXhAw8VkfrzEeav5i6WBNBdM9g/oHhuzOuzChSZ1X+5BSZ1X0VEIL92poO6NL16JJrledBQZf9s2
qs4dIvUTIpSfVAfINVNzd4OuYjyXoJNP1mAEUrHHVfY7rl92s5k4euG13d817WVszDzuSsSxUv3r
bRBUvVU13KY84TnQSyyPk9/21J6P2e/ekGqC1bhYNhxxJ7rddsQ2N5ioN0/Z/rsd0OOCbzlnZIhx
fknaNQAm6xHDHZIleSPmJ8q/8NIEH+1jCd3q+ITM2bGkhdEgxxLp1mVhBqHNC3aH7EGlJ0cIddzp
u/yxfv4nfNJ4/VOXmOJ6QGjr6a6IwdUeQP3tSrsjETS/vT73+DZZZ1PbD3gCcZ1Ygy0tYLiaAIRz
/eMLEece/LAFbhdwbfXZdtDb4fJ+stSt4l6ZhTyis7d7RWPu+W6CxrwZBhEKgugkb2hsLMNVI6lC
Ldk6WDcksDrkPsqZYoM8p7+MyUoHWyTcw7JFQIFWq8AFEQ3d1qDfYfwZV48cnvSPDFuXYqlwkbqy
8S9TLCW47DuLJFS6WhR2/K9yW/fH+FNwOZpnusH9XKMPKF/ExStf2UKcmCClImfYoDq56z67XJuW
QsoQKFKbQUxsB3HdFEuNyiguoYZ8GhrVxvda/1vf03t0ANhI5SqJRAhsvYUvq9QpSaORXr/r4fpB
FyyTsiujolBhoiJbaLtowcjN+dRTk+f5MvNA7XoZr54TbGVtxSzVKwOMy0HXGHwGNN0yYeWaoevE
aDi1PPBotNF+/UzZNnzJRiBWpUFppD/tbTeXC1taMiXF4TQxiBBj2AcLyuI04kmrCuq7FIp4kQiq
bB51jWvweTcq30V1C59XtyrPojiBs9yQmqRQLHiOOaXVxowKMD+esN9LEG92Oac5znogB1jUjiRI
SZF6g7yEV+L1vQKK0Vw4pyJxupgMdsBu0/+SPA4ivN2UWJqp/J9Ar4owTitX6v86k1wXu160Um8F
WiT9ebkFjgCrBMpYf/8FlvDGkGAGLeJkb8PKJdnv+elafxbfjoVmiI1+okRwTBO/QrNcIHpv5wgG
1MBqbIccK9V+3p5j/k6UAncKP8AgmP1LRxAch26rHUPk96IuxvdUfktxIo8Fshc0LK/DvUzCKOZ4
ebxf0kLWtW/H08qha0s3o4ugiyp18fgHUbZSqNRm2UJa0xM+sirtVvReQTfa/BDV/ZqJpVfrC/ET
Q5F/L7fTJJ1qVacwZwtQNq2n0Bxl4koRHqLvrs/Imw/yA6SEO+Po5IyVn1Tq3lkUUaugj9b9PDdV
eNyEjkX8mujVU5Lj73ZMn4akceq8h5Fxp/F8+1SFZXMv3yPbmJS03LnVpsy9oT7X3soIGNh2qsc3
/UZ1M3a11lKJZHDnFrWgRBWPyIjAitFC7weMsjj7gpHhhKF3i+g+yoNbLhJKkcOZ7KiTqDXn9sxb
jCTBKAPkEbNnNp7Zez2Be985bRO62tiH7Gsh3tjau+DIoGwHToMMHt4CsjohXrRYJ5G36g0hYDZX
+dIHUHA+eWji7PKUCR3pWNbeOClu8AsUgStXrjMN37IaGJ5TsnM05UVByft0BZ+a/dVy3dDAvpBL
GaHqjERIFrI8EUwnmzio9ApdC0nac2zO6xFpJg+x0Y3MDWPwhgjCYHzrlKJK7p+0qzEFPieVjmvT
oVefJZ59gQY/UnmvW9bsldSNbIr4ClI8Ug5iVQhkpiLaRsEpOyS1phVgfLl0x1jT0XycvSLAPDeP
b/ni5cWHoSYH7Tb74FcDg16OzVowH+i5X0fNxNuWb5Wl2+wEJKQGcjOrN9Ptf+MrkWzNYo7pQtKN
8lyI2fZpiqsisKRdKnPGS5lfiaEHqPv/MjBNAo10SVUrDI3c4roZiA0LDyqtrA2pZoqBGMRgU8yh
K7ucLJbXJz4ptGa5lbj1jrQ33Gdnr1Dt/EjrSJi3jrCi/HhZgrZfY0GpJJaq+RrDW2w5Dz+sdkHz
QvueDLaFz7JN9HXP8UBSG5ATlVvlhblWjpl5OUbP09qqcoi2897ArlCDwK+MBgLrAtUiPlJEPjMd
rfJ6LIwl+G9NT5RXX+nbDorM4b4HG1Cr/ABbd6qRLpae8NkQgbWXTB6JyuD4rnmEqcc4KrLKoGY5
jSUJgyRd2f70Tejinl96woHDJK5jh25KwTy+72eUV6Qe1zOtHlW8RjHMyvt9tRJyUQPJIK0HxVZc
Vl/Sjd+9NCpeyvV81BRdw7wZR0NbW8hWbOxHoG1lg4uZIDHSutoPEVjiO6VbYChmpDBmiSmBdIUz
WyjVdb4OOjmsFKBAItABa44LbpHjJjoGO2wbXsyVnyL5d9EV9E653E/tbInZQqhInFmaIC/VQj9E
KDdxgvOHlNzEm/fyIOGV+O7cP3VC6KXVBy548WPWas6tUCyN/Gvu/vZLfIvszSbQ5sj5RmZq+mQg
x1CWJu+qEiZiybikHxADo+v64dDCrU3CTju54qT6OSeB0S8RbafH2j5yl/4xuVrddw38z2v2+lh7
wTUV2I33qnWL4tihZdqJEEkuGnVlkkZA1Velytg9iOwkxwgK14lbIk5u6YCOkc8NzRHgppri7rvA
2avpQGAO/Yea95j31xT/T3WDow2/ib6ONvGj4tVFf3bQzdJ1nWscls8SuwR2avtucJynL/cC6n8V
Fe90lVufkPVd3WzYofDWCnmz/ig97jlAKGBrfVoY9HTLhd6ZanxEnNDWdRu+8are0HlFd7Y2zBoQ
FNpbtV2xrV3PirYPJqjn7EmJBBLnoy5YUN945UwR7WBwvRUZjj+HRQJC+hJqfrI4pXAAIqsyZRif
J9dsy2F6x1KeBhQ5c/5uhB1LdD8PCYnL02KOGbSWJQbGo6c1cg70+1o+jZ2tIU/VYiPvfwPLmlJr
FIs9ZxCETTpWbBERS17hRpwFPEpfl3e+Vez7Uygm2Ct1z+GAyqZC2VSRiFaHR52osWpKnwe6JXoI
bjgeTxcOSUdAMykNykBHQQrNT6ABtqfFHHugu66s7Jnu3naxFKJMwUiVzzRZH8BWHgYwpzRO7mRk
Addr6O6ADUFjkX8ayG+KyHhquusjrM90Bek/RcWS0BvW3R5ivWtmG5jqQlI0G0ocPiSJY3cxBaFY
ORCH0DmvjkeW+5ox1Bw4BQLjeVwnW4oJ5I4RU7M/zhUf+bSGA1d/Ah6ytfxPZmET0CMRP6cbUEzI
4Y5OfOxs4QaWGu/0OzZb95Wv1gCCCGkEmiLetq88tALM31y6FbgCXUeZESj5Rigk9EZ238ruJ2Ra
Wc0pu5bsZuayPTsmcvSr2hKpQVBk+tQVGfiqw4g1zh3yPFWhXD6CdH0z1CAlaafDRuV9Yz6ACJNO
QkrX8qZx30RvswQZ+M5vZ0jVr3PYjET/J5YLQGly/fk0KKl5CrvEtuQVYWx4uH1LbnRruF1KiwJy
3/Vf8v9si2iXJ2DYKmJ6IEyC9N0ke5g/cMA9ylWVZo5XYIX+Q7+QDBYJ/SvpuU0Ox9ZP4n5H3u2Q
pFTAK9fnbX19VZnw3VHOQ3I8kh/O9UjEr43Em4A/AgpxRBSSGuXNzdTnI80UGGd48TZ/hVsBryRQ
QFo7n4p+nCpShlHK966ApQxk0Sj2E6SJl2lf35/8S1Fr4wAX0A5ediEtup8VlqllnctpshQKRYSc
QBL9HuSDKXmQ2JCvc3xNg5y/w/Q42goa5GEXgCl/EMOIkYp/ox6uBSgW0Rz0NwoE3WUv9iw32rmj
HFCEsWQhiFZT6pXTVy1m91WPl8zXbkGS4peqfvJliRolxaA3UNIc7NCdcF7Mq5u02bx792HhBNiF
iGJyVDemL1j7ZlLKofwgymy3NQzSX5zuMKjTrF39g2FA2zieslnRmAYrjJ3Vc9TtB5FuD0K1G04W
CtKvIYh+dMSFm6AcsM2GqB+3S241/UfwZVGjczp4IEcwbhsxE415OE2tVNjMR08zL58EpfL+JEQs
WdnO+zQ+9Xm7iEOm9gO2KA2vHaA4ehasdeoxMAe+mKQriFnhY4kouQxEbHBh2ejXxSnCrb6B8ELj
TGNCs5LLJrbqXPxTY5VO5pP4qtYvQnZBcSc42GB0oEWhCyPofwy8Xd0WHM15wmlxHJjmbsGWpxg7
Ol95lGOto+Xq0s95JV21pUYGZYnyxPsUNnp+9bN95cNWs3NHSYiQzgmgdYA+Pq8Em4J2i27b0xRa
phguF7yzkLgIxPUqiwwDqLt8dH8UdPLATmIzJxOZ4sYmWOyDnejdKHpDom5PHt9c2bqMEEo0OCQV
b3N7ZutCczr11T0oV1igHENRxXROME+Wz+oGuTkJEar6XI9EkyINLdLASFFCBIAkOX+0nvJwVMRL
qYrtT5z2NbD/fO1aULZxEFRd3vNU83+g+wjkHx2p2AFgr5mR1+1E+63gWK0/xwzx2naKzbcncEk6
kJHJQ1JFPTT4EH7d/AO7KzRZ/sn0r+Ssmocq3jNDk5El33BshNBkulqq7DUmfjZgeOABiqOnY3Cg
aG5qsJ3wuMVFbJTFjK8aw71xU5tImU1gLUkAyDs8BmEqKVH39QpPoYTn5EzJdxdTLg9cf4PoMNH7
O8Ck/HMawZKhhLc5ioSRgY2Le2QZYeS/1rXJwl6zsDaKmoH+MQKHelWNfbehyD6rZdU3L1fIWyIa
Por6D9vlD03vZnuHzb+Od1KDEQ6JK9pEwMYt4fz5Bi4c8o4Upe3L8rzmTBTjVtgyhbCFXheZEY6p
M4wZd683+YcgmNhF+cN6nFo/QCfVdsIJFshRS3HAJzYTtV4Yme0369PSZ0diuFoMYDbaPYH69d5B
1HUCq8lJSS5p6xdlr/nrAXHGkWXBv9/NlxKLcU+rHNEQvNNddGD2NHyt17Ju77nwcMg0Ui7C4Imv
MxhW03gAikHC5sNMRy1gHGY2l7UdWRg3EtDvFY9lFN2gGeuBzSmtTjasSmdDKYKNo6NgRAKDUmuY
RtYLXJRSqfOyP9DU7gkFKxagxE+uzOsQs4PkcHQ3wBmXBoIgXjErYI+76deA0q7LCoUjZttbACQH
6/UV7aQ+Vf5+Gn+5VmxnxJxndU0qpkiCbJaW9WtrnOMHFLv2ecEjmem0wpgkMlzKnpzIN6Qx8Dr2
qtz54lu11yV9zxnUNI3Iw/vxirdBzykg2g/E8sSt+566KVVZ61P0WiCvqWdQOvYApogM+CkD9nL3
JewSXmnoBLjmY1T5O/4Os8MdezMoVODq2uXe54ynomaSs1VmRgwvbd0E3snPhmHOfBmc6e1TLNwD
EmwuCiHkUwFrDaAreFLuUYhkqsG4xIPmB6ohhkbe9OBs2OtwjjL/e059PekP5vwtsSYGvPNFpXDk
bK0wyTlmEKA7O0y6Do0WkQ5+ezZ3VORxO41UOt3pgWqx6yIVKxpQa6qMGlZv8J3//GbWyI3WZFLE
B7Q/8nsePja0udZZ54YVVPEyz2Y9l100Hdxtc4lEPSgSErZCgzvEUp6V2jzv1Tn4lvoirvoJjzDq
5bnUgyCnDkiUvzPz01eWu2kkbWk3AgADXqKWg99k9DQcSpU0Jvsg9XzcLI4p0FBeYcmvCWJgoubM
iSSUB9gi2CtRuVb02OAO5YgM2J5eYEjVhjAk53npR9dCGXQGvgGlZaNFy9vJz0dHaXR2l9ewZ9XS
v8M4qOl0VV8CUU5Z8a+9H6DM/Zp/Z32lQHQfHrZd/Ltpo9th/hAbHnV4+ZUlImAFnP3s1cvoipUx
UDqqiaE9iGfYwL8hd2o2gCcOkZjEKyPq9LGRd9tzSBbwx7REp5s2kbDEwGiyhUJCOntcodnwqkKp
U00nNaZjVQbhgfX52Vg7OxBzvIO531uiMdC0wFPH+RKwq4RxWAm/baHUN/9I422kVVwl2fiCir2c
AQkxWusD0Y/9aTsUX4H5wY+qcuwt+nlzoXAOngyEDyiQ/zqNUcMCaSK1eS9z48NHh8Hh7v3xQgAj
8qmv+mH8pRdexK/5h5ALKCKsUtZZ0RJ1mlbGtRBzfi4YWRCESw/6rf0wjIAez6bluL8Zk4qRrokx
nWvFTxY/8HLZhmkNVmWEckwvaxkMY///IIKDk9CXnS621FqyD5IY2u58OenkEvJcrVX++XiLuGWL
B23i8EEudiUqydmq44lLXfGAzMOnXCYsQWHv/LRsgJpYoO7EVH1KF9+7gKawN0cn96ExKEmPjjxS
VLV7fU085igNmOuKTFJkkUDen0H1YddnlowthnRaXSenta7lhK/RFwZJhN06FyxHUbyy6Qb7VlYo
fmdPSqTbjC7FG3Q0+Jit4sWzY0g4am6xBfsCULTi2lsvB9QImPBN5b8B/h4B0Kx1Xdza2mAyYlwa
g7SFv+sDnXL88iNivWtoLj0AOePSPWi8k0UZA19RI1gxFzgbzzOzGgtQAN8ULUpXHXgP7WJ09oMG
bUvtd7xB+sceqMt+/BhrhQqgLGaHTMUL84ON4EiOCmdY9x5mifReiJ75JlTzOsXsGjCLIuYCgxU4
U1IDVqkJ65TEQEYNeXLC5c7IZLoQVAjWx5DmzxKuB1R3J3/duf84eugY6BDFa59k0fhDRrK6XXSN
63r3IzZy9Mi77yXhHSlkoMchYFoW/9YipBwxXcNTS6gv+BNoOYks9hm+plmx3NeJroTvKNclRD5B
tzSk6IYWjsauz4rWhBAYBXRWKby5hhzvH9nEAHIIfFpWg0ACr83kt36rR6YPiycD5/pdWY1J8zXL
lSQ/6OSzqFPLRGMH7HwkPDdROXGqlWmgrJvVUkh8r121LyPIjefBxXgWg4AcSTFnn9WYmefct0V6
vImPJg6g1MKRjQKDQPA5J/8GhBw+uifkF+zWPj+DkW8vEk0p34g1CAwiLJkOiXEGacSOpPjHDpbH
Gvg1K93+EeFm9vQ+cqRdzTPRXTM/pmfn/QfZFLQRG/BwCs8x7IxnX5dHiAogolYZ6UGH3iLFiuco
8N4VzwA6/KgttJSAxawGOep7vRhgD4lpsziUqi4JqhAAKuC2ymTGt6YShqdS8Q7z7IOyKGpUV/EO
yvyaHFq7eqZ7fEgGppi9XxFbojXXOJevTE1MggrnhKlrrVb+gn5pZso0EwB+foWy3UYgDvSes3VM
aRdKODfCH1cW9z+lFA+1wbfjEQuDEGsfeV9ZAPcgceRZyMhcKlaHbGOprXczeyNEtTCIX8h6Tw0m
KQ8xHrC7YDaud0Nvm6xpKn3jaO6t638X5n7gUrSFYe1++O4kKmT8xxYCzx24Ry3fNGsy0oLK7V9V
QFMjwS6XhgDqclIbijrsxcpikVMymnKtaRj3U/M9a+sPiy8y8wI74A+B7fNk+Z9bSjiQmO/mkKLH
0/1DxNg4HqqIpYy1YnjkCFvmHx1IpXppfKowduJiUa9HsDnMTTd1UaB11AlYuNiLKt7es9wHq2I/
iKPq81XoOPlBqBkxpsln6ff0PwOyBKZonZidxZFnuTLtBTqZ8lIeotT9FJOC7CX+RQsyCsSG1ZM6
lNLG2AgzyTzL+wjj/cPbpprR5aapenPtVhpEFvrR0woYjgxKarOdxLHf2SqYmIZekJ7kqm3ONI2d
1GhPWmEv5ChbwZ5NAr1YC/0RBt8DQtOuYsSatawePFI6EHOAczONDUco0Gdq+wDy2r/S55STe2EC
fuidPUlXFIM7+0E3xH1ikv68vItVaJypovZ5ag9V7JOMnP7yr3oq4nyomi+xhbX04NvGfkDKP+G7
aFhHyAgYi73F/uP2ZQIlRzwH779kdAl5mQqxOsdl7GgjTpvSWhKwKthIKIclYzHy3sSFZXRxNGlK
wlsEr1vZi/63cyoSXJCZXRws6S7mAV5r9i5cQxVrbtY92JEMJOnoxtOSuSytfmLLO4HdkSYy3vy1
Yxar0vNlyGP6JEm8SGfoljRi5kN0P1jZeOLwrgZALXmG17TMHUOYAV9BcWeDT3AsWLQi9qZoe4Fb
fC6izpVa2pdOin6k6tUHHcZb5ciXLvZkjwvm7yXlyRv0ZZ01IquUt04Z35Wl85E572WYCQU9JklT
EtwczV2toHY2jzPsfr+08bJYkGuz8+pu6Y+0acehJLlZ9SuEONskGGeHsXgCUiOggtjiVAxhRmWi
0X9+5ENU5+OIfO1NvNklWVXdpURbpKY4QxDg5csvYM/QR76fUYBji1/N53gVKJlHizFcCLhW1WcB
TIqhHEzhpnCBgd1W0aKhc4oTELV1HQGjnTmF6zJxp1+W8XQ3M306HHFUmm66v+iw40b4Uqg2jVPh
DHpH2MfUe8iFpEBt4U2SBArKVTkVZvePer2tX2zSvl5PQ0vXMFaQ8AjZK+BSWSkFkCo0WXEkDGPq
QAgQSmevcuOEdRTfKXGCjlPGGtdoLneYGmxIYqsTzfilRlfCimwj8//R4gF7/JgOUFj+QKGxt5Ji
1MHaARf6H4EXp8etHlxDM+3JDE09nxSMqV0I0xcZ0QvV61PZXse3KelrSULyzKRKgL3XdbUeghiV
iOY/ZUk2gD0cC5z/9gsWWD4F6Q3OBzSsqt3zc2adcR8pxFJgruWEyVbcI/iAMAgiDqtHBOGHvqhx
qUVsCINw2RYHN+4WOThqAlTwLyVn8yag0m71Lqd7amGqeq/uqDbwM9RvfGprlSfww7ZzDRUl3qM0
0+3Eegy+cQEne++9XTipaDiceWYUhnpdoAFeoYq6DY51sgmTFejXeJ5RgCv5lK4SHPNbbBg1UHLC
cBUi8Rec+AOZcVyPWc27BWt+SOzhPsvW/v8ff8rGTSJqSZHhSpYi4ftW83pkXBovpHNIcEFo1zkf
v8namMYWH9s3FHsX0hDtkQ/XBVzdoTeTub+UH8lHvBUnYesKEyQ9aYrIWnHby3AMK6fJyzOQ2BvC
l+s6TUGbp8pkRD9mgyWtfSBIYBg1JHMR5P0dthBfZPPh+vVjxN7xQD0WbN/n9UuMtcJyTmW+JVbD
WQsKgYCCTOXTvMRLRC7Rdm2b3RDLXDOcz7d3EWnncZ4r/Sz2vWTQ65+dJTYAxsc315qMVBUcDvso
Noy0I6tQK0xv8d70SDvp8fZR1zBVw/Ord1hUYH3jW9fQevEZSA/7mMZlGAyqLKj6lrjjhZt7zNED
o4rv0ljDvX/TAl9TO+rCon8U67Np63nMafmmCeE1uJmLd7GyC2xBcO7pg9lNND2BoIrhH/RMn936
BPhUM2tvX2nQGcSA2EetoPjlHMs9t11HYcR3E1znX9dyOLyoNXpg5tNlFtQL8zFtC60K3S92lzSM
Hdfq9Pevvt0fZ9aRapAmf8dR9EtTEbyJeBsIeFzpVL86Bq27n76lqBvwH3T1k5EJZLpxpxsBDx4V
RqcyaUta8Gnhk6NFnA8P6T0h3ZPtMXm7EMMYntGjgrLERFe03+2KncfnqQaEI+rQGlrIwC6fCt/n
sMn+Prn9yDY8VGcLFeJweBbrYMfn2Ip06H+KjEwt/oZEdZMJd+g+XLPG8M2Ck3G59c+vgEuQ+dMD
VNpFvzkNb89MARRGma/G8DufKSXhvylZHT0OAIoWjYe2oawH4ppxnlyyH9zSxSoWvpRDFctUkDYy
1/gpWJbBDAnUiZuIlTfg/3nldBCBjB6bu8rShjf1pFpTyfIje0WJflWBUEKhGTKqsrmJ3pH2j65L
RjcpJI59C7g7aneeHj3RjEU5ETGIlXHXBTLp6FvLjkuA4vpbWFvMNfCDYEMgagDCrN0+SnHlFOxI
vOKyf435H0kuwcAgjlQWwr1UuDx9G7/xp4nrQVKIkR/fYh+nN6jWE14BZ4W7JmpTVikxeC8jaJeT
RY9nO/ijpo8rKZjhF1CIEDjZtwhGElRwR2Ud6NBiN9zKJ3qiniO4tw/Xvm90zzmm2Pijc2GkiegZ
154rrYkAWTtT4MvyjH9brAPwlMuML6o1qdIvx47HWsy+k9Cg/HVyjJe6vkYx9ycvNoDyep5O3FFX
Mkd3m/pCXsjbyaztdjHyw22EZPjSMxW3Vpk2rdD66Cmdq1oww7um6VdbLE3vy5GqKgsDSF1cT1+C
cCpc8zlrHDi50ll73g/dwmpViYnqWLno5rL3+Rm26lYy8+VkvFI6adaa0RiAUs11nlHyZeXui+z0
7XMFjMCa3quwCszKP0zl4gsyMv1do5tNlDvsBWbx7uvjiakTZh9hqC7LARpUFiGuZc6kF4Lkok8Q
sPQkr9qQle1SdrcUYOCaqF3GehvFiDoLKCIO8UAXjMSNSsjRpqcBov4dGN+YGddjIfVeLVwkqevx
Il1J5hI3Mc90NoX76KedR9YX3okUeJVXliDmcWdz3NnbA9TIQYVD33AUgiqqygHcNJ6+N0LowK+U
7Ekg4/yfPZdGQzBswjTxskfb3n56ulTGCMMcIuzbO07ntOfbpmU95qGqHgdbeFsx+dTDAcVZtkFD
dCgddye+SscZ5r/a62nLji8b82U4wHFlI3QD6vXyfsEi+jGq+uKF83rLAtb3HfLwZbgNenDRT8vv
PV1SRoX3FTOGIDYCfKo4TnwMaykVa9yI3EqFIRWJ51diJ6PrR7qCqlUGGP2vn4fCw8oAe0jfD6sJ
Wkl2SBchcopIRZIGQ2V9z2hFmdlw0y71Y47DnTxcA8BFoUnnRuMyPWpBsb92bsGHC32pOrG9J3rU
npaAjPliruORyA5GZ+36/GFgPA4aUlJ2Qvnvj4m7WVsFcat8Khrt+O2FyoQfdAkFAHxmooTk/NGo
2btJE2I2KagvlXwECBnnIWCTHMFuknmLb6v4ErIaI4r6Qsl6tFR1bI57S5bl/yoHdPaBJ80vMrJr
/3Efq0xKCbScp9ez2WEprRgxhGA7IYhmF10UAm2tYrZ+LtwgNC4L5WwxhWWM1R/xnBNxHxPOyiM5
S5vRJLIIJ6Ph3jj6TPgn7Ck1MvaDTPiaHtPZul413PoT2X4l+e+59Qf9ZALvm3WH/skaynzknzrb
MjThNDK4IquVzSGHBkGSJT1i2IHhRTkY7rGfiIEHBsZsf8dvkF5dgNxdMMHzRC1mUuZ2f8hhcckY
JJlb6nryyy0zoNX0JpDWYfS0xBWRuvT3bW4DIDDja2Va5vBcfOCL7rGzbWhF87wLa3bmr0RTb5Mq
8tABiDKpByYs/yPfJG59jD3Pl0LYHnC8gRodmMaFSTZxY6g9AtjXZgMAVW4PZPkeX2v/EFrkySWp
kV2JXWdCo3u0BXHdPo2Nb+EVgbqLXNgdUlflEOpruHBWyx/uZbj+Yds1fbg8b58J747n42aunOmK
ADwV6GtUZrdSueug2nG1GW3sJmt/s9pWq+8s4W/KOE0Mfz73AwCp/097aKa2RSf+VRh8Od97RTbG
2fTKz0ZtWUq71N3xIwik3AGm82eoyzEBKmk+LWfnZNc2uIQJL5TaYWHww0GqbSa1AwLZP7YWPHxk
WvUIfJhNapaQFziHi1dHp/0PolGL49mXVDeOeWJnoFhpsWnwC+gfPLPzOKRvRo7gEN1x4+v6BUyP
bZwJjmdvjapso2LaLVN7mI2QiyIwpCdPyq5k3k9Yp8npFW2NnVM/CDdn1mcn7FfHd5K3m7ifsh6P
hltxhjdvsJZkjYd8hd9fNXLiVEMClpXnz64eiyd+UiyJKHc3Ww7X8UGImuLdY5q/o929o95Z1p/c
ilSDqtoTg4udsVVhJl/q6Dn7JTgZ/MktdyAB6fwI7OWtI4CC0KZEcY7aSITz5mFgOoenP0Pz9A7L
MOLfSlh+vrroArgcNlEiN3zi9gNy0AlkPTa/MiRLdsm3zsrMuMxuFHp3M4r5ixpG41cpCsvhCm9o
1UL0pAy0qvXZLNT1pk5ZGztzR4UWAa4L1KzMY5Eof2IarzvE0GvvB77od7BndlTVy3s5QaCQ7wau
ZL0aJJjE3Rimy3t7u/CZPZ8OfZxa6TAR7wWP3z1yT7je/Ua3vzte3jbXbKLVYySjbr2A9fAKB17b
nCC1+cKsukDNFet1+1DV+RTjWGoa+1SmyyXzD3wD4a1En1B1MrDJX6YRIBGPUyWxBK2PDx3eEXMM
zTVn/XfKt691immzceK8fD2FnIHUTqlGLe91b04zIJ6AsVrHlkZp8I+cJfWyCTkxstvjVqR8VgCq
LgaahxSaFZqYA+XR1q81949QKu94JMgV50PPbPofbrC7UeJhx2w0SIDKsHoyyIYdLQ6eljEvC9ng
6JQ9/Pi+BzjdWSkQDblRXY0iYHGWFTe8/25bs5Zhz7HYjBlfWcl8G/9II/q99C80UmPkSreOd+pO
s9LH9nQodAS8q/Tk4mXlBp0LVWEkelwzYYPZ8HM9rsiB2SKqHzuayxIcbGF7t9Nu/DK9bayrH0DE
Ns8+4nHUhWkWxSeWnj+EpWGS+yIjcwG5EpQT5UHz1wIo+WfpIdWYM9OZWDH6NLhwGBMMNGxmCtDH
bv1ZASfssB0LwTNXo1BiXFnco9DdTe3FYPLe16yk4zy5XpfSSvsJ9b8n527AnodyHiz3WTxYW/mX
cTT2bHeKLcy1jZNxw90xusOIZHLECbTdvso4kQRr8Vp+3JY4gvja5L4iVF7AT3O3Ow/NgGdHnNfi
FqY5rA5pKdqgk20ThDDqt43d8GjG4mbv6U+b8XJwPj43zYMdF0mk8a4h3uenFdx3Lf4WScrTEfJD
+8Z+Le9SsIyFd1dm7+rgmLF0JjSYTemJ8OHWU/V69OX+633asWSefWqbTfPRnDYMBTyaqphD5hjD
7knwuAvlxSTT1SUX8uArtnwisV5v0HVQuyBhkQC+kpQrHV7CEPsgVpVV/+9MwZGcZhVUJfcHA3rb
DbNjLhJmnNcPhzvoAbKd+ZDsVoEzmSfOdSvALLYfBjhGqI9YjSt8XbDZxzPWpQuTq9ctsnLmvOun
VKjxC6jAO39aZhoYXcEq5khG30tAsEGs6Jf95xk0rB5XPymgXLr1MKGyajKWEIQ2ui0SIh2R0aDn
+H8uahA4+lCrQRSo3VKlGwUtD9KyHXHvLMBemDMQI++K9acAZ4OxcLt4st5PXTLzJeCv8vV426Yi
0S7qrNB6m5MIXvguF0jUyWsammoqRHm7PgOeHTMNP3LGQPTpiDS4WCO38CYnkQHKdKjoHOcFUahB
yY/CIDOBr6SBVnmAI0xQoIlmDlQPi94yTh0+kbCSJftp14Z2SjxcUDf/Sj15vA/slNmyrVnd6u87
6q1LKHnBGSaQrNva0/JfOt/52HvQjjdccRXFnHkq9YgBQ/0EjdEWT0rD1HVVXlpK8tDeAUumxAUd
LmKCBVAU6x6/fM0J+ZPpM4zpZY7+QisYjA9gbfZu7UM4+qCh3iXrK3if5/lT/J2h8JFn1HhFmtIY
6Ocia1ApGEdc9p7/Cze7a+8NzK+QrSvOgIKfR7NyVNFYx3zQXFdw1ezX9OBOBvnThNWMrxX1pDBL
2c3wBf68GNSFAybVxEiiGljc1Hc8XCyjog1DhFBx5THsxzSvWojhNoh6NLVs6NDV6jDXHZNsGNrn
gCktQXlIce07RRAxPUal8sSYy3fCYIzUp0YBEUxZsViuA81777a48qWNYa3ffMCfR9Tqb66jK34S
xJtizKzJ91FBQxSb6VlWWorCTAi/Mll3C8o1T77EuEM816DetGTSO1XqoWfmAGnxuKQSXcOmxEwZ
S2Bz8vH1YRcocGZO2bCW3BRd9paLr+OyLW1fHkppx9ACbjq4IREnODd9qAcdA75U4DFKfvkKG2Pz
wcwYt8CJNMyA7/0jcwV6zZxhl8xZJfUYa+HOtkTxQ6UaEen0zQXktFDNjSiwtV6/wKXvXxPpqivB
zKh+8Cm5f4Pox8PcZmlvUHscK3/9IbS0SI4CBtHtOZv5sx/NoexrlNBplNJGiunZ/Hmlyet5Y4Wm
KsHIfhBVLkHnoNcyZOBRUmVcgiMYCsDa1YSyotBZ52H+39ZMLMKm1op1rjt4qs/jQ0Kzj9p7ibaH
PGHRzH+tvy7S0MM4oITgXZ8yH4O1FbqgdmFQWMcqCZwIcYj/lsT9pUt4+JIopV5rRhiW/yrm1QAQ
rDoonbjxxIZGYyUQ6d0Ge3CELH8Q33f1suXx1MJEW7ZGJ2pc9bUkWDbfYqMtRJGi1ZG2a7QMTUY/
nbBszT6I/Kg0+PEq+cEuaoEiBmrardmb9KsaNKivFk2ghtzA+7r5p5LjK7zrRfT9Th4CL5KIDU4U
TjVAWMlNHic9/KHo98QNNXvmUv+9UDBGodBvB7O5e5k5nj/XkWVtNnwAoR1qPnheB0GKh7oWtq8I
qwrWVrMdc0yUARp6UVJ2b/FgYVdDq2K2NAZWCFbzponnpMFbOq6DtEytfdjBeqMSTGHP0z+wIohz
TIrnJiogQWfOlxsNHeUlYXbtQv/cE0+OW0qrrkcOKesZxMsPUQC5qxQFFwsedHGHKIq4VBklGdls
u/Cb229HU5vmlaP6/3CsQFEc6QCchAqSndTS/pgmn/hW4KWAQ/NwXrNwqUDJJedELhYdko7w77nP
u1/LO6yynhs+hgCUmGL9sl1XSJzHxWsUceyizWAmairMvX3RHEzNncmF2rLe+Y1JI1s0X5a7u6pE
ZtrzntOYslpIQANCDwNM8rPsb2JXy4Fy/HvRU0EOxe0whx1atdF7QMmn0olJpt42zgTCl4BDmS7Y
SBpciWg29y801t6qTtHMOB8zLNsvMBRSW3BT8lefDuAcL+kghvesk/QLkVhNiF1+qkvnlm2hdnvJ
xQR/aO0HG1MH8tLE3TEs6CUYvQpgqYs9oFs0kPkBxOOQolrQnezp/azh+Nh4tFB4l9y7gBAQJP8A
tN2PQ+K6Q3Dqb9INfr1pFZaMnCaba8P6IGsP7xqM65eL14aV0ZQ5hp670gxMXOg17bxiu9HDHhrE
v0eceTnlCvsCQteXF0/RQhSDis3WtcWnrK9dkSF+rGWR0sC00S0AMn43yAOHgRgP4JvgqFbhvenU
vbLJXWR4Uc/PmdaHHBaMXzkiCBQ3HH1eEz1zmXCeDJJICXye2So2cMS+grnKIFX3afkvHLr/Vac6
I5/sAnlWIeQXbUG6GOIk19N7Ly9Qt0km4VOqnSvZSntUUiPLtI4fsIiCvPlnVA2D3MP2a3LVp7oG
yfFbQ1Quss3zGqaF9JqOu63QBe/DLo+AdhpKVOc4uKvs1AskebHPvwTd1ersiNgkGMgHGh+72Y1A
h4OlaxEdF5+9vsetLGFgjZjRoH72pOEy6ChnTgUGrfMNeISy6tWHyyb4mCKeMfl75o17NcbS8lY+
Zc8JS7fLIVR20KICE3/tEMthC58/U5EVdT17QAxnpM1uREk18bAMG9LYk3L1Y1XIBl1r+ag3EqCR
tERHl3ia7oEzHF+kXtfvoc37QEkbsYvORoM8emS0O0HCUCYvXjuo+2zeayLw180IFFVK10oIWgWf
7KjBarR8aDNU7aY4zZ2egRzPN3/66Wygq+AAkgIITI1xc8it3SLtBPGdZJc618JmqAgZKrzxuTI5
Qspo8YQYUh8bmTuJy1Fh+7b7aHF9fsvDpB5QLk8HRXY9jpjdMo/LVUfc92x9X/uZ4twPALhGJWLD
HCDQm6Yp2KtpZsVDRZYJfpZwrLUe2sQQC4GYPkVeN9q6o1Ilk8MWRefxWGRZe7C6UCX+FhG5w/Ym
r3ilG4Zkw4OFt0BMVmdCyJbligxeBpPKacSqejiI9iSTp2Aejy8N2T8Ho4wEDkjs0XJ/shnVzLMO
cNqj8es/tkENGk0HH9vTrrP87MH69JlAYTQ560dkSqiKYbdUZG3YkCamUqnTA5t/KxE1mtOrzYAj
UA10ZTJHRcMKPkytv/cNvXx/rroyLt/P1OIjenFwo1Xtvu6wcfJsSzjyaQ0u1j8N+gPnHg2Sx4Cs
LhdTvAmw0XWTiL4kBNkY2GoTJ0Hico2HQHyQyosXZQHYGOXyOYg95JQWFosW7Sn9TVcAHn3Wae3Y
LHrx866G2tRQYx/mFl5uQkDUGIZ9MR4yLVLMXFIYuegMX2/glq6+517KhFaJmxboAKJq/AXX8ekd
+GbyehuRL6+jOajww6yavsx2HoQ/0wrnS01nsTmf3sO0RgoCd6hbRJTpDndhKYN8EKlE8sQy9hCm
4Fya7OzQ3ExyL2tqyzIuyuTj31pRNJTdTeC9nJ9HnZwOq6CH0LVP2Ma/uFH39x4yNHqRtWChIZOl
PNy8aycMCNqxDN6eHP4ZAnQKE18f3dGgCgzzJbb1t7qC7C0s1q4nHkT8VxzJR56fQ9KJ5LjGiO5t
ORv6McjYlYDEs/2NQkZmiWw17uUGNp9fEijKQdEr5qS/Lrwdp/TEoGML2KZECDJjWj5SQ9VNKwED
yjO/Fn5aIRmQa9jU6HRiWEHBYkeLUt+3GtGDFWP6IiiObLbo8XZoOJLck106f4tQTyGFXXVYEaT5
1eOFC8g5l5GNOOJX48EfPn5xWylgfA5Nu6qtBWbC3X0YhfVVASy5dke2M8tZolrESO8h/jHbCms3
U7YuOw2LdxgJWa6s8BK9x+N7eRu55CnKTarymF1FOtFLfRDIPz9Kj3KN2JAechiifsRfnJuwMwal
gTMAydeaNMaJBTB5BlO+gEis6mhOCSeStfhsrAu06X5+w7nipK3aw5Xwt91WwIYuKRBMpiJZJCkP
JAt2oAmcuXvVasbThndrBAi4A75ly79+/rQ9brSXV5Qej+Zg00/3alIcuB4gRKs1Pc+MGaEQ2eb4
2zUohSUuN+h7gaQ3rQPbFZnm9hfMe58onZia9I+61WiB+bNLOOX5r8adIrdrYm035X22AeyzCf14
qb4E9UFA7brRnRyVFJTWazxRoabfZbXFZQsZmwFpoS4QbfYLSLsJTd4+rk2ZmDGV5RVHDo503ByO
ZtxXxS5UO+uvWK6w7LhmedsadJ/6oJvn1WaU33u3kVQOFVBM8bG6OJUgWMachvU8bWN7gK7IfkR9
5k6gocSBJrb34fDk9ZvsgavWpjiLSWt1QDqxCEI84+3UgeFEQiLaGSLZsajNNgMowOf7BJkH/4Ij
51j9gn5+oA3ia+Nr/4hu7nJWgLpCG5i1JWldi60HcuPzhrQIqqmZg7h5qKsgppOCKhcGoRKNfTKd
nG6rQeZNGcAlbVqY7i3VzRfRNHaRbGErISHMvzMFWSO7XXeHha5nssUVxFelmTPs1UHNEkeIcLe2
rW1Edj+ujOxt+i3RIOUcYqg4XJPBzjTMFW74YRp+enaLJUw6JVJTLDpsEggdWH1LDK6RhwB/BhXd
Dy0oLjUmF8P7esOQVXxWIAwXzaioaiI3h5ry26dNaiqy7jo9AUnAguRxZIiQt4J8+vNuPlcpyzmp
GUco3n6sfa3rH66ia4+zZLntN2/a8wCD3zB3h5uE5szw1f4jH2LUBugmDUlRMBneD6azPU/BB0TC
LLOXT6KeSOV3oDVW5hb29S+d23ZDhhCVRbX7etvThjb09fwOtyXrTos6zpUNKZuFRlxWrI6LMqwa
fjP++hqVlz/VDL5wla5GKjERf/2UxX/GxKFykWc/HZZjvcWM/m5HcuorqTdcvNv9oeaM2nF3xUjR
0GE6KCyHhFkVPGmvVGwRPv435xo9sVGxq97LbVfkyHsekT/Ti7ckJzLmu6cQmkdGMySdY70TMn8O
THdhlVRBz2Eo2/nW3KlB3XDmfvGe+yOxFvpTymSXbWZLtOkVcGVekAuWC8YagevMi18IY6QUnuhh
CbjxGpccuk1vkRUl2nUaed1ECMnaJHBJCVdE9JUCiiFGHCc+Mx29Ky6PW8Jcaj6e+oveip8hhmRa
aNZhDPINPET6lrAZ+ie8RRLNTtUfwnCBbP2kByP2qolqxYQ4FzrNSrYUR3pgXIjNZmo3/gxeDGcR
23d/cYxU0aBsnL16AO36mKoKVlxaBa3D4t0gGAl2JrFagqYjINVFx7CwQg/FVP0Vly3LCuaFpTZv
sCM3jxZfSe2ASj98Z4/v8FWHBpWuH8Gmy9sq3i5SbPE5zlxif1C0aaTV9iGh6522XlXZ002LlsdN
ygL8qOjm1iN/bhbEfioVTfEeMOyWWxU+llp2B5KVMzOMcP5/XtL0vTr7Dx77sk5D/j6V8EE1U5Ra
z8ZwsCJW3xt0w//Ti47MjhfTZJktHTTbKMKasCDsOJftODsdJ9Fj+rLHL5jdYUgW1vqJ27x5rkqK
wmxrCBY2jcW4/PoGB8lmGBWWBcXwOYwqHwc39McCL7E4XodEIevbzi8uX7t4zEPzl77oJaohL1rN
iwWTK/3eD9hoE9i96M6+SBvu9uARX/dBTIypGFO9HqVaL0msBfap3NhHwvwp05HjhJ8Bx+qKTn3a
u0pl7ektlFnSBYSKPuLy5QLw+Ox53kwSsXhFZK/lYXWKcLNfevN1QVyHlNmpzAFUrNo20PuCUAhP
MsbDOCTmnxHRiy2Il0EhvvyK7E70ICjESTuw3lRRptZ9AAjmIM38AsJ2W6beI8xec3zJjpoGqn4p
vM0afMQWKJMMwruPjL6+aIEAFMb4sl5Kmv474Y1+rYXsl+xwYoYbVs2koFUO8clJIMeKgkzR+nej
MXFOA0ZdflJGFWHtnZ23srZoItFlr51zreydCF9GmvPXH26XQcGKPDtF9dYYB1H3DKvoAqapnAX9
VkvAVi/E8AmSTgL59XhHDQlsRChGZVUqMz8oXSZg7GEslkSXBDImeIQ7WI+v2nNpGzV35lLE0ce8
kpCnox/2jxGEPEU0Bv2JDoPyYAtypMB++sr+UJ1Smw4jRFSOD2ZIylYvXlD1pVAlX3MTzJQmB49C
CEUlQUlBi97tX0Ge8tgwPFE1dD1Ptr+tJOobvD0wsUHz0TKvBATAsamQ8jNLCShOaKpDT6eATq8y
HX4046IAzxJ4irkAT86oVFYYLawcKt2EcM5tbZQjKhio7VHWDtOa9oXJVz6vzq6EwvyrU41wPZMn
uDHwfKrwtSuF/x9mD3VR+n1btK9D3+QPEFy4c+wskxlr7vj0qp2bxfy7vDCBGilKRDVS8Lc9AsH7
DmPd6aDD4KvNXJfSV2toc4ceisAgN8gKAN2mKwH5HPaEn8bDBDlPjF1ZZCTpSCNvkCuXZUdLi7Dv
FuSnDJ4+q3f4igyPN4B3io0+XYzaTOepo8o7aTGBgmvsiTTXExWYqcE3P7lU58Z97nQTkJN9d3A3
G7Nqa/WVrHSPrSsOaqbnAEzfBA7KqQMM2EpTkijKTEBOXHY1pqIODb3tBh3GHJLIzZjDwac7knQh
gzH6xWPpltP+UIWaC3tnQSgdfd8VsuXQc8H4aewILqGuZ+VDfxonYsLLPq2nmK8hkAEgAxg4E713
aEfy1AnS48mz2MO00jZERkHdrfORlvOfLpSdfKNj+U9PQrwyycRqSU+wdAUQ3/uyLnPRn+3kxuFV
DZKrF0l7if0gv/53iRmCBPn9ukquJgJHLKLuUKO9P1peYSgVqZv4lutZGn6Wv3Ym11/Au6IJ16mo
NXwrOyp5OmPyux1xPbUJR5vXW6pTXonMKxg2Ni7NrDRhLuKhVtkbTbYKoiNxUnmP6qFr5X7S/KU1
wX52gxgrmdRR2IB6pRXp7vpAVNXG/0tRl1O8o87aMgOlKQcGWOO1qU2m4UdWbg3s1hFjJlCQO/Mn
xUGlNEb3D2Wax/H2pTfsQaMxShJEUeOWn6UcwsUVZgja5BhZK36APetGPoec4zfLsHbaTu3/CxqR
Kdl2bx87+n9sMhv0JF/RSbsg5lEGtHFw0DemnXxPycSn/gBvnAIHAY2/sK0KeKy/YOXkR1J+tGrZ
+BVp9OvdEVA20DN5tJjMxsVsTnUn+SURDthyeVIJQIutazTdnSxM4qgd9q7pjlTK7SVwNnYbaMB8
lIGpIMMk84Z6QEt4Yb1F80NHRZPh6rIEqcpyPD2FOPlo1iShXHXdnR9bS1+pCEdLHzlFgoHEqA76
kh8BnVCz0NZDerxMs2HFwTyQSrb8Cxln9D7MGW6x/BBdYTJATUeqHSMOzMUga/ZFnhAzL21sSDBx
IwQJQdL7bA02vRjggiQMdcAkGhpa1ahyePnriYi09dh8SbS5XP1c2uP6me7SH9a740oZn5MFbe7x
JhPtn45JgZxtdfSjORp2vObvAy/ujblZ+3tiyTyJYDyFkML8ooJx+2BgK2JoogUQnerdYiXn2WyB
Z0MGRdaaFXvd7+IM7fgr6LrlgqXIoRQb+PuyPoSxsP0IXeAkEbyyC0U8VIz0kTwMTIfQ2TJX/u/n
EAcxARMco33pQlKv0liHHJwIgdZw5suRhVUMTYo69hU3Dcy2dpDvl609rcCtkUM2mSb/vMH/3Sxc
obchIAyjvUAvxBk+nu8X3UUdf4mX9lhtqp3DqWOxF5Wwy6pKJUy7mAqkb66xaGBl1Ady8Mx89YC+
OgvRZTmr0SsH4+j1b0OsDGdxihCNYlLVArUmkHv13wdUJwxih0YsHqTaHFIrVyi/Xiq9azcKaI2R
ndVu79EIXiCmkD/VFvqXfLbb/3qDviVlp36QinbK+ReqlSb4IXsxrIFjR4/yOBGW9W03VGOJY8d2
r1Vwc7n9IbtJp2hsGLFdrNxAOD68yf80RKH+qaGKyhruZNlTp/9nFXngJocx8Q5RZgyB3Os5xmnJ
p+jwD4HFL8zJkgxvcJ26/tpLpmqs765dX/xENcIhQqIb4cuVxdhC1an4m2PNIrONQDw3lVlKBCiH
nJGUJ2Po+CWqoLqTHmLLTloedImu8wjbEUbznr5Hx9k+cJIWFZ53rTJv/DhJVlLAEhxmieJ8Z+Yu
LfMcq100NluMI0ZgJ9uT9Hl0YoN9ZWMiw/fY+NtR/HckhxVYXmaHGrtZZMOfV8VEfIRZcvmlDmdN
Or/1SMx3xx/K4eMrdq6Qn3djvDk+/0FcYi8T54Do2Czu4HNPOANXfDcQQmW8uGo/YMyxb4+3IREO
AdLLM6KkpxEf1vXwYoeqRB15NBPIJ/UHOfbb35YS0FKqkziE2kJ8wqD0sdNOpjbxkvHfM1G62Y5c
9TrBk8QXi9HBkGF7MBQReCKyPOD+7wxqk1sCzs9OvGnceN4eGBoIfF0xjV/aZkHyKAkncVOBxHE0
7Y2CPmEQUaN7+6KWV/wvozLWy97QqOYjqsNGCb6ZiLIQHaK+jUEgR7rpjIicJluBi9IFtFLfPWZn
jqjg7Ys6/TZfIfTMJ7t+EMqlwUkB9VQM0deV6tC8eEbpYZBV9pgIsPW1wu/SR4BUfbfeUhh7snZS
wVHxVz/0P9WP2FwQGN0iKniNciWvTCxt96U0OU1S8Rqw27rkAS2xsLbbsd1NjXfSsG5nHuprQVQr
9okUbCprIk/V17LzkD3QwrssP9tbbU6xueJUPe38CGJPm2JRztdT7PK8e25PXCh8/ElpgjDrjUsg
yPZa8AZAzYfNa+tB1BP5O+cBymohCSHWEImrSUTtW/IeVgzr8pv8F2eSkjS0NGUMfDn2PJ/j9kfn
SlNjhBbdOe9OcD6y87NhiCYR3acIHqlJWS7P6pBe/uQFVVsGLYaEFP6uvU3+sspEjWZMhm8dn93D
UaM9D83NChA7fDnlS/g+LK95Fqf/FrJgI1xFMoki56QKN09jME9VTlrqlMYBihH04t97lf0PNHyo
ZSvHX6yve1H0G2HAG1cA09+kZgOYEJEN4VUHvT19xDu2GpN/gBMEXguE8r2bYVkosGVTmZLhpjOr
LaRyLDEKXQSY/KNju74DNgp2A8AxQkbJPHbpkSYvDZw4I3H3/uFO4D5qVxDlFO9PLFkyeQWCyTDL
gJ+69GUn8gvkTXM5vsERht/DDMZ6n+0hXqRnRsiUukq7n7cLaFDoidhftaXT/28vr/2CKAJgfP7a
i7ZbTKcFYQxccVpgxdkJkSvPdxWOG5bH4ejsWU3BeRt32Blb83li+5GFPYBw/PHFcN1nazOUoM3S
lxhnNjrghBtYBYI0zYxTSMRlIMXH/CgOdFFcH1wHFp/s14xiIy5G4kCkuPwifVkaHt8yghuEVVKh
s3euzFHldljquD4CGRv4Wx6E9x7+xE6P08yzurtpNpLi7o3ctkjOf+9DlQLwULLjuX9cfkHYaGX5
saX3vUGp/8UYMOy9+vw0x3h+QoOoAU0gxXpOZEI57GPnc4gL6Ngkn6t7eShZ1GP2koXglqaNDllk
wZELkopH8r/WiYcytoqR1QKTwI24xwvTGmby99S8AMblOcbe8+xBje4bJKK0lKumzVDKII5vtTGI
VpUUvuyxTl+tQjoa3faDmEoHk1nniropXcuqk3y6TnCn9pP96K7GMZKX9AHYTzRdBjUgXUJDELue
KsjDLJGhsWXknlzg6Ew2m6T8LBRs0YsMuDitVUT8Lc7v4hcxh8yCwIhp3uND0F2DoMfctd565SEe
SCcxH4myVcnpo/b0Sdvg+M+3FgNP3D4Wdinbyl/MAcIHDEtLHOivDp8JCcNZP5JnkAGDdNfhofVy
otEFJCxH3PpUhfEqoRad2IbL5xUAA2+/j4/Y64uM8CJ5KVNJJupHwQqR2bpohpehKycaV4fKraPd
lIXamZm4slFf5RucUmGHZlfI9yMAUdoNlmLqrHfapxIdUXohRgyATGxJFkjAHA3kKzMCm0syZ4Ww
y34AkptMIe6Zrj9ZCmfze0StpU+9e67/yOLZxUyNExU/oacMSmk0rOP3VkI+PEfr171NgJ12Prrk
OMEFjLDgqHVNvrunRy88xfT5ao0ZZiQy+XC5M9LWd9M8qWM8TYI6gclkjc0RhS6B4C0O+QmW2VeB
0i4wvy82lLeqJsgz6qpkyJ6sd2fgAGB3HqI4654+jgQK9jnSFAEcGKsKoeFNQw0Ahn29wN1E1zDK
39fJrpmmrw8lTuA4/9FmSaQ7m26J5J/hVJ+EqDZVXsDoIDwjY5hiVLGqdBxcHGjjSxPSJO0Yl2TR
GFMILyz1dBtgXEdEITtXcCsfAButcsvmIKQDJnRX3shl/Dgdc+8JtLXOx7EzGBglqx9TpEDjtkKh
+NwPiKlbrbK+cNMbzRmmZvJ16WmxtvezY4Ie4d+WGnehZZzoaJUmDwBD1WL4nXL7WZE5dsszczoR
5WSj2UUCH2J2TIx+6uyIayaLny2TQLeMyikDKyOfGMOJZ+Cbp13OdLE+RYqqLR0OCA2zI3bBc9w3
Ds3lQxrvFj+B5mDJZ897YXa1GXXLOyxLNvCy8/NTWbrm9LpvyuG7dqMFtJ1HMWKdBbiUtA2HIP9M
Y2mlNukRvKxh88YFbGh9G1PX/GwYKVzncyHgjqDI0PnLkphG4E5taBz4No7Wd8noY/TzGTZAYYVg
npMW0TDYKNYBOi+r0vMgXRnJqUXyIrEdvJyWMJX5bHHGxuReynD5B8FKSoypad9xGpBgpFgIg5v1
nAlZXJ2i5mLFrRqM1c2u65QAq1IIjQl7TC21FvXB4lwWeVZcVY7eRWZGEYD6XDA/28zVHTeTnhQI
RFLpNT4xgf23hZLR7xv9+lYrDlxeI/24i5+PogjWsU3TmnVG92JiBEZHpUtHa7HOMxmEQdRWBKTy
aAZMcPPAcOOCPHbNfNhjAvoWH83SoPqZIWTW5zCfpCoD92iJ941d8+lXdkgt1BuKq1MLtVatXZnm
G44wnKoGvTJIraGWEhJ7HrXLvVy/7bFE1nnTgD5eZ0tVN9Y3leVRrEmfHW2OWY9qduyVv8DkhiZz
0nJaGABOAcVtHWJUb+xwSfHW2mPHJ1mGVL7hRkFoBDJ0jfsdOq4uTO5k/lo33Y4wATOvQaS2IxKL
8c688X3CjT+N11y3Utimrxi19I9pXbGEf/lrHn/KP+r2XB/p/to/5NhX9uAe8nVBS6PxO+HfZlaV
uOwtN8HmBv/3EQKilJ+s2XvDeDZMQ8XCOFzLiYuJOUR0U1jSWcWhcNx/TVkDRAIVZCis1kaYeUyX
aTk65gu/go4wNYeXYXTjoRTU0Xjgd2tX7tNKKG17xa5s9D5LmBPJaOHd+0++o1+mLLCXz/oEd0wG
6Vx0Oavuk+BV8X9YgnPX51NVmtM12sxfm/hliDtluU8iXcpBSLAaqTEPwEy0TMl9ChiZni95cTr2
esSyKvKp/9nCQfFqR8jAqhErhB0n4iUkxUrZ6Vw+C6jEsw3e2wiCb4Vwpi7qLP3Cx5jyM9wGCfnd
yRseEgq52AouCgF64ReNOuuNTeXk/WDNqeFUYDITDBB36qpvMAUOMGU/pxT96zkF2xi+et2xFX8u
la+TctCksKkAbgoRZU+Gpr+sWXEzWdBfP+rrof0s1Cb54sPKSkCWd6divJhTZc3HSqnPazLKtb4c
GAm6MAGZWXw+4UD8+M7OrspqydGVmmA3q14/cxdgBlmd3V1550C+TKOTO9PCJiRyIOH3HsVwiaDP
3OjyyF6ZuYXGgdOXWgzxOQ6bywhiiea8wzhpQq5db63d3V26fe2seRyEfuWGP9rjBxABKE6by2Di
mcp9SB7wGJp41BccpMUg/vhUJSSwSTn+A8bDpmCZVbnuIPwRgzFyvpFKV8iroQKMGfV2I7w4xSsJ
Zy+rwGovvic+aBPpvaYgmHjdnk+QwN6VJOfB0cBvY68jJJLDPjwhnyecaIACdQmXy2Q9fRYzjiaS
f3ajAtiLdrR+r53W0H0qhSnVXImMnktz0CDEul2oGgYBAmfE7N7orPdS090BK3HfFRkzVAOMGiuW
WDOHzPqDdqgUYlm54yFH0qkeK7B7SYGEr2XNiaX5krMQktPcKP5Ulh7eo61A71jE2hIZR2yYAbfr
j3X++ElSi/tJsADixEKYymKiT6SHkqICjZ1ewcgSeSgks4xOffommD5y+diL89v36fz0O8+qTKaZ
zvTlFsN5Obs5Z/Zr4AXBxonzKgist7JTnU1qKurTDxq+6Gc2nz30/Fd0xIEGHk0dAtywPUA3vYzt
g45y6OOuzkkyN2z0RQ9CEntoXNMzS4g1Dxon8hbOcVjz25Bb9y6Yb/NWY4mb+EnDPVMUAn5zWdlz
DT5Lod6nLWLe6qB7TZSTWjBL+tmv1+MNLSA7c4ozyvAprAQdoG5xlhE6WwmquAC87WJdk3Z16t1B
AE/mr0l8m2r8QW5VWiskUuW0oqzjVJnGoNFD2LsQ1XVvw9QESyTBgDAOFao+vcedzYxSURAzbcLI
JViAjFuIJSUXBw/KaO6Eu4DnYimxQJTpbVDS4DHyc7nKTmz2d2REh+oinW0dbHERyBhNM8iRo25z
+p643qHYQwaUb6tHifukIsOdLQJx7cy2/3uUuIZSVbR7f9mbSUCzbgiKVa/BUlwHREshZ/0Kemqz
BUQt/EMaGLPOU7i3SnMSwtvqjuZXRAcdpMJmWpe1xQ2V51xa4RUL3RDE2mSx1ujpVnnsD3uH+31y
uLTLmOWqrlJwwU1+IZC9ApJoeCNGt+QHn0LTkZW74Ko0cJxhELsBTkdv/04MdfFQgjQNnfYQqqmh
dzpdyThh9TjjSK0tcDZP0oxcjbsIUciqliyPKFD6j1axJLMpg45Ci6lx3w6DR5CpU07g++s1l/sX
oPA8zF9wqRmaIqQVnw303DiLDv8GvVpeUvJQT+RQzaZ+QLExaZ/ddBBLbAeIhmI1OEE/DH8uyjGl
D4U/vyvDqo/GMBGxfTBss6B8GzMklzWPio/FQLWuHeu8hFZBkaw72gGkyN9vhBD1w7ICj5gZUF3G
dqGGAkzD8DNlWj6eZVS45CIdycIzPwOL5BylhHXtaJzn//CLSWTD6vf+5dshy88kSfxIkhVGsYq7
GOJ85UmqnPN/gLJTrnvsS4pS3ONH0GQMtktvndDOH2KGXhj++teJ7mMnmNlLqv7bp9btYtaXvuNJ
8ssToTkXWfGb9+Mm5glx0Phje3eJBF33SNkBZSab9ELr7P7m1PGPyojoFAENyxe8VJ5QYqIIXMeg
MtsZKV5UZAM8mTNxMyEz+c4yRBFtXDmjIHKKBWPmR+snX2ux2qEs9IxuHqNisMgXOWXODfG8XPrC
2YB+ehntw59ydDYVd9HQBmT9sX62kWLVU6yUkqigV62vCpulgoMAKNPcjwV97GBrGC47/AxiHGNf
z8Eai3SsS4GoNgunL32Ly/NuBeqqgxnOVl6cPI1KBzHIVJKAF4AdTERqY+SSU7sUbS5unJn+tRE8
C3PxyRLl7DEHcT2yR0YRveAwYxMezE5/Gvva2tMnu2vtbyf+NgQ+ur1wx59R7IH3CKmXDskc1tk2
y3jt0V1ntdTuQzcjCuIsjDeRwlXNlXFPp+2H0luIjt6LTJXWD7+GTMj6ZmbtmUrSBlVjHWd4YhsF
ywD69o4qfN4RO71Q0PujeqWTY+0z2vMNebFxpE1bjXevtd7LzacBRsEfFJ+ByIU/JlPrpj7vkj0m
fN/N+V/qUTigYPPVWqHWr271IzJSkmIJjQywecyfh/aJJOUy0DiPn9Ym4x06hnrwIMUcQ4roM/Km
lngrZtFem0cf77L5ZchHRIVdZjJIA3jVcU2vCbr1sLDtGP04lMfP89z9ShGE10GZzKojwzlIYKOC
Gq/19ni0mIJG28/Zhdb6ceznV7jKIEMsQOQUKlPUNUW64aF5j+lPJy1OD4fQQqFCPPZ4oSBBmwj2
FKhQKxkfxROGXb73TCFQ1oMwwv/ne5h5Mv9XqtzXFYjafri5qsj8lEK8F7xs4ycHPeseY46f4L0c
BdlyevKPg8nG5Hz4Hi4XLuVJjVIE8c7E4hew/L2lJXqzgU9BRo1kvi5fwlNva1pUfm0vRf1aqc58
mwDGor1fq5f7AVDGjdOKkNxBQIl2ghtkUX04LFJAklVozA5PyWPK1rS4vNEZhY/bFqPXNcYo2xzg
xVVWD/60QPYxnEDnHZDG3mYt32JYIrbbKzUg8FVO/Vhzo1ymS3ENVj16So7/s8NLNCt38slRC7kq
MlBj1I8wuBKs1J2LwGdHoSEwaWOZ9l6K1peHgITRqubQxv3Rc0W8rvN3dWw9Me39Mex/pJSH5i5k
eiTYE4Nuf5eS1wHVagEfZKs5Ehvb+NfAxZoiEm6NdAP+CxgYsIHtlC6DLby1IkRKq6zVrevZ7JZ+
8PteHXTwNP8nDnfAAZYWRY/WGOJXaDNF7hrZ5W2QGTaOLMBCCsIBBtiVOvcJyZDmhhkfbutWzOvZ
w6X22UuEOvTuOz+dh1XHmWtJK2KkE4dbNUyOr+jSidjZwq50v0LoH2vfjgy9hJ0fv3C9gHUUW0CS
QiBZ6pGVpZl0nzi3+ua/uKK2Ipx8euioT8Jl8FwSe7ZuWy3fBfR3XtJmMt83xW8k5zGqNCAQ/f7V
4J7RAAfUgwRySgxKSjj1HopfZiYEpkuC3f1imbYr8rGD/znTzW8JcTwOS6oIRJD/wajFiZ23kCzo
5RGIuqs3EtnhJb2E8fjJ/FXNxrLBIxSdOS4I38A4u6+icvcqL1qYxq49ez3zbm0QedNJtChLBhyZ
zDQt/cwAtQ2I9PM2zgX+EbDkahjbXdIJNduTjnlQ4h7hYroz/8wp9B8O8TQNT6+joMH+bOOg4/fj
pGjFNyptugFlwI1V4al7YO316hnTIeGAzPklIxzJ52NZyU+fAlNLEXrkO3D2kH0gHjz1gE8fJyNS
l4/c4Nmek5DqAV0gwytnqrEbh6f8I7Juk8k6Rrh6PYF/15biP/L8M8oSVNVRNrcPkwz3gpT6tzaB
UC7b7tl43giXS2nKrocZumBsw5tL8IeVmUArh/UrfiOgjqtsLLrdTnfQuv65/MmEgFHqQEsHXU8Y
+fQ9XdokuolEH7fys3ujiYhiddoq4vLopMUYwHZzmDi/faArsco0cp40zveLV1efZGRa1j+uqdSA
YSLh6q3ei3/QNln1MUcv2c5mLYGm/kt4hFU4iYJ5M3duipCus1MRNAZsVCqZZuagzNCHZjfRnlYP
rL0y0p2qRacIaMREpkuKjahp1tqQSo/87IZ1zsGyBPsamdDmfkZXheB7yikeeD+VyCwTVmDHnCgN
G36x1FnisbTQEC9Q2Lm+O4zoE2Zvzu12u5bhw8GCqzVltFIREI5OlmT0sT5vTOLeGGI+rfhx/QZ+
3n46TT6aKa+W+EhDOrfJObdVd5vuLRAuIHMo8Ws5WBfWHT+6G3ZpIrAjY8mnMNZukz9fQFcKvJU6
4zLLWCGkeD1NT7/0JASRCtpubWU1buS16n5XErTGPerJf/KoFYRWGMePHEe3amQu3u0GDdLyVyXN
cOvbC8YVFMzqJ2TZ0fm2abj9KDiUPUusJ7ibldjeNhTMeLuZFlcnuygRByuT5cxRIXL9/0Ky0hC5
0r/T/rzGLFM+3vvKXyjUd6UmQUTdy9Exp45uY2dItd04Tt3RHgbCya4/MhUM+OsJxcnzOmNeUD+s
P30XUeqWDr4MaDIrZETzsJVKgJT0YHjSEtgYj0taQvXWb7ef/biOKfr3oRE02E+Ou462W0VQ4oNI
MwyNXJbpatadMw3lB6L/xFOX8HsrzAmHgPbZ+2Gt8tJHGlhCfg4JmNvIyk6uWqB/2p0X2ubL+Lsf
2LXxCBkuvFF4WZhyqEDPsHF7+YWowhTY4GwqQvrGpN7nQ/RgmUwEsqm6CdOKAA/WbboF7RBJFE2M
WWmhIKjCXG/LaOX/Pk2uns4O01796Wc0wObB9/LDkYAFP1QtMEdTBE3+luWOq2am27Z+fgUrYRAQ
qapj9bb9ynCIh3d4snoqzytroW0NttW0CtoA5TVKqclm2/G+GaO89TN7vex4rDaWjaIPgd9SnX0W
LElX9YnsFUIdPhSU3HN/PTJw3jX1TukbDgy+wo943Bl6KyuvKdMso6/S5uuAxHgixShVp8DfrbFs
u0vlFBwzegMWh2RtzHi7PgYXyumRGSd0oW9UiVEGFs77MJewzlFWAJk0KcXlkMZXjmERatDyr4FW
ZNh2neaLc17xdhIBiPl5knguNqxHiP0Q2qWwWnkz6MHWz9Ud7/ka/GoFfJ4PaPPwia0fdbVLuko/
eMgstRUXI6AlDkCKRykFHMySWxuFF44r7tihv0wgwMk/XmhixDv3/A7/X4IAFVT++FwXU1kxYVX7
XElJPDNYqhH/q/TZM14CKmPvg9TOWvoJu+vmJvgFOyzK1o8glr20zMLjTpkysrKCzkuOlqVXMvrw
41rGhAF/5JU71nWaL2/9fM73ASF5SqBTpZGhBlJehZ/WPYcgRnCPjgib5KGRjoX+9wIVDy4fbOUr
Ia5pVdLWCu43W8EHwmTIQhkpcR3xZ0iNBbuoYN1ceKnk4w4dqonVd9PXNB2CtISiONQ8Zd0GrlwS
4wqYJLIhRN5sG8EjCrifGjR1qW1gRcI6aS/37VlR2AndMQj4y5LWPFe7LF5Gw62EU6nrlALuXwp9
PsFOasUIZnGsmYung0nMsELZAxjKOnUWJW3ykJVTD9VEjMXkZbCCstoB915MNMu+l7uNqplq88+t
LDIQ7JCa+yiDOexc3tMRFgoZX0EXeBrTPIcrQu+Hefy5vvwqpwpC4B8zxEuZ3he7ysxJCssP3fTT
OhBAQ7CYh6rW4sUadfdKVbpCWFzLT+eJSiHqJ8VQZ2i+XIS7GybSxqJztLLlfErHWuh/qBIHP9XL
DCHM/6zaCd6EPHcA9JdcJtyYQqFn8SB5OPIukxHQu6GdPrL2hgN6UAdPUdBXn07mcgMoG8krAD1J
XFfby1zFgR1s31sJxNdYmtaJGdH0/Rx4q3/IQPCL0Wgoc8dIPNZQVAddSgcDnc4lkPcol4QiGoH+
toCS8PpxNEK066NHPwXcVUoOIorsWP+4a4HVe9eXu37ZG1Chg2AedzgypfH2Vd7K2FfHtZ0Wmb/R
OCn16ju/oKDfxqHhWAhAy99QLJQsOiwqCQjx4x440g+CLRKg59AbS+yOKvLe0qeNwNucNfMxkdS4
lH3tYSVCfFqJTNdnGVO0ciksvXC49tw8hKGHDGXh5hHn8hCn7lHjqL4hnoTadCupP6mnWEDw+dYi
SNXoqXZdVCnhZhUd2jc6RETek5cEbLF2sRwy0tH57rULy3oN34+v8XcocqxMEbpuPPJv0MwAD8gM
RPmVXUttFof6hhSu6FSvP7kpDH6HyUbZT99Sh1c/ktGL3kED1qVDIkFRiGcAeWJCdL5xopOV8Rrt
z/WF4+rEZxpOtUR+TBa6y+SNFA/QT74OtNEmFXzvIEbtlZOVIV7EHg5OJqC3GcoFxEw21qQCUF0I
MPZNNArX1LMQs/4/LVGPd3/1yggWtKrX6UirhTDK8ciPWyUbQj2RxyY8vA/ZAzejTOn1fcSm+Gxv
ZNCgbyUhfr+ZmVx7zlZWV4QDOudcgA5Y4XK6Vr8gltm2WDVFf7hFY1zYjWur5juUOuZmOcz8GS9W
0ArxNR2yqZN6Diseid2/uymL9mVcfxoNKYqT7C3ozHNHNYhZ8MoHU+c35IkjIUCmbxxSxnEDz2gD
lbDC7KIDi+8RinBTLFtQ+9EBlS+nKYBPhWbZRHoSMyYp3nCn03WCgCy9tC+v0hid6XoYbF1hv/28
nV6wZU00BlgfESGF1hbEaWWG3QqEWedYm4lcP2XcC72QMhO24cmOuK3HXaZbebOOsUPXNv5W1BwV
KV0UNS0wR/2L05Gpbzxmpc5qmJn2TIBEs2D5haWy4OceJEpCVU5xYlbIvB1eRc7afLyZduIo9wvl
zCpAnujGjPsIoZCVoQVQicx1f7ZGYnGILKSs3mrkqvX/FPn4Ew7Xf2TFzK6TLGRLc1K0tbSMyqIV
l92z8ZvMSfORzCrZ2e9p46wpV+dGFZYprA7CesinLrvFJMG3IMcDQO/ahy3+GNpLmtWwwOwjqop4
yHx2s3QF8RW1T6xsxuHMTwgkq45Z6xxOdfzmhqqWsuwgTNZ1ijaU+GyKZppfCUHzpjzo0MUEHOA/
TdPjSf/b6ev4qvNc9NrDUI2zfORikssaS1gdi9JgGdyCXKR5lS1y9JJxZaD078kfTkx+Kcr6QYDM
uZ2p6ML9fFrK+xu2TVD35uE1I+PqiD3ox/dtusJnyUi/RxEuwsvLrqQ+om2hu6divojGun7M1NiN
jWuOQAnDBQFO/PW4WIRfozb9vQpRVu+5kEIKugpnIzPBryZSnena2kferrZEgFKhBtXtKwi+zdq5
RCw0nhZYGm/Diem87q3/wDg9bowEk2M+2U8BVR8eow9QFTDAWzu6FXErFLmeJgh/m/fka+SAdgsV
4G3GFrAdGa64ZXk+KfCZZnjpIUNMMh3Ax4UWit87RU3KKne12AlYmKRuzz3hSo/426WqRMy+KB1M
rBS8/W4b0jIVuIRzF2EcKwqCrpAegbooHxkJNG3T4Fx7OT/ObD7jMNZbLSMzk5V6ltmzO6LDkUyC
UKBB4AMtv9d1Avh9FODdcTdQB9+0nboJgl3qCzlNkFUgMI9X5lN2jxhBPjdL2oj9Dbf/rSJf/og0
IvsIQw7vMMQTbbAUJhC/Y9uPCQuxbKiC/qxeex+IZqA24FS8L85SDuo53Zl3l3w6cB21r2rWTLjY
uoohshaVsO1rkD++y5Fsh/e6yCE3Nyc1Orv5GCFWtLBwwH9QfL8BFulIa8Go2KmfIVl8Wwu0zob0
0lrqrDMnLtMrg1Ia6/MLPMRTRlU0w5yIo2QXr1lP32lxf8TSRJ/qpBoEnEui64IblKrA2fLrbuIG
paG6Sa0eM+95DHBEW7kgBQCzLBz9E233lFK5qYF3J+mNPdG8beBK3xaUGevvVRrVfWpSfqz3ssGK
p1xr4/QPvuXqJqLo021VwyMtCcaI/YN5IGKc4ZDGqVYXDcspFw8BjTW75sokr7rFWa9MilUQNNFg
FFuExepA5scIQusSrTbHAzX/YsPBCCugObSdM9U5PTuKK1COByRDxb8g/9wrptetZo2YW7uu6RS6
+1dExTj3tYm1Lv3u89yodG8JQucCtmMHPe7i9z6/Xg81FHaSm7g+FsKpIYZD3D2oKr2Zory/F4Xq
s1u2jL2hCYgUuEln5qCG90cEm/TZT2wa4HeaU0xmVG5oqcfzDKODTTDBN6Zh3GqJ7Ho4VQb+3pjy
evHwfFMdsNYRxYPQLUaLlkr+FsOCKaSz9J40eqlxMagiorggfGELq4bPpaqsGc7ecTXjndAT/Kxi
phL2Eb83nxkomzIi2fzNWJza/KPXzhi3lGxIptw1ZJfxqmbZfdN6k1JajOQjkOBeayaUxgSpCvbN
KYewZtsIQTdVQmvKPNcFRtRGAF4u8QJkcHoYr22zzg9sAinMmJfNWMZvEE8P0KEA/eEnViifgscy
cdMOSP/IToCqMdLa63hrnPLXgPYbHwVo2qGZU/LJNlFkhfVtiUjeL2H+dA2Mjf8uyy1yL2At5H46
vTunGE9/cWLFWMkS7hL1Wc371jHa0v4wGw1FYlcbbnTwNNRP8pnyodNLvR4FhhgbaGcK1l1iiUGJ
aovC8kAsNEdnOxLLEIvstqrsKx3GlxTm9oVCAOX+sPtmP9MqOcc5Fha2i4o3YTOumOiTxQiTDOsg
B9NMVjeVVuKLHHzN9+enALOwqIwzw8hBsQsdApR7zF1IXX0AYCLlLZTQBo/wbN0vjSth7raTK6k9
B0RKGL++X2PHXrgPF3dL5t+xGfv7UAdk+JdH8ZpTniE+4rXl4dfZ6Cnx8mfrPERbtwwNL8+bIH/G
wILR9BkDtDlhDzdlyj7qvUuxxzS7QBHEEam2Se+rZOjSFfK3AgxmjfbGIcYghQFRvMGBwYvPeW/z
sce6IAenL0GyBjpO1dKprCuHiQJjAzi5QNHlbx/7bAK+hAtf6OtQAnexBLupuf29I2sjcVUFmHn/
wB3nnjB9U+jycefFT9Np/GdUV2/UbwT3W3h/cCe1MV1a6flsPTGLtLlBj5xMjBH5Dlc4MoVNLHFK
F2KspDZyLp751Kz5GFl0gOwW/S/TybGMdr3eO7jpv234a/2dOeEcT7ayLh0ND8iE0gP6Uj6477au
TX1q+NVkBfhvW8uUp3B8khfMg+rsxa2nK7I0DticmVn1uImX44egGTxzKmJJj5eiJbpDnXVfLZZy
jsoM6/zsj69f4aB4Ih0vx2LoW4bvzoLupxJ79JaquqQrAnL9C8LY0EqlkbtwT/cSB+YJ2pbDpHHX
rv+81vaGPLs+GUvRooLiNuRJBR+C1O3m193zHc8V6B1+LzQFR1cbrIBJ89twZjSYvR3URz8dCL5e
gxVpEdDOr8ebITR9M5sZdu/egBe8mJg6rWs53vB65dkgpd3tmtsQRgbphIPDvfcvVdY+WgR+iNQg
kqUwrMsshHiwOydNDBEcoNlT7jIEWhmWK2SrBr1iLjFnRB8rxYhRn4Id6ffQgQ74dIW1xiYHQ+Yk
KKE8XV8qqdrDtqwivgRckQkY/cPPJGh6qnAUmCU15dN1e2R+Aba7UBGVrIRDC6JZhtTjQIfBXgZS
pDYrkS6mWrWtLi27IsF5WMhCvv01xLZCfh/lqzlAg6YFf9+TCDM/i8cClO0WoM5j+4lTeRd/dgi6
fNOVKZiTPh1vzUBLXZhgoAk3zTWegPSDgw5lmnib14g8YPsW9NJE0vXPKwq5jsaSnBKws0pmK3xp
uI09TUcQx6Fj2B5ePog/XpLY5ihIHUbS9j1QV/dmV0svEIBZ8gtHiSme1HymS0sUCMn393KQiIQR
vtjxttYKStRsngYCgRG2l1hA8bNRhS3tvo2VbTicEUuntWbxh+UfZ22KVbRuGCNRgAwtrRuCLQMd
DqwjlO9vmmeaw5JRelozHcCjJYr4RXG7MB7qnQVbSpWA6LUqBRs/OP96oyR8Tju3lDffhnOO3G/K
H2HYEbfyInQF9xQLgy7tjZPaASkv2Q9WYu59dzqB++2IWp+UIrxVyXJKYtCMqNiPQXLz16YJHMTw
xsc7ACqGZ6Lbm4PQP7OLt8SonVnRQudnYqxozgrtAhxdEoOES5yWXrbV3Aq6VLHgo1A5zXvs0K+8
BFhgEhrqcEg8+x8kpQ8rxGedbrg3Du1d5e5JQn9F3nlItkh1gmLqFUuEQeNEFW9Vha6GzURlNedS
2/Cu1iZxRKK1oBSzGQvzJNgaI9hwyVQWCGiLnxOGCaZoeZUUyCd+t342EhXutGJIBtZD2/RIlxje
3BPoSCTVAaLoRUkiOzseYZ5y6WcwCgzapqc1l4NvyQCit6AyybSwQLlZ3ccRnOGwP9aNxTHUccs3
u1NA0c/F24ZmaoxHxdMyEdEksJ7CfTuR4DOHEHylqnXZz8b4hGp5XGnWE1HnC1y4DcFSqEN4T+PB
lBj0KUlKpBA27JYIakTcTkkqp4zGzeebLNXwdrt94TZfug5v6SFK8c3naWhxP+jUYNstDuIJDiif
h/VL11ziQDxY4dS0xagYY9QXgU7I56HHZY2o4mx/QsgsUvHMLacMySmjuorLvngWWq8d1yRyErcF
uvxLMc5vs/MYXzIpLlnKA8rv12xmxrksAcHgmKFhqOretlDY2wTxhidS+xL2wJxshtWTvhvR+JbO
ihg2Rtwk0SHLCfogD8AYTK8p9nXdiDtLV0t3p2ADbW8QShytfz0eV7tHhhgzY8i6MPYvPWkZZO7B
J86hzpNRx6TKEP8Z6OLLKM3+YN7Qsprfd9L++Hzzhr3b2OMp2a+6OzHJoXcce7pCPSx75cSHqc40
UtWXalO+NNEo4aVUmM2zyFs+CkK1sn/P4IaS/xAwSazoyTE/RkvnDsxGpUQdqp866QUZSe/hN0r8
VpVRr/krnpk2WuqPTmxJwWH0u7EgHbWL2AXvgfJbuyeGIUtpJJSSCHqI4RWVXYn4kDgC7QvFVTG+
jAcQahjIh70d6jt+h4PfJeW48XV3fWFV0DY+OmMP79dtq6c4fgucLOlmfTakkPhJW8uQhxyA2VNV
Qi74oj4U//yX4dwHAMB8lTyaPSlDddvReVaqtM6A7emnSrlBKJfofTx8zPrqf7eAlmYyLY5Zm3Pf
D6Bjy+jXUdt05lBbqbsnjizVt81+7j3yskO5s4fXFiDll/90m5BF8lrkUih9NEkZwBUiY4Gm7xB4
UMnfXe+eYWhSEZtJjQ6/25xCfzUoUSTwbFj6nOOg6mFSPnTw9M3642tbdtijrmxSmnAO0hMtcJ1l
Bw+3VcUzyJWdb9eUxvaCoxPyDN6Tk/d9yrnGeohyuP3Ms/HnlLjalGMwcUvh3PyvppXcZA01oSrO
TQPPKkFgHL7vzOQM5YwYn+4J9fBPb1kYo/0FjY9D8WX8NpX5XTW1374rmM04+uIHo+ufTlpfe6/8
2EzMRdWOXBSJlUKH2UuW8fADjjpHhNDTjSFkbPXj5NQTicIn74NlQ0qKanUi4DIUut374Zb891sX
+HeuZ4mk68BpOSN5DEf+7E/2eeyekTtER+NRsbEenkiyeKAxRYEUQvrPTB5LKrFYOQBVJNboTq/2
niWJ0X0ORFrEFQdyzUBE2D17IJJxWga1FbfGP/DFwcEl5ES33ei1WdP2gzo1rli8hL+fGHU2Rtub
HfSJIpofNp7/4ckVxvox/iH7lViGSFWBX8HDrIVfgv11DBZTuNK2F5D2vGiIUsEBFW9u6/W6g6T6
oo91yHmVzL0FGsif4hPtwPWGBQBJS4u/UNJNjJ+SXq3z9xodmB5/G38ZGs49yG50GYi8+2bGlN1K
KWN4KvDtKWc+jy8XkmFt8HYfarlKKlJwNK8HtU2eifw5+WleMK7H1Y/nXY0pJfU+R0fVqt8pHnsz
YBDIk1G7EsL86ba/QEwewmHMKCQiSEO97dVns7VgnOWT0uTVm6sEoASVZ9kNVPpO0m/olmx6q3ss
lWhZqbPqiju0mj6q1kXPGecMnAb0CrSDTehZshMw4kLTZL4+Pb3HXOlhSFuMcMQ+BZPD4/5nrCwT
p4jzdSVRcapRRNKeBqCbmrXn4Q1Inp7JewF/Me/tU8tP1X1ppUVxFSndypUsMT7THr59iAGSI/VZ
7axBs/CQKp40adV3YdLiyVzXB75TukqvY0dEL/2mBV/62Zy1iLD+Iycm6dHPiaX1ZH5XsQuYKIeP
DaFQ58d5/OidXFdDWItNTk/+SltDKPRiG0O76M4Ioeriwjk42zANXI/bKR9FJrenhEMsvZPvtRqH
vQLBIdcXT1mfY36IfZet/jqVrPurPblzV+R2wgg0ah36BiZR/exNgHRl/lqWEfh5FkITXmxo56Ik
tSO18q8hZRJ5o9LUKfdL/8ukyzAc2IOgh+RNcu9siyH9GUokmeNdFmoJQARnF64nnqjMbWjHPUGh
ntPqc1JxK22BEEx4V1Pt+g99/1lWGXYMX3t0rNA7j5Je/C+5QGUbv8fQ/jUU3EYJiHlVGOO60E3w
eNJPgDxwVmOn+ErjPoPVH/x8drycfYtDgKQ8lwwmbYy1pMXf/scUxwjNP2Gfp/skjNP6z3LinNZt
OgJ+jJW4fKMMKkfToyY1WWPWDhjNaMAnffdVmshvldTDyRNLXHY466j16Q4o4XY8pCNjjMx6zUHY
a7OjZZl5tmvfF1vZZnq9ggjAoGXbBYB6cmffv4xVxp7BfiHkwWUjmP1BG1/5IMXz8tgCWNoGg2XZ
SEO1g3Q52c3U6w/agn5dqboLPPXjffsyqOi6u4/80AkxWp/pvAYZeBvoldUk+TlqoKlA5aRhWUo7
zOhO3wrtNCw9ytIQD0O3jOUdUT1VnBr4i1D2Bw3mXP2lVPMMxCGMqXuwVFGG3BbBbA2j3ygYpc3Q
Yoq4gFKxgJ/s2CoIaHYABsTEVwQILqFfW5Z/DSYv6rMyITRg9n4O2e/2Mlnu4G97U0x2+cTjCbel
dhWDCw3d/dpVTk6V9sSzsJeHZfAg+Km3BEL/abazjlmsi0kKOws9d3ApFw4Zr56nmeoccaqgkcUa
9Y82gBBp9uE0yiZ9i2VLr0yuCnhT24sgWE1qLUzKfl5NQ4DtuSDfxaU26Q4qUITOFsTBI484bEv/
OKEuFnauEE1/J8jmOKxJCmg+hDwP5nABh10cKihWy8RiljmyQygjLtYf0MobA5pkNRk6cawS8+Ly
BDIyNHn3MXgeiiLJLT7lsaTCjsMyKR9Z60BRjgSMl10kApHFkHpNw65pwS0ZsEFEkNI/yryXBr2g
Vr4zgx+g1MhXz5Lq0S4MzHW63FbCrH6iKPP9qJjx7/tIEWfifBfG1vSe+YQJ9RnHYuEEBDmyS9OY
YHLjG1yK7TccSIbNKhBtNpYoCaWb0WA5wb+XR9piDJVA+f6KoQhl3kGyvmfYlYLRDtaXJaLv7U21
eP5ka6ET2F3yjdI1D9DW8+vTDe9KlbBlkbBxxRSPm7Th0QwDDDigjhqi6qeXvh7PWn3o8TmbxQIC
E/ckCSVu2t1br0ZppC8kLzvksZYRo3n6aI5aq6M9YbityHK1zMGulsHsL7Uf4DUpKY49cjeGxXC5
I+lqS1ChHKp+4xE3Yyi8A5pVjfivwC860WaHF1/IkkdwEmgisFDCSOStWR+uqy4hfH70+9P1UBCC
/Eb1axQjbnLQa6KTL6iNWws6JBYYqkPrSsfCbxYOpusudS1bP3V774scTG6ixza7QIUSk6pvkb8x
hmuU6qYOEKFSMaOy+7yY7+VuvmbPRv162r496vgWIVlI+WdijuBVZ8zYvxApizjt/nkJVfyPtTNX
IClxegMrwM/4ZnDsoWQ4auHijR1TSjIsVdiMhuAk1nbS++Ny3Cjz/5qklF1TLv9z8O2dEVVBT9iG
h82hsxUFNA9hPAYeP5hcN1GeSW4QJzBk46lfhuB+JKtwRYTaCLKfrCAj/tAzy4IR/x51fE3TkLxD
vkEjlWtzK+uzhG4EyxuWLhXUXVMYV486OCRwbjCnbZ3/R4i8Juj5p41WzIwl3j9q74ned/oVzNRM
O0StMflLsFVau3E0LADciGX2jXor55vpZMvQI2bVPZUaZ4kIIP8T7S9OxNF2F4LIeuVGtVlflc8P
3LPAtjJvpShKNXm+2fXH8WYPlrYZu0F9xb4XsWQgw609TVEhPQXRS/7BjoETOaZFDKou24+sH1Wc
iz+6RSDrkenWrdRU/I/DrSxr7XO0IN7hRSl/snQLQ2KaaVwfBeFNv9VFK+q4IOCYm5/K1aQvkb0E
N1L4iU0fjuhwa5TvwgaaNOdrAXb2NcekD9ci+gMtMjB3dHNYIOrrBcgALkKXbi7T6xrpuMikz7+K
wrkyNKlp6W5DIwsdHnnxEuLT2LcLcbYb0Ap/HiBslcPgbZXHvRPd82kIkOOH8JEAAtS+3oFLTgkb
JLYsXKCeLRj/Pum5mqG1g5L4X1OUMxe9VzYfC0L26hfHRvF8VcbROiLYc60YlJTv892GwETjHjOJ
TbuIaRnBLLED4jABJ/x5x+MQf4u8UHChFt+ErFWCPcrpvrUHOfkQwuu1160hx9gMZYx3Tit7+89M
HFEqNjHEcrTOl5pYRmws7K4ryn9NDpT+EPBmjcXdc7yCC728rXDYZNg6pibm3VGyydJYVwDnyQOn
I/fVYmU2DUiCsTugL0ItVzBBvjk17uSPagXVActD4wl19mOl9gws+j5FR2ZYs+insINSgRqf8b68
mns+tB5ayBOowYDFYbJWymyqJccrJDNjXruhgWlculD5FGSjCFkCdBvoS1hO/2ykCVkjcrv4hIyz
25FlZ2zYGHSyXYAmEuLUmPpPPat4JKiPGdLrZIshIkR4Dtye8uvzQOYI8xFOtlkCq3hfkzSu+xjt
G1GFHtqgEuCbJaIhonbCSe/9EcY3iDwsWXgmKDs9/6BNf/VKkedS+q/nDZBNsQkhmyQQs5/f+FWP
xYpkQyMR6Kkllob40hJ5SFi3DfBt5lzYdi70+A9gXu9e1VUaV5Ljmtnk3u3PZev5J8RJICK5tGRp
EZk1jsuNFtLkxHi9Ci959In+MQO3RzseEonJsdSIB7fvOCSrue/P3BMO/gPpeV+DHpAzyIULEcaT
HpVg0qkbrnSBHELLVs2DD9fh5M9Qt/X6VvMrng8dfbr5NzhHbj4K91v569190zgMHd+QgioZ1rf7
Mmh7IU2DiYfRNjgLwQxii9Wdl3a1LO3NCmILO6TfAyoNu65ji8N/AQHGxFg33WGMB0CQ1amD6uMu
JNq2melyI9t+t25+ypwFmx8mKqkMsmonZeV2xXRn7Cf1Y0TkYzlD7D741z7mjcS8HyGkUsAJfKMH
zHpnrsve9YxqpH1QYqvQUIc88CjMed4cEMZ5Lako3GotMlbG52F6daMlg0D9ksctEv2ACs/Tn2il
rupBUfdXTF9qJzhn8KriGXGTdFx4+eze+RpYNuyD+bIrYGIgfv6JAcWSfZjWiIJAmAULejkBxvyy
AhCyTr697YwQP7PrDVypljzYLGe15VHGbEUg1GSsOBB3CnZwgKeyG3/SKtr/JWYL22zdNK5vLu/i
p2qqMgPzoJ4NhmrIGHxpNOubzVrcTIIYyG1mziTRNAbAC3bK0p0Q2nXWqaqISmWPJK9bsHVudNQa
Ez7roDeHgYIPeSQprsMzMvkBc1Siu9hMxNbmXHkSkygLvfp/l7OqgoRtmHxdMZ0llWaKR1SGEqMV
nh0N8LE8x2KGxax6C6AP0St8POv1hvEDav7ADkR7/TNSgBdL76xJ7CZE4kjEum/cENyOLzafX9ZC
Sxk7mwZ8FH0Gvy/0ORK+5MpPA3k9kaIb3XGpHakMqeFvySWHFwn1mwTHEhaaT5FZbRBbrMhDkZn5
G3EfYakVg+SWGVRrRAxpJzCfxs7ID1vEparuwFtlja/NdYfTyQXMSmxo0gmlTYFEgSmn3Phf5YRm
l31fBip9P/oyc5Ld3EMZm4knwqDDH4NFue7fixa0umaWO+QKZ2e3FzoYGgGoQDx3SayU9ilC4nNI
HlQXHzdLlfWYpz27aMTUak7Axo6It48ScmP+eZMmrK7SQlSKL3aqXaDWM8o40adxsMW8Bx40wfeV
7Lk20DB3p5bZg8W1ecL4hFEQxgfgEp5MxOKDuuVPH/vp2hhTAYgkwCpPjVIJC4KG0uLg3w9MNn7U
TeK2BSmc11gnG6AOZ4wywzlM6+mLbWtsTocOApuFIL47hZ6mGbgZi8eGLeMm/G97RfiFsUs12doA
CPX4WCZhSvs8G9Qc9ZMaGaXOOPATVLseKcEMzd+NF0uLhpWJZxJXmP1TugHydPRYxJYf9gMU7fjh
0FNJzEuG6/8rLPDBeDuqhF6rwieQi+mvtoWliZCVZ++c40ABrfeJ5bzczfmHPlhRlz2GoOH64RlD
zyqaoYUMmNlYxifuFtxjONyv4cpxCaQ+ChE6FdR5qCFXnD4qoVi2/o37xrtk3t1zfKBO+WT9bACp
9REns+sWrZN3svk91m+nFvjJNhRFDC5EN3KMl0Wv1KwV1SwD4ENk6aVYuxehgDMe+Klvy3+PUruy
61CVJtjQFMiC6sVSA6SUnOvjQ2F19YPIT8bCDNyg0dCQfTXhbpb3XQ9CtFyK2zWr7XsAq2W5vsek
7M1fQ9GAPTYz01/wDxwFw07Q9jhLzKX8plpDaMuRf6+LC/97lYE4Ni2b0lavgAziKdY94IcsjAjp
Lzj9oXYAPVnz1p3m5+RZ6UZDId75XZfPYxBkmAAROuTyA0Biy+Z+hQRiNEs8oyStiD2Ml5+tQ9bC
QffqYPKcAVqvHc8HfM4/+FOfi55QCJb3XvgS13SK1MbuLSwhS+UwrzAQAs+lsLOJGJIsGBPeVvXB
ao6/2jSYBk2PnQHfTwM4VOdGEtDoLuyoxE/rWMjUhN61uuHVp/pVe7lglnGJqlOFYMDhL9KQP9pq
dAIvbR34g5xb2lEcvS1Aj1Ypo3kUJDbgavFard9kKyZKrptnaZutRBilpe7Z7OrR/vxJ1FdgR/dH
8PfcFplz7cbYwm2SUrMtPybi0LFNEkrUItH4vGlwVC+gnY8cKBUgJBEEByzUysW1iEvjq148PUoL
sMYJ3EbyoCxEM4jnyKQpfT6hwTlEKx+7XKC326Wcew1KGX2nZOHQ+pFNaZVdSs8GCqcWnxQdeW24
H5FfS9GfAvKA3cQHCbgw1s9GEMQKCDz9U2wKM9U32/agQVZ+iDv4vZi4mwU5vhw/DmOE6Vr51Rce
YFhCSu1bg8XuxeDR5rfUau1EN+iL96/kLa04JhFiuCU5MXVRMskzehQPgczql9glI3Sqrx1rSWPe
GdnSFPQNVTROQwwEmijyA7UIQyAMXWpohcZlY0L9vRHjGxtmzKsKUpiTHF07kLXWXWUzX2ju3kEs
NEf48j9/2agpBqB/l/rjsO5JTavsi/27LxjUDUIM9Syi66fwQBoWl1dA+s5nf26CDImHQvqV2Acj
1/zyLghQJNqav9xih14t8JdeVuxj1nWqjJoIUuFKDSrONkDh7BnCjlDyMBu1Tve5RH1w8nrqhnF9
mHtJUfzEh/ABCGgeUErLZgO9hx4dyyYj0YfRITwjqyEQIFlP0sZ9JM/cIgoNFVykUIGsXSZzr+S6
+uO6o6DH8tcAtw44jejNP5Tr3FQO8oNN5ZSHLo6CqX0wAdF5XwgE3U8Iyo7/7Tx5qTjKZF4Ur53w
blyn+Qh1flM9xDTrHg0Z6Ltg7wIIqZEw84/0m7VOmRWpYHLMjfHR7A7W96S0NZ/E8J216rVxaOAi
LSqcCPgdvcKKHkUsEEJbm2hEWBZwGsHvHr0ZcG1mgRZkiktmm0FCDxM7NPOo7kX7mz/3AwG3SUZU
VmGKSM7riMSSJ67SHYLGnjLxuika99DZRT/YhXwoqr+qxlGStTh4xPY4x926dBXagZ+b6dDW7n7J
iYusNMa2ImjERu26VyUTLtmlc6BJYrweckon34equCmIBEFs9bPSj9YSxfKoXBvgPT7L4YPDo1y+
GELNqs5eN0r0T61NsC7IwZHjhVRGuBDGIL3ZbpE3bZMOzcmEAtT0udrnBlbMp2EbAyDUMU8z4T5n
m5KZ4RCQNwmZauF45V/qb9gpmfUOFy7+D0W1xEbmT44K4bbzzgmp82WA7XDQfDJh3pv6Y7wU6ctP
q+KM60no1bi17E7tb7uzWkEozVgHF8HTGCjAn6HEGWA+O7IFq1BZOnAvRET4BNXrvdA0jAOcNfTB
cYFEcL0FatgNze9oLtxBZFHm5nfVIyCj9+98MtAHiW2Pll4UCoBoy1lk8s24bCxlxy9pYX+sMbKQ
lz+baueiGNIW6Zo3EsPu0rlRLmP/MjBm2x/a2Lt9rnmyk4Uqnz6e3bkOO4cHQBaxui6xWRJRfC9L
UsJtxEhUG7E+48ij5vNJJRedNW7mNVhxTokBvxcjQ0DY8s8wvjtkKHgBAZUL1SbVGB+2B5oF+0p9
dhofY4IiEiM6WxmWcJK5HzzbFoBpX4s5t29+foACsEzOm661wakwZ0SIogoQ7/9LfczMGt1eiD2P
rCVgYPvt1OMmK6R+J82EhCtt5FrFsCGfwBztWHHnfdi+h+PZMvdIaUaMhzQs27BKSrh5N86u3rT7
gB/TA4yKoj2qHvL6TVmL4r31qa8sh5/1WBmBbGxcsrF4sdKMRT1j+vf54YmTzK9vjAlFulzZXgiA
e9MF9rq1i88umjAXOE6zJVVzKimMIlY89jHqz6OjP5P/3Rvtyh4xiBmUBqrIEpKQutNSAgE/4i22
rX1qMEPuDd8AXUsU/JgiIlu+/PuafPNNjItw9mHWogc4b8m+0Zo56yoZQSRbVrMMrcJKjtg5k3sj
SPBet4eh+8+Ut8awEO3Vs7mGN7cmJNJMPawLFHyNwhpPff8Ltx5eb7MWDfnopCxTJfdmez08fTdB
1iPZQ339uAvKOI1xE3FiRvEx1eUn+rZOtSQCUi0QNc6BR7RkteWIczPfg9gq4RwHCwjiRgHRmPGw
6Ur2ZI5xLkkewNFZ+LoGH/KhijXxo/CrrEUeVh29wkjaXGwu7UIhotp0YVxhKB03Y4/H1dR+n2QB
OfnDLpFv8JjiHi7BNgvZv2bxs3hft1bbeBQ6i8jH20Sueipwhi56vY6vyUA7Y9WzcimpgEcxsMEq
RnNWRCI2Jrc5GSP9q/7y5IoAdN0KIinD0qHsWhBYAj+XrzWTsKqbeemF611CkmR/Y0rZr9cVCp2B
r4VisS7RQibyn4nrWFACET5XRttvHZwxYccgW9MGmROOQCmceneHjXXjk8Gl9XM9G0vl5iUu7lnU
4ey59OPMkugN3O7RZ4kuB+M+CqJ/LghmiRXJgJLuOKYTKeiFQVUPLfzpQFxcKjUHopbMp6M3LDw9
v9AdP8E/m9NGovOv1BYRlX+fKYpKzEBOGI3ZMB3ESbbhLtFAGfe3I6oMJvY7Ho5Wx4CcoUYMOlOx
0XnZcjVn3/ASIUNAX70+yFf+AWh2k6LPSVptnAfBNZc+IFVdBC8ORzq5cAOj5caefglfnztF2wxh
ioKsUvtV1SAOGR/IbryPkz0yYXZR/T2S1vcq+MWI7hmyt0lgakDnFMoYIDonuYkoPU74Pa1GgrgV
P370c42nk6HZddTTvVA5QGMOe2tZYKaGEbzboB3regS3zQNjDz1gSjljrV4n/Hwe0E+tuK3cFbSf
IOqdmztGNkgXYMj82Z5WZ9TxaJBxuT08dEGLZxSNIxaECnKvodnNxgePbtR/VPieqSj6okH6x8QY
dEGgKXRK0mMBa12n8tIOkX4XQJlK9DcROLJZ0KuiNooYgkk8qTAIKilEXSLfm74pp2e0Ds3KSAXP
baxUYV57sSm6+itbml/asYFg3zHTsYaOG/J1Y5qFwZMyQkCJ9O8p0Cm9oUfo8gZD81SUpwJEilsf
R0OB29ra9nH6bcQJXBGHY8hFW3q6OQlpcvaKTyA6AimP10qxXe6Vn97a+tdUtwlpZyjqcb++V4pE
UG3KV9dVbHhhL6Y1sAAqpcD116hgPf50QDGy44YEJYtLEceSQE/htqA1mWXP+SExcFAG9Hswi3hw
XpR7H3a4yAHBLzQ0HZvxGBEagEHLQ4gfx2XTReLoq57USn4PlarcsbOzuq06cXLIEkPbfFpTamBR
M+u6h4813BHU/Kk9JO1+3K9Off3n4U92+kuUnve7ZgW31sapmikVFAERV73uv1D9Eu2eSJWDr6Ij
PALqDih6h0k1/bePqc7RpK40eZji/VpoHb2OfZajElLaJcJzbRj4+SuIKEVyiOApdh0XLCeD7Fmt
wAhbUHILy5wPKIx/sfl+HtBXuRrkCzFp3mhKLGoYTsmAF8hdh1/EsTEUm3cnL2DRoXGVJyqumago
2zMpZSrv2baYDnIQ7/gXWHNmiy5/vZMpRDnNsftE19epnfMn1zXUi4+hy5Y+5Fxcp/UywlTm2pNz
yzJJOIkCsiuW1Xx4vNDntcfJ/rUKnYmuFtDkVeIyMkjk2XD4WEcV2ZdFvtByhWO5YHbRc/O35P8v
DilK4HaBo5D7Kt1F4rjKzh6ZTUeWh2X4OZ8gUXKsyCChi9bcxCnNcJghaD9VVBkNYDyrx4xSjMxh
OlweK73Q/F/UGy9leZ3j86QLJhPueJt2w8FO3BrsHtq41ntbawuTlkf+pH30LJLm4NVwuM5ReXsG
6Byr7JQEz6w35YDvZCZQDs+Q4Py/qBghZamFtW2Ie47XRDPWHGZHnqSrOdXvPGtJQNf5ftCZzYQo
Jlx3IVjNtAIjp0Vua82sIAGoZEVEFUZBr2EM96rYIQqO6YNRoonAOT7q3eeSPdElcFx8o8hAEtgi
FDz5MNmAj4w1Z1J8hkk4HhWveOOKmbxSpNNo8A3Jaeg4xhVlAL3gemSAhBiBhw7u/3jCn56D8QD3
RNBMCpgML0c3GbY+wZO7CY8aUmOJKxaWDiQ4qOUZKM3+ssdRpvN+bcDEbvQ7mebQZbVSV4TGkNOd
K4AVFdVyPTXYBwuEbLkDDl3p9S54mM4/aG1wBXw5DHKzdElhtfqbxuWwzjlxmRvzt5M13uPMI/04
ahB3eJSkXK9iQWI84asXwpxn/Tbz1fxgh1UKeJItut1piIYvUgBqK/OK8BOqWBuzmub6luhr2laG
IOCtHPTryeRWVKpOa84cVJ+788PaKcF5eYyvUFzaIGox8UUTWxUNkqzO49qgobGjibEkMLs8thVZ
mSlcD4TbgN+lZfJ7E377yIX1zcNtd6JNjUxQZ+m5yaD4+XwVUX3w/GFmWTdVoigm8Q63YcPt0v9H
Pzklui9C0JbWi1pUMQyZ5nY6x2SIyYiXM+c8chnVopT2I7tnkfWVYwsWrNr6bnhY8kzzv9f0P3Iv
GJGl7fLIP7yNmmoq9fgTEIe04aSGp3DaO3PW0JpIWLVjzleU2ElwKaziiilSCtIXgSQYlEjWizte
8TbTnQHYWRGJ1EA+znl5dJWr0KBvV46+Piu8GGLHlfaP3zpAJCCOHy2Zermz489Uh3VOYpGK15aJ
HUs/7ldY1rJVgo37Gd8Y+3qWDq9usK289xhOGVYE/OXdfxRU+ntyQllTMUhNhPA+CrIDqTfbrH1m
KIh0yT4m518fI7LrxaeH0Y5+iDP6HCqfF/rWymSTdY4okD+jBDJnrvS8dymOHWCfkHUxVdXhYnJT
3bFB420EwYaJ+lWMebkuAdqaoHcWw92q0oY0UbkRyiXvVjG11M2qX1C0hcTQb2aTdlHfl38svEHo
unw77PLz1ysU4U6bOe9f+uBLLEoD2+RfXkMTKIcUXBCBpmaBrUh5o7bYL5RKfOmOYbbA8TXUnIFC
ognH1UqoiO34wEbdjBgS1T87QzyA0EnhEH6ut+U6R9mX71dthA5nqJPbxdsYa49TjoKrkALUVCDy
K9wdtt0hHNv0vX/nvwK0hVj2TeSf6Knv1h9SkO3ErwZwLBxVjcPzMLo8mLb/viuhbypJscHIWhpn
0jwbC68nJlvLBVSfNm1fsaqcMDHq6OAy/Z4alBlEcnl5yDUIF/g6zmLG3GdyQ4jfJeqOieXd+QMF
j0X7fKYoNuhA6fWIh7J6w/+cg9XIN2HBd2EJNS8icJ21fAN2l8v4s36bN17OOyZN+Sqh5eZCcXXf
PivVuJ+JWr9VYUaxu2isjkcWylNrCymCvUVVZ1FthbHxCCt94wcD/5gF5yfkwgXKAEanSjYLpPQK
xapYFCcu0nLdZYwiOgKZsO9bL7aNPQ20YR8A3Kaa19o9bw32LW/MBP4/FII2w1Pnw5KfIN14qOxl
u57jj9BBasqPOo+IcRakYDJ2SrUFriGXWviJHlvvxVQ4khqQqJrSQ+uRMDakpiykuKgY2qjNtqV+
RqG0JZ8r8vZoywm7r5DiDLHHwxYSpyhe15CuCYYhN3Cyo4MrWwhDz1NVGupEcT40koowX7nwK9Wf
ATmTWC85DnZ4IjP+Y2pe7KU3z7vomQHEJlRnZ6fVl8TIlxeRMY1dDUbv1CtWozq7eYvChM4KJ7eM
MX2UKPYRLOZDWURGHTLZ01qTeb3GmhzmINvAdcVnqrzSgRIrUC2NpboS+W1GEy/6L1OJ+iNLSVTn
FS5nVVYM8BEUqdGleQ9FNucntB+PaG266zSWSpafNhH+uhKULcaQKaBiHNL9a0Zs/lQawrXcF0MG
l7F3hxIHOWNeD9+YBdNYD/y7K7pepksj515Poc1gghl7erU4Pt5SBLZthCJuo6vYZXWFym+qOHzK
+xK6nNpODH7cc8HH8AJs+Mbjq0sd6SNQlls/QOJlQ86KHg2nTcFIDOohG2S9RYrC/a7paY1l1VE8
IXboC1GaMttWiW8VWnymatJkWN6MoK/NzF+FdHK3dO2TOhLlfCafIMa/n/8aYu+yL9hVhlebERl0
hW76rTT7j+QtIQu1DmxHsURP8TQ7wt4zGW2/Qw/P7zRdxQim7zIpKHOHTb5J/tHtWN/TPVpinUpk
Ii/G895i1pBLnb/4Y7alK4pt0k0735ZdtjFSksBfjO812kRW7uaihLSQohM7kR/66z3ybprPVmMu
JRzqlicNTSOmaehfojysViwnz4gcjCsYEp1eOJpDW5GKqRRYBo3II6Z1X7kpJobFtFN7m4UTNrdN
PvX1mrzbpRv7GCUh8nffRcirllOXRE4ODJI2vkn0lS+lRAK0OBNOALyeZIWIl7Et8ptfx2LY8P8s
FMeDouFF9u8wniGTM2nQRODkljBS4EfMO4HzJfVXKlRoOp3WdfQNfH4r806E5XsyyPWHDIqHc6wv
sgYs1lX41Pt+XrLG85/k+OEoSblWDRGu9TSqt8TUacNvTgYFI2oZCof6/F6X5UEmC5JDJpupkFKt
j7xaAdC3w5VBloygljH97MRdIAQ9Y8aA/Njz0J5Zx5c0PaJkOMYjDJKr4RDFR7I0yvQ7f4NicEQN
mk6v7HijjVY1XKK+Mg+G54NXpRqWMnWMhLmsZZRRznknj7QnboMnUltac4ENfmYDkJr9dXU4w7jI
16ea+kIs5VbXB2kgabaP7IoxYMAXQ6kmfkoLsv3srypFP7I1At3nfVBfUUHLW5TL6+eYG9g0alX4
+GcTv68yY9c7M0uZalqV9HvmnzoFI9yIpzNt8KOT6iouQAzcfa0PWzUTMp9aCrn/7Nsx0owfUIDu
kfAhSxbL0Q/erTDStHeHn6hbrRQU0M33XMdBfagInUOkpaEbq/556gzaONDpEfnQPwuqYFill0P0
hcqB91m11gJbjZ0HT4xT0WsQ5InVMr7a1EXVCWJGYRs3KnvL0reFF70YP1Jt4SofPoa91/6ciG58
hipueL+KrQsByducD0cOoy8vLUnKH2fQ9M+QJd9ZFvKsgz6EvxoV59UjJ2tXTp8N6BX2kQ/c2cvX
Bt/uaE1+4gVimG4NJvMgSSpsv8wcwQxwFlXMff+E72yo/v4zaikQhbieG8ezRtzy66JOimak7FXA
/nq1l4PJjAOku1WZfsR5ticu87iMaLfGJqUu6pXlc+PoUi+CWZ9zzYJ2h8rLK74ZS8l/2TFInC9s
UF5KE9oovcyYXqxkA8/f17ht4c0aA8QhXNmRNdDCrJMseo8eMR9oARUWtm1cOwgJBk7zG8/lZQWJ
fjYxfvAx+ji77i9gyLqxAbHAk64u/Wb+aczoKvuYkXisk1g9ZvpW8HNnfMbyydKiPsP9fl1HZ3nK
gTitB3Wp6aVHrVSK+7N4TQ1J2oz8NqwKBRsY3YDEeytktssKtfL/n2aCPgLuBgMpqcP/p302mR4X
QvgF3ND6OF8pLYIW/DTu8exZv0DWEVj6uwMa2eocg30mDdX1oGdnMGoi9rZAckdg+amPihQ0PGN1
apzYXyf65WCBn7H4RBeCaEGnm7sSYuO8C/HZvfSrIXsK3ouuSSqHaopLgwKEHmjqEU6/4mPSs6kr
tqfxdJkWGfi/aTx0mirbhpRUyOXZgenoc1/L3sPAGee/IMyhqI/jPBhAeuHcvnFYPCmA42NHLHFQ
qwP6H2lldTpYl7/+SMm0ulKeaDQ4q/8BBXErwQHvzhaRsVmWPE5QuDHshPmlz3spfk2s/clTv6if
Uk1vzDEImGl0EMdFR7YlCwW7e05beVLW+Wl01SlGNiL4AJMCqOcXQPEjr93T65GXQmrdbR40uQJG
3Rp/m2qF3TV6M+ZONGEbrDzw+cGYiRKHebc/OpB7kcs7XL7iJqieZnV2N0ULW+YRTsY6JWg1V8bj
1H4hXNBZmmpLqUZnlTFx7I8mLItXIJUKdGqmhiGgr4mjTnm6J9Y3iv8l862ePxo8i5Nfp/h8c+/i
7d6h72ObpguXlU4CVhGDHV2k5hSLgPreg8zFuTL4ffUq3rjF0L5HDuOOk83/4JwgjvGOfO02sF/Q
d44RxuaB7d/B/EBr5A5XD3dntpi0t+xS5H59hX0PANmFgCN1BJctF+EO7mF/ijtsR9TlyOjE9VOW
39kQa2dTsGSGUXHHF2mySxQ9x2VUdQYmBVTGuSXlnowkUFuawo+nyiCx9OBJc1EQgRC305Lsu7cg
KLFk7ETIyadeTwmVXR4BvQvHKva7ilZCvURlDWXTz1/MtKsgdAweQyEXalvfihRJyOh79myY3SdL
f4CerAXj/SVOBMcER9WF9JiCc5a1CIsn/svH0fvFpz3HvU40KpUhPNBfnl+bJMHnT7SjyWdvhLz0
uYLCTZx+0Rf+2cxO1uVtwyOwEQOPvz+et5VIoLRiSAzMsqDEWR0Pn8coq2aRneN96DJobJSuCWc3
QP7guecHlS/UC0ih91XJOEfBXNM5XNeAG5sjKhvqn5lU7i/6Is6JdfyE14NWMxgz1cavAZEdzKXW
amnutSJChL6CBya+s4s0vf47hv4YAYu6JmbPlVrvnd44Qlzf4r0cpjpUZjZ9zJp3QtQemO2iRGbY
t8O4Sm3MPClarNvkG4E3HAUFGs1fdPAMGlyxgP5NeUsWJe9i+dEsnej0BbtkiEtoWtsru2DHbedF
UN1yD4oEnWeVC0nN73fuzox61QrQyQQeCFihsKZuLI/XbLucu1gGXUiy+3KJv8uskfLc7L5CR5r+
GkCOm9obgMFnWKf9s4BNXYPf9fY8K9Om2tTUdp8seA3Nnsk9SVW8Zv4as+AC3MZZ989pn1bAJvSR
PFY7bdVac71/zFb0c0Bk6cfroVgJVveh00k18sRLtS+fkUCAaEDtBcSJgvCaYU0bCqG8Vg73yq7R
jCAhZBQQJr7/tkxeI/fo4rzsnbEniC/c/BlHm1wxht8qdYijywl67Pya4wgiHsJFkendHBIODY3K
pzcTPo2tZZnSPN+4clXlOrSNkpku6hLp72yqx1bA9SJJMN1nkLK25OwZgwfQU+V5qpI9GLo6N0We
BvhLUbEAVVuJWrxbcFh2GGU/VnQXcHcRwZ/TWCq/80+cpr9dnR64sjcD3txTOKSEr25Zdi01tL3q
UgtTLhkw/XIMONlN+uazBeePplEkXMS/geIcm/yl7vFk4/psk5AQdO7WVHjprE6EE2MHnszdy9k4
DxtXGH2vmKDgM1oQkkSIA3lvx45tsYSl8FQPs6RY6xhb0zsM/6nIfTu2UdIokoq+Ejh2+2z0m69o
4yVEkP/+x9KO3oLUnq66/b1F3OqScVl3a8eD9P2X0CYzWDMvkae++xt0PJsDCtqxfiLXOlmXaszc
iPN3zdb/Aatb7tgFO6upPASwwI7jjdFKQqs9lGFEnklTmgS2Y4T7n7jrrEVMreNYKWy7Kxi7DHx8
cDiRLFh4yhFpn/Lf26jo/fD0gDBu8+TcE0Wpciy/ETPxaH3PL/bN4pUg40FYEUST4HqAkdEuBkH1
NydenkXSinMQadOhB/mvjjHtflG2cP64/Ef1h1TmZTfoWerY24IjFnu6QQALtvA3gdEUyvf3mcNJ
n40yVWLS94o+chRt3jHLAsOIRTlWdi2ioFSnu5V65MNM9GzAa6GUk22wr/2+U9chyH9Bumhf7cMA
vm4KP2VGOKNeJoRFCbaJqhv4EZq9igFPFiamlgkzGOlAGnPyk8MeNxWczE1SNENQwXGhIh/M70ns
D0KbitQq2h1fbacmPSPbkvj1Z4gwFVytfE72/gasj1cRx7X/TT1MHrwO5CDUunPGH/aoOikQ9IFr
CfSvgeVbfiGKK4nNgFff56MU5nWkeCc93uwILaiWqt0u/Gkjt2AvuWwY4j+f6uIijObhdOSAug2l
KXoKbi5hKTnarNcq3/o5SPS4Hes76ZMm+b1eyocMcba9oHX1xAJOKLVlpVMphmYCCY/dx4pi4cTv
ZnAsfoasDucXsfPNGM1Sl5W8mdHD1tgHYrWDtLDVO46OPwyE6mcDtSVYT74ResRwzmCZ1x3iY+MA
iXDexTeBjSVY/UGOFmjft88wHjsDq8uENSFIGHkY06Yh2Q3QR7JYavRjydA0wyDPUHtmL5aMj7wa
O6KCYOIIBLiTkc6P8WKBexjRZpTRF8BE2slKBg04moZpT0gwQAPht3nHMO43a3hyJK2dhneKZYEK
J8Ye+aCgdzw+vFUsbcgt4r3tYL3sAHj1T71RVazkUZEapSPPsthzdbVM0x2dNgP+gLKrgvZJi30T
PiOowEMrOHUFVEaYfrmJ5FnBt3S4jOnB7L4EdQY9qYHgQESrprrmFvVx5RKYbSXDjrJ2fl0KUuLc
UkLEWtvk+y74HWk3NlM02gJ2wVRZdOCVXwiYTVF9bwF9cF9H1lMho0EM6l3YLiSXKhR6J3/1foK6
tyArNVrqrf2fzVHGJDzZ7h9StQNSBW0dMnm1oZ1Yr2AZu82a4IwN0cmi7CbvTkaKHr3upvcrQyKx
ZmO3/1hpNrsathZM113ppF0trDOJGn4JLtjGVDEB/Q19FiFOaJ6mARfwVMkRbyTkLSqVZQF2jTR9
JeHWR1TGrav3Yllefh0C0HsH9sN6EFhZYuzDrvIh5sRiYtmfDchsdE0oCu5/reF/KYEXI9a8LX1/
tXvLIZ0v2dorwfNFr/wqtorAF7KhyrEn++lduu7WQf6y5Lot+rUXIN/my3WK9KVadW5EHI0Di8dZ
CKHGgk/cd6u85WRP7HOP6JVbBbTq8hQ81vBunrY9ex2bs3pwYspfjDvlrCPJeaHelUOyNtOiFL2p
mvAaphetsCSO6Sc32pT1YgLlnGm2s/RpFzo1v11txJd6qsuX890+mlI/ysK0mXUctVFRcThH43KI
Q2+cFr8AdtjSK+86mLOS//M5ElPTWQUJhvtgts0yo2lGp+pGqrwTXN8ZmwsPaNg5b/cu41hmHEms
v5FkaTnBvJ2yutsRiyEwkl27Zltn/yT87/0o/TyD5tfbRVLjSP9eq4E8IKig7hw7S3hlPhVsgTt9
2JQ342lZv6FuwfH7wJoyzjnxYnn+gr4R7X7iPkEPFFhPfMjNDFV9xgV5yO15ovYvekbIqvbbS73G
hG7N7S0lj8MPqYnn3fsCjqdQZNSJO47wZbCWxBOYqH1Mee1ckDmCSjTCjZBOrhQf19WrxUxhB/aD
v4ml5/cSjlJ7czwKRtRqlgVmIocfZPQ+uR6rTSSF2/zO+cyqy2rLMJSO3umC5PufFWdbKv14fE7e
EJbM8AkkspQaUvFYOs4M6yE28HNur1+sR0zgIOIS8xKq5uSxRGhfzO014fxRwdduWJ4KSqU9TFji
E1GkBWZUxZJap6OTK+p9cVmrWBdkqaQA/LQ23LOOV8HBcZeyO4Ypot0zhbDpkEBzE80K0OtOPsEr
e8D+TTjlkkTMZ+zGDUQKuFphAlLYjGA4sET+JrpvbOiQ1THfbfKdhjP2V1n9f28wLv0hk9hetRty
52PneNN4MraNXaFCbXDJEOfFIBmH1zkzdsT+08Uu6QwyhdXxz+XS9/Ao6GqYw3eH3YIbZiHQeuv0
irzaN/uGmKLzGiRGCRx3h8wsIBuvTtQGsiMdnjFOfqEbvKSCnM8d3EIp8XlyWi69OtMB+cg5hIX1
Tlg07w5ydGNxI23TwMlW9MWrTYD5wGkZ++JJI+wIXe8ynIF6BkKJiY3kx7WedVK61AR1Q+twzyHo
7rGUQBB85/agZZ6Ew2mvpR3+h0lqGh5S+Ok2iZOPsoZpGXKaTdkxVciRa9Gos/ix1YUFdY+aHYeo
LIFGiziEIPqSyOWMIV3JCws1iNd98ZBAv9fRG6nD3zka7z/9c1/Wpr4V3cBen/L7Gs/mynXCb4Iu
YJv+SFILOktUSWFrR4hHR+XMUwkIz7V51fzFrZDcQ8q1moTa6kQXZLzJuAs7prVUrzJF3/IkXURC
J2bS9Ako5w51o0oQ9oP01Mv8WCE2BxrhTKvwTaVRRbwfz8QRsRf4YwFZlr1ullLshr3vF0jcRH2n
clTt14qYjEJhAHb3Q7uLawLF3gmk1MQPtASxdPOGSMmn1T3EAYMZEngumq0oniXp7Gow+SsXJ5lb
6a+M7ULcuXruYGA/HbTjYq/bEMOmSIbp7Z7p1tLX324DOluu7k9T821S7MQRtzjcAKWiqPsznuug
Xk/gz0FjWQU1NinK0kZRA1DrWbPZx3O7YziEGVzaXKaAWu7SlP400qqQy2VfmrNrZdBeuiq4+AzU
MKi1/Q6lz5HrOa+i1XOims7HRRiq7oVClqu/AkThQ62X2bHE56fKBWjpY5Hufp2pj4HM7KxHhArz
eMMOTIfZr5sEuwujL4/cKa+mgcL7sRORO6Lt4fC0wytoKRDJrxniqeY6BCTR1eepyFfYdQcUbhB2
lpWBckUccHPS8TygWe/pL+M37aG1I3eO8AjKmXZ993hcNaqltCvSbMuhAwmQJolfsmEOdxN/Bi/O
wUtXnXqGJAVSj/i8VswNHt6VIQK/Jx6iNPQs+PH8UpLykRbIcC6FGT77AKjHeHdlTmUrlBAjip09
iVnKNTAhyxxC2pk5cZpHDvkPl1f1OuYSmL8BJ6g35Dt/W+kSbYsKWjM2g+i/XsBQbcY3vzEo0fa2
QgNZIG7po69DZDciFOCZjNYWTMj4Vr1Sm/KyLfQTMWONMrwU0r2P0B8q++m8/vh6cFT0JywAquO3
MR82hYH9bPklWKKDcx4ZTzV5J5+yrEHg0fB3oWaB9UGCnwsMYSaRXIYGKELO/0deD3/ozbWabbWR
SOsezFJ3uK9RLNnhTQMNjncI3hfdnIMnzFGdx1eiw4m7UA8HQzHMzQcfGMQYa73Tznumyue3r7yE
8gHZ2yQ/mGjKvX+KxJU2xCJLMRN/ZJhsosjQomqvf30d/OA72JJCg8QnVtzLDMOaEjegG6vqqk6b
9H+8pg26O3J+Xj4xIIFnQPvz0uxQGQ3KNhJQwNBs7Fqh+9Z6FdcP8FFMXJ0fGbOt3t04DGmp7eGA
aydRCoNsPopMiyb3D9ojaV5yzE4uLOLiGBr2W+FT2iVfi69X1iOr1lYQ8uOSdhZ0EZcfFjxHxXnU
3qM5j9ImPTHE8iLF8tJQOqP5oX2YdkpUQnzl2g7E2JijlwBMO65Aobv2oShu4lW4NdYU/IWR5qCd
G/jfKSx9Nx/SUxMRkTopC3kU6kpeUiWhHf2nY4seqHDOASl1BgiuEbNJcrussyXV37xfw5T6ZQ5D
/YaI3mB7feUFxBVc7CpFxvaeJPop3bPn5Hs3qIKNvHT6EnKKkULrBum4m3J5tyrz1ZuHXXrM+AL9
Eu8t+sYg8FGLuREARzbc202PHmgS9zyFd9xIzPNEvydI4c47dVYvuV7rvucwXD6VGjmFPkAF7D0B
FeD/72JOdomHsBAgdY0Jl/wUnmjDDHd5K3wPOxy3YIXnGNB3YNTCliTCYM3vU7/uXPQHzkntmHGK
3V/OKa4/nNJDpO0JAG+RlfutKqzwa434dHViGCgUUkOWNQEIwBeVitzOg5lVWsW94Koao2/8zY4/
+Cm/+FBCyRx/l441xSEK07OWHjJI01tdzllh/bKeHIPwV3WWvkYvCimPP2GYkiZy2djT/IyBbHmo
v0K8377BpNsQj4ynUvg52m2dib3rPHHWCj2QSDSy3zwmYzwpFSNsrOg4PUxgaMWwR5JRIXx/lJyo
wGev0ZCrixu0HyF+A2d+TlGpFUJth/7dfrhxmiPvNQw1vN4DeL/3lI3o+ZJiWCwwMNsWTlMAYTKt
REVq8lKBTQYxf82PA9Zi6K7iDv+Gtr0P/cCkniijPeulcmukPcW8iF0a+fEcQQGZfGlN670pnauE
icK4zAuhEdKzncmKvtX5kOAiuhWu3flYmxVqRr076itdnAv59KN/oMwhOQB/YXgHJ/wnOzzu1xJr
fbnkmvBzxJEq6tvOq90vr98Q2m5B5QaWqdzGi94td+UpFik+V/MYYAEJbSYFipMSiKFiN9QNotl2
CsaeRJDqRT+nvmCPLeDFRJpD2WthyNeToBnWCGTPqzcDi7xxzsHZGKlFFNT7ayxM3H+sorLK1eFj
eZ425j9DcwL+zgJqQdFXBK0onR58s8CyAqGPSd9/8kyt99mkldlItSAnqAaWexbxXg7vkFRQTL7D
nUkhgNSwzMPtpQOJjjEkK/JL2nvAVDyvLs33LSSXNJUY2Cj6VbILPT2LYJolSkqjfH9Tjv/vV6NP
D4kzWspDXsdmPHyn2HrwmfSEs+W/qVxQ1tKXwM90nsQd3UtZn2hjeT67rzPo2hO3eazxbdC7Rwo1
aIPUjHJzwlSWgPSKeGsQSUeyQCUszPdrDXnt0oBCxIn35CtRIlq7A9Pg0+kUYn+AslxFdDTby1JX
4JNVNUrlZhXsXgDUsEpZTKhu0vMNAr0JICtsscTx0UReiGQgjJwQlVask9HtrH+gmWAmK5iJENlU
BkMgeEX/bzF4O3gV0OLkfCmUhvxrW5+J76b5MCIv0ygUmUsJ5rRn67QUjLUgv4zW3jMKsqHEqzgv
fuZRAqJNi6ClDSi2NonUIHxah+s/WgMXcLezq9a+N7686++2UPr9pOZUAEbEKlIjGYXnE4dlY852
YcB2JGeK6grg810zMsR3lzMEkdnGpo5iO7iHCl3W1pV94jEIet9v3cZ8CfrB7YZ4LUCMyMXjxC5w
I3kT7QZUQ7hTPJRs06I7TYyvRWvR2r9NynrUZglvAVDojfsm51R1ZEYDsRDaUZ5JK20wNVDtT/fn
RY+tWKpnSIbuJY+TgFXi3ydLqQaLfa4vfJaA5CEYDE1ufw/mifq/051hRmig/zjWXXDi2zMr38u2
aTBXGuxp2G+RDbHD+SEoVxpZPORuAMFG8ouOdPefm2zk5TyJLWc9DbAwLgG9MCReAank7F7MMhSa
fp6iu9MVfq+5TmUi2gl78XeRmoUaRN9JtR5P2E2yJx2jkJt0Nmoecshd48HcqbnEdDmjPLBJFxwe
DK4EBWJApALdtGfDCEzOjQC1Jyy9mBRKqx2x9rgk1hyoTVLpzpkh6G3abhnJrcsuNWSyRbzmGm9W
cQ6Tyz0WUC8gRZ8fSIKZPDxXA8qIFvscMSGIUN+6JBlfueaYF8m30L0tZtDve0dJPo5crquwawgB
d+GbNnZek8xbUtInPUGCsnA/Hzy6D+JbD3t0juA5sWo0GeU2bX/0/Y+n9ud41SamWshoeILuVJti
XBEasX/03C49OiTEe/WLZN8M175K9Ce5v29rXY7RQ8iSlw9ljHW8nKra2H3+q4n12An0gNulvLv1
qavGmy6Lmh3+UqmDr1pMfYIC2FFVGKLYno+NdpV1C2ZMg3BuBl7O0OiAjWMTBipn5bxSLXJKGCle
p+03T3yIujy+lnB9PCcYo/erbQVJ6CTGhIYzbucbtFxOUqjrtzLmPnmAGyS6BhskncWWyUVZQpud
/UDjYkxV0ixXsIG8e0qfw8S2QNsm5xPqyuY91KmygoCui42e5tWIlOWvCqLwI/zqPmujZDaT+6J+
15PzIwVKfQwKCt9IjfCNokKmU/EKMGrgYHRCgsCy+Tqjn2oQ79dZiSc/s2oVYXk2BJ1dBUxIMmVH
BYPlkEhza4aFdrjKZuLSee+MiIjx6WCKXyCSy8csrgLmrWY6xPBXYPQebdbohhVCVG5uQb01659I
7jw7r5sIrqJziF6LOrXl1c7oGhtqZMKdo1wvJbw0+duptYhJk+3KPsFmMXUHvfKbMxHJCsLTbqIW
XPSFTeKzh05zgXfUCHL7wJk7NZSK+SOMzAarO3gauuCyb+hnS+QBQcRSoo9bVPng8dpz1vGU+46r
OSYF3X25qM+B9gfynhBVGvb2e5Dk9T/vRk3zHjq6jewKRm9b10Suq3KvSGLV01fnEzyGqeYPQY9T
BeidQh8akmJ3JwuZItO6MMdmsAB42mLqViiTE2aEReLDsG3VN2xLKDZWookDGhUVVRRCw7pDL+TS
djqK0QTYRGivrbu/Q3y+pfL7YNHddP527uRN5389pWBbuIP6+b7b/8v8MQpZcc/0t1fF9HvGX1TS
wS7WQKLR8J0yEy5j3QDKiXDQ/6u00xG8ftj5dO4TE5neXpHXtl+GRT1T23YPwwWblAHe/bFfMZEL
BzlGr2WbmkO1bSqAn75PBAAjS7TaODjTkmpF4mMCounio+FS/58kkOY7aAEFDIGmvF5NI3QDa8JS
spCO/C/67qvOqyyOtV3KEDruwSXhnnNi2bQdz+oFbgX4fJMSDBeCY1WdILH+vVD/OW5SepCmlk36
HkkbHqQHZ4O9s1RGJNZ8TfcF2AwcQ9gjSawB1puDi23fQ2m4eiMTj4mL8yIEqZOYEzMXyQh9CjsC
WRi10mRgsERkJAaUdW5n25ld23QxCu/3EENO8sx4nnUnnOBukxKtiS6BdPepKIrkf55/7Hqt3E0A
8inkwEW6faJs+Z9qI2VK83L8QrS9va4wHf/fUEBsICQCPkm1ccqvNeBRxRPfWSyaeOjqHRZEh4jV
3ved4rJELp+a+u+RhldiWJQcncSo5ant6d0KN6B0TWJ0TX1rjkn3RtyBLeiyxPMXhheuUpnrlbdx
XbBhhGDuyj1uUO8UnN0Q7xpIWTJrRvVlaBfsBS4swuaFulMxQjuAbYqsklwrcg8ZUcr5Bj+VMmUp
3KKVCm/yD7SReCd+hJ1ViWW6c87BjrWxlApeFWTiEsn4ex7rf+NMI3eDZT2Mq1NCeWkKVXv6h5td
/wNkksii8c+jGI85JHGpAEhMt2NDFbyRXW+UJ6i32Q5L2BNYqhMu+v5DHRbrFbIDqCZPO37sbSS7
Ge3X7qOYyJjBkm6bQWR8xivqGwA3ugkpl4Mzn3/9qSRfDnec9Ne1lHN4JHTaAD/5Vh+u45lBJqPg
tbaOasFnZD61LMZE8Rn22RMGdsCCPWFKVEOyFsE5cORvzgnihjL+yUEbAJDm41phJ+/O6+Esnhtp
9ErMXrg6yriAhGg7SZ5FFMXCBxNIsVDVuW+RbfWQPvHbWFcCRQhkAjvNgir/gNZl3/E5gFUh74Hj
qgBBLln2BZEL/Ykf+ZmCx5anAVzmQ94hgmEKxs4gGenSw1A31qMcJAAmRhamKZ1jFmZxEirrpn5k
f0TpkDvr12AZEZ0G6EuT5DQoFmvpqk3YLB1GdZuQeq82YoDIcFJUAFGn++qJG7ZLriRc5Si3cJBb
sIFGYsIVP5+NmZ3W3Hv907qlhD1O5fsaEo+2sx4caRvEpr0VBQduuUIz1SVq95qhXvtEUcWjUU0w
Yvb0CrNxta3xI63eOmNUD1iMutwmFTehOKqsARCsRIcxJ9HpzqQNaKC3L1iWrPO1/VndUJE74slo
m0+PvGfUtqnfcGg1F46/4iCL7LtJKcyyIr/RpMYI4EyLzju3tP/0u6wvxr+aoMdpz1GVN986an5e
EmPym8TSx+ArWlRSXASQquHsA4p4+xHaxpxISvogtiQkpIJqMnzYvkEMwiGDKCZBQp30qZOGXIdf
tO+MbKZk5JeB2ySMofid5AXczGwMURlS3+Az7hBaePy6zo57thtSGceIVNKYsnsrEdC41ZoHZ9zO
LHSAWkpguqH6IQyhUFvWB3izCZ/dxEuR4o0RUkIAaVtSvOJTcNm9H5WaEJDZKISFiK9+9XuHugd0
ycZmayXyT3gE2GW5hIewd58T9N8fzwbIuUwnlGUZBba+I66lE6X3KGrxvyp6Yf2Lco8vjI7BME3+
g3muCg/5TcmclMZhs4F7Kpjogqa9sdRVXN19WySp0aJu/8zhx7ucgPUlB0joqHw/wbgigy+Pmr/0
pCZ/j7LkoRM1DTjXoirY8GxKh8pOJmiIRxzmDIbWRRct5m9QWrv0mKIeAmP895B4LKLtj9E/eaCA
tmt/N6p8a5W2xaee1sNc5d6tkceusQxAsk0FpNhiJzGIo3okt9urqr1lgyIpPRq/0arhqf+6pGbu
PHz2LOTo+1XjsuZhSH09xvt6FR//Om2oaXPdzl+m2Kv+cc0UNYD3IOfNE35hEci0NYCwWENsaI+4
gZ9GhYGZU6T0vQZBK3yE0VZXQeHVvAeMAkirZ7OUVYCOk/gB8ycvu7TFxTh8IFRYfychWUKjuP8S
cPDcvH/4zz5fBhMGbBw1jtyZSA6+e7QPFe+jwibqQDZkAVHS86yaloJSkMCVoybNd0/YYnllVrqC
w/D5Lb1UWAsDR+Fh6AnwAwV/4dV0yIDWO8J+qlYF70vcdl8PQalhT6yGw7wX56JbFpf7Vq4zoVzU
KDU+6HyGPEZCIHuuwcYMfHinJES2UE/UkATGkfF166XGK/zapf3HeGM9t8BqKHfgup/UHBNHmnGO
UYWLDz8e1Hc+i2PCB2joSCsC32nin+cwrEYhAXYww4K/9hpGjzH29CinnD6ZfYrBmQIAZaAF9SMz
Jg5tYyd8MxOHLD0a/xAR/Sf/8/BfONiHhbp4+K4vfLchS2M8ZWIDPvI7vLC4x+46pDKPDJUbs6UK
mBLfHdE1Qf+WTg1+IlKlYnaSOYCUSdzP2Jf0qX73R+J0CbMvMHKcflw8jB7/+b1JfSNnhTr8F6JG
nlFE1cYZ2phzCSOMrGBg0pBrPh5TxMUGb7nfs+7EjW6CsR3zEKGGT2dnw+Jc8ob6tXi80/8v8ijB
icY3474JGKHbwGBF90+kAAiQWlFg9GJ3YQA8P3G+PFvAzkYgCk9x8K6B3b6FfqeriXaELDA3OCyl
20/yi3QwIyxazobMAAFH+Mxj4TWkAKaHwjcRXrhmkTXacNKEdOHBhC79zRQoM5xoaw1m0yjNUpwX
y+sSPHu2Qw91PBLUCfLAnGtMoGD6Nu70Dsz5/rSdI+dmwJ8NFNzRCBMdRGARbfIPiTjzcCn0Rkqw
qtlZiB2HpV9GINRaZ4esmceJNfcHSH2mgIGQPZcorUU9xyRj7feJec/lEA6r+v8IusuigBMKyJnx
9TNyBomDTSdBn9efUR9wwpS4720PBk6Me1btIDQpBKGNBGhJvjBIDmstcfTtOWoP3pYEBf4Y0jK0
z+Tl5k3G4qma/5JWlRN1GnPimgL+1sCuwcBFh9mk9zzsVKBeRHPNqmYeNkbBj7Hdl27XmarpUBpj
hWQICbeuIVyThPRmxZ33j+RHw7jU4pKi24G3xL4wZjQmiadwI0QjcXhCcQccIC/7aemFpBnKWRom
Pf+l75G9H/BXos3qK7N1UJIiJkhqHnId49ONf4kTfMHTq1U66PB/xooQyhChyqRZZtQbhtzvedkb
EiRII6qR8ql9oq8DLyyGG07nUTQ+gnE3xOhtGUqdBw41oAVE6FEFqkU1/6k3yPhtquRsTsR0zHwP
pZWZwyHbyGQHzLeUNmS2FdbA7Sp/DwoI8QrLL3FoXkykzAaGifRW5/LJvCCKN3Z0a6SHG57CYw/K
dMA/1TT8chkGEKy9DtYW7RLBCHz9C4x+fgC5Z4MOt9YJMGFWCI4mfVQ4BmwqI4i/L1O7TmxQA3/L
rJSEZBhPfr9ViiaDvRv6UTePJZo0uv0MJOiNV354fl+vxQkNKh9zA1LqJamE7LYko5Y22fGBTZyB
VkYE4ZPhC+RVR2oZom8rGln4xgfYYB+9SvLPRCH7rqIeT/0gwgMXw27qpOvao3p4F50H3ZabdWbm
Z3NyFwgBW8mjoPoZUwvM7UHGBNYvzZ55Xz5MDa8MqGQSp0+V1g1oJHI8zMod9obdWzhB/PUFChb6
nhhl08GZXH41/jWivvxTGM9cfoc2f7wYMDiagxHTciYrqWLxm749gcfgLPx2Jog8xyHGl/zYK+7e
e2d58s9OVCeFtw3yUu+and9H3dUhIvP81qcTuhurQfDfxwflDYJrwm6pi2Q2p1IwXEyjZlp8z4Zd
aHN1K4ovmbfYzkeFklDxYoD3SBLURKmzpEgEomIKLKZ/rAx474SoAJAlfxBYG0oQHdfTGOSllMr+
hMXfTtKzvVJlEuH37d5Jxrb426wFE4fKyIHVXgYXcWPQQ9d+rfEvrnB+tuHRb3VkaIsluavb4fyB
sxdfzXTs+jmsI1aw7zdN7da/Mt92Vy+Z6uMBJ2Plsu8Fd4eiq4DW7ie3yOBpI8MKJ8sT63DUg7Wa
27GOBmX8Bj/Aj7yhwLAMeqRWTUhxdj8dH0l977rCC9jd4KyLdJ/IjLmI+TTp7apwyHPVb0GT14c9
RxRgdqLAMn4J/vk/HYNhGcJ2MEkJSkV9uaq7P36okhDonTEzXZuuCREnjC531Sb2InVHm6630gv3
8jh4Y73/GoSvHxGuM6PdSQU8MxtexZY2CsYlk1h9DLlpCm9MxpOPUtcCh6jTx0a+xf5Vq68A3pnN
qSX3T02XwYwvulULVDxOGJTgY784DrPE23ClnKEiyWx2JZ4rX2MrQkxRj4X1A4VgFdvKv4Zy6tm5
bp/N90DyMjmIzTN83+ueX8eYg2DWX7fEz1lITkeOKcD/q9L+IahQvTzNFh4DViafRzecz5Hqt+UI
ZgRjk3Kecj+H+w3/D7K5nu5bDlzR4PB3gSZrJcc50tckbtKQ9Cj56kIUkTz3hpnHGJmKlH4MlMwV
u9lZRbg8rTpNJJRJGAEn3xIzlQFmTNJlhsmRE2VBQGRvsTIcMGYRZH2+FREvFNzfwchPzQqQcY1I
OPSlivrIBsbWQPBpdLJCxO8K8hVHbXuiD/+3k+08++RbIVnmO6Ti+j6RAx5fieaCuNSQZeEYJ3wT
NjKftp22MaKAJNgS6II9cc7ObcW7Nnlhso/Waco97YM/hQREGer7IPnQj4LcXStObR4veVuGPWE2
huXb7h4LeOtKHdbkSe3J1AfWu1RUYw8LjYHbQbtwCB9J1Vqfxsp+kFkuoG5E2Eltbg4ldfI/hAH6
06NGCilVHuY3fUSwXkBIsju7S+e7ujrm4r+s10kBs1GFzaBbHLeRdIoqXG0t+LUzZVGI1Pf8XdsK
i1B+gck7WXTCBN43uozQpy7gGrxNs/Kr8f3j3IeBozehnkKShckIhStP40RMZDO3+VWZu0tDnO4M
7rN6D3snTHCv7cOsyNIKSggdmQ/wFUHlcJjlEu3TEuOamQ/478IiHMU3kTtBGyAMgdrymjq1r6GT
VFj26B8e1/zexSQiDGHCL3l9uSQBKNSEO4Sm59iQVN2aeBJBdc7hKdcAHU8tht8ynQUYV8a/+jAl
Q45WQ5yxdXASODS1Qd1cuDnEywaFyV+70usKqpuX7xb0ExzVP18YjP2Tw0ikb049+WqOoe19ixfe
Q6JqqaD3BVdM1ZKjU7cvqnGGOGdalWce4QiWhsOmruFY3lYTNvrQRp2lEFADoRU1chv3i0dZWjcd
EOEQe6TthT+xNeW6odvB8Fw7ePTH/2R0lT8MEkktyhUvft5v7vY4IaAbY3Y5EFmaeY/RtAKVxi3X
pWxB/GguiLZpzOi8Dl+bsg1pv0Y16vHfj+k7IrTB0dAjtrKMWM3O0oYwkDrLytmcVs200foWiKEV
e3TWCNC/te3SH2D5fI/OlyekNKR0LclfwPPV3YIDm3hyYv5qSDPpjyHSGDgso089JGE3hL/KQb3a
AtKwn0SVogAeEFfZ3yxsOmWjzzPGvRinL23vtoEtGhp2cmj75ROCv2aTcLzj9Ut9n1NBXVz3oPFW
bZev8N5CxVs1tf45hKbC92sfFN/O0UzcJGpK5w4VDb3Yj8tYILFoCzH+X0JjGFSVtdHIoKkrWpHB
dleTAahA6vIabklpnpJAI7s6sJ/c/TbH745fL3s2J9045QDVdAdVWpAz3pwwJpKxpV+OoHj2OD69
Sv5I38ukmFKKxtgWJcfu4iRBKgdxQoIN4DIWv+Ay53uH1ocjUHbizaBd2WKsCj8sqzcXYzMx54T3
8B9p45xGuUS7ji/KGHXMVnY2Zyde5of76GSca7NxQysY8O1wemCwm9cYiEmo79CLq4/n+NhtvzA+
DpGmfNEbsIyNkS0IOY7SwdRX9on1t0bhoyTLDUGPwqy1TFI8iU6dRmNO1P2r4BbSY2J+JnrD7Qc3
i6Fd+fYBud/6/NAuMhqAS/G3+YjMqbzf+Vr5jGZVV9aJAKI7mQ/wWxyzvIlZjhQb+lKDcjKfqW6P
3p5U1HNdMUE/m8RZNBoPDnfryfMEZq6atShAoKJYAU29b0094ykKNk5E2mgvhUnDfJSmFc1z8D99
7UJIDHZswTsTeRAbeXhwrLydZQ3n6i+A83eoOiQKDMicKnyW8OSCInGhgZ75kf/UbTiOzhkCViF3
j7dzC4toQg06/+VSpfCk1sh37C5m/AFamPvwmXq7cU8QnY9e3KFa6qI7V1CEt9SMPnY1sHQ654gP
51bW8cPDfcjrzkwnURGbup1yAc0b2PTs9Vq8sizLzWDxpXfMxOhVZD+dGkw4JSXCmhAArap+AjdF
t3NA6scJcwRIXHemO4Ak8xdu0WXQC2gaaTTqyKJDl6yJx9VXKPjCuw839T5pIhNcrOavkNzNGiM1
QpiQMJyp9Dy94zrdXEsfWUSTqOZ0vdKc4gJF2IINdeEti7RszdTlx/kAeSYJ31aTpBRDI0eidw5K
c27yC+G+S0H/iIMGKcREgAexDQiFvGp2XHphohXuSAxyHhzamFTj4lanwqx3jwpNxnirHtyhGVNj
wy+qyED1HihbPej+0+MlfhxabML2JA/6pYu6qa4E4P5z8IB8VpREIIL8aVhheAhp99eVp0zq2ks+
Z07W/M+pB5HeiSFwRkFc4fzYwt1YvEO2wIgvM+5UlN0YuyrWjvhpZXGTC1Pnhw7aStyw4/Cva3az
5CvIWJ27nBwKpUWJar2UvqRUZqzGamHDnDmlc+VgDHBbKalnzclykkfxDhuohgHGFG5QaGv/KbZU
s8khyJVDe/BLXidRxTojRIQRk+LlBP/LUqDt3D/Oxdf9cf1kr2iNUlEfEjg5dARxbUNMu8jT8z2K
vKLAI5xyvXkzQA37oUIYaEJlVoN9ew8uOsn7aaoOqWXWUIEhHmtz6nOTJLxU8V+bhU4QVBA9Mer6
PQxMXXs21szaVDcOojj75mNUzySWdy6o+nENKuROhNPJx7iywBsVXGlHfHQHsN2c27QrBGsqJqQo
6XfMfUv/96GzXLbsD3KSn11778hM05H9TiKhbZDuVRLNgh8K7PqtyhuSJ8nJ6kqn+AWwx8jK8I3Y
DktGermcFT//7dE2DmepKKh9J2THknyxOWCPrUvtvh2Rx8VYDEq9XrsF7ovfzYZz7kN7YXvGPPSG
GDLl8X+tKV5jxCGu3CRiLPkor8kGZO65yPBF9vMqdV1x1CxIq6wam+RZu2q78zXATiMUawdqTduL
IFk7X0dpso6LFJmKtLT7ut89sn+xkp4ktpv21ys1n1HGTvYXeOE1n/F5n0aRxcoHg1W2LtXrFRTw
DpH9/SVa5pxrAb4apct+BPQtTrO+5YyCOEE+t/mplsXhFB/Fh1NHsQXKr9VrceZYXSbSa6Xq0kY6
CbuB2XFj22on8/Go4ZBtdVv6JtMG0wIpQP8jYxPz5U05wxMkrcJyb5SNbv3PdcYvnnaLpt/u1FS5
YSCQoxrLHO1ocX/9V5n2y6a14IcgbwhvXMpJSeJaC9VoRcHMGT11hHSRVVyi1pbbVWwuOUknwl5N
RGKrOnmS6nQHGP8ah2mWNB0VqrrCYYS8c6CndxF50wd/e2dPFW+RYX1n2CKQUeDKQ/NeRasPBjlp
r0859c2aDHxYghHcbLNT8oHFgRt+fR7U8mQFTolsd4zn9j6i62yL9O+XelghhJgs1FHHcCqKqcOE
cvFyLMG9is1c9c22uHVuCfkuV1GgUnlSLm5XpsmbZMvt014ZUrCrqY7pVz1rKcL3TnkT0iCF0Kbb
kaDfq/Oyz8t+DcfcepeSMOlxPQTguG9P+UW+bUI8b07AyZFRmNv3FLq+yQ09TkGKUGp6NVWYZhat
PhTW8QRRzNL8Ytzm6qY6bL5D0gJFYkOvt8ofHekqTPOW4fb7Vv1/3+3+3bnr8ucHtzZH+cT89F/Q
l1j9uloRuHG31zKIpr2ewwksdoIHwpIQ9IdtLgQ1So4M8Ypi+qc4/lwEhua/tjVzBdJjFjbFnKS/
RTf5uZfKeScmdZpcSGVPICOqnuJSH6YngVY/8J2dKXsEIXgiU+51KQFa4vZgqf17j3qfG2RNQ4Zg
rX5k6/SRy8JqCrRA+z2az5/LW2H87WtO+dYJxHT62/LZ3E8S8B1YNL1rpqq6G7v2Oyk9C2AxjDW1
Fqwvxu1WaABpz1ZSAcJfczRKl/YbmX1HrX/9M5H7MknTx93SW48E14ONIHUxCX8iPTCvLExFaK5g
uJ8z82DKucP4tRwRW/Dfq0nRkNdge/f6GYaK5mz+UuAC0P9EKd5vV9UKy8Xy0pp0wT2/dQL+j8C/
jbXfZKpraZyRVH+AgQin1D57nK+HSKoSkMeK/OvCkG3ZB4wwZZb9sZOeT8gjfLVJaR5x1qS0Wo1K
3xo3tA5CX3a5gp3mXIH9w60q12OF2Uqznn8i+TiDNNbe6vl1CgPHfSGbuwRnaFE3G61I5JDzIjIC
0ZkDPdxaZ1yTQbgB/xF+tyzlIbdvvzGn4YB2EfVSoM25MxBAAfZp0pBide4W3OChMAsvFDRxhzTU
3OVQPqZeza2vQosOutN5EbRwdaufFCgaP5K9yCjD0VJDgnirorImjCxbfZVTvbfc7Z7iM3uaImli
xdaC97lmgqCs7mVUV62LE9Ue8EEg14ketR40wVnfgb4pITZWGrgGy3+kbvXd03me4RBrxEgR9tFa
dffcHnNDHKXwCofDzp7BFjxvYYCYExVuMiBNmCJFzQ9dqAbH5yjkIf4uYSSzP8NXZf7r3bjzqZ9g
ZQGsJB+LeGzfYY3wrT6bH5C2KG/XkykkbhksGTA05/dQPMqmMgtf5a2YDInD8nO8B5Ig/je+eZ4U
X43ZTGII5x306adbRuKXpFxchdxnC/aOd/U7KB18J5RbEtkhtEBYKvk5fYv1WgKdE5SS+x/Yeo78
V8kT29INsSEljJx5vfT/5uVORn0rfui+b5UPlCdXHsjXbgzdP1kjhL55MI+7vMLaAJiyalkFAicG
dazJQd4QknqrM7f4ZgCelrIC5AYBgReq5A86m7nNUzP0Nq4MjDpnbO8FixnKhqUQKq/ASG0MQI76
AqQztLmeZKeJynD9/FFXN80R7Bsl4bbzcYvYhJkr8g/nuQv1jW31nT7hdd+leNhhaoMawtzZnJQO
brGkf3JHFiIE2zvNpqgwsv1rhHTZ6nupIb5LU8dz5RA1ynLJ8uY2BwGu0WpNVq039V6pk+vk91Ly
6iuMOYMfhmZqCNZX394P4R1VFoi4p+X0mjC307qyxu/CSxmda8wxnemtaKE/rcnEyklxbhjSJZYg
0/gzKOko2Wwga+YDizSQMwB5ESfTJvnqwST2bdkrt13eIGXuTqhRd09+kAgVijZlNNAhmMjyqYoI
Vkad4XExjH4L+rqJsOv0ZmMMu0seOpWS77YqaL34ybS3cnZAcutXzPan4V3mw0p7g5iRrGqDVz4P
8CeT0SgpglakcCQlUB74+pO2qullTy9ItEi61V/YjVjRL8y/9yR0oIJrr5BjY+8A6Vtl0m5MJdRz
KXjI7chykNLmm5mjEzoy/N8L/fPbsYjsZUKDVXgpFOSgpgptW9X31Bl8+xjkFlb4Hy8Qb+dVEDgj
GvUA888NkbDiCp46oykuXxjJVdIlvre2kzJ6I8acgdueU7T0S/1AEwwBWMs8k9linI8T97HjJoCR
ykqHZ9uCYrOrqUdfeH4oyXc1SKQtKTpijjt/aIhTbM3Pl8xnDagD6Y94jlMZvWIJF3aL+Ozk0C2Q
dr8u3ZAcxzi4nrtrEZ7VgeWSAHLsO6A6slQIb139mio8ecDZi9oBTF89bY2eVAays6N7UNc7Tvxj
b575+Suh11uQRKe9Mb29jQerISKTyTXkTWdMLr3ew9846VCW0BhPn6MPyK1RI3F/1bUmxbLDewh2
wnCauGeIEmX380XAF2RJh1GfAjBiU3qCqMbXn4nJ5jZUw/cknvjXB3ids471MhE0zJep1K9p8qxx
sjr+PNDHJkPffaBYdkEQ0ODbYxx/+8WUeX2wV1GXigRc+vAB/2aRDRjdI2bPyBJL0+lBBEam074J
5KF+iQsVUzXh9QJUtArWXeR6uSywql/I+GYbNsNBb70+Ud2HC/7kvA2DANpiWNVRmMfNUFDULfV7
h5bIfqaakJJ5AeIx/KKQ5tBebAsROsGB+nNg4JtdFEo6UjD411OlP2lH0EwgJrK7MatKng/nHMwP
2xe3Q3gAAtA0EdZj8TkFI9accAXSuXTcK71hIcbGFqYJfffI+6vsVy1wl2TNdCqv7y1SFW2VSS0l
g3WcnIThRynvqJ3zQgBh9XoC+cNwE9vqdgu1J7rgXVduLsxLEM2AzRjnUI6o/f3reFAubmOOXTXP
vs+gh+KqnpX1v7ThLZ1Ecywv9bS58C8mgibAuHm/yCSsJt/1BVKxROmLy9z35IbsbVJQZn4DGQdb
0R024ZaHII4PsnjjCWRqJ0R/8Vk8/ZAX2qS8rm3yD7NbHFP3P3WdRr9rBh9bC/dJ71SR9DwM1cZV
6PDA1en+I+OFUinRpAdrKy448GILBT2qQwficNNpJlLf2JRPtN0YKdBmEQXB4sD/lHF3Nupz7Vq4
gcpFt1R6YD5onU8ispmgSGFQG1T3ZXr3O741KiJn+xJKtynSFSQzGJO8AimB+HrzmKl8Sq23Zhh0
1ytSkhzFGoFkLlT4i7IL/LPBmygWMLk8GzLS9sC35Jp6FKhMdIrBwR/4/kddOxfdHwpNNwzaNkGr
5ejG12sWFWnIqpyMxQchFpupFHCu/NtMsHtxItPXutMqD1d4tn33wnAQmxoYbkdaORHw3IVghbsK
aS5UrZrk8B8HBrkQZ6WSMldY91O0ypZc8IGa5+NASmNhqfsWq9r01IPgjHTaVPi3RwjhtpzcANCk
oTUiwtTeq0toW/uvmhF76pShYd/QwXadnCSfo2KdMs2IoiWLGYqrL8LvJ8e11U3W4wfomD96xm0a
8sGDiAqrx1cTMiKxTX56BjCgu1IpCGOqpJj+5qmECrc8uu+mSywR9pE1c5qiaoPhoAIi9TEgBLLP
muFOf+DWMqv/6ihQlCyUeNSA6wIifvks6d53+J8glH8EV5bJt5GzhI/YmP7WIPwqM9G1D/e3S91t
PXlDXXct5t8HNj7jZ/Z4JEhnNPlcuaWiZy/HSV17sxCtRfIKd3wt9fyVtCtKP9Bx7LLzsPM80Bqh
ptvMWnDFnWlcpmw+ExG04prXRc08IT11CBhMb4YdiurM13TaUR2RM2uWUxhvhlWfe7HATsOLCrsZ
Vf0AUZwPcgWhOxlAQghaGioHayacZqmT39q0vVTjhRes8QFtAqb4wQJ9mNWdzp5uyr+uN4XK8PLF
51JbiF9kqBQKTkW4yJx5QUhdZVaDdRdK9rYerLk69sG3icAU4Ga4GaMRuququJfRo9OW7fJSBVcB
FmWPhfzfUlq1Z8odEH3cVk3nz5dxUOv2ObvGSjAXzdPHfQUC7Gqw2kofhkLLPVGtMsKAlSpj/tM6
CX+y4IDEtdPFZpzJvnFY/QdNblMBJoFVZ8V0IP32Wlrm8Wf53ceVzR4sCzHYZDeZgeEXNPj3HwJt
o/NyB2Lv6ffao+w/5aGf9oHBS4gw1WQS47OyalMyqIWnN07osO2OVpNb8+flm5LhmMMvcOMXjnnS
9cRwdhGQe2z6fWiVgxOlDPcKJl6YsmY6H+6YGiy+HaurYHlY+Bl4PgANaJjWPGq2XaoaJ7HjhC+G
WNhq7lbJi81T9gTPiGGzWlSL8zY0hxx0FhCs7CTf2JNwc7zvj/FjMmeCsv1dDYapQ9VPRRNdPbHU
2PvG3IT3RHDMQqsM+HGlIphbtxJQItyex/hxyBy66QMUfaGvnTBVjhPKW0gmS5tf68IDVqwZvddc
IrB/xEc9NggI2O588dlEwz0qYhyGikrIhDMUavAdzWWKpd01IdVufGXr7xNDfsQ0Sc9mRn/dm2oQ
2MSaAHU5BX1CdNe+fKqGYDYo1VYAXU7KJ+XX3X9VGLIMJvOCf7g3SfTaGl9WH075PhyW4Z5jPmbv
4liJ1nbTGdk/F5gZ4DDzfw0E9nBo4P1jgRjtG1SyqjwloqL1lHCn2zV91E/7uD8hJPt0q39jwHUa
5MezBm44O6OrDJ0XZ6z1pEWDs7qk6VTbo0BppMJ/i6BGJQC14otfWR1rtxuZxe01dPOHAc0MmqXP
MSXhlJpf9zYNg+LmrBErtykmpqsIrUuHHZ+/qIb+F0/5iuTDHY2t8ihmyTHbyyLZaWdvLEP7zzR9
KgCnW5R8Z/sSxIn+jBQ+8rxisXmBbtGtyhFoFhL3I0bsDCfMcxrb9tYlkyzhhS2C70yfzrRy6UUF
sU9RSfdrYXhZSJ53nvXFBnuP7CU1GoBNhpwMgzjPYKmeddmHMhKtOdKAE3DUPrrPztMJuCWjKATW
VNCRsJQGjRoztXLZAmja9CPcOSw0rUxAc0KjXbEbQtVF51jh22s7nyTG+2+qjipwB5AAY6UAqj9x
1+QhkzJvJ5S39CzihxNdiMUA5ZJ72gIIqTq6K1/TD8+prdKEZt7w9tGUlXEJYf5+Q9Ux3K8AoGld
EXc9E2TcOURzcA7NoEHotTrUSUUofXGLEX8CzgjtKPPvx3vRZMvyP6evdBGIyQBuWnzsDqF4vX1L
HUw/pSz7ibIn/YJiN2LPhdSr87uVNKX3FCBGXPVLysJsT8HHSgb+51fyGLpMLtGw/bQDI1A9Ex3Z
aNDk6M2X96Zu2YGTeYKC5lsQvudAuLSEktXmyXtyUErnAYuZRxqDGlVGQ/8/nWHrnEnVnU/Ng8mq
xULMsGeMy6rzTj+Bn0NLS49FAgWUMdryr6q4PeTFzrWOaqbQI08Yrug0GvmHa9YSy9xVOK2xDXSB
rypW8R1uVfaz7AZa7H6W8WizcjAf/an3PmaTWHNFh4Ynb0jUr0W9zPHggpiZ9QN8XJRFQtj/BMwi
oEBtk0M2rJZY10LYLfL7UbsvXSLM+X5IZfzF9FejIVgpwCLjc1jIxX9ye+MWRV+Kt88B5pPSTXzp
6+Ag9YYbltgX0cpGeZ/xZnZUOinw8QeHyzRL0pnfyQ9AXJPakBETWQ1ZYABeues1iEKCTz6uY8IA
OXtBna2OeNPLn0dFKvHP3JBOLmxLQ6bIvuHB31PucqUBVeSqw4fTe8zEmYLC9Hrp3DJ8l41hVqTz
2Aa5pJc7tMLvUhPaVeVSfBM0VdKvvKsBGQj/LFYhaMfy6PTD0gfk8gqZtagZXYhEjZ5KBjOQaqsb
auwXZGenoov6LyD3iKRYBoOv+fX7dWIaYyG+ee4kMHiTJYWin7pftX/tqGp9l+NuisiqVfCg0Yv9
zn04G28GFPEe6cCo+SctHxlZS2PT8HKSJg3mTCWGwRXblsiPt+jF9W+YVnti48YD5VIJn/b++1Cp
b4kmKWYMOlL28pWprYA9m87OZnp1vlnOH1O4XXy/wb6kU3wagdyKllvOOQYZRweSVy75okDUSksx
cLFcMsZSeA0eVrG5+GW3ZrF+ZSyTap9QG0tD9c+5k+jax9fKwO4D0JSt3vYrm0CIu+EIJLLYolD2
Noo3yt2CubBdfrFvzloS05DGMVCfZSJsYcLPJR/p28IttC4S9L3OkDSW1nD+FxYrpPJvJ6Ck9GiE
TzyarU1/WQorFXd9sJ+AJtrrpGqUPvbjEmMPQmRyOzSmH2bbM3t6oHASYEd0iu6X+xB7U50dTwsX
QTi9Zozwnku0eL8IS4IJolWPEyl+nKjTbUkDkYb5d7lN7P5WdxfDrvSinTsiz1WwTeMXvbGwQoj3
P/ewQtc2i2Rtg2I8GJOTPjJ6hl23ihiDeNmJmMWn0Y0osRiktfbU7ypRExVsOB9z8QYB/s2bQLjl
wUBxITGlI3/PagDfNEtxXAKj7fW9iXHfFyEAusuYwdOWPzZp4/twTMBQVpddLfa3iCn6kd5xOpbL
xGxrfsloOs+eLPKq6lYu4xKQ8Uou7mq4O1nmebH835uTwqFsJz+dXjT9ltitE+y43Xj2IOQlFSp+
7jqB6Aq9yuvQOYCmqkUEGitWiexsx5NSy/6GS3xIC0CfdtsHUf+BpBgFZwK3KR7n7GWkJ9Yf4zP0
CGWVBkAHGMlOFhcfQCcTcTclUYKMBWHR25xMcBuDNFppGD32cV3q2ZZrs8rMybfZf2v6el4bxxJo
td6bqD9P/m4DhhK2yLViJkNqFjyGJ6AFLVqHBAmV/iXUAb7npoA8gNldadZLks2QF4J4b3jpzJMH
07zinE44PtQlVvPaOuZ5VsYT6lQNxslbfVdbnOO2PnVgwQk6/IbSsUYIzoXBRUsegGALSFTsHm3Y
gdJ0o2d4kLc3fM/Y4KlUlmjEFEThR+4DKvVg1TrUdeg6oPcp6HeZAtMDqarTux/Io2g/QT6kpNF1
5hc8jQRSjYtff/awb491yr6XX0NvEFK85/wLcMVEWH7XktlYupNzoc5OGI7hivTPwfv5rGt20hz3
ULdM3NBr+gdE2z/qy7avSBfN1GH007A5HeCx8ExrYS1+NQdJ3bOg9UUenYV1t00ltYqyupC8WY1C
PfGM8oaDIEkezFabsSldapSc8wzzX1k3OntzT7kWDiIHRMB13tH14wixDsW8Bx+GoLX0jhJEfT5T
a2l+lgCI9X5rp7/LjUq5SlWRlQXTJr6fl6YVk2awb6ryr34BnlmF5To4m2HNne6assIT4coOf8WI
ZKT0OBjeqZ2tFcWzMmwGxkJMhsNeKKFx4rxk/Nt2X8UYMBCvUuP2gIfuwX0DVEcq4e6apwvcBxcZ
DDXfomw0nSlPN7CRwu3QnEd/2N+PhuUYiD/2EJI+855jKO9VHKa1djUIKslRJm5mLZPyIUccoZq8
c+Bhx8eMcdnjpYTwHfjJQy8SC0pUrUC+6VCSXt58mOWLgGrIOPGjqdKa6ab2j19bOBS9tMwKfhVk
lA9bX/GPCnBF297jXnkTGdt5/F7zS7bZqz9Pfrp8hr1UrdXbSquKTYJCVWmsXHPO/ieii2yvHoXN
ujWQ1x9Jqxjs86V5DIjTNuNBzM9lZzTXaEle0nViDlQjaRNgjR+dcBA4tuo+vXH471/zkBITC8ZC
eDRxcPJxfpw0heiBWqGZVxDlTpye+Htg+Tmdw58Nw8lTNkRzBHUkWvGekt6dUjHYMi27zyyGGTZ0
rbakguA4Mwv/bXca0ewNEtzYUsBwhoIPmgvnpTQ9NNiObEPKhw8tUQPwwSEIRpj0KAgNGeJg+SVy
AaVucjAPMC2f8ibzWhPfgQOPDRaQwyEvQqnr20PhfiMLiVevBgVGMyx6r73xuRlnqdjZMv7jhv49
mI3Hovi/gPmWSGjy9cr0hinDaPUe7l5LOkGbDbkjbm27is6GUMqn8YGuWQSGZuLFYW1oWLihTiVu
gfDffq4jspGIf1y3ehFKX+27lU812dzFvUSngHdzhXiOUVsSyw7ZHrJlYWDwN+T/le6wNbMpfSjW
bla+zKee4j4q2qDJArf/BUBVWbduApHVM58J7O13B/Y8Ae+4qPCNO/IekGpQmF+P9Rg9Z8hslbaa
SD/aJeOaihJzS8x8W5AMHJWvJp7n1fW8yxz6JWhhCoRTtJ5SJ8FUZLQj5KeF77aQKavz3hZ3KteU
h64Rn9O3KspEr/Aua6PZ6jlPOH3KnXRjT5tIKqE1fIYZ9rVty6G+Lc01yBD1Xl81tgU92JwG+0uz
1GkGdErIb76N7FVzTB2AXcBkWuq12nM4iN9DzeaB1f2/r7QtyLpjpnzTOhtPPqAaWGIYRz3QPqKt
1rkSFBqx/5qI0/fP+yFclP5BoHS5OPlGZXIYGcACwhcHYqI1AeHgGmtbS0lxn+fpvQ0Cunzvcuza
vC7USr1BJLFjk1LlIw7KNVx4h+sSiK8fnzUREFsqCUsYyEumstnYYCb6UlEXJmeBUzhgbwfLbR04
kQ/uJu2i/ZecXH+ZvbUtU2QTNtyCaLoOydgUz5jCBDZxPhgHh4z2iKVW10GoEbOpY1K4nsfbiT9M
RB95kyWiCBcL/ixfG6atWE3dNCN+twp+qmf4wklp/c1RYkWWeebYFPsyXwIofmFPYa8McWOgmV3c
bPyHxHZnxLRGxtw8XYtPO5oQBAO/nBbpTFzFjr74/0VCjA9NgfOhe6HR6lrBh4/Ro2cSX8qehE/l
5JZsQVDL39EgpZN9NXXeGEpcYwyN8wHm17emQDxWMvzRW1hh+8htqHhpvuaPLPLK8BHFjoEMAEjC
WG12aosgrazpMHkl92eh+K8zeit5/zljdEr2bbQvpfks6L2E/jqQww2oy/oNYQ3xn4T+djfXdCPr
5PGpk/Aj2fHLOrAUPz2RU/XGiVOyPPQeJVs42KMmRLnH7M9wSJgW+oKdQMf9u1Aax2iFcQDEAWZt
bYKKstrwQ5CFPMmc+XkrZlIdXhMerlC59velslvXLEXrJsPFB4IkrnBrulfAxBQtw5jN3bU/guD7
IJqCZTT5OGLsUs8SDNW1WGZT30us9pO8UrFRYqqa4NBrSGO+NpSP/x+dQSGWAi+e+ZWqjagXN4Sv
y+/ZU/3djsu1MDyvUWKTEKsnXsJgNQ/LSAeBLN+4yqI6a/lOdHXi8cNnlxdk3ZGAfymlW9A9HfN9
JUI9oBbbKmICYR6cteWu62goQN9qBHJ9+O4vc7mMkTL5IwJOkDxycSaj1DZFYSZi+3z9aOvQM8SS
eokEyvngCTfuy5/mJ5hI7lXf+A8uDrhvuSllkOZN/+egRg7UJcTQ8Age1XdCNxAfQDHXoWFXypBd
QwPx6MMfkSYWql5VwzEbGNJmIbtgxlf8MAOxAe5A+H2gPGyzfqXEl/6EistwAOM0BnTEjd2s7eY/
Czbt6A2t0CWe8bBSk/5NTX9Yezqfx0k30d/rlkpJEL4BpEhvzzVTYMKdJQEJze/q81Rn5Irso0gG
7INwKQNsKud4x/eL47VF59WyLutolNKg81/anzBrFItdHulxiKU/jN5ADowxqpOIGRMhKPSyzkKA
M0jgeEBcq5gbZYO0hNOHyw8QF/iuRqIrxGEhtVM9/WsNRcrkrimBErp02znu1cGvGSEd7sfJ1h9Y
pKOpo6Ma/detdN9LvHWpDpOJEW50MXA1QDVYDokHxiqVSJ5Ua7LR6VLxfrp/31F3sZbkKhjk4VdM
sR0zpszchmxuspiRVai16h7K7DHxPo9u+D5Gz1jqzLadQWfftR6eZoaiqnshUOHdF5Hyrt2NOAUU
XCAiMQ9SRo8jdERCHybHvk2I8ul9ISpdTeUQjlChyvPZQ8REfpz/xqMtZtjAlBWoYce5FAF7FZ+j
gKizvWth6jNXqkKImG6dHAOzcY7TrClgFXRsIlRIWBrIIUvDDvN9do7O/i+CNRxaoQzsfPbzDMb9
uVEpqyICvEVhuaqr54VCjP8C4yfyxj2I+uA8y+8GbbOqokVYX0C0U0NmjnYDQ3H1nOrBiwa3KiSU
5nPq+dAXDafYdfi54fhtOexY8TYu1UQHU96qvXT7/73yYvum3Qw/G5r3I7BHo2DYE0duRhf55WZE
iFxM6lQZXFAwIAW/lcJOM3ZgzGs5UDjMQWj+TEBu/Tefig4PI3vRUNVa8rjsLctuGlDArBwh1IKe
FlOX8sl2nTz//aS+ZmKd2at4xrBR74NfOHbV7iNYhu3njqU/2WPWTDb3PBIxhzxBP/Egvkc2b6YR
DEV4EIPu6aCPsK6PBKv9I99/UicBNv23juftymQlP7NnS2GxzALx0Q7lkpd8k2bQHrQ/wCZnv0YE
nheiGShhikmH37QpSQrhcraX7yAHk1gXrCFo+CVo48hFHTnx0bKcRrKjp5eKFrzp75Cm2YCf113w
V4j+NHYU0gDf42vJUocpKoOOFrVMzE5ONiPA2Nw9YqKLT6zTV5Q40YVB9HC4EwARpjXewGTEPvWV
q924pM0DW81hIclPvy8HjTpgk4yJQY4sGtmnT/yYkM0ZgifPayEYiCjiV40gH+rArO3PxXtV+/Pg
ZDQL9e70G7ZXtAP54/2zzxJy8dQeMofooYCqpu8WieSefyJQ5wJmHBIuAcO5ccvPdmpBlGBY4dNT
LNyuE7NIHhl24b9Qz82e1Z6BQte8qlOVQOxZFiePzcdF3z81hPZqGd9rNvVuYC+N6JSk4XJHZsYy
6bvooBCZ4sBCtpUJ1rdhhOE3q+Csyt9NOjWdriY6SuqA95e1hxAz6NrAmCxMnG6uCOx0ArMuqDBG
fj8GAy0FBEq285b7XurBIZXrncv56Pupja3xdswCO4WCIBPX99OSfWbQGo4GVAJ1JnT2nOL2Dw5M
lRF1+QHf3LO3C177CnAuIfbqNxzSuQfg75qVMcD3ooleU3Xf/TP/+J/tLhuMBtTjkrZuB1ZRxzqg
g6frWUGDlNEEfJUiREyEA9r6IRA3iO8Je8KXf/ISOaSM4hRe0NhSNLPBV3j7KhMVj4/8Li1I0sXF
rcq5CA8x0cmsr4pCX+cGEMagJkf9cFn6PDw8wNn4zOg9xuPh5jBNFzxJGGIr/0ZJkFLhGWaPHqdc
koisfwuen30kEWMgCH9+NT8a/zCDjKcPdaag5gdvCT23Y5rkNs9xPBVP38uegLFi+FEAlO16EYZs
UPwkca6F0fajjR2FVNB0oYumXbQm5B32f/ZUXsWVpiDfA4/ddKqVC80SQyvA/W+wmN+GqQqb8IiC
YbX4fccuvufPUkFOAWo/ahow51dHSPdx6m7ZE6Wm11HpK3SNDf4J6xk26F9wduWD1PbrGz6QmZgn
dFlWU+z7dDTohjPeRp4FcJQBiBQ0sAOqgffkwcYiVAAVymGIB8dRSNhgDbztGfZVr59fl5+VLMYs
lfa2ulsfVKvO/X0/jOu8KvJr9DjN6hfa9XIlyjIP8Kw3zx2YyOr/GutJ1WYDVAuE1prn382rmb3p
EapHiZidUt1syFpRBnIa1HISfeNbN7kJEpzJSaPHXdL2JK55MXL7UvIHDWAkqvATI6p5tOanEdfS
Fvkgi4IW+79e4sbfTcdo556F6XxyENw+nq7K3SnCUuwthsqsmBHNmYxQRphXGyQapj10ns1xZ+nV
nElznkZLEfBtznzn5RttYKe5GP/Nsoi6pqjddjQdrfGvfo730wKrdNDC5ONTSdW5DsERTafqAKQ6
FrkzaklaMe5WJrTC0MYfCFWl0/+oqBumcXFLz6S3ZUgnh7PMAB7ndLKTufZ0HspnODNlbmy2uO1f
yJcD+LaqesNb9cZssV+LFs3bvg7NZWaI0HjMYCRV2cxlDmxEd3xbrdW9aXOEoh3Dzf0hOVcbFPZh
eMZa14bFCzEE2xPe3FspjU+G7eP8nnFLiB8Xkc0vrb6QDfwWzoXAm+QYeDth1qE/1kgCmZzvMrVz
S/cw/RATEI36ih4xnHCWPhIP4ZsdOrXqbNBftqxiQ+J3qH1p79/wlexfxidAl1nueENabyoqim1o
n3/Xk7F73MWUbldSoGLb86WEjOu5Udyh+W0v0a9uW/sUnhwhCJXvylYQnHdaogE/ySkl9IkZQEzy
28KvRGCc0SgWOLCmzJOcmnd0VJBQ6IFiqWUAfQiuoEbKioXXW3fX+zNyRBljNI6O81GeRzYs3zsA
5oq8oj58lFFdppzd9U65eI3oLu8iuZAIbaSDgUgzuePZ+L94cHbwzqF1k+V399UBS5HCl2KAZIC7
nn3nyoAfxT8BEfJ/VTw8AT6lW29xcQsYpjC0eOMW+FN7b1m1NTWVDvk0zAzXPfteSlXovtoK0Mnh
RZ9ns3wsnJzK3SJ3BGQMAPUVYZUNScN9VMMxNrUX7MSqdA41ChFyAkLcKAnapdzKFv4+01tZ7Kp/
NYOyX9gN6GOuZm2AY1aC2p6Ig8jtP1a9XfLHibLmbsmK7R9GSqoKBj8MeE3P1DoTQT5cqrD12W/Z
UvTWi/hD5Dj1pTs1o4Zuu91RWS2u8b4LWMitiGtLtrugelAp/9hmUom0Rhur2i6BFF6XvWE+cN3n
v5ctCntclO6pLy976Ie7uXnGpHOoT9vATw5Mq7vRcc6aTIbElbABDpYxvzEijf9SQYMOElDODl2a
JjrOaTtE55EE143V/D6G1jGWrlAUo5DaXgSdxJsKK6X31pejaAWAM4Angp84Bk90oVyG7iCcP4T8
niQG+3dQNsocd2nAxuZIEN4LGKBRqBJg4ctu5DgExVOXPUDL576mMnvVFiiOysoPvaxeNolYPCUS
QC8mpMnrS4pdSvIr8xNlOe/oQraHUHPwspzzSOKubfEUQdOWRZYNHfYgMpLlanbU0hxcVIVgATFq
xSFA8BAoHOSY9lFACe2p+FPFkOL9H55ENlQbUSkIMZI2bEXASWAFGTlb73oSXXsdywIv/IeLLDc0
K73W7XSvX7wRB+peKTrlw2TnAWC3wWU5sO0LetThu1ZIyw6Y5SlrVqdEniSdnw5F44oXAGQ5BQg3
juBApgO4JEaKVffnAq88ZAiOHmOlkazroAqHKJZs89dyK9PM8Ae1IjgpU6jXB31Dg0NNxp48bmTX
pWQzE3T+tDRhGGU2BlNfg85gCTNPsGVdjG0mVAzUgaqFZpqbrFT+DsA/H7KFyNk3zZXIXxX9kZKj
440H2YRA9zOiILhWO5RaQouqygx6To1JWxq42uIQa2YCsf2OMvz7excvnlyWd6MQGlR2926eGkEy
2hSQHNlJovLU11y+YripOPthrUtvauvF76QH4KPmjTYVB5xy0W6AwiWkJ7usWtUeXnVw8iFQiQoK
3BVh6ktbl9HYEYN5bBxz10y2tbDL0ng2dcqN1NSSgtKUUN7Kj2fo0UYbt2/PMSsFUXmRaZvLo/l+
vNk0kGJRd+zNzOm7HBL3ogaBs2lMPAGaP1aciloNhIGueH5w4Pa0WmAnOR1I1yS7yeMPx4ExcyL9
FgVBfK6Z3gE0MsW0N+aeb9Ohk5etnbo/vd0okZVsXOGnAMpcLCGLJZ/JCalntt3/pBdu7tNlBL3+
cL/Vbd7woQJWYVT/2bit7p9GrCnBQ7l82QuaZfNxsfi9UfSgoagbRpQKvEGVWfZ6hcMyv6m7brsz
M0OJryeVCxfmaAdH9Wx3E7tYT0BecspFin3HZRMYnmR/yiBWu15lX9pzFKnCepiHG9YyVykX8cop
O44Lg4vJzM1WzgG90UUNihsPuV2CTxWUhpq1e60RIiGOoOzhVaGnh07W1XzMim/Htrd/JFIpvorY
n5opcXm9g8AC7iQ0STlGj7MTYs+JNugaRDvgxPLhfTwZTAEUFbz7PzlP35bC1y35BFJ7a3NfhzeD
AcmUhm5Mmw1oEqdMAmXEu0GeCu8WhM9qiwka/HfF9w19mSzjck7wKrLi7kyK8LbqQkcHvcQe7C8b
8XRcOjyaaUTbqwnLHS8DjryNlEEgyQOeLzVjUeLfRdwWipGcPJgeVqJB0HJtZOCdg5/q6P2ZHin4
d50P72CV5h9/+ubx6wSNOeZOiYH9/kWa0/y+CUhA6T4xj5NJRXoYdB7Xz+rzs9h3LCEKMVt+sZ3F
pioUo+37wPCSX8aGthOQdJfsjbpCNdaRlR4OuR65msTy/AJOWEMBHY02AM6htqXjq2oI3N1Gew4k
s+gfu+CkqIUmHPv5PNx3p7N3I6yOeTpxu5n8xkQc1mpZdqHOl/8NVu6z1Gwejz69kwBmeN+lfRAC
ECjgnCdegm/eobwHmA/ZKsa7h1oeou8U7lPKBG77+dNWPVWUjWo9YDRUzLWF2+a3LE5OWW3h05ra
X86ZjEYwMdV+hMxGsuHo3OCHvrlv84/7P+MqDO8TGJXwIxuPVqOl/HHM63m0MOyuXL/gAZnOkhQ3
qAOrWsMqgmV54XbMLRklHKZn/lHFekkphbfR1QswxXzllzqLiMew9KmMPasHy9dFYkLx0k18tFOv
Z4N7iL5U04g3ZzDH0j4VdT2HqwXR5JslBPj9Bxz6pRocN8Y6eC5X+FXcDaCtGdv9am8rwZZ2WD66
aM1+ahtEv4VoyBW1O1mGnZb6AeQFDFYm9z7z4yqSiGRUKPhFcMl86p0c/Upy1G39KoYW54N/wQnb
rDNo2GlpUHCLQtWuHDT+QhupP9Kw/c0CktM8KeSwj5jd6ZdLHV28L1aAR4nOK1kEfPxCBDA+OVNO
mWx40vjLwkjmLkMLuNqw+Sv/M59jjjr5LX+64lAdAjoa8QL1QyK4lBt4bqYCOBy71FFJTvXt3Wr+
XdoovZgVHv1365b1u0X5158OXf8c6V2nPHnW/Va3WsCJDmz7Dlw2pTGv8bWWY1foGllIWruWbD20
72t7LwAKNTNYjYEyNSsGJM9dmtLiYDEYslYdu8nOU91Jrz6+5Bbck+jBJYtUBMg284uLMG6C6xWz
VepDZRsr3+bqCCpV6oje0shhxt4f6xMP/sSKEqt88UmB0P4uJL+9+wNKMmgGfvUV6xKr8z18GsRq
HxfAFFGClwDMhx28PmhmgA6p6tWZaMP4zMA0jAXMRJwnh3eglyNuLlHhZkRGHXKa6XcI1jaEffjF
a09TF6ZVEqGLKjISxW8VI5yhIz+axe+g7asf2oXnQq6wnMGk6JdsbkJpw5WOuz4jdhK0kBDLcbin
V1dAJVSPLICsgoXbgwrW5PDrkbb46x5Y5cJVM3Or835sYrMkLUKHbaLjZGYb+WdlyIK0Jai5N46U
FKBL86hzwt50vQN8SYVvJuj1zorhwCfvEhMTmNkQ97KSQDW1sMiRi+LejcdyWpuktnLJDF06iY8e
OAgtYwNi4EapwVTyn1K58FMy85szK8KKKdPwuiTD27vONA/RWRycwJVe8HW6CAGFfe2zWFbSE12M
53DjzdlsESBdBnqVj5yd2Kzz28FRfWa0BI1lZv+RnCPcAemXz0wnIY7i+LmPILcnBJpEU1a78Jfa
2Cd930m7Ch7BEB3lZrFzWfv29Xk9SI6qjDVbiMMJQnqaKrZnDPviM4vZUvRVepQO6xo9r9dBIcMq
tpVTMTG3HGRRZ5x1FOCIMO18dxOlWKu0bCYOK9rhCoXV9odEZAwnz3Q2gykQDTHKREJUl+ilOXFA
hRPb7R/yPxnBp7p4wLyDxb/pK51lT603y4nAAtfbGijucFvvV2qK8J1f+6DkGQAyeH4q7ALsrvYP
OnwJ5M/iwvybsiqhJtlRxosfr/+nO55A7Yyw0yoqSqJ3pR3ROVaH4LnNgMiUoodd13evVZRndMpK
O7n3mqpi2D17NkL72/MY+yAsUXi47Nm9MHnvfNduwVTRcg3Ek9CHbcd4qqyjsediCyyqjyhWRfa4
pj40Q3yyjxoWtv2BqyBM86R43TBkC5xMLJj9UvizjdAdnNUr9iLvE8UUN1Z7gevgmv+0hzKc7vlx
+N+h3Bljc0cCpqJDTagW3/I5RKMNJmdKgrC60icva0zJcXZ6PZrIw6kChu6j1UO0gd05hNQSEQts
YZN7x1U1QiEbc9UXqKLURgSnNSRzxtK/tv8ib8wOQNxq4dgW9FplkQCGWorQYEJ5UaZD84ivEgvS
zPHBPEnoJsIu6ddJSQKmR8Pi4m1M9smWxJxEy+K7WihOxNaBGnTAtFe2JpGfcxUWfc0AXCLmX+xA
KoMaG/cUKrr5tcaJ6N5ACO1xzr6tAmTS38shWSH+2OtkFAP4QLTL3ds9NgTsHiyBtIpDKMTQfNfZ
+Q7NCBTTbAeNx3EjHquRboF4sbZi1FFEhsu8xJmsmLFVy81zc2NK66kaMdONZEWfzC9GLB/IjrN5
5KdYOJkTxZ9/9EvfDPZAjkQk1tcoCVxWgmQjjDQV51LxVtFhggYRXK/1PIwP+HAAm12zZvCzahni
d6pozjIDir/zRKMMCqAwV8k+BUMFDKqepvA3XEj48jFcnZ0r8O7+0UpSUIRteJSBt78bPg4GMRXd
hk8j4nTpc68h81lAdhESswgIb/blhIjAjCKQNa4PQNeFg9Q7jkYdra8RCbYnebpccJAnZse0hvg2
kSeAv3mcmoVkQsQEqMDKQ6+cChEQ2CpYkkWNzYxVnDljDulXquCKNjoOnMbT/rT22qODLKCtwCHP
Cr6kQb15xYDjWFSCBPN2PUd7u6tK4NvNb0LIwgHem6frhBRq6/fyvuwkb7YqNP1mqrAC/nw+ZWMJ
xt+0nAosNMBSAzb3bnuXFtzYueVPBgeKgOWQs0RJYh2k9t0ozNHqsYFrWE12SNH1ci/CMy7at5jk
CXvsFhBeSrp7eKL41CyJJu+C1iyslPrg2uPKibk1SoIQFd0zLH1hXmx9/u1NU85mkLa5XbkKWxVv
yQgrgoKjMlJFC8KT0zQAeF7eGMKHEf3H+cMD6VBJvx/CbPsovis8scSaLlbMbE+LIUEoFTpCsy19
YNf3K2Q14m9vKdZXcKqEOjVgUyT9745xeQedlgAojooJ1qCTDqVXK4qcr0l8jVMHn6wkuDDWBH79
A8uD5IE8AX19EE5MxjRNC6CxHuYagwkNBuN5G7s4oju5mZCampY+ZtMf+jcmSLrGK9dMsk4Bh1wf
DU5F6pfLqMjQgFgwKm/foPksO7sl3KsjVp1ZrIchMen6WUPVimZIFSQUMLZ37BaYEcie10CEMvNg
FtIwMpI0gJsx/OLu8bFGFMM8RxkJX7qJlNSyrDST9ehdvUyQbaCRvYP7WBTKMBL+cOCduWFSCrC1
kuU9Bo+8g4SRLAcAOE2W4+QRHdU4quVee5v/HmqQWwWCXch3i6PLl80Zel6kYA4kiRtMydFcBLeg
4S+fNbJnXGb2pOOf/Yk46CFiExNibVutXQu1q3xdhlX9a1Fp6wV2yjOWzDNAI0lkjbPX7qPRS18X
Elcd8Po3gMueGhWQqvA19zb0HUeDRcPgz4rcHThVW29I3Wjejd1iT8B73kbOj3kn3dSbLp/S4Ciq
DpaMgq3TBKIGlnoVpoT0HxaCvYq/o260jantgy/whtLlyCgjB1KDR2rpq9VbGIOJo+62PMu+bujv
UjykBJZWL0ucSKiAPNDP1WVYOg/dbU6KlX+F9VpuKlz+t8K1jrsqxBnFHV9TQRRzvSYfIprmwMZt
rgpv+dLvFQiAe1PpAdl7YQznt88Kkv79m6Fv4D/xudYhmHTjzKG+pIzekLnfsgjEpEqUIZYG5N9W
kU+2hbVJA34SfQXLj9UqVNiIqDSbS38LXeOJRi/k8xibFyU7R8+T8JY72P2BRSCJCEtXzR6Uo1wH
QfWztewwJFYsNdXw23XmudSB4Y8TqWfE15YSP60NjXP84OekYdzmOJYD5cxAiKvdWXmXvQgFduhU
CbTu6AajOgrm04DvapyupbksEU5J/Edw+xvwx2hRVkwksIwLRizwYVuCFFD75Y3ve35qcidL4TzJ
5YUlFWLAH2GJfw0LyFzMLBh0uKIW2YX3kLwxNB8ANb0mdGBDHPhp/yWPSd1j/popWlBV8UAddTXT
8NxrrccW9Z0sygjrL1SZ+odstTwbPe3ug7YH8xTv37PPAiF4AcgNUfnW6Q9Qqu/RyumhOLQCsY0H
QVwRHe8XdUbYJRUHDf3Pe7WLxT/CenRTIKRpzOk+JTTVq4d7zD0+BsbZdhcNW6bQzQVXLdAmKdJP
+O7iU2NhLl6kfLsrNldaeODNjkf5BeRbKcGgI4EOLASJvMuAayCJtaG/TYY3rxWDOeRMjtxa+FJ0
f7/HFDM0Ln0YjQGTFyBTvJ/75m/0qfwHeqmfl+evI/szNoH0c/7Vb0vm8ZfETmnF3I4OjxU0rR3u
S0ABmTW0zinUIeyqaAzgElR9uJ4dE7mhkB7Cg9L6iolItn9wi6hAoIwGaZ4IMOAyHjptEk/Iy8xz
WZEgKYdvRC6AKNXeJL1seSnafIc+DU1Mx47k8sk/6vD6Iifl4v4CAeZXrIyuSuQrYiF9iUyBQRUh
X+rKLVf54X/LHicmin6TB2dSaX+H2pVDQy7HiND4qes30K64U618+k2NlSZWL6Apu4RjvvzZHKYY
jwdZiWXBn2+uFD4EiXifpVeQMfPmABjzEnikA1qtuszuUx7AvoodiDQl/LxgmMq8+g5JQtmMOYuB
0Ds2s6mvRLQMvSbMJV3b4+UizAOoiaNaNOyUG17gR8kn3qPsgPZPVdTD1udXh+bZP5xBUzXDGfNb
ZsBTuNpSCppXTLnv9LhUm1ia2EVa71KNvQiec5PJ1lQOOa2tg1BH7kNaIn3UpGf3vKZoHL8NzB9V
bR4iNOTSWMPcnQzX4iJnhPvikfzYrgAjWZbFisj0cXVfw1AujU+L97SdxbmxsFFgw5oK+vmIytzw
U0WJdwLDuEyMXFlc3q1BANH5kmhSMzVE3/HWd4vHSzaJ4MX8mWBh8j7XKOqkhiRNIQoMNUE21t0o
G3ckW79ggvfd9KIp5Z8pS9V7Cj105DDBxR0f4CFJJLVBFVeXMfCwJVhMMsrjbTnzEP+GLMAqKTVq
1E98I9DPJ9t+ub0U8hFH+bH/sisUTSnDhnwnbu89liVisTOnSaoO8k78UkqvaPi8dWp1ri6Vxd0n
nieldEMZ4YCuPQLjEddPwOy2pGSRSrpN2MHWL6gxeamjD3ph9yte3Fjliqq0j6FS2Xn+n1yQ+C1N
DIH+77FjTf6lA2fVKitZ3VADtU0wLLMji0EjaXQHTAhLzk5Fev9Ma3YymeYEKCQ1tu8uKO61sUJg
pn3v3D862YONHANZfBrmHIT56ojoJx5PY3QI5ixR5dnolSpv4f/06nG8OmnreL7+r2Zi1xM6S56J
uL6FB47GBa9P5bEriuYiCy+5nSCsCvYvq/+M4nvEfR8Y+cpdflFALC/OHiA28OW/W1u9SIJujucT
KFnQq2W2sL8zL/ViGe8dm+AU2NwExacySe/fmUIAvdi0dZWZe9W+l9wa/KiVQogA3JlG2Pw7Ofa4
AKp1yGXyF5v0bcVcFh8KhYPhVdliffXphSoOK/ZaN9ii+GrFeRJuO4OOOXSmigW0vyh35rBMHYdk
ajbN56xn0vsVcbdPbMZffvVAHp7bjm/EY/MoREc9xihv+DU/y06MtwGJu2+PEXAXEkOXKT8Pd/vy
+jGm6CCdezw5U+/iCzgO4kpMp0cWbRH0JcOlgOZXXG+EoFPS/pGFfN9SYXSaC/yLp4npyKxKbysg
NqTGcr/ej6dll2WDz7wrBxLCGuXJKmLWL26G4wo8SHCUc4s8IUdEztcXqFHndaSeSewJIKjzYZ/u
W7NYQPZegBsZb1n2qOn6rBeVDnUiaZk1mmOoGhEBanJkpf42bo0eRA1mB1zJTRePtYIe8DrvrT9n
YJqDBEeZtTNfVh5OMbSu7U3+IW59M/pjNcmjqzVYzrjx/F9B8JoOBs+JN07joUk+o/y9XbZr+lJf
7nXKGWwrWqXXWkVXbU3cHgGRbNP+t9acUYzmRi15inMPgNd+Dxw+bngE+crHDuM+jofAqVsDrRom
sK6xy/T3Ry/pGBMHQqkdY0xcPhXxUwYt9yGap5cqCTk1jsMGwKqu5m1u4qbllUNhVE8DAOOlLmhH
eKRpEU5I2vElx2/2zl/vpzqrvVfar0YDgYB989bpJNiGWuD3OctGX5akw0y1FeBcYr3GdLc3GSXi
2PjgmhWtc/tOkdH9vSU7bW1DdHvggcsb0nknyy+qW2YERkFuZnJZUg8vn3+yXx38DHxJr1mCLsC2
gFNj5IE0iP4TnNIsqB1/d+l3Pax7fCLyVTA5jrk3U6z9Bex/qyJ29a31hi47zB5kE90tHi/qlN56
Gwmvz/3j/UOUk4A8zZ/vr/aLViIAs2MpoYTip5DwDZ6kayFofp+TatkuiaKq5+uMQ5mVW9AY3/sa
s6Wvj8ypRCJCp+nWsFcQluAiwz/x4AywwMPlLgNcs3T41bvuhpktFvVPussE+Goqac3gHMYnPh85
sNw13k4akYxFACdUYSFM+N0hfEa0VQgDAICmz6kUfMY7MR31X064VrFbjTsZc4PCO6JWoEzBCuyO
PUbfaO8m5mpWk4aAhITdhAF+W2VuY+ubKFziR18XFacc8bSLAJDR80fUE5LvUs8FR1VhVaLFnHPX
TBrgCd4jP2bIzg2Id5dTxdB0W/iQobpzfoYRAUgOaW85vIl2eWbXltKRfHsL4LA0JbDFDhNs+wTa
JakfZ5xcjIuHjhljEyba9WNcaPKQZVKn6wb4jLAIm6JToymWbHRcta4+14QntBTTXEGRxVGDlgTa
M/oZat+U6vDln8BMl51EUekpBz1o5m+Um9MAVzl+0B4R+QFc1UOQ9AsdbJmpNWUmq6BYqzNDyTvI
AkIkPIg3ZbL+E8zpFgEMztdGDZL/L9wXGOxu0EPvb2Q24G526itD6TjvhNP4l3U6Zq9dkCNzPb89
1l+Kn53n/YgUaKXde8FnUnPsrbgEzTLjUCIr6ehJJW8fO6rGlnTLJSrIs8RNX0kD0on2CSZROteR
iNuk++SFTWAeirFTJDM4yDn5YAnLQl/1Fsp7Ag5RzsEJqb0Iw5a9pJTyL2ioZ1rIuX/XBGSqsfwf
rU9WOlYKqcIkvQdan71xfFOSq0Jk6i7QmMpvW9sebaVIq2cPmq08DhLRiI0EHfKIIfxZdjH0EJkh
/GMt0CFfB8VYSug2zIR+BJ7Edga1mTL/6dG/meuRzEevPliaHI2Lzf8lHZ+tlINoCfwJhmC1/ewU
gAfujmvZwezjBvXfXPxrwGFZvr0RI8C7NT+QmHi3wZLG/0SklT66jPwihZ9mopC4WcYJeSXIccMH
d/wLpbR4uE+f68VpjUafa13bXc80KQKWp//to21UUKkbMho7NYqNuxAGGEzZUdgDeOL/Yz4c541n
ZXjDEOY0TVfTghUB+ttkZYzGW/5+c8xvt/zQzS5Dof5VRGp94sQu40OiGm8Zjgl/Ugqd+2vrjkxL
vdG65A3VXrADXbkxUsXZG3EgweTetLHP6NW8ayqqn2eLwJmXVMI7tW8u32CKllpkFNseuESIh7/5
0165W/67KCPt3RcRuoAsDyZRhP98YyTTSsIdgGZhTPTYcgVzbwtf+U+WVzKGv42AAl2fj3Z1ADzL
jYkUNiKEgY843ulf090XQDaBjZy7ZcGnH6fklWL+7F/L0qbGO0qmVUKxQL8M61djQi5Sg34Q2X6c
if3Nic8xMhSv5BFHwtpodoak8IMYyEQ373wEP+6aBv9AEvmnAq12ErTtAlAXu80oNMQyAygS3stt
TdcK5Ixjt1IlAGs2H2f3Z7WZ4q/fCwPxBSZFq7JraHJqwyX8BT2b1Z81az30zFgPhBLiOCHbcMBd
mICLpdP5UoLIHrdsX1tof8ZEoF0NHb9q6nuPpJ1VTPrxKyp9Lc3bIohlNhe5S+yI63W0eEd/A/Lu
gHriJwljfZdGjjTVp9q6zCo+YzyhS8wLpgIZShRX/yOxJqs9zn2+zBRNQ8ux76BdScnSpO4l1XxC
IqLH9RMQ52v0E6UC3/VJo+zcCq9ol3vjKZQYA+vtfE5mHbsdnpaNJ3d6EXzoMCOUAN2s7dviatkZ
Rwdr6yXDITFPYSyUv0Cq12Tzly15A1fY1tMonPxA61A5e15REAts9yDIaiGkLoHHHFQkKV3gl1DK
aGoBJ43okV4lMKYKGRr8ma8BjRtp+Z0HEoGyUwUZdA4b6dhCGF0DJB/LUb6pkuo6oB7ZYlC4xCyo
lP0FadJ+o2w1QbAmWJn0m/lckEAeHj1ibjQEKmNV0inlX//okJTGR1UcvmZnhhtaIiHgS2X0PJk0
Ng70C05/VN7X2WiW/CKPYq+bBaYqhQRQXz18y/Kez56hoa+ncxs8GqnnnztfgI0PnBluTTcfChde
fmRg0wBOkG6hCls6pQqfFhr4+vX7aFRMgtGbafEH9LGwRISiSfL00mRyc2/eHTBt/PLTHakqqtiX
pkIrUovKqH5yjAAaGCon3wNKA7it8uciD6mYQRmicxyPhH0tBvWCW0vAcd9LeSGGCo55ncPFa/8C
gFlcmUIRuSJnNJwVMFHgNQd+KKuKZFBahOG1y66EMEDA3H5BULUcLus5VjIK2hjlkFjKbBvxBdDT
CTjFNvia1apZ+ioBpcc58gdFAbUthXNappKF1jTLZaUVb0CEAG9ozy+9vx4a4UHlH03u84vXgZwI
V3Yv07SDOT3FWxrKgm1ckX0D3/8HoaILkwFkTf6SNJQvmr/PGOc1EtP56M7FbcFDu7CTQcBnexB/
hdlJlJkENYLdbHbqkkaB/XDxxBJfgOy77j8T0G80096ktrAcJNclJIFnZH9Z28uHvbtCB6uaz9rW
tlNqx1mKkhankqJGpvn5+QvDj+EeupLRL3fNHmaELKrPm3l/N0X1I4b6bjArOXhKNi2LUBm4PGbB
4ewL7eLR0q3zZ5kKOZAeXKxzw8QG2slAhHIVQVZ0d+GdFEPV0WvK9chSmJF5dZ/gnM1U+40FoVkX
GaJyLhf9+YMbMKbMtU7I6pMm5vOWfhLOsFvETZBWbgB9XusrRUY/FuXCyirjl9hbfd1iaT6HO1nC
UDYyGLtE+bpZweOkE8r2cFSMJVmMK97G9oL2lu5NM8wqPMcm7feaF5fWPpGqduW/76AqUSKTWgaf
YY1d9rFDOW76BJ80v4HGnGDaXbfluLYb49uzvoJVMo/B6oGFW+tm50H2USagDWB+r8d/yA9JrdlL
fNswBaDf7fHpeN9LvcdQCpXBKqRcFT+BTCsikpRaEAXEMWfGNyPuyx2rSU5qjN/YcdPVfDvjvJfX
f86fmsN2VozehjRBsScMrMS3AoA7W2I2UGYZLvM01EBxdp2KLywxVTr3d/9cH2jAq8VS0KDVCLxN
6mX/I8k7IDc3hI06EeVtAa9lGYTOSsDewy86MslPFq/oOgWBTiFK4uZ/fsVjCRkombmx/csk6R5b
GuG1O07WDi75eUH/Jq+VOgfxSSwqWGqXuJddUYuRUPHNJazu96WgRUkKMPlhbi5lczUtFuhSDvAe
J3VlX+UEvNiKqSBeEa6xwvkwYPPCGyBkUthqs54wDE7nhB+d0muBA2sO4d4GR3fitMv4CNieWbEa
maw9DOQ/smsK+SotCWYv34bLk1s9c9HhrPZEAzHDnHXKg0jIJxZ8yTEq9v9dO9S/Tx1wIeEh9+gr
pjYjjFaDuM1OncOwiWQiILxbawppA1theQf1sgtDJ9y+Yyuu5nzWFY9y/Y9fLXfrNNT7l3czrJn1
iyLhNQVoLDx6jOkUuoUH1Q0m4KTP7ZIiS1f/O6ZKIy+3L5Vl9hL+Y5zIZUfIu3ScUcM0IBZ0WCSI
xftYsqjnHVZS9Caxpds59Ivc01J6YJT3F8DJkC2aGMYgU1tAgkPaCzzbpuGSLbC9HSzJ4jzZYPjd
YT0auPS5uI/ZUyQ0nBSV6BOL55+qdz4CrQJygzewiNNhH164xYDZgm3ocygACiEovumjTdjGpXw/
yifNxNsIrLvu/+xeALH/zCYdYTXvVclBUIqR5/bxffIAPqu0PNoqr+XSi804Zt87oNMGQKkwBAdV
tB+QTGx/fB4ssW7UfsazocuEL5KlTxBquvrpQI+c5TzN6CJ9XiEoDAVs+HoRKZYWnVg6SDGRi8zJ
qESJUBUh8pwPWB1f694EttFPQ/BwtQ1ii2DPs/Y/qr6crHF07Va8VYoPErDjCPxcEBkbplgtysbb
szeYF0jMTyTGPXhKPs85YY5fqLx88jmx4WNcgySGxp3C2Oaav6hsnDiYNoF5Shb+9uXmB5pY8xYf
ErZR5mkFzLjgUVPR3r4oPRxR12K3s1rMtMZUJEUme9SX8tF4A6OcDXdHj78x5X1il7oxSVSZvtwI
dSZfdntVubJyLsuSgC8gujs50bnLtD671++VAVjF6MMdwyNqukdz3TWo78zwQLgv3UgvEVeiK1Xt
2iAFZU1l2VisXqKDc8Va6Kbp9bov7VLO/InBBXCI0GdiFysBEvN0YH39uA0kV4ohCL4VAuj92dEv
IG56HC468GSAvi5D7LrY5qWdH8YLT0UVx1GiGK9G1v/bDyZs0HOWDbDSgsXJ+BiLj8sopCsM08Z7
FRUtZxNjbI8PAQY4aJlukI4dMozjon4LlFRckGVoLJnWxm6CAac5d4LRRJr6cvk2CBqqBr4Z9x89
RllsG34rLqXnad5yXOikft8z/FOvGn80fDCJlA9+BEpBySawp2CFfclWc/B4pysuTvGihFWGONPw
ug/ZneqvZNWGm9qWcQoOgP4bhglw2hTa3aUvhErmFFxMAps3PvGg6JCRq+TQaSq0m4LfER3QOVTN
gL76jZV3R6ppHRlSBP0Og87DvpfI+i7/3Girbpv+LjKJpKXEwxPmAXb45UND0hYee0/T7DHhBwGj
JrG/aJo1EFEaRUomC6IE1uz0zw4VAvNBXm+7sU9a7MyvxukJgipzvr6Hm/yu2SpKHwx7c3Onkrjb
R4J9CynpeHryFRuwGn7OU/BNXuQfuVm1KtWcm2aNYipS4DW3VK6mZT4Rk5ujplOBOsLie5gU9UI6
PELxVhy1noCI6y7DEHKUMaaEHbM5nrArp25Xj3eedqLppJb61mdZ09SK8l+mv8soHytxqaxPBbmf
mQdMbzwXbtpQGS6B0vVAGzBBIpfYjIUVDNcBzctdpdueRnssCumB2OQtL5jjDWq7+RySGwLarTbq
d5b+FgtQ71pS8rpFddvpj8PZREUYUKTe+U7qfx/oRc2h/jX7BXmmOTdFHKV8N4FCMDT7iPQd6OEy
tV/Ze68Tkd4/XLoRJ/2BNWJKIm4lxkI8+t8XEAWCbgwn5HMk3w/aJa9ZEXUnGPAfZ8fp75KpLziL
PYsElk+mbJ8VtGhoENWs/BFVZ2Lek3C0tcjUEXtuuBNFRZeosS2QUUCRTMdboBKkMGu05kmlAdSI
Y4W2ewK+HdpwfnRvTsXFn+W+WcYirQTcW2Lk6+sH5t5N15Y8vGdvrHMKfOz+dPh6d/V2/mKUNLIq
aKmgY7+yPiS5UEbQSVjhHFd/30Gc8EiCZaHYzt84bxfPw/FM9O3FGzGyXtyt57RDBxMMsBAvU14h
RwmzmFGNH6Mrgg7VvYGuacO11wkIJrR5H1i/UnPGHC27Egk4SMD/x1ynGrJfTFjiF8Qdw3v/AOKQ
emhrQdOL5k2sZXVg8GVwJY9vRk6mIGTx+UZ3UOuPVwEkV+J5aY1jYjJW47Xy565Ma9wZL+fjCq/G
SdYeYfNR4E8IoSbN9fudEA72O+HH0ETwZIbSPNRKdIk4ypxcFk//6nO2tAPhxkRX8t9SZOISgmAp
MO1CJSA64rZbAYOinU56pj6YsMD6OZKsKHQIlLexP51Vj0bGzOAvdxEKd6zsuYWwkAFw3/XRYnd+
3Orm9N3/mGPSNcKucWhIQmJihF+iIz2ZcA5kccMOJKhD1tMvNMOgbZnd1akT17ZFepXx39VZ13xU
azJ/H0od/7H7sAttZCJeb2iy0ALv4IKeC56RTgHt0V3pwnQfQfAdYEptPHjxUFq+MxVlpJGgH2iR
/88GcO+URx0m1SIyfr1OSao+C38x0VXtAet5UkSdjrcvj0fOG1sQy9N0ibNF5CgCHmXD8dfOKZgI
ROG5SnerQTdGFoMSdcpqV7QsE5lKVDYZ/GnPbsgXfXZSXfAod7zsdWpS40IAGPoOyoFyGBCuNDph
tZ+i35KSw7pGlFi/vOrsEK351TGvKOag2KiPVa8EfjUOR6gyNc7v6LZqjMZ5zhPEB5WyT8oxqTC4
+9UbGxxScGsxoBndC66kIt6ExAoBxwJjHfRseGwsBh10tUxcE9n7S0tlLhGakK8hofujEJISRrsn
Ssg4hZ5r3RCUSiCOs+M9PNjRF98zYJZbCvpAcQIZxif+YqRXW9Il1BotyxuNPz9Kh7uN9nq+Ze90
Nr2GtLGpxAzbFJSPwE2sTzB3LW0rqhUZ9rQ54IhX9Olpsk9z8LrQejbNj5nZBeN3tTQmumLyKyUq
CQKqKYXMPj0e8da8GUx1nG0p54vmfBH6g2LbCuQM4z7lYwNso1KZvQTV+wOykuXgjWiqpXSvtbi6
i2TuTkJdd+L2ua6rjQJumg3vU7xNIyGx7GhQ0v7lON74y9tM9UTrKPLsnuJVX4+TclvnukkVVJvP
nkPTlj0zUbwCYWhsnB+d90hgBsJdd+twCLbb8bnUQXv4vwiRDq8044YKmAuAs6wOPgNZBlqVsHa/
JC6QjKTdKOawWZjBfUkXX3jpSydOPKXlTpsnA+5ogyqxoOIvOKdVXKjNgy5D2Td2v6il5fcrb3Qm
i6gpfqqFXxhBHdXO4hnj3+CZjCo0vX2uQ8VtHNMbZ+ZhXr5b3q09BGllH87iu3U0FKK3QkeolC1n
LZiwjSq42ofZX6GyJ6z1LB2o8/0r7FlAzj1bsLsbr7m6Xg0C4CJsNrjqyoB2YlNjMWvt97e7EyyZ
sWLzWJLTh5a1s7GAq/vB3I45UCYRNHLouAXh3EK0bIgjQqE+LNpLRrdgO2gt9wyz727RFuAYTXjB
vuJ9ql08MCFa8a+bNnIu7luSJlWUJvTvGP/eBALiwg8HTN+sT1Zww6bvHRrz6UDR+NeBV+zQ46ys
4TyudFgMC1CQP/wnGb0eAWjZZyjRC3pMR1Lz3dwmF3MbjXmyZLyyfXKvGbCNn1xo9e4yu3jVbKah
A7mJ3/9UeoXpkojPEi70gpd0PqZQEGe0Fr1D/XtnIGG6WOLeTBtlcP1WUktr0Q3+GBzdN/86M4jk
XdGaF5nAd2zzgzrwgfMLL0/bg7c98jkdP1axsDDfXamzpTchTULmz4gkhDHHw3tPUENfcD7qvGIe
jkpqHY4xKlSwtjm7CpR44q6i/oqWQsS9UBkGJ1Qk+mVXDtrruBIJy5BQRFR84j8RPx+fC/1GbcQ7
Yvj20KinwaXfGxS2rzmbYNpH1UdfW1q4TizxRE7+zEouozGmYvroS5ORU+qq6OktkfUyLKvROx0b
mQ0vlDEl8aStERSsmdwwDTrX0tY3u2ixXdrLkQ4lBd179bMvN+SIKnlg/2GyWlG+2uuk+9TE19pC
DyAz2s/thwqkAFfg7NLB7fuOcz2Wxsctlu1gfsqWM2eyoIKFS7edBK+reUSrJDY62G2vBvCeFfx+
PLLvzngSpcAwx7tfF8U5sysxskab9PX+HTl2NM63D5U7LWomq3VGdCnf5UglU5+b86molP8GjgvM
xO1qpfP6GJLD+ovBEIOegWlNNw9L3oH4bK+6Z9F4cKTsi4O40FXFBHCE46VOUjxQM6BWlIeRev6P
ciB0Lk0o27pFtOlI7ZJVoQeO7vj8AmA0p2nLlFkpvTO0EYMYbh+trZRX2RhYpYx+U2oMAPti/f2P
8n6Av2WHHQ0jH4sbyvP6XQ6P4/NaWvWggZoOnSOvGKA5C0qsSdOvJbxiKa0UwdXgGi2cq/rSicom
EWapwqsJPQ6yMLvUQ24aiGE10Ml3zsumL/foiQczWPmKUShHcepg19Iza4Um1MNqMyUwfddO8i5v
ja8mZJO4UylzoWU5vX2GqOoRLie4val/GIkBfCVZRQg/7RoC0E5XfAkM2iwl0FfzJgIovH/90nmE
/WT3bmEiszr+IEQqlDV6Q4VSfvQ+LQYKkLRIeoMI3hivFHzxGVpiVHD1/LGYtsn2JkKleKf42C5D
8UWs0Sy8oo6IeRLYcGy1mnXYUs1iYg2IK6V3xrHbeaHQXd6Fw7nXRgiOIUkN9OUnA93MTBJREgIv
3amVDcWI093RYbmUXVIZ8Dhj0/hyuOssDO4i+VQ3JDtJZFY7V7hmcR5sR5nRiEB9IriSem2IZaeC
NuU3Akl1hAzmuF9ogy5rXzNF5ZTuirQpQFOJ89WpuPSVMGZdAJ08wbTJalcf6FQ1HJXR80PHDIbK
1NCZf/B+3M0zrx29vzIft40M+iFw381x5h6WTWCA9uROOMO08FmkYekZX2YPsCUu3iwucG0qrMV/
M0yY74ch4z8UnJd3Ig7IEK2YJ5q6DNlIHQ6jPql561Q/6F4PGjjrbYvYY7xhwxeISan661q6kD6J
qS8ycODOGu3SdDbBPXfUgB1lbv7AV2/eO++Q8NPLqKd3Fz5IFtHcDR7JahpHo/WbekPqC9sDNqiK
q6xYMQ2SKVmqAgo9M0ar/XOOiaSlxumpvJRE16+pEucviqjHxFROLtnhaS1OkZF/ing18C9GO8B9
xmU1ZmpOeZZ44224qiPmhdqnHwr++G6SIcwsTHqLkUUZSsf5mIrjGS48XxLk7/fNsD1l2HRASl6s
RhotWb3Gv6AuaaE99FByM44XXL5zGdIkmsXh1tMMjMg5bh72SuMA7dghlL2iuPFre7H1Q8nUbaTl
4Y2V2gXz9rJ7QjitElUy7jlHstjx1bHoz5nVIwWPwwQ9431g7MXe7tPL6czcBg5zvbaaoj4FaGhx
2zygt9Ha+y+9cQie/0LRqFv9kyt8YDIp3+A54pkFPXtcc6NaORgkdyyUcEzDcBGQJ0pAne4PkQd2
ILTo1AX6MDfTJIL8cNPrY9VmueRN9C1TlvIXK5RuitHmf3Z44N6Bs3XEF4hga/nHkc1Uy8ajMZ0V
Q70wzJT+pnv/8n1g/sSsP3sDUmiW23YB6DsdsAykIe8ndd21fJZuzkeIRT3IJ46DQDRdnWy4z3Oj
ljK91yGARY1tgkg4woEIufu5AtnjNi1VsXqLg7XMt4Os7L3zC3Cw+gs9MidypL5h62pBlNen+MaI
YOwVnFAZ+xEAKlxp963GU7FtRvi32966ye/ozGTE+4p5J+mSgZzxO+FHuMbA1a4gMjCszZ/cmxpI
C48dceF9oOGAYBmKj60Lqv0JyIbkcm36sV1mioOXG1SIiRNr3/uU/SsIlqL/vEjQZJckpwnke9TW
6jC3sJdcqt7iiYxIQzXYAtag3yNo/2Mbng4rfwOW72E5KGIb7dPsJT1PHouqmanpuExvlfXGJV7t
SneAVXkYiBdN3rEXTGzHDif1yIiQu/TisebhJkgCZN26s7D0tjv9oTF6eGnqh55TnDKuRvvXq4rH
gHGL7NgWrHtDtzD1yaxK2v2Sk4rYCdNXlrXQJKmaF37PEy79shyh1QqQMZyQYWmgpJAInRf7Cb0h
A+FaTlMm0t6S7uzc4mYyB1XLYB+B3rRzTrBUB4f5M2ewMoX6m2mv1aJs
`protect end_protected
