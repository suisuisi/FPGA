`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iO2Bdkfy0dqqValMR4KhTWXpD0gDQF+kyoly3tZBTZTVs0CbWJ4Owhu4jxMCf8X2gbWR6iweF6Ks
B5dmLHZTDA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dbcEbgyZfx3YLmYpvjegvD9sRQCV1qBv0GqFBvCakC3SMR/H82zqo5uv5MZldBGUVmNHnxF3Vejx
zSqxUKfTNc90CS6quuoQe0eeq3T5XSdgwbNtjPZKvJuJTmQKT96yB3CfQOz13fGjaLrn/8NBUBBh
I7OEoGGg7ADph9V3vRg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bD3a4YgAnaoJx9/hljj2C1rODcUhawTVE1gtdPkNj8/YjemaFM6/sF7Q0CXbDJ7a+OBrB5pUgj3O
Vesi4yVmFp+mGmFarftWat5KmZiP3RVWrXwdzMj+f8T7p+lE3iD4njqUxIUz0TsUaNvFeW0xVNNb
OwTEX04nyt5HrU82dltJCclpFxE6yrP9YvI7l328bphwnC63xxk8T3yXwCrvj3VrIYuDT2yMRxrB
TBCv/Fe2f07JQyV73J7+DGAeJG0B1dTHeu48auQT63g1HsYaUXREihEUKgZe70QlOqlPbrr6Quhx
2LXE8LSdCA+FbJ7LlQc/Sgasj3ZYjM5lhEKleQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GCfR7acMSeEtOw1DhZKkUXjh9Uw/vUar7CGDRG9rZcB9NFDtQTltJeuKjFg8eaeKH9HFBMryuX72
/tmzhtFaiSTjr2na4ncL2XV3QRXe7nQaiHdc7cKBcZDvdSSMzOSYcIxLunwLwQTLC7sCvINmlxO1
NXnYzJVL1xb9HP8QVnSYpo1p+gCXcRBZzrOjZjCUnl7F2t3ZZStSGjBEyXVLnV+ouU3+247oJAOa
kC7v+pOtG2ho4KclIg0MGijjPs+jyOFU+b5C+ufQp/zL9GiZ5waCjb/0Y1vkBc9jZKR7YRnv+ASG
ju1uP8oqEXR9742kXRnW4HkMKkCK1MLDgWYdqw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L+AGKmFZ1zoRJFd2cA+zxJhkgQ1R0aEjGQCGRFLNNhLHZXpzGDIjdSLjralBVRJ2rD6UcJutapF5
YaMoV9kphGGG2B07dxBuIimVjOxS3ZQJ7ru59ddfGBxUe9EHrv00Q5hTwoxig0lxqnmjSSnfsDeF
weTIqNnXkG5kqqezKC8a2FvUD5QWQBibhK69OAdmhhIOwZmpfvQKbEKgLX70BzcNlmLnttRL7G+q
XZ3fabZ42+JJHDLiIfveB3Gp2Lf2tzTH1u2xx5aEUr9154pnC9PWIwL3y3VBAT1oHR7ScdoGDOEy
HoYUiDibldOidIeKW0KrTeAIuBNmtM4R0R+RSA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V5ClnklUs5Wo++EDemG/KeowZlAfqB8SUrvSxPQGrdIwGfUvoCajhuABAWdS/L/pQl7Eyz51aiuw
KzPMrWtQozAEITf1xzvzgKbWZqoi4PQD3rThywFsFq60u8DdvHYM/kEvit0cZVFvG8rAbtlseHLu
0vU1kbrNgxb3bxjOovg=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cRqAgScIUeXUwYGfCC0XDtpcc+mFNm3p8oTcFdtIU1nnlMagpBMqRm5ELc+m/Yw8jBwvcvt4tUFv
u/ypEEw+y12B+5Pr6SmnLJ+NVB3Q3Eyh4Q/d7p3jReIIsUxrlENpCTi4PVXMKr1B1Htzm8F8mXDq
y2UV+0SC+4yrBIntsdS0S8jPBERhfJhzNC5z38pPHANtM4wGGIUuKxIALLz1aq+2AjLbEgFHNrzw
2bJiDwRSTwrY4Yx2MSzYJk3O+cQBUe8nJDPx+aGEvDzQ4ZdJMNg2z+iaiE7OTaqK492Jb/1jvU0j
wlI+n35s2rrnc9QgfljdOJuueruPuYDi5vTTxA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296032)
`protect data_block
31mVfBe/eZtrisFXB2TA7ana2RabY3xubPqZRC5bxb9nG1czggFwWkspMm3jQ6vY9nt783sTWC1S
WTPG4Coq7KHxzEblyd02PpsYdxGsGYTiwzPP8SaedJau+IFc2PV5dX9mafMorlLNHdewvFHa8bLp
B1uaX8P/W6tAyAVkIWKzTTaEDQch1jswObiorCrRN8kaoQ/huHBpwB76PBCFqZCwEjj0lJBf4B76
pqlXRw3tN3NCxvx8qi93/flBmyRFSe39vgjaXpkJvPMAFc19siR0l5R17mX57NwpC/IqnPUubT1r
EoxEz2w7C9eiBylWYFP6OBtChHOiwUPPfePefsTW4m4rR+izXE2MK8RiRq8ZOMd17jMp7rDJ5Hzq
LtPevR2pquZERgH8xiVNoKa/1WzauFnrehfFztfeyqUPvwIE+7PIYMZcoovebeIKJYk4nD/wZDM7
DB85NqhG5zL7Bwh8QNn3u+nZmm3jiz7dACPXKumdHuB3wwJHTCQnje0cBCm4326EEqJrDXGxDwtk
RNTGHOx2/X4Il4N7VhuE58WKgcIiyXcy0PAVM8c/Esf11DGhhog35zbTGp8koWD/q36dj4stp3Kc
KvwJ6SQvYvDo9XG5a9NBE4kFMNJDwwl5kRmLyVPFQZZMaq74/FDkAS5cRGWh000tvLRWPyf7WeOg
SfXVQbSOCotXHrY7rEHu7f6pqYT57f8tMNk6Lr106jD6zrtrX+eJ85/fkFnrEXyX2SuUBQEOmGpT
hZX5L//0siSQYLXwQKZCzwAxeBNUqnjh8VvAat7K4z+b3DrLTDKuVpG8gjVx81/gDfetR+dncK3Y
80iosZScnYFt7OFBpVwpvlq/kf95xWOFetyRlgGaUwYrygP45PG2QEz+4/qFOGby4iz/EGlgqn0s
FBswqapGY3Sxpz7UDjzy8l653rGFjCYjdbwNw4zied2/Z0TcT0AZV21iflEUBDeGABMCr3XbubBJ
r6qgBLUV0dONToEqY4Bh9EWZhxLGVoTjWKsgedbkhGtETgjuEM9T5KG+44GjPyOkG+znlQsQgS17
+5XbNsp8zVl8n5zvcnLmsUYtSyMF06O/rqYCChGLJfAVkqwGOnyxXNELnntx7nTXXy21JV26HOOY
JX4be00i467H5fh3+aEec6LRPYy95KjFQtDuPcx6w3iCNYBBz+j6Hi5Blul4X9+IgsqIqKD6xMMh
mVpxFic3Va7kMQbiNOif7wqhxjUBYHIPTMlZchwiGA6Hej8oNAFPRdLMo1OOtGtGRDO9Exjhmw5i
xwst4JROrK9sMTN6+t+7e7ziQgPCnrHlVWQHmxHVnffeUTILzFiyxu1G8WCNC3afFxqK3N56IjvU
p7OzcP9vhtO4vp2PpB5aIx21e5hX0f3UM6AF+RZe8/ORBSPKpsrwnzoHWC4sbYN9UHVqD0fOnCRx
STKtxdvnRzpPci5ORPjeEOk5h0p6WRwxp6YivNaRys9R2Dj2i7J3lyX5nklZ4RSNkIkqtyJok1Oz
SplIUgX+2LDo2b4kzCjdepW/s72yn8kobaHHVW+prz40Vq7XmVw9lYmSn4leaxuTAyS0zM0e0Fgh
xEXzfIQqJX85XaFDod0bdhqn5R8ooPNBubmjWAMrfVbAuxaXI9B//1CqU3t+HA0pX/5cYezFSyJy
/r+Ya+FojZ0/XjIRN1d7H74bcsSwe30+kgz39ubbl1BUt+zqE83ZeT/tnL/WSHuTUgEPt3MAdcbR
cCs3/rYFbOxqhYnV40HM7KotLI3wYzjQYiV7OfQZJp/YC/1xWVVUU223NL2prN02c3DrxwGCtx4K
QRVq4vS0N4cB5ZUq/ZLdLg9gTkrWQLiwUbE2hjetxO4nnJUtB4nTaO+19KVknxP6xx/NKFnaqgj5
6xcPtROMksrMzJi2OCBw4VWGamwYmhLJFVXtJ909I7Yur01xCi1/vL03cbpOHYUMcV4IOBQDTiBq
9FvH5sxWvDVn9CrtoiOiR/CYPUj//cvP/Zj/Ej5QoxwhXuajw8pp2KklfNleNs8kGII+Lv/dQ9cx
bdnYOAvqWerFZCPYK0tCH1f1Y3B8OMgHEvwBsZghcPLhsuSOHQiBokTLlUr71fopgGyMx3kHTQ5e
jHVSgauVuz7t4HgXWEVF34kaGZfTWAyXTot3us/XFA+gayJnNMDqaRoWk3jd/gzLZYl7Hyk6XXhl
g0/bsZt4Nu8E7ntfJtIm5W2sgdxPyMVIg+1fL0As+xBGJLvULhRVFhRTaInHSz3BZoKDHU9LMcxm
lTlhgTaL4lciZ/DB0MmA7mrccxdK5jQHJaO7MbWTETPjDuigLehFmsMGwSdgyDPzwn0tuPdUJYBN
1aaSC5/IUjg+i6vgU9ACRu3+I2QpvORclu30MB9rfrJZ9EFFEmfsAjz5Uv9YyRl5REC8j5N6a6WP
zDoWkLOzLjS2K07lIkWwRXA85j8lkV2gz9tUfzRj87BA2I5UoldyNv6iDUiGEGZooY2Gs8bi+9d1
ZXTjll7E6LugrwEQ6LqoNmTs1VKYuefWq1R5hLUjPc1mRYm+lA2gIt3xRcQ78vNvS2jzPV0qC7IM
9b0QEjw1ZA2QLxoDWwNBYCGwGsj+Vbj9FMZx5Qshsk4lDdken7m0sVvSYy6ErdXRZDjSfQTuQkj0
GChuIlpWC35C/mH9/ew4E2bLUCX6zCHhN1ohyFRaqAtEsbMOd7GGuTZmMhfRxGOK/tdH3X9ymnm0
/Q2tka8gtybzGjouFOI8OZahlLNIyp56FuNDtDkigMfyC3Unrt4JPT3rhVcMc0vWb/r+79pR7DW2
sZDmQ6JJk8IUny2KQRtVJTvLNrRxTlFoh1K2tHrfrQxQv7oyZ5is0NppFWIRu56WRff6H7z8U4qZ
/xQI2jix7itnlCz8GjzIVKHxfED0zYnyKsOajuBEev5tIZtnRwj/1AlmW1/TWZs+UwYNSliQcnrx
Ko3kdc5NRyjgQiMBuywhyXVZtjjrU9+BlpkBoGXHGSzF0kQS1PsNZXcyuGXAVbCnakOt2ZNEWUKJ
xz3rrJGxcBoyxuMRonK5+QZFmN+7wwItqk3X6PvbeJC9DYf1/TEk5hho9/GFRLniGZUObN7FGjPB
84GHfFOR/G7n5KNNoIM102kUmzE/AmQZ0Dbfc/3rMBss9oy1lG1yHCzeicrcCOmRZzpdfPOK3zSx
TvWWaDGhC5vH5Px2f8LlDcHxBnP8smA6dZNnYPmVJTYrYdmqBV5Xupuvh8GqokJVjjZYkCM8AWeM
6bi2ichIXDmZsBe1xiz4uo0f3rMQRWL5MEwloyIAyDQs2E48uv8PIuNqzSwdtutaE6IkdFubE2ui
UTJUvi7z30W23omWYQXAX8BYvunQIrQekZNjzkIR+yl94NNTy8UFdrnQG8+vuVwUUD6qMKbiCrdF
/gWkoVJ+CrKvE6Qm8px9EPV1RoOQKtvsJL/YayhVjVKwTwSgWe91U82V+f0/MHakySG9KTxfVFrq
MjQmSW8jsZQ+MHk6USUDF5VRsToEf2w6rqPT+Ga++G9icMAXxzzKTnx3CBTi3RmjIM0xp6CK2vnY
vo0ZDmrju8+K8aE5we/qfDcIu7273ZAs4jviYRoCtUVgxCuwSqovrXlkorsO51IvX1+/SD8hq/tf
B2jQrvOTZCPp4KRBS8C2uaKr9zd9kFLp24TO6mDKANK8OvlXavySjabtK1RJjmYzCM7D/yr7Tnmd
Ze1eZ0WiKe/PWNUw6/WV/SsUn3hWBCgf8bCqFsysecRYVE9O3wVGLBtnMFcEoByIbxiB7F1fRcCI
dIU+xbD6GrOF1507CW45yTH3tbD8RFpuSLlrqHlY+p1oFBgyCIDcI8wjCuU9Y3QsulBw3XQ9mfgM
Dnf01Z0lPqSP1npaxaq3M7k9nPrcqfX/VUxZE3uYB7TF8SDBqwv4/FYhAvafL5VnYJBI4IwCOGJt
qRZEpIumWDD1q+Z0NGq0Nj0XwtHJFH+Xmwfh18pSOYixFOTnvkABGCGPptATJ99yh6WYytQjED9E
YW9w7UNlUOrE6znwdV3qCDrc1NOcfEZfHoBmJWdIbb0bIST9wtYEHtf4xeFy88bL1qtxdVxgJSgu
cmZSvv0Z/+QvflUvQulvuN8KwvIbp7hn0xday3bG5uyTDg0BQtjYLg5yGq/hJ2iyzR3WsBvd8dzo
ylfUnLxTW08YrqYrEOHI6HDjLz2L5pQCq5s4f4gwBGF+RxydzocKlmdHZPlBhG8gE4fAxKzUDPQj
yx2McD2LwdPTME5XRPCS8Pfz+2cdL5cBqG976TRWASiHhZdtaguoOJVeIABM9s9hZFEx7cTEI+/0
pKdgVX6Rvkjg2XyaGhXHPenNa/tPRQu82It//uxgsOn11r3Q5Rt0FVSfq9aFfrsw2mWR1zhddYMJ
nVQdxDpqBXp0ODLAuIMYOGNz4DGqvyadqiIq/kdWOvfw+sn4WKgIFp4G8DtUG6y+QrkT8avflhZP
bmLx38R3Y/8qX42jSpCyrWKJTR1+hh+oPG9ykvZrTnqwO+me5f39j4AkjgbLJgZ1oGe1QoJSDVOS
gp9gJaTkwSgrtLwKAt2Ycsm6WEX0H1Fbnnznyh7fr/vkDyODh7HEVQIaHJ+PLLNGG9/C/WPiT8JO
vbcRKZpAnN2NcpWuQ15s8aGiO45E+NM7MXxO1wieti+tkhwG/ScXf+8ZwDtr13Qc+UM3JwloJ+ks
t4MNScC5s6+Y4i6zz7vy+dYvpfv08YzxVBt0Wgh6pWnz/v6pAmUvwaDYgdUFePklqpFvP8o8C8qA
CQZKuH280afeG34NuzFYxs/bKAkB9WiggPDPlt2Y80/SQUtNK4tmcfADAclVG2CbBNUYw/SfgYJx
vh0JnhYM5ItuKPrk0HXGuIHPE/fzQ24EjJdfzqxEOjej05buAI+qBR8ONyBAIQySKEoXuTaLUdl1
EvLE85NsRPKDyMxPbF2mapzm/l1bwLtURJfWmM/GJxda/05oQ+VNTq3NKZNZLutcr/Sm51W4Wp8S
NX+5X3lpcQOdVGx/sm2d/FcM0/YRKbSBmusGoL0rVcI4JemCLqYRT5Xr2vDuuDTbLAozn70xgk5M
L34wN4CAfJmqPN978rNqDVmbp4lG9soXI7i6Eaqn1rCNSt71qsUC8lpHsVasRTrgdf0lBZDdu838
w86/1nowpSe6sQhYQC8kiWj+3aqDxakCroexafk22WvA2ATMZ9job8krs4INrB2DJUiq2iDztiro
xtP0h5y5HsJouJiGwCfTdLWOoJipmq/lq0LzLXHGKtdjnR1B5oU/9dMMhxUL2O098stH/mYBLnAn
OyNQhFKu2DcVfbZlN5H+at6UL55jHVvxRz/5CiEy+3VGvdgShOM0F5Vqyaw9C6dotLq6Kx6Ek+oj
+Hce/gRoert1mqTNIctRnnvCEUNqPIz76qPPOX5XP05QowGesDcD3kjlpts03izmPtxHLpPItIA0
/hVbaCpTPeSyXyn/SvenOeWRe1J3JWbrnXotlrGg1CTbFtOTw+FBaF+1S8Nz/HTnXId4QzhmBQtz
sWKQEDK+XOgDC6/gohgiqp4AxD7OS8/S1WRevwmsvgABxb5zp2DHKccxQ51l1lyQBBCG0RV+9/e4
u0PomWZmq7jIn/RW2DWhtH1d14NvvYAN3M1J7TtfdLTAgDGpXIaZexXCVVd9BFlHBGeM6rM0t64L
9R931adQ/bBwiDulGngIUr/YQjlne2wXiw/Wcr8ZD2d8x/zGEO3aSUqWWkJ12LNbFvQBUJHuSACu
B3VV0IYpVuWH0wk9Yn0syY7j5LoP+IPY7dx2Zgx4qNhTjy1NnwC3cxNQVgFfKxnCWygxNb7ywKca
vGAf+1QQLC9GA/Opb6t+o6rh+vZBHqDw9NTCdOB5DOan9Jrw3P7cNFjhEgDTuYgjzwpu7B9bZMLN
7Eg5o6ZGRyky1rhBOgLiGKMuayDEFOkprEYxxbxQns+7QL/JqAiok1ViU9NqpStGk0tcSXJTyfBe
1dE8CENeDYO4SFe4uSiRTRHGk0Vhki8o8sxkGhTqQauPCHBwn6f1fAwVnBNIP4mTEYneCWBQfFJ4
JYZaWIpY1MjtwplM+Hpr1Zpd/I1YGJpr/6R/DULx4Nv1yBXzrf0OL+3Sx+G1NcQsLCR1KJhD5/I+
yBu3Vy/zam+1dYw8SglsA4GFcya2gHsI+1ye6cBwBLROmZgpTr9UkFknEkI4hfH3vl6FFxZ5ggqz
OsEUQx0it18TVHUj+vJfYYy7TE/ztBrxoj1lijW5tfxoNb4flVBOz6TA0e2lfmWr47645VV2R4DZ
Biq7DbePVVKVjwwadW0aHjv2aDTpeWsUV83MX3ArNwpe8d7pFuZt6oO6LHBEYxvlVTNu/yonaRBX
lCRG30R/aGZRRL00KUP6Fv8luEYKJIByIEeaWMkVGY5uCSy9FMsaJJ2tncQ2RFDR6i7OHLpHk7Ix
IFsQCBn+Nrl19M3GLbAnD89K8Qm4K9py4r6HVtzhRP+c/BawHJ6nU/rXTtC1ggYtDeTXUnzPCxZE
jU2kkUO+voyGRuktfaNrk5oXK3loLOS/c4q82hHbAUEtCNBp9GVuiZEijHHE01nxhwsbk2a5L9JK
2+G4sCsif/cmHA+bNH/5IdODkZPOCgvwL1C3BVxObNIVxhVcVXDH54NCqAY6USsb8jYy/VWwsodk
J1mjMybTOELnOD2TMnDvk8rmL3ZKaXQqACdsP7/xowkpKqohN0FUZQKpcZQ5bOAyWKx0tXpAAP1D
HICFtX4igQGLdtsijl+fuEWQwxY9mUWugXNvVIs0/r0h5V7VP5BHDIezj1AvM5LJVmju4OE78nRP
yhLZkV/f1yddBOHOqAaSm87KRBkdGOwQt4BfnDrkhYKGFErR5UvLYseQgfv8kxjEAbALhz2r0YeB
3VFAfccV4s55F/LsqBQ/jr9CvfyQ6PpQ6eODWJI+/aa5dcbrHaWuLrInqB0qXLRoBxbg8OKLumy/
uweDnr8wZepdek8bmDa5yFe9Ovcik+o+f2Bq+o+fECVBdhq5Q256wwi5xeOX/8mBtzn74iEiHfeN
Y0f++0FDEZ3h71Q3UgXxkOW+lLUgaMtIMoHF/EL3VjW3IETof4nqy02LcTACEpLwWtgC7hm1qg6j
dMBUiTy5ZOZHXoDGp6vuFAJX+GBr5cYHj7VnvqCik/Zac+pve/oXH+/QIkpNnFaJS3JzPXXg2EfQ
epV3seEmNG6aMDv7ZvzxK1QlwBf5bL7ya20HAl779bz7t66MAK8YU+xB7Z3lMKK4fToqFpksNxAU
96AN1BpQ7GUnPYchWIIvgEZ7um/qjTM1reqF7oxF9yfHoGzfApTdi7pVMrlgIFtYAeW6qhUsghOY
esqHns0eSNqFsNx7wF/rhKLK3cEDugAqshNXaGF6bBjto2KAyf/x/EFSQNpo7xd6LMav7S+yZB+Z
lg3cZbT5bc+/HWeq/bp7cokHfOpkLpvWfIpoB1QWXqbDkNhaDQRhTeWvDRi1Lz2nAZ2eJnlxMhyT
FTd+lOV3CIOODunEfEKYheiOfX3K2QU9V/aHJEV0a/NdpeTZGdmPB9y2QNuWu7XfgrarwfvC7fn4
8zHlsARgsnnTJeDJlbfa0yvqF5r3iayRw7JLHpq2nVgWa8hNAZG+oaxhqzGOC7h4Vx2X51lBK9ng
99z/umOcGzKsF2GAW2+S8nKhmlZu08oeEapUOb02oAuqZGSts/T+X5Vs653iykaI+Qh0fKg5WUg/
DkRv0+33e/VN+uvOP1aVMaqqekdFX27OZJyLnJ38XgzpPDQpjeBv9gA3o1roHY7IEcpMozv/E+z8
mjnQfvQtoHWj47G/EkxcIvBbZeODrXE++UIA5+YzMZpcYrAKCE4rk8rtirgiahiHJXSCsoYuoPA4
5P56HExG5l6Vuf8tJDkeqqebFU89CyC4PADfMWPbjIzX832+kBWcGG8Xok3WEfFP2xMsv9DP6elU
J0PdRTBD0TrMK/rzsZ8SSPAPimhg6WlJBG4l1n4ijV2s98GDfaQJgb4ZTnEke7Ov5HwEy7Are7md
SK8bwMhI3yCxCJR1tVELHHBtrEWD8+jNvb2KbFOwp+WdAwPv10VMP3uisamPuaAgg0F93P22yzIE
yUNIYjvJ3F3B8+4jOAO+Mh3sgKOHAdftoX7r577/ChhA0Kx/yyVTGuSxzlhn/kBybqRhtWUcaMHw
vbtVdTQYNHUnO4jg2iaEUFIhVgI8EfbptEvoyIK+dS/MuHA0hs/ORjn76aWzZCQANrPUuHFEXOKh
el1ZtPvBdTO7EC+ZDQlOPHzZVZwhj7eHZRSeJy12wzr7UsOmcK7R/CJ2yuZWS7FZVI6jpfjJMeWe
+yXkK1rx/9xyv560GbsrVzMF8OptytBUoWQ2EGb2OpUq/e18EoHGeJfFSjBwy4JfaHCkYzKgs656
3oS+hQDnLkJlWj5k9IqHTyOeqCyyqFvKFwT/Hv2SjS8M641YsFBTReVe9+WEwTfNUx/UT2dhrIrK
1QopI726QJEQajh91f+x8ZRfbEcI3N4dCP5is9u3dlV6sFJOmT2nTlF3JE20CiLxNmWioEIMDgCg
eq5OZ6RR9Q2t8eQdAiWRM+TNkXv7JqyDaeBdrRZt+I/tz37MrWLwhXwCGrSseu0eN8alh4bIlsrV
s5GgJNSHkDiem6v0v5WdTbvPqPZtINZ2sUaOIzvEPb47RR1UEzmSwEDsqUWzU07Qsa5K0MIcSl3U
SDI9SKTNrDlXEP834oDf5A6vZGE+3LyS5qcw49q03M2GmcooigvzBVI4zpfo6KzZEPdS/tuIHpcc
Jd2GBA4SZc0AULco1U6QM/ejobknorlWvudvxMSr8bJcRLmSkeJZ+6BVzAyQAKoK2oHJGGnhoisr
q3Nle2iW0awp/XXWImVBHEr5OaJCa1y4pSgyoLKchdHFnc4zqAnSLgMd7tXWU5jP8wuRN49IWyZx
2ay4G+1QmjAOgxdLTu32MAp0UfCBKDda5ESekDR8VtYyY99drnUBwTnjNe9Z58qxDT25p2qfNESC
894BrLUoGH1N8QtCyChP9Q5TuXxzYiwzuBNhiDXFg+JeqlLwaRXkaHcelEsUpzzfaI0XRcVyZUDa
Wu8e/sUGV3dGsiw6OSlXoVrqydI40Zv8vUSODo0HeXFXTdl1vu33fbwtYWT0kVbUN9nptHcl8g9j
tMOM2tcjiNIuxur5LVf9FhmKyw79XlwwuHovOURMiX4VEGwjejM0rxSc1dAzJpSdKl3O3iwTzuDY
THM/LQSINgGteW0mNva+SOF2MWXK4wAYZ6yahoWoOTQRz6gocvPEvnicKt17++4gZiqA4xD/dY/t
vKRSwWcYfD5v/q6n3Kp58d5CuEo0bTq9uTKwalAatXjdw9/puaGEkZNoTtJ8yoL2qwaCsS08hFaZ
11kzro0rpnvFnLrwaj2ubxr3eY8HqXY1p2cQM3j7EZGW9eMl12nFf5Ts0uPBRjW0JQXgiAUjHjcj
G4xhPztOQG3+m31oWnjPR9cHYSKL7yTTjuJH7zlRLi6jfRRWzSW8Y1eVkynC1OA1WYl/JpOFKpRe
8KesCo96ngmtynJs03DfvK+vVwYHQXJ/hG9L/K46FnGmHV80Bxt/685obWYe6I3jnahSMZUxjTpP
8pzI5r/qAt3O3TAREA5rrl2lPc3basxvzv3FbDZnZJ7bhGcVwbqqFNC9dPJQgCJC5jwtVc9/Zr2y
/N8SoFsA152rgWWxj4i4kedbkpCeS0mj863EeNeH19RLfNlDg2Bb1tl90isxecZX03ttDdDrw+yK
2xA1aorzZOnys8Edn5LAn9dRoDc7+slSw4zA5J7qokFL3htBN4FjkjDLTsUSqL8Mm60zfrSXSpnj
RZzsX9p4+SpJY+6Ob7SbCpabG5gEkwwG4zl2qs4PfEXcvn70t1ONn4lA9K/zk6TE8xaBiCfMIw3L
ZwS3F0O6Zr5S+SdTZtW0PzuSCFyRypjXPNKSXSZ85KM3Pm58mHq57iK56/3OBq0NzqRwyA6aXXhD
vWnDOJ13Xfa/obIourvWoVGOi5Hx6d75OxWm8vTiYQ2PwcvRBrlCUAPvZFRH9J8YUnSyrPtc+T6x
P7tDHaAY6ZxsHpF83qgpZN83GCNwO0mJr/XWmmZUUdUNSVIToDFIBoC0Thb4SalATl5p9WAJflCz
vJYmAuIq+EfjUPX5+f9lMnKy7DSdFNP2B0vf9a5o9kYBWyzBtouRmOLTayWy5jcme6F7bH1ohl+G
RJ0YVPuSgcdrdkQ0qIRUFNDUUmpcoQ8IU4OGPniodUZAmv/Osc0btfWqowadsxoueyKtE4w9SKtO
D7YVEQuyKBPtIRh7k80SRkoShsNeOm8kljnpfaW3nw197UCxNUspb9XPBTDdk5ko1NO2aIjKp/3W
qOtLccCcoE/N9izyluFBp14VPi06HdVL8MoyiUmVxBdhkv4juF5PP+/YyRnmwQsBemfnsw+DsRDN
tDRgJW8Mc0UWm6k9T9O0jKmJMOc4dD6LAqjLOGHlRAIHuLCWF6G+NUwXRwtMvK4QPQamqNxwhqik
3WGinvN9FL226EsLjkhJU4fr/efxSuZJZQrimvPSslkmbsGlUCHEO5GhdJlPdATgc3W+JTu0fPc8
praZxwox4p+AoTm5AqTDnC6ZMKdPr+SskIU0xXhKWjLm/JJwbXT2b0YI1yRSJGcTDYsIRH3sqTqB
ck6Z2wbInRYyQ0QpSgYwgjN21sii3vNORcNWSbire6YqO3nm0MGUFNvBQUCzVtWSMIf688BZ+nsT
zVPhg1TGPZYRMNxLbl6C8FK4XvGPhu2f5pMCHYyh6lOlXSicXQ1CClZh2K9BV9/d6Ca/t1raTiRk
m0Thdi7KYHjuS+4HT6pG+R0OPHojC10BYIZLWvVGHeR/Ris7k2H20cRIDnXknRPOexO6dHvlhRsU
payFWY1C/QVdYAa3aH8eO7pBaIz5eTQB4nwOOmvrNqLHeHZJQ8Bka6R/02t7bw9NlKaccUix0Btk
Ig9ATrDGJ01bQmyGDA63srv4cGMl/ey3LC0qV1cxE6Nfi2LacRQgLmUX/ju79G2fJWT+cAeEz5lZ
4yS6X01c/uTyrS6GEJQlV0nuDYv7XPbvM+UWpCN3RzQFTKr8haEPvkWAkVNHB0QVIt5kmwzRyR5G
ekMyuwB+BQtGTcMsZSUR8+ulTXZu9sJJykApgiWMbCyFCJdrSoM0iaeX3gBomeNcKFhoHP9Ip4+z
lMBITc1dbk+hTYptvoz0SQNAHy+hWX2CZfgzaxaXkTcubTYIR/HIO2N3+vAu7fMHc01atzMo09dB
DVbfVyRDcEKu4Hc5TM3Jip8NWZHKGTBmwBzWpGUzaDEp10sXUMqeBKFaJrnSn6F+QRKoIO60QK5u
RdtsPqomLB5WHyLPgMAoAnfLxz4+h5rFptDHJpFS6874QI1KvkJn8b45dEYec/7N3SNMaT7Sj6kr
Z2/pDDocM9xAeuyU0nS7tDURyEfKphSIAdtCNxPqiu8xPV6CETFzdH5B72IUgzn6DrocxXMHL+PT
7/xGXeliPs+TXy9j0liJkSJ/EsRb2ACcdGMeacL0nsR+WnrPrZbpA4AAsD2tAzoE/5sthxKHgI4J
RLXSUco9JOFMYIQavKEhPf7OQ4OJNiISD8iQ8eb/B1nWPy+J5N55EktoFibNIxLVvB/3vf5E6QwS
BgLU4jqysodLYTf7k5euGJle3MPPnCGdcOs/lQhS8ILR3cv6nWfEfJxInGEe+JGSpFQo0taUbrB/
AUZXqy9W9Py16p/CoYrfVZ33FNmn8KPGxGema3DHTGIugCHJtPyWCTqlCccigJJ5sQfN7cEtBktu
bRKdA/aHlWSdekJzJM9BdXGww5GgGli0qRnSZgBdAYNZM+UQNjje8754lUDL5/2rL+CIP0ol4Pdd
tRm04xZ2xqfdJ1wIn7uNsATOEcRyWIgY5kOfn5IEvO/6MoFWo0zig2rMaVuk21QpLNOF2ebyNsJ7
4hPJ2q2hwva2NejcV+Et/96kRhr8E9YkRS2aKXdNH6Uuyp0zzEHdfAe6+v1urfSqISQWkiKhuLLB
mYPmG1fDaxV1iB7lxEGx+t5wy8m3wO+7jY37HKlqQOtGDBHsB8UMOXrXYezTJ9g+Bu/pRS7a5NAz
LZYTFbUcXXol9Zi6xCg7KofRQQuwgVDZ5sG7K2zMLOUoeB41KWFiHTlOJn43ym5dfASJ6HdPqfSR
Cb6BJFG3Er1fqyjcHmBokgz/pverOeqiqoynDPr9/qIMYeOllxxBmYVx1kgG8lZkJQUiRK5XkiFu
Wx945tajRvh4NJWDTPkLwcRFdSheN585S/F9u7Bd3eOnW1dRQZHz5g6XaF4ykgEggV8S5vIYBxRU
aomOLE8q5HEhmK/INwE+B7qblZ/JDroFtEsJMLZ5Z/WkLTCWM41dAzNCf58VWMcuJBjAl/n95ml3
c3/75Y7wRi6WWdDfb70W2+VI08dCU909rH5NgdarKhKnrCFcm/Y51Rtp4M6auaOgTzjWRPr1r18c
UaDvpnVAJx2NvUzG1iQA1fsrvm1e/5AvLylkK5C0ruVIswFgNDgJngOa7aJiUM3BbP2rAkci1OaG
vqOEmPnPI206q4sZJIeYi41A8rZFaodUuPBGR1ACW+8Z6fHF7pH7nxi1/W4nUuxAhFzYYGznfx/o
9Zo32wzFJpZxpBpgT+/ZIuU1J2hUfOZspgutrSJob3z0nHgS+v5PpfZaPBZlaZz/KYLbgkNmhAKQ
RKfNH1tB0F4tZz0T6LaNE+TI8oVYuRoVqv+fhFxNcZYTsvB8X3FAfksiiEZ/ITZW6qRc0aDGwG8h
t9o1GaNAjbSByLuNTXT2fguoCJqqF/zArNkRSWJfTHX8TtsCafDZH+P711eFVxN+6CuF8RSA0iLr
df4sXk6+OTIX5D4yyNb299v3iHRNQ57jpxQsHomffO0xFM+zWUpVq4sHC+G7OuPPOANCYzmw/WNj
czWt1i0NtU11k6qN+MgcTby1vRUMlYrPvM29MdZOkZkY0M9AuZisnZuwS6MbSUOb5G4eti0iI94g
crV0duyf0rpJnb26B35xUDR9T41S+T/5iQOiEROTJVpfOFgmHsqNfIcOqn07R54c1QUrIvsD5f/h
83q0l/xcNuVLvS+TeuKz2cXd8eEAIx9XLZGyEhIGyOQiI2IFkO7X1j80Q2BDnFuQBaImogMX19dc
8L+I2pyozBNWvLTvHNUVR0f7Kv7K5yJ4xS3yrTYMzwRaZtS3DHVyg+9AwbOChLTHn6eLsFucyPIA
/JOFRPsuOPTfaeFb4cQCD9PSZSDELa1wI9yVmgOXCI7Dea34PKhKFXf5HrCKZVInQQVESNOJooYF
v8uO9rTtt2URofBEjZ0K82rKQ3ulsO1lueNziUnMpyd70dtfYnpWur56mGTIyxb+KwIL+QV+Jv7k
+FT6IufPDT3IpWaEPDQ0S9pXjh4RmrYeGKNaiB6B9POfK2QKkZ7wp5cYqwN548ILuozkeI9rI4QN
wdl45qPvT1EbjGiBNN6EQd8B02zwUcZHC6WVQjmqcPh+57740v0SNmWm+8zE9dp421a3vCjJFpR2
pSUgC98k+9dUuq5LaVVEztY55+IrhW9QrFWVF7SnBXsYMv9Y3k9v0w64YmvoAS6xS6wZCI8rZ5zK
9A1FowVYM+RkQlryYu4VZxcYSyWTeOgrcKa6wKuF+hsQzzYlnQzoEn64CuIk8U+niDX+J/Xnr6PT
P9MkAuMsfJy2vygv459eXlqHl+pz5jg9hG2jZDkEkJEvB2zxsEGOD9uDmd6mgk3CxlNagfWug9y7
gYBlLD7HDwCg3etQPC0Maj7LMuFpbwXJZG4lIE9sac2MU3uIWMynnoxfJbDU6+f2UKKQLOo8+TzW
vouSfyN3p4TIu6vxOBkBoHmityf7n4WtbKN8nSqLLX565IUYPrZPM1ljexASpsWFupx1nDWPBaLo
rNhj95lJC7ioY9rgz8lDctvbk/Bg0n0YTRSnTNPNhj/bZhM0SCyaWQPKVFyk7j359Pd0Ye+K0IzQ
8WBXC96MwFrw9C1ZCxfLOQIQ/NsQkZc9WoV5laH7ABxw7SocKjwKnnXdkMRxn8ydIrwZw9hetJOO
1RY/OkK28+MbHtcgxiBdYvZJ8ycBhaX2SPlKL21ThQP1duBZju6GPdqvBV5kIXdsA7AXe1HGC5hJ
x1XGAz8nj3g9uPK1eVEx47mc5dn9Ysr1uBmgv4NHOiMpyykBNLrK9XMe+BWyFzCut2l5eV7D9NSf
amhoXqa9Ns/rS2kfZxPkEm64JHUOLyzVtA4WUVqniaAmh0xrYhy1PZYQJ+pEGBa2p8nOTGv6LGIP
to1JW3o+pQ4FEfAhPSQFNZt5jYeIUe99PurUCP/DtOE3Y8c40pxLzJdDDODg+8uQmnCCYc+ASXnL
YZY4pG/RDShmwDfQcASGtG8lUMZHY8qbf02hiAHcHr1K28WfZWzFOmi2m2Rj/HD5vR38aLZt/e4H
oNCSIbooVRu31lZNYkG/kwiOQXZXXdyQCX1wEjnFhmOhV9shCpjYtoyBLgnfoKkp/b29nXGt24fW
cUS8cuJJbbW9JIJT8x49mIRBRBHU/OlSqQtpKb3gRL+Zgu4oGxUsmMVysNbTlfmWpu+qHDMdHZVg
FmpuR+v2nLQqJmDZEK+QUHkgQrr+PAOsZoG//qrVA0t7vwSho0W41ImeTWo6RowKSiXLoW5UrD65
8VqrqEAH/hJNdyxObg3DuewYb5GOMkuiKe8v743hq805MOO6EslQJHlNCFcuT36j1atsjJEMoa2X
fSXWk/KvMSFqcm51PlhrKkf/rxUsJQRZLJe/hhhyWKu3aCTIBiG7mXVTOmhOTFXl1p4g+yGEz3h5
yqT94KwJMfaWasYigrICwnGfONqR7ljeRPhwu73r7plT6l2I+cNO0SpUHxUVSp35iJhHOHwTIe9d
Cy4Uovo1iyTo8VgcqD3dHTqB0UVKbUV1Ydj046ZideXvLY1MzGOPB4Bq0O6lQOc6LdXCxbURRUSu
Nxo67iF4eXGaMGIzMa2eshOIS2BBSiYPlrYPI656x5EJx7jy/6GOieo1XElsun6LiRCorlfGR62E
XHhAYE/xNCTA26S1WcHDPCdTdzZAiNlUM8zpLg3f3dsQDWuxL52zB/JaqPZTccfOj/9J31RFPkDB
makwHp40RKlimu436+6sZCSfnOcpJ1wHE0L/Hbbcgm5ERbrWV+4VwZsfbzheLJr39xbg5ihyU0ut
kR1+6p0VkTVQLooFOsCd73VEnIH+DNmyFNbPpVf9dJSuMAucSZiF2tEBGGyL8yujpWdmoY6N3TRU
5qC3syBgFN51bzUy/pAV0dOhJEtcnj1/dKHPUlMY5nTFoiI4kPu4dGWDKO62eTWlu1tvNH/zYQ+d
WXQtw5H5aOlBeaxngBVZ5gKWX2svGqRy8ixD90IZzNThiwrE0Kjtoc/QjO0v0+djnhX5sP6lDIW6
WuOvo9qDcDKeTyu4c35f5q8wfLrD1J2TwGISDJsQvHbhgRY/ZXFAeI8dYgqYeujj4wRnxrsiukEP
eUZGIOLTGYFm6MW4XpxizOu3/jnGewBzHvKTUpBolBZywPT3nudyAvgoHs7ppskfJwX7laufh944
AD7OhPWT8wEhNWUZxwT+TPWUmoveFMZtiygOjf97o+k6LFacIIgRdMoN4MST2fHatEL/m+PeNUR3
SvxChgj4PoFHyYFDpENzFyADN4VUDSzNrg48k+MV3O8+fGGUka/4u33T6Ykjkit/J3zVBNqbVf1J
8ub8p6OqXj6Jo4sYumfQjoEpHqr0MFWy0MBtHtxKJsGgsFK9qYYamW1jVx1TN2yay8OoOGEXhei/
Z5/P1RS2lT85TkA6/zeup4AgfkIbGWx2mp+nWYCDvIPpo+u6l3DTIofxZjH9sd1RpTTfA8izViK9
042hJbmrE9CfhM9W+gDWMPzJFa3DcknuX7cXFnzj1aFV4X6h6QajYND+8Ti1e46a5zOldpfNJlW7
UmEZ2YeZ7dSofDgSnVd0kcSMbSHiXz9lLVajHaM64FuO5lCgNCM7Wks8lC/tSDFaFRhVK8OvlbeN
bkuJ80e7kCOMf2UPJSxfJs8T3Iwag1Tfyhl/HgCMCdoCjdwC9IFBB3g3dn0AJ4uhUYl7gEPwbucw
cmui+avNNLQC2tSqXjTCBZPe2pTTNkRyUWErGL2swklxiLBi6FOZw7Tk460qcE0Mep1HCogv4ARs
jvycZJkUKW9+NLEQPIHWoyRvwMyfmChZ70tgRNGSMVSUcgmae+NsiSVzvfsXXhTm7s9JGYlZGMZP
baW9eF1Jyk7Hd3x/HJs5J0blcH7AIxv7YHnjmcaxZAPC0FHALWEgKUsF6/pQWevhfxd5KuAahlnS
cJESvOMT//0sURXT5hf6ONO2i+CUcfSnvdQtS1GMY5d31nFhMypwWV5xFxyTdoOsYGRLBAsFO1u0
Wke0JhabfpEPhUKdBdm+QAjXLCXKCu/20zRF/MjKsSnWFenBFfhecpZzeqyIcqWSlIDpf6RhFj66
f+gEyUeqFjI4uVM5Cl/RKICQjZ8oiJJNuz6KLddj5XvurrPlBaHMtaZS+BQSEaycdIn4Ia5U35cl
RtSIhOVc0azRNmQt59InEAitpmMSCJO+IzevE0K8/jq+q9T/JJpThFb6cUTp7JgpagYjVIPJS5by
n8DoKWUoL5uGDDrVGVXSijG6giaqWJgHTZkEIEZVLh5fnE5JbYTFVayJPR0sUzZ+5VOdCG7Fl4+N
Um6PLsbLn80GJr2Ft7jYBwu3AgB1QckxDpqtCMqEEpQa4Mun1DzJf7RG+0GklC+MmaDKgdvraCOy
sScsBA1MjSaKsfIerw6s75U1ptcbW4/oylijvFN/+Pz7rRwbS0oKTxIVSQJSwuH/Lnbqzq7pJ7CT
TgZ/S/1ElnLGFQxs5Y/d9IgOlEncIV5n4gUEhAkRfyYYcBeXYIlzkR5wh9J5nkgnpoCzjSsehBKn
1EDT32BT2VzikHzwE4Y+uF70SS3XB7+81Ny1dOAXdFldLai4XbuR7b8Vo5EmOofaLKBpb7JGWGR+
Xc6Xz/lMsdpxSJJphnCH9teS8HbQH8PQb4iz4y4GMUNPHEZbxSA9BXsUGvyceptOgAdCiwuyKyjW
y5+BSyI2QFNTO25WHueMRii9cFJEXpa2XmIUsDh6WZDsUbDXOTIHun4jRcSUUnHH3E3kBCuBH69n
NVER5XbU5ZNh+74ZwnqVovSyaxfmh2PAtW1AoU/mS92nWL7mGAZrBVfwv1HnIIDQIDDhu1HK8xhh
ThH3oio5gOmUNQ2AXlM9WL6HUEP7uIkJGcOBgYuI7unQYeRNAkKv8pHmzWGs/v4SYT1/iwGqBhbo
lTS2pthKElEEwHBZj9/AE6y2qzANPVvI4dR3uzdyZn8zc2ywbOF3VwpOJLiiU/lgIywwnGS2njC0
TfQMaqQ9GF/09b+R3mdjv75KPc/Ni/20OP2B/3I3lk39VVY1v67MhPXyUs6zxgdisGDkAaBj9s94
yE55b9hwCmKpcgvkTSQ52Li7oStAxUWanw6Lnai3lv8P3HS4EThoL8ysVj+3Y/cggf5VLhVRyT2B
t2UdlwzzZq+Wf1HECBkc5H4kS/EsHgz4LPzAsn8+fQ8PCktT/pYxA6fGNsfw/UbmhqdWJuFWKxsW
znoR5AaQZ7aLPhXmuJBQGk9uArHMqnfGOXiuAqQOopp+zEMmwLzre+NuggThTb+QTZ1oPG68tjI8
CcDJK8jrd+6HfETvFDYOOPcEUvsDVFOIj/vicc9rw/MbufiebBwjOvpaqjYuiggkJ12vj5CKHM30
Ig+BRg2Xbqf6flKCFqZ7WYp+p3d2G8BBT/uAtZ9RIrlU9EDP4aGq1wL6xOHGcWtQURzdUC/ibb+b
n6Y6Nj0cz6aePT/Op3Uj6Oa2Bqj3azHWfr9sIP3B6GEti5QBeHcaNR5v2VGW4NPBEG9pxEymjhRw
0Lxb1y1wGFTu4RgJvVrsp25+0vLTGeoXjKJCYlbo5zTa1IgtKY2qmV60dz4UW+hkZ1yOmYyT17kw
0f5izRJ4a88D1/UE1f71RFGwU/7YAZ7v+4VID8rW3y664+CH5vCZSiUFxLSAL/0ggETtnlN5KGs3
WUt8U7DdG6vEVRGRqJRctck8lCLOnaUyCramBoh3PO4FFEaEWzeAMSXDM61bebPkyUf47Cd0fX82
HIev1/FDITzQtiNw2rmzCvYX0IhfbR6UO5VR6VK2v7kdi6R6QrNKCugp8786zWb43xPralMAsfTR
g0pSc9YN3qT2z5IX4yQeHivx3T9v2+tSwsVFEHZ8Ko07GjziTx4dFd8TQZz3Ro05PLJryF1apUuQ
FmXzALhGPaYsbG91+VGE6XEnxLUGCvOKtbCKq8c65xsVwtBxF2uJ0sO3Es8rbSh1ZvKSNdvU7WAy
yIsRRRBMl2PIFzJ3g8FmWA7C6kmcIGRlu92JNfsGh6bqf/iqAVP1NTznr38R9A70GUWhjqRzLiTv
Pp01c54OVMywXCh8r3afKljnvYdl5d9tEh6858gPBI3Q3NP/ylCGwURMC2UEOUouG9vfTLEbHI9D
vtQnP9/eWim89nlwwAU+ASAsadMws51T3VHDfuHfJkIE1rxcctI/4ksiBg7/SWgX8ww6VQoepDua
Sq9n3SoOol/R7ktVs7Prf+0k8yi9Thee2+QVTIZ8GsCkg1ja+byL3mIn6HiDbucULkTYpmHvOSEa
PIyI3jIRZ7JT92eqDY06vqH7B5Lyrrfm4bobHK9ZPrQ47AngP92NhTJb5/ZHgpgV6WWtzUwVZ0Cv
WVsLHiXWgw37E3hfrgTA4iKgjdXEm0UJng3g4zizkQ98b1vyI7cGzlkZJ6OFVzVWohbuHF/9BvIu
dI9jY4IpcfHgaE7vVqdCHEzRMx/3wx/J44661aUAj4Nvn3yO3CRdYu1V1QSBAynTS1Ma1gVWtCFa
JstS1L3+7Pa2zpLzX/dFeXLRr3EsTG91z9XEP7u7GAsV1RkeTzUc87uhj4/HHksywVweOEi25nqs
4klFWIn7YP/epbEBrS272CcBtR/FH8UkYetuVcUEpWiFr/EU7PRjxmtwUlIoiw/sioUUKohj4EPM
dTdTfS6w9lhZiq9LOP2WM8SCkZlyspGp5WixV0m+IpK9ljR7Fmb+FUtvZICzIOxtAidqDRewvO2F
D0oj/tLnUX8U4RNdedgLQAb2nFwG9oik1Whz5VZsudgaro5xoowvpp4wKgxy6wi1qs1uJ4x/j3nd
Yh0vJhDQ2+wt5/AiExEYvGdiELHYCWYSW11JSYdSbsmsk4n4Io2Bv7QfR1C/4h8T1INHxGckGL2n
rpnXHRt3FReiV1ozgmBTEh0r5LBAvHhJ1JQbLD9MBAMRg5KYMLgSA9aJXpXCVHW0ZSJurML69bfL
B7MFGH7XEaJCQ38+visnAdTWaftKPVk8TTdjs9jQfKU5LSpXl2QQaS/XUmLhVAig09Oa3l3jnlRp
DKhgkemk0xd2NYT9RzmWCE5XUr0Hd2uHAdZnqBfzFFlBIokVlXRIfcN21HcZULh5MlAzbXpI+dDz
lKWmi+6k0967MmBHjCvN8gfifeDc5Y6scAW2FHdm0sWpok7OjyqjKMohXcEl/VIP0CAbWphTt7fM
oVPcKQajZqo2XafX9aIeOCknMDkGFX9RQU7DcpS3evt9sLkgR6CHXFAR3vVYPlFuYRl44ve88/iX
Oz8h+6FZxgqbY0J1sqizIBMNHoTWzX3ZWet1zIyf7wJv2ZKF7sJQ4iILATarbA1Z3Ia1+KGpHWJN
YNY1HxoNyy6NhNLA8fRti53MyOJNUwqljUnAb3aimFGLCzYQ1w9t7COO/ux8DvB1O62UYffXswaX
N7SD3TC+0A/ZEuEDccaqScn5cDRlnfx8mv7M5hZkaZO8Km/WsrNeDb0QpDceonuHsJy+wJM9RGI4
cqlOAtcnB/Yptvx3H/nj7veoHrUhP6lZ5h9uDfShBXaWtaPPVrjFqOhit9VXrMvGhmH12SoT1Y0v
KRvCtsgQGB67zDBIZNKIcOL8D2JBvhV1Xo20uyyMBOQyCSGw8SjNDn83RzjwQUZ6KdRFXt+oQI/4
jSL3bLoFHXs0XpOKO6KgCleJ8FB0QmT+OoRFDLJoxnHypGkPWwiUoddW2bVyWAMehOHWpqbaIVel
a9eMTmKcQ3OS8pzeCUmSrYAZSvyJk/w+Bmb8kDE+mPJoH7vWUGQBxf1gUcBG/ozv9tbnKpfNf1KM
CZi0Jw91yobgjEICsY+IYdC5mNdaVr/aqDMb4PppbRHlIsTen8oD9O7Qpb+kvcmjmShTyyP4XVN8
tzVBsHcLbjVEbQvJX+ySHjIRRGHK0oGyjuubjlCKcRGLZEb8dY62j99BzaXR/B5PG0xWQ9SxvS57
jvVzyOJ691Sngv5DokYSc8SDfUNEJZfe+SzQ0lj3KzTEvk75Pdd3CTu1yspNlCEFsQqHXTOWBbWS
uMVrRcal+BQ8JVET7OOYysm3nUTXl1mMkNTeMsciTeZJAk9r9+SjjAnU2WY4vl9R+zq+2yTGqNGy
ghiOJlV7yFfELvHoGKSfwg4+SxRBAyVdzj4q4rgGLQN0fagJjc/Bw+vLB13uEqJpUYKpz4c6P9pq
8Kv3+TC9HdNxcWVs5EyK52tXS9O/pW5XwrM/mUidTMkuq4lSl9BAxDsDaw3aG5jiRBKUT6NHALpl
HajRbarDGjqZPowMpwsvnFX19suVmUPxCkmWeOfxrb3tglBA473UVT05KFMQSvAvxGZmmJk9VaVp
GLmkmvxEMNnhrT8sOl2lsOroYsd9cF/zz8nXQE2ellBTPaqlZzE9tU4J/IYZTnqwYlTGPflCn4FS
6FKwUnpAKczo4lBdNGiii5MGagMiD5pzgXFKh1f0D8n1Ybp5py3zXcG084JwWoAu+2wZ+dWBHf3C
aBe63LBqMdvW+3ukAZa1LTo+Rsz2tIlzdnBQVAQfA8Hyp5xBq6G7moCAb52E9n+egILIXew7LWbI
pTVVDxJ1QVgXRsz/Blc7DGi1mJYISXJsO5MLSyBib0YZxF8icRpc9pl7QFQpxI8dwH49sr5sLYyY
/HD3TB3U3CE41vUO1c5zKLrLwbA//mYyOX2rAJP4cog7UChe1KTQus4pmfD0daGPFzDstKDtzFc4
7QRW5VksqWrrrR7SVManVRxvjvpQjqeN4ZTqIjt8llUxR740FPdkcP4DD3fkWEvQRsQT0qpJp5ey
5Wi1mFdTzSvNEM76cN1zV72lzCfRXUsU18sDl0ZznxQwWcsSVZCkFnzYDzLgKu0+hh4+wrKiE5oT
SFRj3/y5/xKJxMjYqYnt1ibEs2aC27122F/zXG6+/ZkSsgYHhiXEnhx7p7DD5/88k5UGrV16jn2Y
GpOh0MpzDwiouTpMtocK6uENZYgRyMcVXA5gH5lsIYnOSh6K8H3uEaOQd9GQzyGaex0QSeslvE0v
mowgYu+CoBlG0shShr9jmKMmHtKeDkbUIZawOj7LtWEVnNWpjMOe7XHhrKvN/n91EUqOVMF2k358
4gjWgGGI6aSSRFCAQLfYAKC5VCMzzlcga1KsGZI9fsp3/9qV+fXrNAF76bWEPQqGKGkt9A7v/RmE
YzENvFrNR699mjumJk5+ty3z9LmP7127ChtkN6p0pJI1Uwa8QiM92KF4S279XVkxhr0ORN6Q4It4
cPCyQSKZjs0KY+29Z2tSH4CWIm44e12SEmJXXiJCv/ukDLolu8pongh3R9VTIVrvZCAbD92oETMt
WzBFZr0wC40DwWZMv/JcWLdof6bYO4k+K2IXixo8ULKltnkc9Cugo9sdjgBAoRsOBgh+JbaKt0xO
JEsd7njD0X8zzrsSkMBqUXztn82hUdaEaTS0WUhgT2GMjZDD8X3WYVPRdvB7eBznMX5psy5p+aUg
+276QavkOownL3HpI0MvG9kkN8frWYr+9e+hHGpbnLnUiA9nQONIpLLrXQ0vYxbT4Cu4Ghez2YWs
b3Mh6XwVBpm2bsTILlmGRMCgSeWoPLzs4WpcGchIzgF5BluStAVU7Btnn26vtG9AaSuGDdboo0ZV
5L5wD8BUedkgTWtU4rGTrqVoRKB/t8ag0vgiUpYQN4tH3WPn8WIj6hFeF1UtyQZLH6ANv/m6ypSb
A1w8Ar8LEXqgD10Hz34/6CWB8EZbcs5vuT/+LaIk8cnLQpIG/PYGNMyx1o9XIb/VkURZ/YGPgZnV
8InpBungHoWCdhX3aG2SjPx4qdqgwxRybWA4JAcZHuXAZCReixV/zbj4LtTUTxal2WTGwXwaVQaB
gJtNuP4cAjBAxhZ3WelmMiSb4GBYdB7mkupDm2lTph5xp6n80AbnalKajRrxORrmMUXSgMqq3plM
pLgOPqCQx4nlxviXYxFrQiOxfeCkmU8i8W3bCgxAUCKoqMExdNFosUrb18FwlzAF0NgVvvpO9sNx
QZu7Tpu62ZrAiLcIW7K2kcdydM8hmuUx/mn9ac+MnIWWmd35IZJgSlUvmP0o0AHCjAFsgIro7wM0
E/+7T347TvRiV9iV72IeBlTn272YhOROuCLP0kSPwN7tjz+wWh6AwWgylmN7m194hUQmf8+Ey+dT
at/32lDmWbajzU+dQf9+A37g4YVc6PUSS6NUlYsMQ77pXRkA7NjhssGdUC7x+JCBaM4jBAKhHqwM
xRLZzWten65zDAakVlENPHqPs26srzExHiLHoFpYuNISJqs8iML50HGG7POdtVodJKCuwe1rb2h/
jbeCv6MCYueP6wdYGfEdvhnlOHa2axOjb1oCrPzh7+P+yMmrDm4NfCneCBucG41Drqb/itJ7NNRf
Lr4199BF75aODcBDpKjelMDCQXCfRpduP+UvQ7vi26qvOt/CN4wBjR5VQ7V8Qv2bsVvkM+4j/0Hz
/ZHwmHBlAKPO3koSxL4ROur5UfutXlm0XITQdoNkoVNNd5Y6eScX2mYYjYdwoX34ZZXV2hMwr0DF
Kqda98OYBNn/Cbih+bcnSKHXnofmOkiWgs39CbZbxWr/QWxPSPmSHem9Czx8ytdx/zRNL0y3Ij8e
fvXPev8xXCJpyOuP1bjTgPinmR9RC3KTA+ENrZhtS728F0JeMRDzxC4NEhz2+l0THKqnKoynKEqG
FpeG8dhw0afOb3vRbs4SiIBAr+p/AEdw+p4gJvZTJqkU9BQppnI5ZZ5l3HKYxiIg504njn84NJZG
BBf1DEfnM14Zo2hPUzeGeDkcXBUxJQKQRPyNVb5bjl1jnQliGw7gqaAZevQFeI/sNE43ckmspsht
Jskin3PFfmkHa+LfQvFJNxn8vkXmGywZdVxrQ7HD81JvX7HeC3N6RSDZy98bjeNhY89dJnbVAMSt
Q8qMTNrDW0YnLKjDS1hGcpQIobchHPpYLOCqZHFvtCKcDJz0UnsKgi2PgyPDXluVHCpdtR6h5xut
VljcoPI8IOjYw0hEv5dpJgbUPumwPS4A7EwxrCe7bRctXQVqnwK10kXUvdayhvquDkE22gqWve1X
L//xiLcAQ4xaKT1RH2tzGpcVI4SnfeaZzmkI1uT7wwMfYqYPcacokI7IURKdc4O84mFstCsk/U5N
AZf9AHty4CEt2ZxR1FKiiStaej4zpdFpzZNPkJ4D0mAcfcDEyfCzI62hZGluSEJX/fkZjCmcuRj/
CXTZu2ALASc2O4UqWWTkYuX+soMrdP27DdTwVT7ZlAdSaEJ3GmdzxokZkwo4YxV4G233afj0mmyB
wAk3tn+szLy5Cf0D2Z/awdZG2ecXmqgnS6OsPMWBKaL03HXYpmYJwSfBPlYDmUUgJth/uKAg+cSU
BPGFMFnusbdiSzk4omt81RxyIykgXOsuLQLdwDUu/X+xAYX1fLZVlBXMEAw5mrWvyUjN+oTWYPrW
Wx/8Mbg8AmyDLln+eqDTfqPpAPZ9vqcW0GH13j6iIGW0ZbQNF7PywAAUsQ5ngA4kQ3djJT44ST5N
siRmhWq27rbr8kNYaUFN2HxdCNdlhz0xAAmyvThf9fgCPp8EfHNOC3r2KyOd+LVy58rvgfXZOFpR
S1rskjDDILJINSZFTstC0uv2WituOsRRREs5W2CnfURl/uIv7slxh15qwYnNNgsOy1Qt18oDNdtn
1k+7i/h3pGU4W8zSTmGKy/VQ/734n9baU1ohH9zmQDng5UPAWzCdpOzQ9KAak+XvkHdi1ZO1T19g
ZQXlZ0pRKmxMf3I/Db1MzhhoRHUjt54A0kt24+iElnKWzHKJoSfqOr4oieK3lSKrCE9VLQN7y86+
rqt7DYIKWUS5hQJmQg1e1u5M/sl7hIQ5ccON8eZVf3+8kZZNRLIIpWExe8Eb2Aer2BlEW9i57WFj
M0oLFIiu4u8lOXh0Q0EzOSCr1kDMcMTthGVaE+US20QVdXm6n/5x1ZXUZhYX/2tINR6JzjlcENbR
aUeioF0WrYt/4zKmahHEOKqZN9j4J2PceVP6g7ZdSqfkee35VTct7CVqHxZcAEq4Un4J503hkJ75
aKXtcif0MhyNsPbHOF2CykcitQUtk4YN55CNUt7/tPbUdLheHaEO/YGTYIzPzC0g6TG/LJefhb+F
Fw8MCEioLHpQXkUAcXbzbEDrYscO1VvRUAsjCUCKIfU0dWHmMOXXZOGCTW4pu+0PtHvoXF8aE7GL
X5TlKvjTfNNM1Pr43zoK/nyAYwRN2VpMoGXYCMhW1tc83MbvIDgIQZCQMG3+FkmeMN5FjFqQyMI7
53aH7JLTAiMr2wRGktkWWqTuSSwQn0wanHEP6kGOyy4/f+YPhR+UshobrfJPxNwj/Ub1Jr9A5cG6
B8vfg3vw7XaQxkiP/d4KMWEvVu8xrmezBiBwLmFMTiX1GtVTtkzjTXIc+JMTiSZQuW19vNcnBa+A
2lxVJbLixL3J2bg13/yKlNeY32iTYiPAlSsOydQinQuf9hlz4VvIdU3DGZHMd7aWxVY4ozGVqw+P
AMKRzeKWC5ozhCJpTNLxlCEQ3EZ7j4Uz8teRUXIH5QqiCvfXmt/sMaKBRL2qkj5FOZuSCZEIMGC6
x5wvycb7C4sjdme8UC0WtITKvtcbI5VSjp7jy/McntbUno16oOc6XAYvcgu2YKGAEo5ut07WurL8
doeELD5UbIXGcYPUmOhKbdC9NB+jFDk64t9sRKE2JDtliy3tTURzstk49cv5u61eUmAHh8ebi/5i
hf9zeja/Eu2LJmmwhiPhlyjT7+BSwYinceRrZL/6XXk8uGMOchQZrEwLZ0/27mVC4zbd/KsjdC2o
FK14FazzkI4+uIc3RYQr6q+dabkE1XNjyMF3onyCHyCUZ6HZw1NM9AnOjk1HEjzByRMqMXCxpF73
cu/28D88THIxcbnYYGzOsaaDwuY7KdtD8/8v0b/W3omF9CU5ckap0cheOl9sOsX7BoSC3eNFxqQc
LGwQdO3E0eg4Zivt3gm5Nc9xA5rgtVxKs1ydYO/i5MSQt2sWnrh2ITVcI3rKpqcjVEShyIWvaLdd
JP0WA5OJBfAa+QK/Tm8suqcSKCPpZ6k8Ztb3+VS+n+rRY0qNBNfcKY4cfBIfTwUeEKZOoyPXIqm9
veYvlm0GusaWjEO0a9Xv9bNQDdNyHx5iozlAVPW/O1WPCdWAsVzjxT9qHMdHf6uMixiDuQnFZp29
0LrNZhsauf3AzZqT6W3pfSxOJTX2UkNmTdyY5QtWUdIPGLIzDGgkBsReFcWWz90SHLXWaqjOMcx1
G/liAwCEMv/BeNWLoogFQKbu5XMyZ+NXvqVzFUW2Sfn4wp4ngEXqPxiI0hrY1tzwb+zEyyEJSoat
vyzHdi/EZzkF6OTuHQ/RHvBp21FJyBKQwUUnS3Oe5Z+YmB2lVStlzk8gTunT8bxQMtlJkaTROALh
W4I9Qntp+sgTO8ZV9xGjxzjJGrUVFI33vEjz+atS0G07GRkolgs9+R/cxVzRVd5pAmlGd1Gwf3Ii
RMpRDg+ZojVwzdCQG7Gj+bDOJpYfDsTI7K0rkSx0WgZhFTe4Bv2/MIxCMed+4U4vz+R4NzFT5h/I
vCFaT2hTOrDN7nxqQ9lxzMnGUscRRLuDQ8M1yHY2/VNjvD6dO7Q2QUwxNY6N5LWbgMvivSCpt0WC
3lURO1eM3sLJwcWh6I2S24XF61v5DLfGE297QxEilGAZpeChn9Sd3DUBucyRbu0ymB44c6kBdARK
EnHLNk+9Vzder2mvQxtYJCEX9P5dxgOkXhYvVUTL4pP7cpJ1RymaLKgRs+cwHEkwl99ijVGR4+DD
fFcJw04KMoosu1wQi9yFqMfNLpOKXlt1Fnm2v6rS5U+U+gWVZ89+lxBJuD79fdwyRcUhl1gno/57
MmNDxyLYw6T4gk72jkPPRcezufWu/J002ed4dtOvywSTDawwuffBI4xxdGG0fq3RAzKFzX3SlELq
arCAoA30rg9pcfCVutT0ms0LBese6Pbcyl9EFmOLbj7aqTTZwdhslM9xG6YbUuXdYMZoDDNy9g4g
pk3Y7qeJVgSRTb6CJuWJ32tZJFYY+/14RVv80s7Tq0jp6ErONLY8A4hRdEF2CcVbmfjsIWQyWiSa
ziCLdeFagJweHUVJL7mYhin44dSxLyZogHNkiF1CW9mW2zojnDmSYLHSZjyOHcZwaDdL6zXyzZZa
oqQD1hLKz/MrHuJRMlAXjpBnlx/OzrKlebZCMyvLYEekZexeeFCty6YvvNVQtvKLvKR78k/+S/y3
/fou0FLbwhB7hUnFdAa2OLr9UIHX46ENjaB8qYSI8z5aPxjfolYXBkvpWtFHliHKvQLCJlcg5Qv3
O5zSouqE7sBbCy7hkB9uEs0tuiCy1w9VcyYXWU2Q6O8pnN3NhuGn14JFVCLCy/1+cCmVjMadFqGI
RoBAdryeTsarLUIf75IYXF6S2tMH14gj3jz4CsIH6lZ1GRK7Zi+M2e6zip4R0uhX9JL55AWe1I6f
vcrHdYCFpVMWy1SqLOerIYyt98Y62CLr7FXQfTkIX+nE8iQh/ezR5J3NyGKPTnPqbnKJD1HRGRmX
GQzNFa7NvncbsStOtukwNeCw7wBMIkijr4zu2rtFCBfQbd0jDcnzCDccw4cWLpt0IpmWEHG5uurf
twAaifGtYj56GhQE7W0t0FDtJkfV8XWRmk9Wxk7K9vQ5R7Ll9ynIkFPXZBlBYXJ8AgU3wmrZvn5/
W1i9al0KbfME4rsXP0Vh3aO3SFr1a4Lo2/dz8zJwlOokWITdJLkEF4ZkIXgOPVu6n+5UbxuZnq7Z
oFldCYxFqn0QQPh/DfvhtRs6bNdtZNClj+JbV8j6FIcCHsOeO5tDRHkjtK3MtWwUPVq527Z8si4k
X55haAzhCPJZnSr9o9lGAcr4ByEdi37oMNhz3C2x+xs/FGzDpOmMsSYVj0BTN7efLA5TyzXT0OWP
nBhLHmUfLoxw/qu+3FTlgZ774WCtEIFgZ1zRbCee6Gje4Q1vMYjpiKbfRayDzVf+EYuyobw6YZYH
5les4fyl7cC6Qle3TGcAmlll716r6jcrxtrZr6Egft4hxTOmjkYKFcFYf2oGqGxMuROUAeQUvuz5
jtxTcDOAKlRMH0sCqhXgVgRSwxBoTB4/ZxpiNbrPTDh3Jkso56fvqVjtfTLKM+mJKKUWPMa097r6
zH0qQgIKvVkDuDB0KjYG7GJeXOv1zjRAr3GaE0cSJDixhYddqTTVZnx/WEVHguMK8bar401dsOjp
syilR8VT9shcstQiCRcHz+Y7LNmZL1T+TJamQalUF02RQiX9qCFRMSf54x6OGKM09efQUwTaG2mp
0+FkNByAViJwxKIQJxXvM5Xh2UxRD+KhQ3jGuuefYv/lmkgFjF6wQDIgXYWl6uKea3uZdd9m77vC
jYYcOjZZnkyL55tD2Ho3gjrJfVZofDRxAZ87Gq7w98NOaU0MLVJlehXzetuPqSd/RgwEGihKH6tu
es4a4MqupVKqgK5EwlVqHDXCVuOyHWw6Ph5CFYP9LkqoqW6Z1yv9PMaepnRiJ4x2cG0JA+nJHWZA
fUYa89vPydXxxhaMGWhIpOaUTrNnaDw1BQdWBb8ANlPlh37+J8eSFJXXVuCEUptlb2mP123XDB//
qflpGAjWjcmwQCbhGRTsQHzrVKZoVpIFpcrlcOCellG/DKnGuCh1f8sEweYj1+JdiqrSxkkAaGmG
GCYUTNv26OqabJbKP1kZfUGg72aHAkmqbhEbH1x+t4PKmmEJLt4dS81jqqEM5QBkMbIQvvSiEBHI
AGE28di9J18CwK7m0LqEBgo9/xBFgvSiVHxnaZRwgd38Flvc4vtxSorBSrukQDOjJw80l1QT336y
M9ufz3scucCJtxR1CdTsY/d9S4+gONZQ+mdl68yHebGZBcCGYAuY9el4Psoq9rLvyXyLungrltOv
xfUIMFd1anWFh7DO6TfQ5z7sHhzb2/Dav1nPGbMkzUDGqMiC9lEx8skLn45Zud+H2E+w5X20aunm
u3CH8H9jRu2P8X4h8Hinc8QEMesLIrBCZbXdOGEHRmTI4nFTKejeC2z8V+DUkaKckt9uotGoL+WP
8IJb1AQlsW8+0tsWsNVhK9xh+lR7tFDzBe9zmfov1oungHFwwxNlRuSQM03TJHIXhobTncNMtGOA
pVp+ub1JUvAcaCkC4Sw2uZgSwFm41U6yOUDBkAY/uuaiXKbpPA/OJLREw5xakXy6yQczc8nca4qN
7eL0zxEO1E2Wl7+1rPWrCooU0/fltruFh40zDbvDb+CUA/WR07WmJsFN9OQDrwapiAuEjJdUAddo
pIsVZ+WTcalJr5G1Z17tjYtMT6bgBn35e8U00h+1UD061zMd6bZnV/HgdvjWpa2xMBsZyw4/ULjd
p3lFsH0meH63bupiZ7+nsD7I5WTcZZILWARNfBpt6NxkhVr51JWhEqO/jB4VulaFBM2AXyZSZutZ
5xJHm/UUs/vBmXgoj0TxLfBNfDtchSOTjfvD9njrc0vuShik1DIiHWnHeSu5p5HCya4LcAYUI80m
7aQssS+skMZ3z8gJc+3lhv9QR/trrO8BVSgCa42bVwfwbbO2Dav3S8gyig6SyAyjI3uFO4jZbNWZ
iDuIo08vErgIsum1BI2Z+gx6Nfx3l7C0bZ/d2WVVi8QPsVdWJi2djNcLvYSbKut648qJnJ95LoME
dSCjlDKr5RXgw5K4H7npqfw4KsMQFJvTu/M/lj0pN4MkmufhkXN11xjaVweWBTDSzkJT+O/OWFQx
cGJ/HIt2N0uJAyUDA7fYDeU6kE9KNizMxjRtH9yW961EZruWYqH43IEs3Up9lfFunVKDahJsaWTv
JJD4znpSp83SgS8k3xv1dE3xRwjyDMTDONQYPsKE075JSjWg6/0u8KtaLvl+t45ivFFy341G87H4
REZ5EV3FTpmojlWB699JnEIzywhm46CnZ2PUyId+SgB6MZY5sxYYrUUgKIt/wds7HJ+U9EW+0se4
cGWHTMc4tnpNw4SVa9QQz3udrxJlMy0FzA/1imxo0SLe/n+JvJdpRyTdto5j9wsBKdLpqB/bzAkF
R8UST+FTfOTZVm/Pp/q6M7S6nuCuZwS/tkCLQ5RktkAURGvcHkKtHVDQ5WmDKhibj1n65/Q9bz2B
HY1TgB4g7nc/Idc0/0JJrkaCCvPrxju+xCQ72qsdHnpvRIezedYKIwjU4VkerdgEleTlycqcMfOm
Ut5ACNzahpYwOAcVwlxk7+nkSZxs8Sy7dcQySAKyiFnAKhPiLUUQ8DuZxjaUtEbBPw59pF5NFmlS
JJJWADikeUy6cfU00oIGFcTzGmSwRmwK6EOPue8wLjNZX6MGvtx4+QXcqh2trc7HEDO16MPG4iBK
B4jqmbF6mga0hnjylFSiGfgFWx3cVTa+KW2nBLqQf7IAqLF1DHfDcu0RXaOzDUUIURPjClMVnX/5
NXG3wmxYtx3CNwze6o/G7jpldRnpxt62bfsR/7IW55Yj3ZseeN12FMXc81XxD2FIHg/+nrSyhxKe
kc1hLJY6qyJal/3x2KvqQ/YXfw6wELGn+EYo1zq0NyusST3hBFunpKHTHhJvMQxaPkRGiyJWKxL6
NRHaxJHb9l7A5i7tr9tvFrpVeqNO1BTR8gLBWj2aw8n4k/qPzlXBNq44i+PwyKUjvBSk2Fab7IHJ
m1boFLQwMLimBW5WLx+3x3TCwHTC28fWvZlnTkfCOnTZP7yYTLc6KULvqHvuKCiVCLITvAsJs+3x
HeIs8W3OxLrHRfSd9DYKSL8FcWD9scsWhBBPhNwJnlPXduaEfp3WujMbkeRd6KluvZtjb90wywhy
4gBWjRPmuy6cbmVrANgbIKFVFRIrH19ina4LfIJ562/wb3G9zfL2BU997dNbzWTCK7JXCYmo9ian
pxpqoGKeMAu/430XopfvdJSLz2otIC1v4nsgviXDekiwin8Ee/kJeMN2mLqYb0TD6nV2peIpMwoC
RYt0TwcYzqjFrHBgxEJGWbJcNssm1j88YDvxNSKSs4cOw+fsHizn8KB12gX1eJtwNG3dVR9vEUg8
AaPQU8Vre7OUwW8o+tKkxbkcGdlgkCifTjWviVr8xVKgaDN63KMFnOuMeMudSxq1k+JPgbAX9xXn
H43evK4QiAyDFkjaZXQPYqj33N8FCiZSjTJmSsOxuMnrs2i36Ny2X4mGRPW05wdABugcQN9y+Xtj
MBRJW2xoDI69+d3J3ali+x0CCkUAgv25a2NcU4pbAa/Q3eNC36DRmgKuephNMLkMleyceoniTHO6
ex0vV79suQecEsoQN3/aqSOhWVpC3JG+D3TEKny3uQ093hKjVoSgPdg7U7ELRdJSxN2IHAtrvy5r
GmY5woTsbpqVuAnLBGzIggDDvhHQplPebCAi5jcl47x1h7f/rJwx4sKYa1prs0oiNYGIbEFuJQAN
CKpGom9CVKM+c7lZ9j2PbN2XLpuQ52ZGlnqFIqaLm3SctzBCnYHQ9JLMn0soac6s9KgVNSojFPB8
wlwCxZkb3cKgePs2D+tLy2DIl/lkkSRsF/0JhQ4DAEkUqFzFtcGYivE+LOL9RCwA7i/YHoLAac0+
GdMpTuwcL//Yp+Jx9R6KYbyhSKKd5uloLDviiKB1Nrt3BzlRGh34SibklUziZD3I+wL7vg2giYqW
G9v1fYhoCubEcfaUktkVx3I4r9YNPhhN7oYz7Pt5rAyB4t/Q/qgt2ua2MSNP2isp41I8Dvx4G+3n
FUeQhTd1IC9k0Ghh733cuGt2sYiEzhd64NeSdLeqdlOpUNnPgVevj1ha7jdvaNDWSB4RR5g348JN
kHxRIBmByQhUW8pOqmkeGSW/9289nSZ9Wz86nAo8Ool7iLDWMUgFsjw/gdZozWSXDYMOSQH9f2Zy
V6np+q4C2ObZHHjvM5PkneDQ6RtURbwLoc8q7xfJKv4mDtYAJUmmG7A2K1NVpn0JPGIKTShk82DZ
UHUaK3hv650CSwhSvg9282WBqst4V4QM56+uQbdyzzBogIZ6b5sYSQQzSQ9WEkyo4qRUlb//rRv1
NmgKzfYrK6RdQjVynPDTpfnEC9GJhs9eDUJEljYBfJ9s1gji3C+tkWBIrfBRFCGh1svHCC1Vwdfa
a5sKPltUXPWFsiE7RkCgwVteEqeMvTWCfm+eTZJkweGCgCGaucbZBy2RkQA2sN4dLe0BrFBLoQGp
vGWRcisIVviMZbIaOGs1HmA7ELkqEZbUZ1DPg5eQscs3zZZS1uN8eWI29uGXngHnYqwyJfo/db//
Tny2d3wMzOnPk7MnLQqcWyFGRnEHSNAJ7gd/viPeyzlasRijHhvtDTKl216xE9Tj1uGeHZoMKBAH
5dCWHHPMOkfwIxDk4q9aUetbfWYr7yCDJ9riJ/X3SFbgjDSZ4QDWCax0FlAuOcLBrsllqYh2Rt4F
2oWL6vxfdJ+45VG7WSunBHG1funzu19/DS8Qh+m+vXideJkSNhHM+mEbR/Xt5OXAX5ZmteYRm6wZ
WN+n3+zmnkF+NYiO5aXhI1/bWUkBfC5O1kQ0Q+ttZ/8mbidVn5pRHhJyJ4m3vxvYYgTiIsTKINMQ
7nqyvkzeEyMpmgL7AAMpcr7G84tVEU8nvsj82WS5/VYiM/qJVRjknPzGsXmHsShC3ql65KKMCas3
j4JlLF8yXGs285JxedmEIbsoGaKnnTKU6dfRZRTkpn2o0hoyn0I1PqMKgHLZzI6h7yCIxFUimuhF
PB6fs6AvVJ4nFnsKVJiUlRsNR2GoBrfyZC2Dkxd4dBR7r118RvM3qwUnJEmj5O24jBO7tdOjJ6EJ
N+gYt2N00lTYvVYtxIGj8/4T/AKGSXbvdN0m72ZitLfRHf3GR+rTsGqLegwvI8EFoklkaCqEzV/8
U09t3gyudIAthXQErnCzOcrnZ7NyY5Hljtx8hvvc4XSvWaC8nNev//tUpWTvIe1XQcjbUcJD2yB2
8cI2MxnPivCREUH5mEMK/3mWTVx3uU7LWEu/+rHRsATVRvJVlMIsEfSzDvxoAWABP804VLDwzqDq
ygkuuHpRhSRshmTHYfSh9S/pMUeI9dejLGTrmsXXyDFXbcvBv7L47UmybPW2HOFOv0Fms2KxYFVn
53DmlXGxmE9QiofH5gxU4mlTRMdNc3gDRqXqkyrYSQLPD65pph8mn1zcMA/phQrk9wUSgG4PtvNB
J8MXdDGHJOR2ai+x0sv76RC/D484Z8g9nh7UJLmywz0DA7wLG5BnxPxDnGBZ1D+jFaSuqiVpB1J8
enyVlSMvGEI1BCADz092voG7hhvCq0r8GbaH4Djutpk4lIgdCbzJGyAVbV6Kyr9+M6zwWmr0mpSS
+ZTi4I21ZFaUOjIXzGppqhGRIH1xFTnKQLtHzchg/i0RaPfNzwcrZ5kAg+wwZrcX9aJ9bapPDyUg
FiTQyT9hWsrL+5owK2ZCSEIwem0R0K16g1awm/mJZIvRnIW1Nt1kwElvsavgwow1on7Q7/NRKKRC
TJJodpVEb1vteUebOjkwnUvkrUrBebJ1nK95COuMcTRKULLR1AfA01WwGMi6NdKmlZjVESfbPkGQ
vfNn4lw9Ra6Rtm/9PXX156YKbirh0urg996bVAkPm0G8U1eXYDXl6ChvMwKolC+9O3Sw7aI0b7mq
y4WYF0HVruJ3SBDVQ0d2PLlGdmVghQvEoonkVIs2/M3pBvnF6oL/kFo1eq5BCyg3RQiJrYo8Nuc0
WPbHBZIdw+Xdxgh56E/cV4ePFAyYX0bvXOFSm59/MNqbAPXx2LtLBv8KHRyAhK0LEN70f+UH1sSj
icFzdpPYMEjFhzYFKX5GV3yReIXd7GqyK5Vwy/C1fTSsQhKvwej6xorWTRDHG1PX+kwUYXQ0ng9C
MMHfCZRrywcKgNs/Ts/JZEEMpQpipqQ1Ze+5PR8zPVaFiNoxqqPCVX9+am6oueiHU4UsSt7IL6o6
N8oUvmti0t2dly1C0Ez69yUsRKSUY2ersp7CTC/Gv2sCQZWgdD60h/ufLhvxS4YZLOzTyRUkDf5N
tev5OpF/d4rSTwjf11oxMtbP1zs7znXRTJ+euK1Qv5ooOs75zT/7jR3w6uiySfIk1kviE04PPkhy
PHajyx5IH4hMXjdVmtcJn9awX0sgt9wVBi7fVCuv3ksV4usJqJEqQL1NpQGr2qQHRuL1LhGFsoyY
pttuSahMePwcY5cwVqudrqSqfJKXD9XOkM0s57a/LLZGYxaHZEcPB/9JR5yoDCqjxJGJvgBI9gnZ
YUDq038M5duhYR6LuxRIaqnYOr1O8fAFjwymsQE+YPfFnn6AbLLiwLr0CGxo9yWLx+pLKjQVvx7N
6I7ZuepK5FTsHtbiAyolWoL8CKRAE9m96katN92346HIxFqfUlnJQRjdOmNwdewTklhb5xCofa7N
0pKbt5blpsyYATtNX9V4yW9sPs+FLThHjXY4bqzmeCtdsEK0rj0VNOiLyAVSCbjhexWq6PlHMpsl
LeME1KdTfOWV8MpRh7K2LWvwU/oiWcGaZz1mKJcXeOv985GGUx9CgVKBwtkqAMQZct/7ek6p0197
wZKNaJWfFDXNFV015UExvJHeg9FFNkLF6AWgmxEtIX/mGIdMLqwnKDVS/1zzOXQ9Ax8ypqQ6DTOh
seMXalcy/L3zGFrjMi6vkK440Zet7+i2I0yLEn6ozJc4JYiDh2lvvy4Ui1kaRF7M3Z0paPLeFmDb
yXK3yiNLGN1+BceCLVrDZqnx7pcAxqXsrxqhOZVVXg8wfRZWkPYofH2wKrzfxSCjHDK01GhyjmcL
00ccmxtj5n3w0mgH02mVNI/WNJZNpnljlXbXypFd4z00OzgWQUxa+9eHEvDoeSvFYkvXiRz6I6PD
TLkn5uGp5cYI1a8MefxvayZ5bWV6UPY842ToJgvhGZKWYtHV6ZYgzm4xhreBeNPJ8Dk7i7cmu5PT
nDN6HtyM1JsDMX17UOQqkDljw0MpKnqFmBDgOT4auem6QqaWQVC6ir5Cy4UQ7b1gzDKuszDJVvFT
GXcZi19r8+SYKOKUjoYUhkcdVR1SvH4eZfIWiu24iPuNN1agoUhbWzquV5S2Y3R2uoa/DN/RceiB
5gaxbo29ZkspI76gc6JmySvhdeH79ezM5ehjHrCKuzueNLQk97jqOkSwdHteqd3sGoFKIhRgQ1Zl
UV8zzRsluFzNvWwDjlUp2K/OCwc2c1hfWBggy9vKEo4ORYUzwd3C4utsGYnYpOs/7KGc7VANz/bu
WeHSGVht0hzOTVLJ/GUavvPammdckMwczNUvh8Siijfi2iCQ9FaOpLdVf+QyOv2cTLoSQZ5NuGZf
FG/tFAYaOEvIGHXR+YA7gKOopDHnePdSUsRn+oUj87PhrhIrTh6apeI4+eAiSz99yJiVel4uiZcH
wNwymrOkOeVVxmA0ItCiu1vYbQdsA6FetlkhymxaK4iIKJnWMGX3bt7fLprpFxUWULsPvk7ZRZC8
o11PYvFSpPiRQ0VHShaP2VaceIHOVMT9UrVosjb+52UPD7EPc0GbDFC4Yvb5mvMIXsLFC2gLi4WZ
SUkGy1ZcuQTEe2/EOVaNixVDC4bLV3+YpT8yR5zH52Td0611Ik1lJ/lPxPAHIhVs+dHQvuTTr5bX
nptZmUA0lxqb9Z98ODo5g8sqVpapxAyloowWn/c3kZHGR87DkcwP5drOWfq1P6psjQT4aPDGUmNI
GMcYpsRFged8GsdXFD4ETsobrfFfqMVrDIsvND4/bzBmEU8lt03Ow8M35Kb+q8maUyY7Pi5IM25U
Iz3FOAye0a/2UQZX5NZQ16WMdLyzB3LEUQE5AMvHdv/HtnVMkWPLJD3WomWMyG+BDE1mzurMGN0g
QTGH3DVP7yE4hFGKE6+GsDW92qR3r6U8cNaZU+8RM1doTPpRE8Oxof8byyKChW2PkqvesukG6GOI
8jA1Sv50Z4IRq3oFZUY70XAkRLtF76YhLACU6d/FGSsm52vbiQfR1qLmc4/U/eu/2Jep9BNBJjsg
z6QHvtceFKrtQTZxQiEwfsTB7H0q8yhqofWCWFFihCJLkNPY7nOdKbUii26vAEkMvBQBHgUreNpJ
rs846s2TF/xXX9e0ryoQTpDdF9TmYf6UyB6NawMSfuv5F4+SYwMODYHy8uTIywX6BDP6dPjvB+DT
d5S0zadIfk4bWmuFmh3QsWOydbFIuBpTU4cVjM+L6+bKdJq1dJUdU/28OP5O+T2nCzgu51GwIerK
qXsEvIod1OyhrHw6mD0pUYsc7aml2Un2V+YOawBFVcR/+ueG1cyTE5biEpfYNASC8BOW45y2vM73
6HC3bkWt5UFfBJdVq/jEIlxVGAm1vN/weOMQR4BnqTTSwAAom/UfraI//U+uhEmaKBcK5n3f/G1L
9JybzgCPGXc/OHw34nHdkn6iZfLqESniTIdYvdlWVIcl1Czvfoif+sgBTwK3U5zjAe5JM0y67XJL
VEpYfx8zcCRhIhyhtJySBGCDeGNNaKiNWYo735nX4F2TR5bf6c+yhj6DDNoCS1isVLIRnZuc6ZLE
KIyrwOoiqBsy7af517zndqrwHQKKuXTITd3Lil3vAJLlHoplcDI2T1SDgYs8vSKTuImeBarpUDW0
fExnpD34W5OB/Ic/UMx5nBqzk6lZPkvF6g/JqaY4yqT3rETFpRDue4GGgRTNh33RYyFfe8z5eYQy
4PoWYR3VeK/K0sWbpXKyTHRUbPw4JocLWiBlH0CUiPzpSFPhzDxJLQEOmfZ2eFJKWY2ufyMzf1/R
C5HlxcHrPNhZ6Dc6u0GXuQOfe4nR2vH20ioNQP4ZdbIZmoRvVYx1S6qu1qvxCQWpbIfY3C7g0iat
nE1Vn41shjvKxNL7S/yUQb9O+eTgZoEZnSZ3zuOoVbBOu5LvONe5JfPPG3qA/scQsd73MwVJXm9T
NVTE/Qn8U6QWVfiBxm9FxPm4KD8CeIg1vy0QOrwvKkXzAi2hiV5+6d7ZDrc7pbrioJOHGhIwq8mP
+8/nNqyMPNHk7yeItV8sQItwGEPvSbwFnAf6l4xtd3mG2CE4nCq96+wvzBxxIs/HRkD0+KZSHxuO
P9m/ZYkO3fCobGXUzhFHLMPTor+O5Tcdmbr5e1ckjUL3SvoYSUVXvwUOa+kOJRktzjf0+icpCgh9
mML098TMy2Npk0yD1TMJ1MgbcZ5piTIHpE4Jc0+HmiJklNRUR6V2cSjEjz0ioW5K8MqKGthKWNpA
KFe4uQL3/0B6VJ0wUwR8SB92Zvm3hT2KAcXu0Fb6E1ufKBwDSAXPNoaATKtw7On8VUILkGzkI7Q1
jEI7W5D8X+m+cWi479RkXfCHuzEjiDJyXU3FfUqDVVIeRrLX9lO/lcnI5Zf28NZTz+fwxBV3fWLb
INAwWjHZMEGFWl502CxfACrGFaYSh2TiJmkBD4LUtsbYiDnjRo9UMaT7zpqLBgcKz6zG0cV6iqeq
KB6lw2ZekmKIuIrP+spwzfQqxyX9erdLu1l6fse0VVqLPKzz5URxLD1PuwkrqlpkVVtDKkpYdw4B
X7QhpBMZ8BjAdjOkQTulvPaNJubREDs8FSjSHiCJBxcpQmpCAZN2eRO0ezIUIeQxC02cWjEiaFrq
z61H0KManvLI4yXecHQMQUNMtVBgFMUt1rkY1dAvZZfjjuA8Syrqnk35N2rk+4MCwAHY34Y5Ja0G
nBGKWkh009nEuEpPzvAGoA914U5hZsegGEH8HhD7m+Jf6KogjFrDf0JUB7vrzdy2/LVym+z4s+i0
GaMcO/cym4iNsnAZZ9xg0FWQaLp0KhMqTBmM2de/rUZSW0Er00mHZMnlLKy742cKpc7tor5zDGmA
xxIVy1Ne6X6SUSPjXjg34FM/3K8PuzlAkV+7LhqV773Rd0hGMbHHA8eLJLNsbEoWmJ4lIs3FFg36
OV+ZVWlR5Trewr5ZDTd1X5DtuvvjtFlIyK8pvKX1yxZZW5Ju2AjkkLJMHFz7VjD67xofZjYtFL6I
rNpJXT90HYN1TUN4+/OjliXJoYluC7fb56OzQ5k4WzgQglquyM1BDjiXQsF7CkI0B28qJEyrbJuK
ag+WB5wdppvlTQZewV0XDnAYSCDdSMq++pDSWIi0kTqrT5cv7vD8F05fm2MiwrwCh2HmfddvuSCP
SGv90iUK8/KmQMwljHum5RMrBbBez48zkzKPISWfGUY+NDrQBuqVmhfAQ8oDa98pX97Va2MzJIcQ
b/K8e3eoCZjNFfQVl5r2EtPGdCDVA7BrgtZPKsjLcxPxnHFqc5izSUGJy3ygkUUnoFfTlkGOU7/b
do9NDF058QJgRzFLXbjCzXecdDpWPqNGwtx7X7b2wGkaJN5odcOOITIoYoSS0FFaxmgfUBM4K4eQ
4zgTny55LGWACXIaq9Zf+4119b/ReFWRd7pEYTwV/82UJJ2BdicM+DIHnzZMJb5Lc4Ukl5meZNTw
G2vGA5blOB4H0jvDXe7LpM97kMZ/7Ovln+YAEN72PAsKk2O91RuHDM1wkFXGsjh49FzEn9wP/4Wh
LnISgOokyV41oNkUURsrwqfKDxuXfdPaJ/gCcoCY1on1HtNb4iQP+2w5UBqXGuAu0Jxk1j/V/cQ7
/9FafnOg0KLFwue6uZz52McW+Mj1NN7cgg++Q+z5xr2hNOHzB96JpbJdiHa4/hT48qmoAqib8eoU
Mx2AcdT7xDB38UZRmZKSbZB2pZQ3nXG5dP9B3P4JskpyJCaTU/y86JzW9KnXVJInUruxv7bhAGu1
zJS+uifqtmctY4MxGcRCazC4MyfG5r+pdwZIRIjot/OOao8VU6m8xuEvqsmqUBTFeoqZpoLZ20oz
yLcoC75qfoGs1Rm4/JIvRIwrc+jBaAjt6nJ8NR9REjxjPqniZGbMgC9LOu1IU58kpYacaoKSiZRa
CBr9PQufFBi/ty9FpoF+eLBhZyCc4bKOKfXyxo/1LMDuEej7tnAw9wYZl2dsyfRRNuomKrzuKEhe
aWP9latKYUU0B/JDIgBj7pIJZTY/LvUQi9uKH33Cs/98po0aCvViFoAQQgTOnSVUQ3xoiiAprpMW
TC7RWMYegaxcvPLvCns2EZl2ycAlwYnEZQSHLXR9DKyJEX/WPvNmv71/XwlfNtOoZUi47AHNsXC/
rrqvM9COK/237/343BhR7Ivh7L2duEfLZK9KUv/pqiZftgTCRpA8XmzbwyA+/FbOTZhYX5YKZbuw
xZskxsJim7xT93LgDWcuGavGcbaswv/f0GxC9yAftXZdsKJNZ1G5V+uhfmszs9AgD+rd+Ykduj/k
chCXyfa7QfBitKQkXd6JfhjYXK7ftJlAXjL9tCprISrWMZzootTnz70tMRAr4cKkT0E/6BJBIWUx
Js9heNN5eSWW+Of1Ym3ojQxyZ/qqbVdPodEndbSiDWwsUJcOACXzVnOKWDaoijAxNnKPV/nbrZrH
YPOnKzgFl6WwiVRQvIhKctBjXnjALr4pHwMwRnWV8fXcUngGqOa/dD/JockEDx1DoDpjJKBGpiBX
73H0UpApJh2tSm76nSLzQFRsiDwb2jLSU3n036Ju0rrHYpleowSDBhpZfFuv3ROvy66bK3FyH9AH
IoqeO6dPlEqbMRZjyZ1BTE4S0losJ6FpWfR7FzApVrOOLKq+SZCDwLerKuUmVcS95oC6sXTFHDZF
fDsrs/JEFOEy9NgMhbHXjfSfBjBmiNHIZz/gfG4Hbi9+B+/zdHyJYbMxSLpqtqtFOGjAt6bh+zeZ
NPwQ6ASSBnFZyfwTe5++4tpXvI2RY6lITwQAV0qWHLdiFw6wn1E1p31ukVXzRRT6VPbs0zck5YEG
5vWU1Qt+reGJbdJC9d/UuJzAzXML+JJ4kO3Y7tLxsxrZnJs2uP5/FDh0KKGER2eNdIipLrtR4xRm
h+U8IbZEsh81+c5lG9WEuYSk7Y23hIGF1+D8KPWEF7A7/L34X6V+3ryb74p+0Xv+YqqXSkOAwWRc
mvfEgpfEpEO+IiBEfk0DsVoO74MnDANqt+pgupY5Lv81jvwzS4ANxoRJfGkJuePNLuB8jq56/Eht
Ilb4rztV++YhCxWP4ZRuETfH5qKuQskRJVVnuozRYxnmyk+hsOkDe9+vqcJKm0QZcfmsitqQIO3z
1RwWyh5isF2RGgfsF7oL5SXkQtHbrvDUH1F990FmykckpcApHfipCO4OF4OBPKf3PgVxgC9QVLUT
MKzAoCoMnJLs36e5gOXyQ8pc0cG+5/CA/ol9J91U954XnUaLLLzUxAvwKlWjAX9kZksf6QEYCx5w
jjqgBpUVu/sa2h7qwdURdcKALA6PpwbRWQbPR91n9QTgsLDj/DftkxpcgehJJREmL71eDdWy87rI
BkycRwsk8589JRcERhi+ECxMKyPOJTesy+uuMrRZVfgSFKRpKa74qV5DrSnI7unYjQJzRULmbAcE
6WIL8ftEXtIgfz84YFd27kYasWwGH/dt3+nn4Ev+93z62/ez08/la1FqyUTlEzwxQDNAv11MvqHd
SiiqSH8FjLvoCxpJEOel6SYivqFrSenrwIut0kEbURx/o6yANy0i0dhO5XwsMH6krcnU9DP8NLLW
WawIyoK6PuaMavV2I7kGK/U2Yxalm3Q5K3I45oJiWu0LriDp8PktSP/QxxttEBIqz/yNWUHLDNvr
5cp8R4wFaeYw0Ur5Tiql8LVaX6Fzy5pqRev9GIv/RdelETr4cknyEkI3C44co0+98+3b8zmuY1iZ
LSgQ16NRK/gq5ANPssYVtOzCCShv5PR+8T/dgG2DRIgWKHX5To4Oyt2x4LojmdHmma1cZ6wvyIFv
C4BiG5t1KOLDr5i2ndbvT1zXnqAaPb48kQMUk60u1+KOy5TPym4dlCAWIgEU0YbspEb+CLxt/znx
BJxC2+lMuuyt9WCKW6C9nj+NGIzjLice3iEFYzTNM21T7tKocGyrAd2IDsEkF3CxB4NFUhoRxAua
o+3a6skFdpJz0Xh5d3YzHR1a29Pe4aU7U94NJm9sgwHnDkNHS3iO8ADltwgwonSE3yGNt4ui5nso
8epbl+dvxk9HlqkUWS0fKWLm9nKQIPvj2YA0TXhU4eHLYLZkN22B3/QH3XrncWGIvKqGfDLGIPfg
i6/H2Jnk1FALM9sqkTpipQTeTe5qoU8EqBu8pbN+WBXmTYYbav2JsO9tMrdaG7WYXSHifiPYMrmu
wmK3RWeQm5FfXpLMcTW7wCLtFnGTTmmMuvTACs1oU1CdDlQUPVpM9qoOedtf3A8o+IoUdMb07xZb
FH74gnwqzvwFnZTc0x/cIIOPYspQ0KlZNFYjtWvE5lZPjuVOrR3tQ23jemA4cUdFMfpGzIMwRJbq
lEpzYcmQsWaOwTpAReZcnN/iXgKxOD2gQx8hvY27RRTD56VwI+rmOvtN2/j85UKdWsrzPNsrpNYA
K0Y8Ap1ZhBm7UMA4wMTEghvj+kxldL2//+DKzp0GkfdTtIMADTyjb2C+ckZWxiAah3zgNKgiFl6P
J3e5j54FIaudF8HssuMOGTNefjWFrajQM28pUutvEu9jfbdt3BOY5WmVeUDb0eD4VFB+hoUAEW1r
Kv3XBK2BbSQSOZ9rEjLBlOVnldk6TyB46TByRBcnW+KybX+imJvhFqJouejiaSBHHxaWcLqijInh
CmMiToM6LqWA6rdmnVGGHegkTU2X4V3tGBqvQW113hRs79sd7vl7eTLjHiMAvMgR5M8eUl6+vrzS
/obFHFsWF8mcIbi1KDiLeVayvnhdMYVOSQHGKOgGccEuJrDSLtoUQFgYOJi5YjJJO6gNx0f+nYLs
UR81cfu3EZnqVJ6AihPIJ/lVDi9eXFdYGURblcBu5yQB/uuJg3hL0X6sSIljiUH5OEYAbDPaCQAq
l1JKFRj/5ME1M2DL1DXcXMcj1wXmu3UPapLhRpmnEo8/cyabdl/GmQoiKSKcgSfREVnBm1g8/Q/Z
9AHbZJFbNuIYhLvEHCPyYOG14l/52rZlZCS9X4A2utxi3cAEWtKDRJEJ46vP6HZ2c+eI4xgjzNYh
jqyLN6j1Kp9MrHoVAjFTVfrUth6ONqqNv3li74aAMe4Ag50+eLn9Ok5ZMVbZdc3cJHrGAzseIxcq
+oL3zTUuQZvB7lMmy/+dAklsLbwPSFu2wX1mPVUG0Rt8ixg8EwXNVrRIbU7UjmDc7GmH0gAmY37q
PoEUTqyoxu22k2bUc7wV6DzcQGjQ8UpNLrpJePb8y6qsTtbGyeFxato5JB6KU2vlYjGKQOAx1x9S
ck6zDInVeL52ei1KGx4THUzF2tw2yNB1zF22EpL5zPRQC04/hak53RSvi68/J7R4o5sv6iqVfIh5
w+2Fs9pBT3zfi7HNBqV87mUgEWx2/XaLz0qALtNFqCe9FJGybAqxDAca6IHGK5+JRcm3h9r0YgSB
EE4FkbU+2ECUgTYyk88CK0EFFiwP8l6omNeUGMbdSOYFSwzsJfjTCCjNwXMAvpaF4kLaGCMtoCEb
Mx6tGfeaclWmb2V6j/f/9M31eOUK5QMXPJpAwdjjs9cfESETfMauGK1s3djC3KDzIa5yegT67PqQ
mpnuvV6sSIa4nvK7apx7u//5wYzfPr/Y3Owzii6PL+s9ugtazroKmpdwKsw0pyTwJf5iV+GX4Frc
YHRrZSCrKnubeacKz0BnRbOeN7ty6MzHse3Yj0m0Yf+o1WnnEeazIl6OiXFzndkTHu5Dg5O/YapV
j+CFvf/W4l234gBLn78MgrvDnYNiagUtZLFifDPzFUT1rwzIGZXnw9Ra88QksImqE7//PmsE5w63
ZB6TJZZ5bXrMLjSdERIBPiKaL3AD8zeO/hl+kgYxW9QyG/AcAkjuOHiPw/kCaGuLHzndBhS4+YyT
PmrLYXstbwK5EciMaU3SqQ1QSZPw11wlAS/FCw+389I0XSiPFtOvbdzEibthpDnr10wD8wk+0Htq
h5Dsf28b8tvDYC6m80rh6Ic6A/z6btEQ8O5ewmhNH1lBlRl2RFiPkEvNyu80QbqTpgDFzZLeWQo6
57knUrQ3zbAJ3WhLuDyGtwIeULseCLdrrraYZGLM2AdHyTL4WVm7+r4FPXN4JRdZSE+R8KbnDnBy
gL+PKIiyCwPpaI7CJBgSoAF/3ubOnmWsaBONrZ+txjmoEtQ8Hb7L+zJz6pBQw9/hDZTIX3uf3U6e
mLBi9kx5YcH39iFoCIlTYmkp6uV3/WLpmNcKbIxJZwI0/PRLKPamNIUrn6ajzYV01ET5qduuHNUA
jAXPcBj6BT1glU1cVCisG1KtX6zsN7SqyGvS913aXmS8+kC4PtfqlBb6aa5HpRIk8VVwc1ccTddY
OSK55RT6sFZW16FJNhn9+AmDTt2E2mZu3hIPxCkFUASam+fYVtGl3XTZ+4Owhk6RgJRE0nVJfz21
eraWeuOkfjIjIHeHVT68+TvhsddScyvSQjJdXfDY6lt4+xDBGeig3vefv1P2Vkmu1kZVkkRgmLIu
ykXnaprXDrl3qxcdIo06lh5s1sqldFq9xSdzdrk43Nav6g/zlbZi11MR2OjFVptbkA8N/Tu6De1Z
gRmFe8CY1SNMDp1dmm1IDFsf72ADWOywmq1cvl78G/8OWx71KxYt7PIcJuW4GOGb72D966x7Os5m
vva4z2nHAGsplJwxwbHdCLPqXz6jtH3c9UDRfyDbRGem46U83ehW+TXT+Qt4mTda1OtXypRO8iDn
YWvhHV3PKXwY1tkDc61dPA1d853lVfojkLAjWkXLq7pcjJ5uefCDNssh1+Ya4ybDw4qzmKzitDNg
6gxDqd/2mi/MJPEFSQtV81trs51VMCWtEz5P1M7Og7pIVaJDJvMEAVa9mPO2f14On6nvd/9YqvMm
hyitQ7cNSixwdVEXMHe5lfZqtECwiiY3a2w3v/j+g+wTWonzK4z807a3LZMg9/EwWMc6jAxEB3we
rNC3WrhgI7aMvdBymBrcelt//a7Jo9ESdV3VFsG4BXq7US17KORHL7N3Vfs60JLeH04qgSp6673T
7gNYi9zLiYyGFe2vuElNgP+8TddPO4kIu/BY+8nN649WELtAbut0vamaYgY2Ki/bj1VmrRYiwBLf
+cvKMZt+/N+KkADGsAHvOkkrf+iHZHWFjz9Zp3jxhvLWZfvtqnfGWpYNueZBBQCLnW4YklU4vmOz
aK9PajC4LDRLbxhpaeRVKZQBdUnYAm6D5bXgd5Y7oSZAUmKvL8bHSmPQoZjnMlQKJH0sB2XNg6WE
g8tIIBtGtgxEuDlaLMRCWWY7xkK+f0Y1C3RDszKD7fnqp6TXl17+yUNGFWkDtbcsRmhgHs2RNyxJ
qjji74kSvWCE6hUGgP8VIKiFUdVQleaPWs0GZeJS5ZBFrIiy6zUpLGWRXofCXMDQVel3RH2lC5Tv
GLmKwKD+HoIfkIFRw5R+q/oTVll0XY2O0EBx8dDsDPtRSmHts3cy7EXZ5RcRXqlFssT0+8mJOtMy
s8Y1w4ZLdImcYWSd+o4XqJYzyLQnMk4QWX+SA7NlQvSBTnA+zOjQCJeZj5AfFCxehSWOjU/uMpuE
pIYyCDedxr+irMluD9xZkRrIYvBFyF5+qytpy2VG4Ipsuk/XFv00pWlHBjfpZaqpkI2jcxEsm7HJ
/d+Aw8neFfId3V7sEqmgQh5lSiSsttKInGrEgYmRABNsVwi8eK0Oq0GNIZf25+pnKfRN6jF4PklZ
7ISje76aU5j6jpRZKL+dsyBcFMcV+CTyuT2ujPtrsxGCNBeW41moF3fyBLbU/grQboOM3y8lkAKK
E3R3Pom0gwbw7+SyHIY75IKtefxgjE1HXSgm8ourqq/PHH04jTh5gWxmmz78ESfeFwValtiV3W5K
7wDiddEZ7ZOf+RPy1gf38JjMCJNxGf8fRbCrByFuAYVCw7iunGrdR4SvxskgCrgdDSOJM+DfU69m
mws7wv6hu2G7COSj7Wk0uuITPxWz4Vwl8rpjP2xIBDJVGYPRpf2Ksy3J45/nw02ybA+q2U/s0E7f
JxMqkAh2AIWa705RsaRUo7myxHHEkHrOfgamyIxPZ98dIbynjqYTcatRdcByObJOQRAqpK9vVeum
P8iDl6LpCdEqwsaz3MCJLOm2bJDXAgq5oU46gEy/Yqly8VzHRSCQMRkAuliZX7/4WfNAO7nYwaJX
ChlM4SPAt6xhgWCGGnq8sRLp/TeghsFGYCwRCgGaEmjFNMRU747QV/bu2SPp0O/WfThtd22jjArw
sB1WJrjfHi2BVpsY3aFETZoCCjr+8eScgkovgARFNvxqNln7Qe5TJZFw/nnvJAhxUTy+Qxuj43Q0
BN9cqC/DwG2OxWlMVNGgVL63WEvzNnZfk/mPvzq8DAlvMLPLpgzQ8nk8jVS7PQO4v0b6NhqVsuT/
jBrZL1sm9grWbEFtvXwZlfmxIHTCfO2Q7/oix05GvF/pdS1QQUzggph+1H04FIdzko3h74X1PGGx
294M7vMh57WuOblWU+jseJCN+PT7mOm+nxkxH6Qy0x5bPKPvTENi2JnghAIXGKCmL0nNTmRQddIv
RKaM5zWcXjv5cJlavhWbtThWn/kMLQkO6lA7V0vg1iTB4rxusRubWKRkdWhzhjALynlz0ip11VKH
IeCCK/5ORJuLjumn3RNm2oklgVhZCOoQ00FFjGesyUHZxQ7pVNT5zlvJ8bqucqjnPLL1w89eJhvN
6NO8ENB5uQ4CuZn6op7FzB/thttMYzkjg2VyGPY+tXh8/pbpl7tdmfCLHA7UuZGiM+Q7rkeYeTWI
AXu6C9hTzCC0u/8GvDmxAGPCF5thweY4tzTxmHyJaIrLzqUDB6Vyi7rDqWE7d1W2Kmyqev80V7KT
G/DK6fMKGyMrddgovCeICAnbprYkOwsyTHNykiiWPTr1Qx3FfEnNyUfOhjDSDszxCL1JqptkPeZl
8LtkW+hLTj/IyShINC+TpxHjvAGo1fuwTcuvB/zsp4w6534Jf4PPBnr7GlTpu8yFndd60XyhLYXa
2cuLtBJYIPPHVRhoihx+t318BZ3Zi1UfzfnXf6HUEuZh1fSr8xZi7TD5WKzvnZb4aGjcong8n+j6
f2Vdh8p3fNYC4UQ8pVOKnRbFPF6mj/Ei3UDvdoHBnTMZB5oUeMD/c8PjPZM7xNTF47k4j9nD5tYH
PCf3spsMv45DP026kZMZfo+iwbeDaRsxpdg+FsapoZzRHa5Ets03slvsaxwwcZoIahdfY3NjNHEo
X2f423dZ1SNmrO1UaR92PoZK1dMvc0+hhJjfJ/5kdQRRWQHSZqvU4NjoQ51ojVAFBnh6zZ0MZYc+
zGyOBX6Nhj5KsVOw9U2vh5ra7N+AwFTjresxFYkZUKf/yDGIw5AEHDp1Hl2iIgoKTn9VJGT2ZvbH
qWBGANu5PlrW9PUK5IBEw4I+/uxuTj6uJ1FNlKJNC+c1qdFju1GQ1Ecaj1sgZX14og81BLjHbmF0
/TrCgiEGdAOP/XdYpV8g9g4Hgare2CnAKYDFfTmZhJKjpWAvFJ2Fagf2DiDTYZ5lqofYNqHp21HA
8W7pJzo2MRVjr9cLn8TGGQKwSVlUNespp+PwPMTWZfhoGdigft2r5BS88geIaYRrhc1rXjVPL7XL
qXlY6wQhenwbu5oWMBqh5ls0QwCMcxdtpt9IX03PwnKzRuSDtiTgGCRlRWDr74rLle63hYuLQQXj
q5Lv5VYBF3rz3okFlnaTGp3ZgUQzaT7MHWb38NGSDHw2K+PRB9om2U7CWWfEvUE/hSFVgGcPDXYV
H5/WoiExGQDnqprUgLV8qI/VYToqdE0pKARmVxmTz/PTq79HYebM59q5cAqcJ59k13809JR7OkEE
fezl3C6l1zyRRLGrsIZWpfn70vl/wMSrV+V74eMJxNHaJ/syxyEwXhvcIOEta864yzMCtmN0AO2J
liVzcYW11KIxZE/EYKorRPcC16GMMph8tOPsLoWlvKeWhVbDFMaAtdDUm4tjj6XT69Q3MAbFuSc5
jRhAU324/SXmRGTh6OmzPy8M+mRaFmymGCbr/eGoii+j1oJXGMH2yCoVJ+55v/4SkQdKWl6Haik3
ggtJkMTmIFk7ARKL20opEysuRBdH1nFnaf7cBOA3ESPq8xUn8UUx6i0P2DtCnA5NLnF7+AVchTJ7
DOCANkJUPWHSnoW+7RicmRlXok+wGzjwe44v4V+dcsMYGl8fOVdD0WZsmNJufn9lshKZm2xrzc3V
UddQl2nmEgBkOSUk5hl2Xski6x4Ruas2jG/jjldQYC1pNNMqgDU3wvqdnYRR2mY6m4qqODed3i/r
oqPcO7YLHq50IT5Sk5+b39gikRBd2TnOnBexisAXJr+dafNOCfHiQZc2zL/Av09diFnhGYc3Ep5p
/q1osXRsYlapxgWnj7tZwJO0lPGyHOKLsrmWYrtq1iBlYZOvkB232YqdpPpN+Yim6PeeJtMuZluf
WsdOIdlu216tpAo+Dueu7VsLLTNFn9ZkFTXGun6fkRlVtvMhGDC/a1z+SC3IjWyxK2UhYgNOhP7P
F+DA4hvIZv/riwu5wW8sPPEEUBBAWxhTf+B+TpPUB+jAFo2Y82PZe6QQgtiCSEb5FXCjhXwjFZEj
J+YmnYzYqusyYBOeip3cl+l4/SwngZDMTZiE4bzTskN59a/I+Wp2OxRch0W7zL1FaZebKngKZ+I4
SGKKfkH/JbquecZZbDpIIjF5hWS8tjBSSEQJx06SGhJpFRJp5l1DT3Lsj9VZe09t0WG9i4DQKkIG
LezQoM4jUG6V2khPXVQeCREbteDF/y5LZ2uD0/piapFQJ1f1pJVGRZps4/E8I0Lji67AI/KA4nmS
Ou7rOO7u2nTZpzcThZGBtC4BnHEGEXEZWqdEipbzsCqnu9sWHku/erFc6xNPrtoodo/5Y9Zmp9hH
qgXc8O6Sf5wsiImR5P94BhiTB/IwThaiq6VRj+5u8UIi6Kkt2Phf4XurQmFJ1WsKtViRYzebkeIr
R/du8aSvMEWgmaQ+TqZ5675TRCHbr4EgZuQI/xsz8mCB7/Th1USJWqtN0MzriKF1V2i8mOubTw+y
KZOFq4UuOcNSDiJ3bsPDI/neg8u12rVDoyOyKVAgzNTg5J2ULWuYGNwLDf7tYwXk0BaKKZkGYHcs
BdqkPAFWZwbZYyMyN/W9P2yTj6SlRqjog0gImV5Qq4XlKM6rzdBfsgNh9bUUbm6wH6zeVeiGcPbf
dcgfraAZiR6Rfcyq1gZSQOH99yZ0I0VnGgelpKESvq/qyZQ8FNsnMSRZnA2MMB5NRW7LK1q9K8D4
6iM433lxYk+Tx1Un6vUxQii28xI1eHEeb/D4E+spjAembMhbtfJzozIXap+s/UaKWsX1ehb6N/5M
Vg9WkAW9YkNkcI+IPeus24ST8zZD548pxRckvw+DStWOwMoxaW4t/V16GAldgGpGSB4WDEKACsNG
ULsw2zFptKpa07ZbWkWFE+XRqNjasbO0xbKEPYbeXNOi3ewI0KiNMUKrfGjfz4HzjtVcSjR7BKtV
/mMSnIPhKT4k26b2S9wkhKQ//dZ7hLWumm9LRN6gebrKe9kvFdPBizTwmL5UwjKcX557/HrZiNl1
U2UeuRXojfmM2Xo3WwYW5GiMVZ4+ctl6RDmXrFOefHMnTZgY3O2vuQAuXInBL589+rknokR5u7nt
AoZWS/2cpMXbSFBA3G89ucZari6R3nDGkdRf6SRDyrjnQouxyQ80CWNHCSqHJ2q0kpSdNOd5VvqH
DEtr7Lpsq8jpdfBpgsrf3SNQzBWfnIWPiBZzhr9DNmZ7N0VkstXq+EENngatXySjv+P39xCEAT8W
ab5cWZcVJLxEMHAwj1u4smwCAM2n1+oKlwU4I4kHhspV1n3TQnG7kFMh5EY8ZKCFRRP30YUihD98
qti6uDHHIg95vGWPUaU1YyoZqQoZ7mzP8qgSBZY1bVUgZ3k7/brR+d6Vk19Et2WsuCLxMxtj1S1J
JpABn1a8mRB8XzgORh3wSrfVeaGrTW7nBJO+MU5ryuPUxJ5XmQbZjTPmPkhlt5pgZjlezDcFPsgP
rk61sFOhgziPgcdkz9RGqbvy3SjOukZpFSe8BsXgxC3cYSKPG3/tPpoctthjDhujMLasVT91RxDZ
xJjIuNFCknCO+ZTdtPWlEtr8msjfDwdrIvPToGwhARzThmQ9vZ8cAcm7vcS4bBpVHgThDj7ox5t7
NHxoz4rEqi+5NGLTfWReojA2SXuD77Iqqu0xpY5wo1xx7ufrCdGzWjAvOvFLCXcej7crPKGqNEcS
N328swcRBUwhifCVOPY6lvkRHTFXQq4GNppKbo41CzcVXV7HDgJ0g0sxLB2EqMpXalxCTzIrmtrs
Trmv9GAIa5pOOVvMu4aIjSkJKMEhwvMqAFkhWKyJOp53gxO8wo6xDJHTFu6ane/Xu9ZKtYkqlN/s
yIqsATVB7UhMk6uUHgeY8ewNg9eGpBCpfSsy59daLN4TOGIzCNuHyBXARP7cXNvuQpl0a+KZJpsR
EdI+l9BqL4VV0rsvfYxOD+9jhet9F/Cg53apJCc/hz5wborVegJ3o8L5tO9csna+MPIJf+EJyTQ8
k3CzvvWvwnGvZNOqyRSGYPMuPzxbXQZuiBIat8NmOUiRazk0VP5dR+8IePsEuUUoV/p7QPNaHg+V
YRzUzjhVv4+KGchamCQpLN+0w+g5Ld6VBFdvgqdnOMVuy6C/gZOwc3G+oxcogKkF5qo90syoOEsu
tXwZF3RJw3lqXz8lfWOvEb5V76AqFLupYdl0K10yqNKnoWgG1ROpbzQxoqqIGW/wOCvCI6ZbvZTV
6Elufubw+SjANOiYI6xzqzi2yr8a3yeMsk1NpUboS4yYAT6k6BGt8nJ7ZwnKdIw4I3SLTlc3YNW/
BVVXndLC8EWomlWnbXhkHwzG599Bs46MNDFkbNvXkDKAgvdzullRdAVJ9xjOD6HSPN7HY1laZM2B
ZPxMDh7M73vEX+mRaXe0M4EJJj4EQrENXwt2e5XAo9fF2zi++SnGwXhCyFKQOVK58DbJPHo9VDJs
fyJE7JAKPf49XcuVLyD2G21UKwX9HRhQGd1ukwh/czvcjmsYjwjpwvpsjVHci78w91+g7fIR3QxU
UrtVKd64Vq8FcNwIJAd9k8g5X1Wc9SAXzm2gxYtcaC4XZ3iNtVjxE44xmjTjCOD9z3Ne3Bnv6j4Q
rgLQi7K4/yrAt1ysJ5SW4J7Kt8UGQc3M0ym+ok+hHQj9LK2W77rkpNR5hAX3BxY4EffIKPC4iCI1
1RrXovod/tL1BjROo3fr3yS5rur5yzPRJHxWHe4OvayjCYXSz0ITRCcscbHiqmtRc6jo+2ZYtIUw
G1pMof+fFvcHzHOh+vtdJ4CWsgcTHHJeftuvNtyHrK/qchAtjxSDZZuczqW79nrfS9A6Qn6hkgLx
JsC888e76EwYU8V18esGrEMvFpgPAx2D52CjU5j5Y9Ce6v4e1rLGlM7BEJ5Ensyk3g0gpTo3WjS7
cXeQnuDEKsUEKVnazUJr24SNRLCgtZGlAA0ersV0ScSUMX1/Ryix5+x/z3xRKobMLyztTlNPlJjx
TFPFu2xKrpAYoRSyjwy1s+TX1jnO1D/EReNW+1rnVYkTZaRpe7/9fITs8+XskK0tFBkfWtk8m0u7
GkTPbwUUairMuB+ZqQAlslBnRO64r/ZQXb2PzjVnUdPmYrlyfiPOpynjQpjf8elMsO6tZQdTt+2v
wnemYEEC0OLPLmEEnI4iSWt1qZQjtzti+rdxPg03ElvjZ4I+V1jDamJLsW9bURXltY2//9S1IrmD
iPBmC71sFNcM4td1+Gmr9RTl73FnNeK07AjXYVD2Hau7NVJZJMTdUikVK03JCuzzMaAr6I1cQOsy
GclD6WadUOQPKCpwEFno/1/vkHNvuToHzSBZy1LYWCCnRPDRL0Xf8vPfTBufmEGU1uysbxM9/ZDQ
sYoa1m4iWSDXHjNWpjJakw9RyTC05D52jup6S3Hi4D5vSSZ839xHlCTnf4xExiFuoyVoY3JWPYLD
DHts6y/EU768L3DUkpECnfBw2X726+E5p1pHkYDJ3mSZEzD8MCCiRddV69/yCiuROQEZsg1rnlVr
KdUn7SGemESw97Uone2fKee6w5/UAn0Q7M3Z9Or5IorQ179RxbextZ5tDDOGtm9wkCttZvJ+EVc+
FcyKDQfjLRwxVukCVvfCfJngDL9kzXdR1lyquu2qkfVF1E2XYIMMVvETn2alHSwSCZU34VkhlDhI
84k7EdVnbvfZXguN8W9VHz+dKgYT4Lg1k0zhNWBtMNR2htk8x3f/LjUkvesgcdYzOPrGVmUE3/sZ
xmbeETYfbuledwUrn5UifMzy/OfTIhxJeAiFiq/D9axEzNztUEgTKX92nX7EEipdiCX/3DfohBlg
nofF5Of0GVXQN0zuAqlDKWRtxl4KGYpPsLlFU+H2KpKuWqOpefi72zXl+ayoO+K7ilP1PnMtl4M7
AWZzzAbhSF6Lc0qXoLgW5qGG0yE09zJBY4O64npijh5TF+/draFLn5TFn16acpaMvQGkeiVMasxM
HatnAfW+dQCUYQfQoQOqh2eZcE+04GLs01zklbd7RnFzNozSPdmIRofDL9LcRVeZPlZU/U0KchYv
ptFL0P7FlMmco8hT3DrWXZTObha9+VW0CQO+quB1hxsD7Entq8v7ZkD1yLTYuu1KUsHhjKKIAV8R
cfpTAe/HUq3kEQHhjhpjsnqk48g2O/vPjqNrFtSlSh0HoU0x3f8J0CpZoyu6ou2E1cHfts6sntoM
pmlH9jBlKRMMLSvbZl7r1gF8aa3q9YzwxUrvIeDTlF/+awG3hm7RJhc/LyQ/GMKEgNq4PfUVDyUc
Et0cRnzJSbAPxndSA7+t9/D4pWL4ycb33qNxZsfHFSVzHKlBN+QsKU54rFyiY42hYHpNtbeq3CeM
qGSzU98XabhGSCtSi0eS+Smszv7DAvBKDclcfiRxCXQk4TZA/zXBRGmgBwDZ93tExOWe8mFCgwqq
I5N8HcgAJ6jqat7K9v8G8RExN50TeqY5oshZdEfL5ro9eCrbjOk906UGDL4EWitsEJPXb2xfkZls
XKqB+fR+5xT8glAYo6dEepkAfBcPeWQxE4cYnDoeWSq3yCPlU9uT/qQ/83nN2bWVtwHDsITJ4yCT
oktGWNcMiXdbtAz0KDKuvabxV6XDDZxXQddt8AvrQ47HOd+Z1MjVewNdbIYxJdJLhJvhUZpcgFAx
YG9VAibA7k+nVt60K7OnqW3ZC8tO3xWhgu8dJjvDxlns9O3v6hRD49thdtb2D4oApER+TW8PgcV7
RgOrn+f5EAxlLkn4XCmP8suIOD1k74RusdtQLMbO65GCnAyLgpl55UMKN9LpKBPfsGhh+0VSiCgv
VpSo9mt3tPqjUFK9JFPFwedX5Rv1EvtGyjgG3qF+RZKPTL/d0PXChdqxKJopttgKDqwJpCgI/qxE
IvGle02wfN+b/CCEh48wrRNj3kRA9xwCI2wi98HgdabnPi0xNs7qyFqa3sSz94gBlMQ6r4mpT7mk
BLaFmmZB0MhIFPXzoBb8my11pleZqqutBrTN7LPFNmmzevawG/4IC6I7gY66Ix7cHJ9Z6roy0TAU
lNPgnVt6mzJIe8AqBPyLTaAra56NX5Uzbbw238wctrvYlShL/gdqLC2qs5BqEkcbU4GQvlrHyIbT
uK6jB9auESFvMGIY9aI9n7uSBUehG/aqT8xQGXK8n1aYtU87KdWRY4Q9SvZCs/uJzU1Nadfetz21
j0a0I9pwOumqg3+91XbMOCyJF4fvbHYeAZ+bxSMZcQ6Uns/Mvn6Xt09vTkhtnUn3jKBBR+zPePcK
VuZ6trz6OIZGgXdwgzZv7yNJOriFe3i5Gvalc3DbW9TmjsjdS6jeDnbHSH1Xb7imqadW7287BGfw
lccssMUzTjYKwmTdu6zH23TOWokDurXSxjsd6TqRO34kg044ZAv2Dr7vn+RwOIAgtOlnX3X0Ud69
Ot1GnAeTTDHPfqt7+P8hNB84Y+kgF0crsxlatixJjOgHlAlwwTRQhDQelml0STQXzXGzgjjMom5v
mNfvhf4Nca9RGo4qCYyYCrwEyCCVoas3TrmCJug6tf+ajAf83wJ3n68fCwkLyOpxqwU/pPE4y1hn
by3cjZZ6jb6gR+ejWJslf/QhX4sgXGgwYinHypbs59281sBH2OyBgyummq1z3V/BXAb2I+cQY/BR
/oSUm4fMG7dQZ3k8VsHclRhWa5jv7V2ZWm9y+vyYmPvwki//g4Hw2Mt4vyxfK4P9jI9RbiXCKT6Q
jCXxrUw5016SCrjoZ7l3qlyz8ukhThFPATuQPCZNOdPehXOz6U5hxamgV8qPaxduyaRyVHe3mL1S
8zdg30vX85V3oIbIhHqg74NIXPxNQ2pzjuZMSaDH7SfA7kZukJQ40J/eSAT9XacONvkbYbL1a/IS
fQF6Ks9T89iOF5gH94upeZ1gWL14AuyuVdPTu4jLbEu4IF9r+rlE1eOyUgXIYiN693zZf6IrLH8X
73fR80iiAtfcTo/fW1jnb2ju8e8pjoPquSonUgnzGwI7n96wVzgb0CR5P/B529iFbJZgHXMz4l4T
vIKBRILibvLXRoaIG2U5EG7jCnI8jyCXVXHUREYdfM3sRq+/oOBWS425Xmo+DY2LhWARey3MegI8
LvcYoXW/K1SgJfATT8S3m18RDRm9+xX33qz5T8EGfW3FLvbduNZxGAqKSbucwqhwl5LJCRC7jsiB
3eab+Wd/33MrCr//eMzcqb9+R6tjVX8XMZ2kwVBSnQuOBOOAFnNTdZlcp4nW/vTL8fZPijT9uipB
pJ9SGhEw5oWN8CnOMQ6PaujFGORGvfnA1CCaDYNTNzRMXaX4pO8iacNuzC9nNwoFaREgn1RM9cd3
ICjIN6OsXzCYBgSjqgDy+bf7s9gC0tHqC8Kn1lCtN4us9qLGkO0cT14PU921Q1ha3QHITC5JZRws
E1Vcho0fA3+gOQwONAwsDbphwVmgd1mzsbXPhqPf/ZVcNqenYygNdELhkJjLgWgNkqFcZaKK3tOo
2wW59TjS4522l2P9xsE/rQjBvhng3l1maK2g6fb2OvQWewo0FVjwQwDzNqbRtsrtozCC9e/X84q6
QaXA+/dI+phLyperwO7PZwH8EHHq+w+LC/17RgU2MePjq9B8TitH+o3zib4kXdGZ0ca/I1LRn8x/
FB0czuDshxWZgqe8bgwKL2+gqWE/2KhnG3vk4FaiwZAPqP5z/zvOSiUbuYdpxYGbkVudMhh7buG+
QbRN6FfxXhSSzqfY+GbuXScuO8HDGPHqu1GfWIsy4e4EnmRew9k8qnVdLm6FiWmRY4PUDzIxz/Bf
8bv8QflDBXx+40xNITSIXiMFV7zCaPeeZHTVU8XvcO1zWwZIz708HUR0xbzdVK2q5XpEmlxznH8x
iAmDuEz3b+w15smD0qYDI7VagzhR4WD+yfx1cuvKe48FOiUSHBL111eLjkgwzh7HIHGpHp2/gskd
8cGthX6ZWL7tUxeFK0F60NeLepbH2FbpWXW1Qcq8sfU+WKx3P2qmP5JE5nc/l4qE0ON9FMErC/RK
OJTRoVnA98/pLfB7dcLiL6Y0h02DXP9tb4KB5sSqrzuEoFatWD2DB5oGGxob5n4Ti+P1m9Aq/vWk
M+4T2h/DQypBT8Py5uU0iTy8QdrdaGbIj8w8BEEbdCRB6IAZfoadw//XqyZ0FwCieSb6LQZ7492+
KEGWoyLwVM5ItQxhrFA1W0nImppLvr7ROEAQEkcPJACkV7TjfuYsJbBjABf/sPNQf8CAPjLQQy/B
l79uXrMEszcXNqH1vJjD1i8QmDtHsqTqevx8sX6LIewRHZZxGg+A82LXycHe+q+P1k5zJzuA0irD
hpPC/Ce6LMD2H4f1xddefETWLE7mLNh3u6TZZF3hMUsjQesk2SnAVV6PqTChjHLj3N0i3AzfYaIW
9xUsBZg6/FoeYI0cAVMaWss1DRPQDcYaXlWAVuuSqvVN8fhRELsjBi7JrpUNq+naOx0tIBJbJBDN
0eKjkHdn3b+kkyK59lJbs2jjKfWE8JghSx3YFaSDLChImeexpHwwQaW2kWaHJYsATVnHjciUpBy9
Hh59iH3Xf/y2+HfJV9VrAKPOruspnQu4GuADsXxDx7idMbRBY48mhd5nzJDHjyQm/9Rr7rGZ1jIP
yl0yE7JTTqWarLESRaDA2dbl5S8HGRmvOK002Xbrmk+fBMe/ryuLRqEHOdbe19heDw0ngKsPUC4g
7qgYX9i0Ab8G3f5v53zmAvwr9k4C4DeSDZjHBzakOb0Lyf7uWRbBUb2KwmGft59qoJsC+EXq+agG
thCcvXUtemEH0pQkI5B/hdrtwUsRv6aI8gx28gBT4IPJ7YeXeieGuPGhy5UO5bRWfzN5RfVp4j/t
V0PLl4/RkE3D+Qa+VBq0deRG5NhwkBtrJPRGlN7IYX2w99Zx5R2/zwA9lPvnvzZy5550zPpje2kR
8hwpvHEyLTQce6cXUgKfAKYJpkh4VbnD+xgLO+6L7ZzVBS/7t+VY1kYM6+19l6QZkWFUTaQQ7rSX
Kudwg9zlpY4IUoXDQYkobtlD/sgSbF8WNFINfMAorwOlnr+d4xt6GxMB4KOGh2HwqCHwP+oWCx/+
JoH4iF3zG+DsUNZ7CWOvdAGdga4OQ8AgM+trdwZKeAncYCkJqvljjPV1mBA6HZG2nYUgAnIztPRm
/JajMdLdqQBu/hCvIcZDoHRPe3/56ed0DQB/n1alR/y5jZCeI9hiYC7EMjfe7lHXyXcqD6c96Rij
8fShW05maunuVpI3/v7HsYFsgEVmv3Pn+i113OrexDuY5MAGI5/PNmO7YdQl0GRMSs5jKEOcluDi
BWdnn8jOBKy16VmnW3q2rVafsNfAMf9K1roLYkkgJeXCfS6U650IHohRFQN5KYX+PHA6lsE8rPSk
8Q7Ot3+CigPn2/P/oObNpSEWZFckTHv7VKITZty8s0ChymcKSYltZxDpyRUVheAKN27cmdKuC/cX
t6D3x8zRZ7JtFX+V7vT8GBCYcSknl00fRDrRJpNADTQqA+WPMEMyq6d59CuMrmV9/iiyMy3RB9yV
lB5di3lOphE5JlIk51mlRMilwreht8J7BroxDbxvea3qOMf6jYrSM73XRx/CgdV2XT3BwomL/W60
nFM/ncxDu0FWA1K1deDgCw7/OLYpN0OG9gWPditD1Sc/PaAi1+E4BaA1oRAqyYp4LO/m0pj9QR1H
bKrxUaJdwjpuPURTwV2JHPOpXlLbKj+1Fkpgg1jXu/1tVjLqEkl2zBwnVLHXJZteA5HkRBzXxi28
Ex/UD3nKiHD174vKNO9AxKkYQTgJG/YxA13IMLBf8+bbp/TPt8+HBo7FIwxL0icf8ykeMZlcEuAc
2v0ZhIDM4hd99WScZLumPwojsW5g8dM6Im7dDKytdOH1N0Tw8ED7MepHWjQPC9mKTkxCROWPuJ/x
DxC1mwwxxCZbhxGPY1TG/xypEto/QuF1tXVAYlKTmYHft2ckBaNDfD+X5aXrf38SQXN0iM2sUNjh
Hneme9Hgr/DMAO/6bz+mMAK/4qeW59BKziYdPZoFlPHUOHjTssjOmUZc3K2d3HW4I4N0qPIqZ80Y
KCptMCi3uz5WIXmnDFscU8nH+Zy1udPPD2z1u7KBSV6b1ej4SzqHx1WVIOdk+7ZO+v1L4d5hOkv9
wp4NzxULk8xVubLk2CF9cKGHM4p5PjpdUyHI3Gc7DIt69ijexzi99GZvRVVLCW2UlhG0zW+pjEV/
loAqCx3hGZGcTmtTyqDHxLVQ5cETez5zgpl+ZpHG+V9QpNsbQZMH5Hu5oH3uaa1Jq8jgqiC+fA7g
wNVZB9VsoDTDK1ipOfdaL/irWnRULqPyRN03d4dZ/oAd3H9CwdwwP70wcb+mS0BYZGc7dGVXvPIw
bb55RK90Y7RZbHf8wrtXKRADcUjX/QixW+ZeUK3yTvYQW5rR+FxQyi+5C/fkch85KzN/BIICZgLK
kNw4TSn2MjMAke7/n3lBIqgwCW7vHaJUqG2OOBJ2PaHr0Jz9pjwAKs9WVQ4Oy+mya97TDehXKVyf
Y3jYRjaXp6CaKdsdqgfjIpcboUGlddGTof1v3uPol4OXsJ+Cxw7Bv5NXCJvBuF6U1GLVD9GIxM/J
UvITWpuraedp3xMnYPo6Q/jNDw7wvzyEhzy5eo/g+3qrZebhFqGQDFANlmxHAfHVFUKaUNuwqew/
boJlRQqA8n/kUlJaFK78h6leEsgiRfQCrKyPFAH9Esr0WNI5GNzLmE29tI3010vj28OOrjeph6fY
yHGMwUjd+kM5cRhslrwEecOM5QPF7/kxY64JJWUNWZu68RoDnS089WY31bFq+ekSFrKzMlAdLEsg
R3CnlrBS/dnIhJ2Ul5WPOd+pZjp7XuGcLKIbgDxzyXSTJK0GKPgkYg/dwFuHmUofCfSdFl3U/3Qq
sKEaQYrN2JoA31HgrsrTZNblKACOK2KTuRLCCwbe4vTvC6MgLLFRbpLRQFR0jd9tManL+SvmmvoE
ElBrLj/Rfi67Mf1hfyQjbHKb/4R7EJ/sgl8Q6vWgpKfl7yNFo1s2jFyKl+ZvIyLe0NPca04jITl1
r5IBzf5upHhAeKOroZvqjtY5MKtsOTSKf9E+r/iIdsdoHsvylWrDNGK4+9TMpDtHVoqKmz+s4FS+
AcGxIRIsLe/P9Z9JVtfH2rgBEKfu7aP01wIm6JpAQHLF+bRejNvg5D8cBvOUSddlwyQHhYlQ6v7p
lRlHRRqf8LPnzTytKJRYO+y36o8GPUE+sY2kO3MDwGuKJ15Us0Yz8zXaNlzXPbA34qyR0jIRo7BP
ni+UiD1bZSJejENbutTHUQcTARPi1b9NMbM9meVw12W+vaZWAO0cXzuN7NB+52KUTLOdONhTMtxG
Gi6j5AHLJz0A6MIpQlHp5UnXXoTuDoiIqydRE9kD0HcO0PgWHZ7MlghytRgHLhtjtSBE8uWgZsZs
srtmssY4v9b5FLmtLQcvahZHXHDCb8UPjoPkMmdxO5TLtT/1X0qYJhDMc1frnXOxDqkzuF+ZsieG
VBL6CtWGOhkfc/9b2SWimOM1E+tmf/aMzmtlNZKW+0wx/ZhccHTQspb0Xg2f9Awt+wX6ciLIjC0D
kL6lil4rvasul6ISrRP7DUx3rduoYFXJ6eBtGjdUd9FhlD9POCeGuEAAS2g/g+fQH8wv8v+hfSKX
0BD/x4LEiYd9rL7oo/3DfK2IgJQeWspOze5GHOd6pKDHy6CAFLTYZF+zUEsOPckWHaGkIQDKzby1
uvFhpPPB5Uvxij39P2PaNNv1BEoU/m0uB0jAMgcHBErHVDFaLzSPQZE450Q7auPS3bXiONJH0gRw
oxl7Lhiyaliwd0rPIkdM4rw3x/XBW5AGjNuWyXiFpwM0PF8WDQuoS6tJXfdnZ/82XAtviDj6Lme4
TAcrWZ8SuDw6M+jZFxrJ01vXTCIFsh43svZ2IYPAqGbEO6253fzayMDRGfNhIcRe6iqIiBcRBAXi
uv8YSSaItQuzSZoyq/182ydIL+b4kSihA+33NcT3++VcobpCQgTgXILXp43i8Ee2wLAzsXwJyVPj
oYeLmzkOTdN1N7zXv5JRJGHXOtICx1qSyskDLToPYFb8FKi+kMV1jGBUM7SVh1Om8bX8UrCjkW6y
iA2yQ+q1WKKt6NAf1FfEF4oPJKEFW52LoS6JAVZIOpFupb8XcxRmlpBECQVGnQseiATRoLRLNfbh
rJ2qBbYqG8Lhtma3HmAXwrIK+vP/sBidEm+S+zrOBAEOUlJ8hOlpyTZW8WhDSDPp/bzUA6JxgQRt
eDM61uvjx2OaP2my6GvSU8rXpgx1dybyar7EwcnbgXfd2QWdSPiBMQXBHeailN3ZvWk8vSmpJXHX
RxP1wcbCR/kjMGEFhXRx8RUW/VURiIh0MstDB9yI2bT6HgwqllhtXoJqwwLaFjcSlArNbBzijGii
inoTkanP0ZUCr5sOkcDrcgMwTNExHbSdf+GwPX2EpTFM8kkfsEgAHxYAmHZqFuQygK8dpKGUc+1I
sR/GS6o8OAhedgDp1brIzSxRrrC99qiEMC5YxhFJDi3/Eskifj3Hlxsxt++Mpu+fmQmOok50+0D/
/qfGfLSWbAkW+xZaqXbSyOHGLKiv7L9iqZPQk7/NJV3jFf6W7UqYwZGjllzS9vYctFEDQF1UKbUl
+nAtYpUc94E/qNdbhlmgl5hcnSJ8OaDFJMCrRss5QAufz3+gv6GfQ1+uAajP2jPAZb6f1Pa6vFxK
fSYCAE29C2lGKI5fY2cqD2AfgPoli28jduuqDu7GTsjKai/7B/vZd0k7awkYUch1qNiybhczaxsc
6rqBbhJ5oHs2epYtVdF6Qo8FdXswj+zD5l5yqAHEhDJzOAu03nf9WvVOGbSwg2dUoMBdF91IDjn0
8zKN35arBPNcg2Og8lqgxBn5IUjLGjYdCa7qGkhEkPsTixZQeeJOTWKP2kN3/MSmduUnKFfwJ/3a
RzEgd6rcYx1JLn5hZwcjeGznmH2HLJWjA0pPh1fOzUeuLtQUJwlf2xjhL/RHRGZu5AL9GmIDwRBu
0zlDEU/23OLtQ97Bw5A5hxx+t13Q6uO6j7ZbEGSbkSPf7+jarofnRzhIBcCSx6UCmhD/3wXH5h84
e7MVtqt0JJN8XXsXjukehKwLgMOeJn7OAZj6NN1JAauUkV7ariaS9b6y5ZHITUehTlA/FxPH3e4N
FbBcy2hsVpC9+JoJ+K069YTVEsd2vqEO4WPf+tBEay0L6DWqPlES6pl/tEC0ukiok5xoWH7B+PPU
h8H/MAg22p4bZ0VQ0cyW9IGwvKw9FMVPojtoEQwkitC3CELuzn+60qOVYafhM+LBcGTJnLsNkkYn
cU5KMcrBg05sfVBK3fUNGVS3Y84aDfTUi6krz8xG+v5tikffQC7w4wrYse5dVEj3ez5gttaDtp4t
zPJNFb6zsX0EjrVchTFcgS+OfqmEq3Z9piEMi9N/qRjYRrZ2BMDq2TsLmzbWhwEuwqwNerWuZD+u
ENaMU6Qc+9uO2KFdcYOboi/VqbCGe0Jl1CpM2jjuJLXirXlYACWDL88Jcxma5oqr1eOoYTj52dX2
yqDr7/YY3g7sC4b2AgTqtRtmabX+C0hyA1PWLuamn/YdJd/FxPATAvR9NFc7VuVL+oLD3+wTwxt0
CSnT467Zk5s/vWmy/vJp2/f/441yxKKk/G8I6QWeO6a5RXJfsp8v66O+ZPOLjuf/N67GcWPmVpz3
A2aux/F+xhK7asBu6oH9UPrst1ZE0p9ruPa5CEy5mg5RyUV0VuLQe0otY76Vdr6kBMjBnXk4WOlb
eWlkqk+J1YVj2o7z8INar1k+ZOOfwfjXtAHnEKmKRQFbdMYyPGoRwqbFJaf27D8gr7itRznRdqgd
fmXKZXbn4AF4Kslnk1Tiv5u/kvQTsO1P6MUlXKT5NicQl7TTqDFLSzIeeur/vfqXU2z5KEs8+sR2
lW80PDbQdBBjf1wcGfkMAs3tlp7DIkST8Bbi1YPKf964iTRjY8DfjOOUOQGltgwB5JZojZKoNtGF
GkAp5Kv2Oo3iKXNcYxK8Iaodu3KSEmFTlBGTPirIONGGAGnCIQe76CiprnruJ46M8f86nNLQMSBS
GCXUravzMefwmBclAZbbQVGkcO1SFkthB6LNspB1RCMcap8byUuwoyxwB/RNIwfAA7khDKGC1z4B
rPem9hBxh8u+f29sR0qDRpDlAETGNYS7mysor9COWgYaZeDgq+zWkbXNJhDHNiyUclIxNSQsamdE
klJqATdJ4J5s7HT5mFM3aUl2gn3n/6f7zZO39EdlOBpEyANHLyUGE1Cj2AAZimiusEA29W8UU2f2
g6ZIQnQM9xLESwvwXxZkJ3S1Z1T6Dn6ybqFGk848VLzuqnLp1Z4QBNmCMJ2QkGqbLhra2rYfFfHm
YCkilt0UbaQpy3dww/JUnZ2FywnPDORWkZzNut1dsqsgnUaDUf21T3Umad3n10cvNQxwXN5sdJB2
/m2FkU8LfVIp2kPZCswJxP5l9Nsw0jkLehG4eh8ph3gXCl26zqmMEl1Qap8tPBuOqbQbPMy3wLf/
4a9XeZIonEHu0WHeahVBK5xS6GUUQia8lwXMnkNrGxewFlOj78B93z7WzhMTP4H/oDaHScuJkYW9
EUqIIbujh/B0VqAa7oUUxg0v+3Wkr5sb6dpr40Nln8/i2AqdpZ8O5+u9z8llhbEOOWL3IyA+8cf+
+6i3Wumvhy1315cc6Bs683/Q7qDXz4dnBT/Ft32CEDt+A7m6hPaifdOpaMachve9JCk0Tjvhyu6d
2YNzBSkA3UXACC/A9AmIe403FeCRNnRqOGpd4FbODh8Ld7sjRxIMbx/cbam440OGsqcEIs9/PWCw
a3idHC6r+j95bxzFCx99d1RVEh4XMLGQFiPBUXSdx5DdhQwrJ6eFeAVZ/L4P8nvEjnZD7wSPOAja
5YmemS/jlZHM5nWZbgioos7CHxKEj45hpJNKFyORfNumFO+VT9pVKooxaVLeocu2XMRRPK+vGyS9
E9L0TStvyUeegTeRr9c6u0jzeFg9V0xz0TEA2Z/ABGNZLpVWJ1/YcE7DPmcwx2JH4dHFHl+RC53K
78PrEDEGWeduDKXaHxTRm7s4DOS2E0to2sBB9o3Gku0hwSvdsdgtWLRGGXi0WextdVBSD+al3Jxj
Xs3GDWgOWpK0XDqqas82osaC4IpkbCPTTpUuNFCuhx77+O8IT7nhVNzOWeR1S3yzWPiqbGbNjECx
+NLcbIiWOLfZMVWzUzxMDffa3CVOh4ecQVrJOyLBX2a/xns6UPne6CRtFOdjUKlIgFoMH5p3nP0p
iaSltJOFAjhl2cDaedVrnb9k1fKOTtiL3AJgIlrwTvulFWzp70DIku23PxFhwbLwVyydesAdKtSE
YjI8A3AkPs6HP1x1M6FnKJLlHlNGXK26EZzaj16yFXhM93sQcgtzf4jHoDrdYP/JREmqmXqq4lNu
oI//RpdijljYXdgiEY5JnHY30T+JJ1IEYuqgitiL+66FP70i0V8P+tIXK1O4iFD9vMjWHkEM6hlf
cBTvrzt8dBH6+F+KeVZ/lMt8cIqb9/9qKobTFL3JlL3tsAe7s+pY7asKXlDGXQzK6rKeq+WOCZ4B
KkAfQkK9dYuxzvr3MpBXQzJeUu9e4robPeGcyIE9R7scg7xtax88eTUeV3Pr5dQ2UMrSrpq6+nBd
KQC/ND/T3RbZRSIe58TvXIMqGCLg3b2Uv9akqP2whmww6PU0ABjEz6k++ezGlhi121ZAwQThLua1
3C1IDVYpmeY+iv59CL2s+v35gb1msSUVpyG4bH50sGACeysAQdITTs5RCY1fEoxPX3ICH1OhEI6K
usfaVejk2Emy0sxLnjX6lbz0ODmLWjuysi2yTWKRqHDYRCoubO9ORc/uZ++e5FUSzFFV2jGe1pJy
h3TmYjZ3lu/RO2SbdflXUMEchd8SPElwImNQ2BQKTx3ldp7lvbQr0kKn0WWNcz+hvJqYC98vk1q/
TWyqv/U+bTRKjXYA6kPsIqmHFcG3st5jA6O+j0/1uBkU8a0qdwXSn9MfSotDyUyI6Kq/US/wpAey
mYl0EAK/R7qzj9kpLZKHhQEod3HAwDrG+X2WtJKeVA8svLuIP4VyNcKhuFninRaoa6VBeHoiry9I
ybMJd254RJn3nG/IRE1f95Pu6v3D2k6Jf5RCKN9vvphYy3yPjhJBqpyfXGbzIxy+IhCPyZ+M69Km
w1xZ/Tpfl9scj1Zk5Hw/UDlI+LQwJwNmmeoWtr3KRdKr6I0RMzNc79SUlMvu1dzBv86tzscy2mnP
2x14Uy3i6iFqIEnX06f+OlEzNu8wvS2jIJWzFwBTyxoLWUFZsdnjU0hyRPGKwcmRNbFrWIKK5dhC
b7LPgiSAja5MwvfjYtj/xMMGjh7YyvYwJdfSxQhEre3lFWSJjSwfzNo3+yXXDDozloV0rHe3iKaj
oKrlTEnoqGHo9a4CaU2ugwdE2zNrptEVOS70Lx55OaY86k3uYF8OP/a5hObg1HRcmvQwh14N4Dpl
vF5mCmgJPhuXKLPNz8hpYA5mkmdFFYU7nRZmnUcho7lTn0Q5Mj9cphIj61Y9IpKRIQbOH0hSBt3N
dzZhKDBJ3Ybc+Pbf0Ca5V4LlsQY8EAq8RV3qbr/EqoFguWGmAdz3mSY+O6Z0V8OTadEYvAZUMrhj
3Zu9yb0pgzGco6WS9LnsHpIHREPPkuCowmin8ZnAv0d8uYxXjnf3XDbr1ekCmK2vA/CN72HzvT5e
eAQ4EpIGF77fCYOW976VWtaCijWEHdy9tX3KOIMMZj0FjX6KJCriRh8eCUmYie8R7pscIU/OksBQ
jzJOeHrmGN9lMu1j6e++vjSiaAH7bs1yhftFTDILV5pFbcTiWUg/YXAfQwTNzJaGD/G3Msr6/wNG
neA6hmFYYTod+F+wh4IYds3H/x0vg9ANSssBjkQ8Msuw7FtFDuVxThHmW9EWvD8eKLLcXAoKT7DK
XFE4VFxOhy/AXXJD1hkQ5nom/gClfaVLf5wPKCTf1plkP1khAnLRyINUE08ElMdgZeEraxuOFSpz
om6uzZQyRk6tCk+k6QvD3DiMOLXEHGj3nDlOrBop7dLF4SaBdoX9o9lIFE23/DJAzkvtHRuDwPor
Wm8IRyl1I/aKiaTyTr3hVR0WVInc/psqjTYikqq9xi7jzvBkvPYEuWibicHoZysQa5UL4cpSaoHT
nLLoAc453w1zQXwgDkuSkfDMFMaykhMB7AhNRTp4LiUoOiSaSfpLaIwDpXPmIAAdKAyJ8zDRzYSS
CHzoSsE4AnUcElTt1DHLAyUByCtLkYzEKdOaGcKqDpQVH7hg82jRJd2MKTTLAT2sb5GStQy+QCt+
iH3VYbp+PmvT8iP8mYPYfYm5RyRxgrwalZaXIj51/oV/9r+rTNSta1ivjv9Iu6qfrjAkJvAYQeNY
AVFUshouU7DkTsfZBjAqZllEzApKZKLmwGWDE9DXO5m/gkAkmIoGm4F8c/1mfmbf08SuFkf5Oqcp
ELn1zW6cYGjEsyh0yIdGJ7ZHHbmo1pJz4gZx27YX40oOqJiLw3W/qXRB3mdI8qtxF+xozqK2jjvs
HOyF5FEqwroDVvYkKQRs1jvfkufzItL+A6Q2H899OVF67xNPs2PDwNuP093zo5sYcPS+2T4o8qnb
CHVQizLfzckN6iOCRvdNhMDdDWr8XTNjfDiHG0vOcfs98Z9XwY+6GMzMGj1B8cIVlnl652HuWgv8
PnueD11NELx/T+NrcucfnC4CYYVRpgQnjwWMd0dOLLhMtiI1/eLlbWFqfDl9bF4HON61eUHPCrA/
cZF6MCLReGB5io4sZnxP2mrm4n3nTrI7AprcYIeluBRHBOdnxLSuxLGWEC2GIVarbukhG2bPN0M8
lzppqObNPdCEWxn1b18NFg/LHNo+I6jgax8MB3w4c2ET01RtxjhPASOrRJy1qQf2SeBKvDkiz+AU
XfC0aEZcI5r6NAY5j9mkvucN4phbegJptdR7QlpNcXjd52U6LwuTASP1kjhCmi1dUMDSy+vMUYdg
0NV/GfCdbwcSD7UEccIy/cMEpVbGDsif6kokhEjGvYJ6l+6kERmel6cTfyP4fLsSG1Tm9d0dJxi4
H11ySfjo34+wmWyWOpNwfhZCiXZyQFpTy81Jszwp2HWklis/H1jseRtC+xkPLLxvdq5Vrz0dERUk
+wyIksA6l6jkUh3dVNMKx5zMiPaKLQlrVO6RC+j/EByqy1xccT1YC85JcMYQF2Ko+2i0Y6gRezPR
NDYDjrYYBLGX0rp3+T14zVDBpq9Eq3Fh9MIXvOJwJGRC6vsZrxUYeX6m7wOWS33HdbnxmdJcwavf
JcVDsJ8FjFNUX2D9Qp2xqE0tZ0k3Z9V8x83mfVpnTFhEVYjqAkiKzot1hEqgEny8PH4xc89twJ1X
3iqASv/pr5Tqubseiys1gkB9BJqG+gxpclXksUupaSe2K6/KR/Vg2pByYNfCNzSH+K2kOsV5tnZg
qOfu+uOunzjT4SCRiVc+/o3X2AHO8ONP5NnzRAm2jEPKn1vkOsV+znqhOZamjgrtUHgBzP0BUrh+
jnYrroU6zIJbwmScgjJqza7p17dDtJMZIdEheq25TVjXj0Oo2kNu8SHtO88mLDq4+ztcBWA3lE0e
so6Y5KjkJTQSqY7dagYAfiIuL8M3xHLITgyvpje4okSNeI8ItRugpjh9IXOUDN9hOB1QWbQkreMY
rc0qrUJBoyUdMIg1Uh8ZEogs93OkBYKCcu4G+p9MPQsosIdmZu8MEJmhtjiroW4mPopHGBthj51K
SPcklrA5ZzMEwluceK+0B/JKSqyoWmRgfcSTYP+8w33w2cFn1eI3puFOqagpslMTOE6HwlK6INvf
v5t+d9Av495HcQfakv4/cMBhzxsAIfO0KArMNgncnR0LRNuEogMOeCOqfthJQP4vIwQp3sUuUrcy
c3Cx0i69wZI6D3Hjeg5pW9B78sqyYR0/bAgLZTLEGgr3zXdCdcrLLNRC7fHHtI9HifNo3RDngYeA
cs85NvsfvFEakWSiPEko6Hzeu2OfTBCEFo+MPnzjcNanu1IJ4LS76Xqq3MCGNPnqDdRLgJ8+3xbB
NngKyfTNwBMciuVH7PNX0+smGh+2QLftCyrNQhu7IzvG7UX9YImjGv6rUruuAPjHoyoBY2hUuVSx
+v0G1E/p7OyJIrYZIDieYAhSn5+nKrZnDIcrLLgOyx7W19iqVvy9iNqxf2XKOxsLH53StaVf+uBX
SbikgYiM562af7JVdey3+b2ySq9RvjCisGkE5Qo+sNKuoA/uGAcU4ThDdmYtoDEqp9xcUQwvEQkx
utTi8hZRWvnWkwX71GYyUgOGqcJoKVLfkFrUtkSQRHJBi8EohnUW0kkzmZsuazxbH2GHt9CjaM9b
8EwpFG0Rlqot03jUpJK9MPjy93iZjfyAP8fiYf4ui/3YT8ic/L1pG2VA1EIoikJhSAApnxYdwdZQ
NuqzAhevCvo7X+GaYd3gIByB/RTp+gSHqYmgKRrH8i6jeeGts9Ti3weXn3P0Q56H3nHDgoqm0AGo
74vGlnwCkkDqMmZL84YxfZgjP71+46Z/SyEn+53wBP2FieTo6+iyFhlG6hPti4Gaq3qJF2Cn0gr9
rR7ZYkPwuJNy7mYDOocnRf/leUPARSSkUQU4TsYDB9C2hC5/phv8f5clcAJwRwK4A42T8N+FNuHX
2+FQahYbpfZy3oogihWGQQEdfIkl6lMF8n3twvcKcLP4lD4wZ91nRCngWkUXrW9yQZoy0cDZpS6S
0zGdUmcFmdXlcMRrbQD86ADQbsZAxaVq9QLyxoscuY1DO0kyBFUL4wBLPM0kga3Y9x3OARIKEXp2
tUUwFDRl6Gm2es3wjNO4EHnLthcCfrSQb26dN+Uc0d0qjySGHLjxUAPpn+3rj7qiE+fhDB5RkaEq
jQUp5y/LM2wgcnkG1pA1vB6s2Bd7/CORWqQLzYjge1mxXVFy87jyUSJrwAzZ882E3kP45ZNTJN0B
8jdTnNWyy7GSgCTzjR5Nc/7DzIdweuhoEhwCn+TDdBZeSoSPHK+Zc7Ci+QSS+Nc1vhQXC6mWnh0v
bbUvBNCo3FNxiQ53tEP/GZzhgc0BX2Q0XgjKAH6dgsZM5wU/tLnRlv1+GTU8bul2SzpALxfupqLo
OmuADFV9X5PiQFjrNM6ygvXW9ilGY3H1YEMdy5Y/9D14BsKKmb6xTMDAgjTtSeeImOcMY35zDf/w
cLTr2seweTpDoPNZFQU8wMfBUvpfrBYpqemBJUk5Gs9KbEE40i+fnlN+pgvTeVPhJ8NV5WzPBvB1
7u33fuzLWeGm2/uLI29FcS5MJwjsex2yK3GuRIH78sRmdIFssJ3abfaQBnk4u76V/XKYgrAUZGDE
1LZsUk/I7ZitQLh5ZKftcufasDPNjkN8U7kRNiW3VzN5vWKoUGlM1FaIAyekMKQYTpmjwSHUP136
zzEO46qJOEhi0k5DybRjJQde7kzUp5olF13KXktWvYNIALhcecUeIXInRvXkuu2ASp+72eBu3pvB
uTS8zWEmC57bt8EW/eiZ3AdDfuuk1sFPnYs1hCZTJztPSSyJU2Zt3bkF3lVfNxN3eB9bwFTvDShm
TD8+Wgmc9lGqo+RhZgzteIpw24dsGu9oylgycSIcPw4lCUx3AnIxtljyb+Rz2rw/PVpJ9FegHqBi
OrejFfsFCynSilHD0EwZPVODbKwuy/2GRv04AevTewJMbxWypqCZb12KyANa2DEqxRIdYvZJ/65+
P+bhrYZOLoJ0lyJI8BxhGB00bka1/JHDVljk8Gq7N+xt/jznio/FoW6o9FcJyfRxx7/JguuEkYaj
YwzDhQfjHg+18PSFC3zzrHq07KsMgyOsQqroQHuRVJ5rxuG943PzhJQENTaE5VVQ13IIK1VCmEJ8
8A/+LQ+QqtcziLDhurFuBf2K5ZfUGCguuRxcJhviBQH45VAb+BhnruXoxvSCSkEWAQnJiQRMhCWT
6TVPf1uy7ZqvA9oucvzGONjDtxbGqXNJpsSrTsnBcl9c8UqYbSs2QiaysPDf5zTChbwulQTfC401
ICxvD+TcBEy/AqYm3XhZORZXq6st80uBJxJ6bw8239c2MPmaIbRnS2LVvdLduEk3vJxlNrLLgjU7
A9xalzB3i/3ZZ/kVaZme/W6UuVa3eflxBUjA0CoxTi0dbPufxQ7f5B0O2HVz6wUEQuHbBTAcc7zA
9ciIhekMnp7Ofs9k+BMURtPcb3PVEpvYIR70qCXUH8sIKsqGuwpzauM/+H37BAc2selomOowOMyg
i1FPTx6PtuYVsnMDzXw/eXyfPU60FgM9u2PlwcoT6RLbEuxTAxUU04rqqMzhLRplcRyL7ZCRHPyJ
YiuGoM4USQ1d8SN4dvh0iR4zYXC9FgcQmSID5QJ8WUDpiao0Y2U08Bes0Arq/UG5MSJq1zCoq8SA
0I+Pgc2kjzZLvL2OCQQE0ymk36jKJZkunClNkkzxTzd9AZsGFBez+4Ij3ynv/aWUSCU3Yoxq/v3b
9uGhzsJRk81Rq3/26ztYz+Wt1MWXngazRDtuykqb0oF72HzVApIqy8Ikj5zmIu7PlgLOWDid/1oY
arhjILae1j5eGxuzTRIdid8twm9KXuvsk0z25xnGGwRewn/bXeqkHIBAp8q4nI+uniBATWXJ3AZP
LACRtc5tbqpmv8xCwflAOzU/HIg3RhzK0CB5HyOz/NjtuVdCbJD4h4lGLsW7V6+HPvziRXAAcaqr
hjGBpuYLXeG0qkIk4RK8NrPjWBh1yfTx6cHDPJKziKs6FynEJsPwA2nP2uXYU4nOI9KvP5yu4m0W
A0i6rnaJeBbQcJPw37vCKlLf+Xv2F+sQY/dSHI7fjrdDuzXHWEql09BuElJzFeBEa7rcFC2U86+2
dFMCB5xeH2ji8JYxAmLriwe/VwzfQ7W5CY/KiO3RN1LP56bNq432ugnxJRHdS2/Do0XdnNJkGH4P
daNHzCTVhIlRkgwLMVsPRcm+NLvUZLvn9mHIQ2uggwRHFlGHmZ7CHe2u0DeN5ycdmeSanzgq/zj6
NbO1MpEGxXm+HnuDecl14ycdN5UO10r8VO2mXieOpTGA4WrHlasjYWrZu1Rf9c0wZBGERQx1Jr2X
VuGSyxTelT/NKZWO9KVx0RN77siTvg0YAh0cDFmKu8SLcJvF3wc/RRhuUD32FkEIbIKbWkvlQYMh
daacWdQRbYYBdab6R1MQfJohUV5M2ccAL2Ri7AV2twFn2d8Ix9c7nJjKVAps8Gne+LqqP0GYjBHV
TahwSTPPKv6pBXFd/qLAC6bAiTfUNkJXAxZjQHphhizHDzVgEAf37Z923ZXmubxPozRlroTAWB1S
wigUqCjtv4I1Ng5ONNl6PlLe84e2Wz3VZYePHrim9cijJphw71w1oWMPqNklU4DE6XvG05Whr287
zmU3vFcArTXqzWnA4MpbYl4Vz6jQUSQra/gALkfPdPAzHr5Jy9wa/FEAz1ZskxDeVL0rCi+iqL75
GceSdK5wI//a/WiXx8Ff/u9lGWCAjw9Flmh0+18VHt9TNHFbzTOykUAk1+rOtt1/GNY76G9dEVT6
7UFMF9XgwdCL31nW+xubm63q+Ek6G/ewMVq2G+O2YH+m/EsvsT+EIUHJddcP+bmtG1LQ0WgX02+v
ZcTTE/T0U6085+E2etIuhZBJ7N4VfaGRqBCfhDEQKKK60z1GTCZdRjqZwAARQvBNUKWVutCf3voE
GbI4ACyTwMVAuEtU4n3QbzSxE3cwvrZbcfJqBxjRr8cyEKAWq5dpGwRHytZlUlskmb3f8S4PesTH
3OTNjtyy6+/cs+OuYuXfRqmN3bmFeb7wAOG/7UqQzeJHwPtFyB/a4kvQi6pZUSCzo1qdS3238slB
pwtAQRnjh1EKfyQlO68pNAgzA53FipdqIuTs4mb89q9HpGSCQjIj9ksNniw1XdE6ll8OvewHvIxX
XGy0yWHX3faWrw8eJWWCT+HtP2h2JUZtzxFthr6fYMzeN0oBb7rCVFEK+m0XtRPImRMBiVVJkXb+
UPE8F17tLrs/2BL/GX9VnV6MiHtIViUhpKwcQDFJ6AZrqsPNGU93p5XQxhucmLy7T5d4e9nLUuIq
2aQPidf3MuHLzkmvpeYRj4pooEKz3jjZPkRczbdRRH/KPxN/X7Op7Cc9MR9FAmX6Xyfu5++ZzLlB
bm5CxQwjrixM7EjfYTKUEsABa7EYJ3OK/i7UYF2hFd2JJiKCDZ97bDnJ4Md8ftcoylXDNqX5Nrey
4CM0FzyC55eBQFHQ76+mNm4sSsAtFS8phM5uaRvy8NnFIHI4jSDTUDid8dESSL0iqUG+G81uM2/U
vWMuzCCkIDEK7P68bWUptY7lPTLFNIQVIHhNCc8nHjwuxZ6L0dOw9CCCSMK+0xYq6czIJxO8vqpp
rr3mipsHJPwQU8zr03X+Efc5DVbeoOanSFq6kmFMgGQCwR+LTGBXaiVhl0MDs3swSyeu7F+qNXVB
7ROUJTBaNI61L63tt0erzCMb7dD4+XfVCcfJphn7hehRyWakmYoIpfL4svG+qxrNgKf2LoCMNqJb
37uoiVOJZjuiTvG9ArRP21i06do9Gh+8pSesfkNINjuhUQG5hkdIhvQLsmbNPPiNhKqKJgD8ljp7
+i+pY1AWX0/p8jb16mp6jwb4ulCb5jROXaNC4f1xhrVM7Tu8vLqiqzJWf/OPOL/Bcd1SKYP2xY6t
OwFqQlMHxkCLo3DRcXqVGkcIMUMf37K/SAUjOHf0U8uqu6kGtd5aeeCsMb+LYBUOqgtT7UIshzxQ
v8/OLNdtxypVKebQA6CbholfNIG7ul/Hemw6dzY+AjQ08l0jXHKxie1yTkYZlgnPzj53+3RYIZkb
P6z4sTiye63nAMa+XgGYzlOMojHOgLujrJsEj//bwzcKVUONJpUI09GZX8VD51m+tJw6AscyIA8a
mnB/BlnI14E7g97sJANqxCWo6eB+29ONV8iT4B+CtrVMX2AnH1xvwunhT6gxasLIj8UHgmClj33q
/NW6z/qQmattFBZKDBCCrXayzDVNHUFtR2bAR+EZfcbgnp1Zqya6z8xiDNxUTaHjC5fBD6mMLcWR
gdMyNouZssEW9EEqmlROw+K38WBK1c9NgSn7MFs7J9aXSF5frAFDTWlsJnGDIqMBa+qekBPNTZJr
Twg/iUiHkW6XrHin2DKu4+B+oJiB7l5m48iA4IGlHjKUoD589DiDz3ssGsV3KpNPUPK0YzqNV87H
dvI3YkOu8bmwFhaGuBmh3MuiqONxKYls2o5oypjL8DE4JRZElFK3cCLoTSirkxcHuznsA8pdg2QG
hXX/q2Ii3U+Sq0VahEf3ADGn+bhMiclaiEIcFletI0QGEgtjJmgEPk0a1eIGFpVUmtjj/KqblTQt
rNw/XJfSIfQJvO3kNvDAp6bYvmck9PeA+VmvBfOCR/K//l8fHvtq0hofSSA9dU2KIh2d/45Bm3VD
LlnNWwK1ciG5XdHBC76ieaDonV6+oPf1QQ9YCgO8cm4QLDOKZ45L9gS7r31HsRlMA+OP74kMmq03
Z50zfbyoT4pXN3p5Tn3vyySeLoWdDw9aWMQ5HzfR1TdvswJc5zHKcPQ6Tlh6TH3+A9cHJVlXZ6m6
V2ngnwHbw6j4rEDdQ2xpg3HdstVQI1i7xWrv8Unc4MOchvHNHF4/m4B64T7HikvCwyBctUv+ibUL
ciQ1NTBj6Vr0LjjGhg7c29zq5Wou8DtXV/w4x69pJB9684E4B9/FBCiII0lHKGKtrbWf/xdu0+j2
MQDhdbKu63CMuwmxHpXJsGhmYc2lFn5awN1PeJuj8l6kG3HdWQdfBQ1oO/c22WJrK8twXAN7J1TF
7KpP6pcXvvbThGqWF9/s189fwU5SErzqyDZey52Ztem6uP7CbtyX6MPj/xctMHlSXf6Po2UJvnmk
n6pWKsFNcawAHbykhDXo3Z5XvXwmW+sXVR32SRjNaY+iu5NbiT7dCLPToawfHdMxCPnbxQp3C6zT
GdblSRnUDIHmBGEEShv2c3229XWNpHnGgFMk8DjpcP6bj9KhZFLuRYRFHlb+OrkOfi3md0Q4nMCj
H4eXaHPvdO7/gbZP+pqpkDVeb/rTxevnvgmntWSZlWk2zyAZowWyB05OUwqL1FkHLc6uqCZstoft
fdYg5F4KaZT106EHnad4u/SJtr7etDn9cVv1QSA1ApSt2KuizsusYik/D4ImzwZFkA0WHM/o1KsR
kHHWVQMTIx4eGrFJeUw31UUW6i8jYjeGBKCXy5dlTmrMRNw4B1UVgfuAj/K701/bfuJe696jxxYw
nWqfn3AQOvviFVqKYQoch2P3RG5Vdni4X15AcJ+Wlrd8su18kJ5mVW1oRLh0ZgnBQmF50KAJLvFx
rO5MgktfQmX9V8xetlHkDEF46SQ3JO3EGNIVYZ8vch765AkHYsJm4GGGbosKTq1HIoODu/eT3mcH
yRnwx5Bej/mjxUwQ04myKNGvMU7ZsFoPoPpozQRgqkMnYU7t8OjbqkwXsA8r1QCjNNAzhNX1x+ZM
FeU/8kNxjSHc3/RoKM66pK1HhjYZeeWxqUOBYitQlEzNg0XRc8xMa9Tj/Stoz0L+dgp3BwUDV9Dx
nmhV9+eQu4LsnWjUH9x0hpFfhQHgdqXGEOtLhETv9ps/uZpi40fwZCjOUrQst/Z7J3UwSKH0U9U4
LcX6gFck5K5tvEwPEMX8zb/ty6qAzguF5nSYRDjymybNzSSxwIrkdHFP5P//fHHUCjAq15QeXpwz
1Yf9PtzUetElE06QoOZ3KZot0OAvnmJYbaQexalXxak9yDFR7x5RrIupGq62ugGxeBheh76a9lOT
vbV739zJd/OjfeOnT6ygmFfyyXclRoeArBaY0HfJzzMehyf4U3jJt8VttQzn55RPgYUG8doViw9F
M5rcNtJeOpwqkrcxIWSwDUpVMP6RmzY/vPdM134sM9AH5MJCfmMEsR+D5y7kAcay4jI5/8kfZ1fO
X0hsECnWX8+IU1jlQ6eFS1InpsxBGSqM5v8Hlhs1QEhPNOohyUsDV/7MvDIFXkl2fHTUwb6xaE7Y
RcZ9rK8/syh63puOK3dyF4fUs9QwLagOBCy/hddLAxfmcLZsO63va7M/UZ9FBTOgs3ZJStA/juuQ
HnKbKIVcfSS5jVtrAyEE3jxJTIFrh1HLUk0OEV1T+JjkJpwNLHVXj603cDIc7/50m9VP/6rWXBP+
erXs+S5rBVwj8D/0ySXkJie7A9Cyerpp1jZaq9FIzDm5LSQ/c5U2WhdAsajehqyvHYv/MooQ+oAU
Z4oi24s3Ap6p6yUhVzdDU4/GdD8/NMKFFUbyaXgVKPEMvAbKpgRwjjjaO9MCXs4N4a5UNien0hA3
7sIZJpA3x2v9h3l0N09+7SyURK4zXR6l/hpniTy9PEsPC2yb3htz6KjGcUMabv8qljFtgg/5JSXA
5JtAZhOmXFhYRbge6J6S/g2sV3Ol4v8ZFs/I5rk51Uu2jbPosqsRncRLc9ekFcdF0lwuBygBaCpD
puuGka6+rD5WUznNm5znoI/Ple0zWFS+BcR5QifsN4WkzNpIaGfkialsXN7pSqprZd3RqdEOo5Gt
/Gogkv85hgYJ/r14eyU0sfGr2CI9BOsQ3oMuAye+ITCVmJbkm4vrlLru+kWUj03lxIYH3Q4XDWyG
To0Ju0s/1N+oVh01DrZDiB6TbaJRRPZQcXQxkO8pdFv44mGTvPgh6bdJ+1xXPVA3zNNw9HUE6Clm
zd9hIbF8hrsG73zF8/uVJ+jLr/8zdolUTV6tnN9f76HVKddSNbD85L9SsKLEOHRf4MpF7f39qm63
ARQNBtiasOY/Iyz/NapMzIvPUsSbe2OjvdBpqXbE7mX83foSPVG2+cUe3F0Vp45dJhMOSDw185+p
SvxCyiJqbM+kpjPMQZj+f3Kr21kx1n/65ZMno20lW+ayCwWdj5B+KJBxjvf7Rj34hFrMmxCyMFcp
GOQLeQqj27Ajdtel65atyC0hv2Kt5ErW99MELCh6zemv/klJMwX8H7sTnNZ3vuNfNAFfHOFNPsEO
EBaQY+z201w2goTjz6O+vCJRO7S3F9Dzma1Xerh64mYfv8EhCrR4n8fEAHwl9s3mSDyIututpDx6
Q1CUxW4m8sLnnoitWtTLZGzjQnz5bVFPEvWj0iXwsUdxPT5plRs2MZCuAPN8zuER9UXZk05nnFLs
Jq1zo1O35WwlR6br96Hmb394HzbmP1lsC6yVM7Jied5ghw2mvonvtGBGKhI8E5tNUV1PyauNvv/f
REtaT9YaX3I08wXi4h8rV/kk5wGDP3ShlRMhn1B7kEWhE1y+luKbSvGEywQh7/M56w51iUkW/cKT
TOchavyy895WeTGyzE6uJU7dn7n+/Nnw/7rFgT4xrFMRHd3/OBETmq0alHerI3/oZ5MN4X7lRFMD
605fEU7+9PIIKrG2OMoR9l6rk/HSzUyLxEwEMZJHpJOOt6EZuQf8A0tmptoVwg+d8PUuzurrIMTC
YCmEw21q7vwi2mKNwJgzxNMzn1jsX2sREqhgbvin1I3xg8kp17TEQz/fZl5uQMPMYQ+uxQ5H2cHJ
ZUsjTuRchc9dJJFqS+AwD+nJgnnPDzygdZW5GbZv62DWauU9GiWIJJuChuJ0fRO7z9dBKbwLv6f3
nBuT0zJuGUypts/U692U0dBUermY/kEzWUs6NpXZL5S6lp+mQagOENjCVZouJl/UcjBxQHUNXwjY
zerqC3+tIdxXPDgmjWkLR7bxNfqbIn1raEZ7nIRcBOd+meCcZ+AL3wC4al50BvBatmbEUIYFgMNH
ZAp9TcII9YYcxjUyRXrQBJzobdyo1z2htG8mB2Jq+C7YuQj9LH8cRjo6pJPsM6MXyoJdByRQXM1W
k2qtFKYnHDfxl0ovCBHtfjxXm1itGA9sgf3fy0rzaLJ1UXFMnH55i/bOh6QIWOtD7pZ1GkXaP6J9
O8HMrYd4kw6K24hAtCrqhBPDoL2IRtrIiWKr+55y31X2ux4Q0pWrN82YoUOpk0+TzXdKEdap0XxU
GSvx1+ZCAtaRRc3Wv+fC6DSrul8UNS/JVi0cSdZoa/JWGELP/LBpycU4JszvzotE52inqJyBnhnO
AXQXLPONzlz8wlVxA5xlIxee3fMliA7ckItWXRF/cMUZ9dLs2dtxOR3qQHbSrMnZmMXq+tGtNSCf
OcQ2YErXdMSLEck+BJpvDjdOmWJzNQaFPJ4julNjq/WU2KgAZli7mdPnaqT/oiQPLUXOghq9ht9W
A2c8C4K11zLgUDqniz8pXg1BonB9p1cqoMur3XYLLtTrG7haLsMRP9kQlfswoAjHwggwsr8tsWkg
VqpKPbJ71RN804Xxz7cwCUmD5Zjaei1PMYSo8wtX4Ssis+AAK4FNQRLX8dgDvibYu7qn313j3rbJ
9F9UPJy+zIaT7kMX2z7Y4B5/wAZvdiLMyjluWa4JYuNoE6KrvNAfCUAYJcgT3cT+pskCiG7qfapY
I/nBPynSG1zRVQVCCJtMnP6hh7bYVlNuiO65AWmaRV5u/8zPdZIoPh6y5kaiPNiCn9hYbDBd7I8H
D3InU6JdVuS00wmQQGeNV1sTZ4g4HT1JU0xCRvuE4U+OP+eg3JiKx5gQJHb80TedZ8yOiNcZspZU
k2pjDuj5fPI6LSnxcNtu5QyhcByLW7/QOTNdwkE9It/1YMBUFprPrONkLJjDrnb5AOH/JV7Gnoho
Yn/ElNyvvDMt6Q30ZUOBp3A8OC609MqkfhiRM4SMRxybFVQCVafBTVizJoestx1MKADLS0ShNykB
VWtM6A7smDdOp9ubZsATblnF99y4Mtn9/jtwftrgewhEsmhyag5F6qd2ADjD/hk6dTdAANPRRb6g
7N5m97xoUoccoT/zs5qTyJUSVAS5BM9VaIr0g+9hR6uOXBnIgygsHmQ+Iwj7d9qDbjM9vu3/Eugh
IOuY93FUdt15vRtBjxq0soVFzISdn0rQlw+I4yX5T8HFgbCz9EtGBXsN4PjufQ8Awmn3MriysZR5
llqjpEuIm2PGevUGfK61YVDwgYVkmNo/Fi54PGjkl7WNotHRGksFZrgLEu6PCW/F9HwtissxH6y7
dvXXbWNNnvuyT0lGAf8lel2Z1iORq1Bl1DnYnSm9E0drHRcBW4xMA7bKaG53hp2A0GbYyjegJGzw
0jOqlJXey7Oi9dUvPIBvuOew3YYaWA2oJCsm65TNtk9rbDUH2OA/HanUgmY/4yxWqiD7n+BcCCA5
bBBsXcgK0GUvEBYUZ+FRuNMoTdsKD3qDHXnPb6CitUH06ENhwPoEnygkRGwA4KcnT3tpve7lYDK7
t0YmLohfVLJTlJtY3eilu/tlgeHaRdrzDUd113a1RJC0fmiiP/XebJoCHNIuKTAzomGD1PD9fMJb
tTQDPu+m69RDivb7fcp8Qhfi3HqmbrxZlhlUqlDHqOdKx11jM7vp6RI5beQBratdHJ0bBIBen4yh
7ekgJxVlOkXEOIbiOHd3eejWFGm+TenXYOIPWkLIbYOjtnAVilL9ph2qf660/uiV5iWXdxDVMXvi
t7bXEDVtcV3+37Nu8uK4+gjo3IRR1GzmqPa07O7B+5Nps/v9VJJrgzvlUxiguxIlhCsylGEkQtuy
RPb6dWta53ADLQLGvCFWTHmvD6z92bnxCsTJePIp+S8lcK1mzZq9T5/MLER7VscJU/T2hbVpjl7o
ohunqigeax4WmWY78SDFl6FB+bq/sSSbuEy9DwSH0duQUAQo06yKoov35AtDyevx9TA1v5Mn/Ygr
NENLgf4v44Ar44CvtTJKygTeMPFknWpOZFDfNmFw3TdEdOccz2+it0R3OeP12/wi4J9P4GEh4jOZ
FpeIhw45msXERSEk3zbnMhCCCzXRRfk1ExO1jRfNZ0tulp9LtyTrGq564gLBonhSByhDrdCEOxH/
0wDUiL3CObEPdnXvej7PzfcsLKRt1hmsjPqp6ue8Iu10TIhEDhvt4zVHOTj8ys7IeQ4Mq8wk5mZm
T2Cfs67GOc5m73PvISLzNeoUn/OWv+YlTk4LhgNJyzrAPIEQNdbxMP3NIuWmnqesW0pBBwC+6AQw
ZRBZjeeUoPEDRTyntJWI6Hez9AIMno/QIVGkKbEAYcmzqScB4hkpOlCfR9NFLjvaV8O9Pc3stPFo
QKor1Vahlde6qbg9IR2VCyPV1gB7N3UDWDWaj/qVcaKkhnvSw1hwjXPANRErWkJVNwLKz3kZZXO6
V3F0atMqB0fr/iLkwvdyr8B41yTzcGahzeTYmFVnAsk5ubr/HH87vjaS9xo2qqfChY3WsDWIPFmX
HMRluprknBuiWs93cBio6NzM0fNVk1NLxI0jMBMp33dIYUsP/wOJPSZ6pMdIn/whRXwEbD7/I4TP
zunk1pop32QEyKGVDOYp7sTRBKWr7T4IJk0WV7szpZ1Y0It+JncqCTRlWxwI7DMGhzc4koIZRyib
ugJJk1mzYyKyuXNFibzSUo8nzviW74WWCfQVYXhGgUo1/vYdUgjF5dhBi+WCvTqf9DkwryPTCV7s
bJwjCa2xpJV9KiDD5ikrrJg9G2gF9GhNDLeirXJbCMs3jzWNBvsknrW5Sij69cIUQ59XdcWo0R3h
g0unu7GnQynI7xgFQG0SgoQD+f3T62ePxiHpW+xOuxq5Ey/1eK8o5NufQzd1bPHL1r2TsrhLsQ+9
z4jR/GbrJybGkzzmTFY73gVLVNNfB/TA20UbCXIiZUeHpB9LRDXwObS7I9VCH98WtmGI2h62zyBh
YZbyv6Cwpl12CgKFNaPBjJL+R+Lv9ft9CYJYhsSLfwfzf7mmAukz6yoi5KdYjDCSnPDXmfGqdMKy
aWrUXh0dSE0N0VI3zFSIPp7BRv7vPIMyMF/qhgUP1goSkqWmKVFukC5N5ZSDL1NTDq8D8WDUdbJc
DSPyhqP07zjbJjjdhCIadAb6GehXV7KbpJMV72jKtiL9vgFd3wCcET7THE+bSPVCiok/HxvZ+Wx/
nrf6gJsK7fPsV3z9YI/a2KHZHjHMbIjapqvr30YfGqk+JHHJ2Vghg7QtwcjRhoXozwLeEYK40riV
0XocS8L2yPujXoai4EqqpZMPJwi8uIdAPugBzAz69p+BwCimmKBl8q4qiwSdM9k6ZyVDuZLoxqe1
fKD2TNrlEGdrjBbT9xnRHNU9tCi05HTVUUmiT51l9v2kCI52i6cE9Jth7Fy/44da9T20Cb+q39OT
73jEFpe35XVc0uuzhoZkI8FGavECPt+sr08+RsZ20I9Y/a2D7oP+g7w8zkiLbx3zRrTxh83YWNRM
V7FpbTAf6/1YfMKSWJaCYcrZVYs+KerGd/be99TCH0pVhKP9g4UvwsZZHcOtjPtwpwTPeFOmRmzn
mqRC3mZMg517fxsos6gCtsQqFoJ1dlViyTkHPooaaA5MoSUjpvpbW02aEgs7BzrRnpGju0d/6n2+
VAwK+EPOGTGWYnsPXJyAlH0l8wCRj4Vb3iWV/oKS7v/K5VJQDuejOh3PG7qfMSNLsuWWHfN81alc
TEguhpdvtRG1X2YMu4edVX9jvHL1oy2WCdwPL/J/Tc3O8syllUcLOvJ09nZq6DdF/eKC+F5mQeZI
p5d1s6lR2abgHUvHfexnicgBiUa1JkBcwc3OaPLTzc/SlSjhZ+o1UxZIWBUXCrNClIMSjaTr5s+x
N9WcooiHiQKQskaWP8FW7Ti7m04ogp13vrUzowXgFRzBpnd3NjI9ND0JaW1CM1XJ6MD+hAsWJG8e
aDoZ8wwmHShehpcZJFQSesp+rRZtfMsBihuhtRjkKswc6QZZEoXLpOwK69DoESaX1nRx+TV71qqa
XFmblncW1G8HpiBYbeH4Sv5V7gBk5N6OpR2RF9FLBebwwrQ682qx5Dgh8KCNLz28Wl7hcCIlaJZS
yY6gGckc8YYPM7ZBlznQA0Bj++9CtsuN+bHLNUCaLjsZnHp3D5HyMMI8h12Nzu9fam4m+R9EaQgW
DuwEvwDphN9CxeKQAIOZr8DpJD2JN5b8ZYfSRLyRPnwRIEpvfH2hflMiNbEMND82PhLPFDIcGkiC
kBY75TffQI36DNSgpO6BTAxJqc8aRZtG9N/5JpCq3mwFxNKCdjWm7iadnyWsOUSzVXFOD5WSLN/M
hJGc61irwznwGbW+j5B+xRTzdg70GTgZ8xboqnhvlWhhwbbQNoEthL7BJM4KHJms4fukU1O+xxwP
0hb9WAaFHZPZM/39uTbXgnVZrj+pqHryac8jvdEdMbdFIbeiqb7Cj0YYiq3qeXICY0ZUSqOJcgT4
l687VrlpfjnqiQ2+f3W9P8hE0dAdIUkS9FRop38D/moIGx3JRS5D61+nqLRwBS/wC9kOme5aTo8k
xK3qkQK9xHFhfNY2r/Tzg1IKL/TDYXEPybAnAYvPh13SnMAAw8boDFblK04TZHLzgNfTSBKpby7/
7geNcm01nSF53xmViviRrMNWp6M45iUwIeR5jFn0kFtAt4IALrSWQiEKjoK7ugjj77+QqeV9h5NN
ehEgB715HVG8Hr8TBFVXnklfsNQWDxPz1PFE4GO2rLnLYOjwQYzh+mvujl2vZmJRwuJ9lEe4uZ65
2FxQGVtowJMB+3mvqOYoAFa9blINBFl+8GR9boKQAL6bfevzhqKZ27xi1Hh3HCZ6aRBHAVjA/VUa
mnU7Z2ueus7S/wX3qU7aSC42CzTz75rQnmxREA5+zgHhd4x0yfhOXIgi0Pe4nuXtOKnlV3wRmcSh
JM8Y+VQ+5p+5Z0VbZLCyn2CPsEiW/AlZkumMn7L+gtRBXNpzwrT9rQ8qzmO07VTFWcYPSfXHipZM
7He3jCUM1CTuOwOLOKbAnuqO7sTsbJTJztRVkeFwxoGmYnUx/H2ZWFbo9BlGcRpmwayvPlgwZgkK
GvbKz5pHtwN3AMf6O4BdywfVGrIWuCvrnBKJKRzkEB1TaKLpWYkKsu9yAYPxcWbmaexJiN9kJSpv
zRUMEwjOng9HlDyW6re1a9gaBukClrBx+s2BdS7Cb4MF5xFLRutVTTiRP4YBx0RZDsHHcNUxNlHW
gXUSQ+6mXpXvd+TB1eR5tvRQacFSy4cGkviu+Q5OEaQ4RzohfMc2+rdeNWk4gwkUdmrDzPmo7oGS
7enDxgGpc+zH7Xz6l01lPL6otehjs63IKMFCPl29NytBnPEnNiCifZcJPdrkRVCvChijXXbsiSCx
TTxK2HIDRkMl8a6IA09BO8AEiPMSFLjJY9LV/C063YXJt1RiB/X7Grj0fs/T8bOtyONhKsnZrzRO
X1elcKalBb/z59l7jG3/Oz4WxMh6wEKSZKNXhTLBCp2Bo2UjuXLpz2cNN2/HP7Kr2mwycaGnIA5a
nf/Ekl7gWk56ngE5emUWj1kueAkDDErAI6J9QHr/n61fzVJM5ScZR2FT/PCCirsqVBvsduvz52xW
2Ps5vlf4aluK8RH7dB5b5VpSYCGWLs207lWqlaLsL0cMxBbw0RdVMDmeVQCJcVU+v0KPOra/USJe
QwkBRiFyIG06rHV4GNXz0qbMERL4GWO0FmXlZGAzC4+PR2uLVVz6hCECwTCSF83nPqIZtIoX7oh6
QVwBYX66gSpxBsoOK9G8bpdUAVWYiY6jy9c6Mlyt2KOUUJA2eGtCoZcRjasReyCwRTAaNrhmlfiA
Zgtkrl0t05Z3vrkF/nqBBJacSg/hazJy2tv09u5UyS5gIFNhEE5vWIlg/R5fjx+p6XfDHTXq37Q6
+OPjeFTyKMR04EJzpNe0u67LPHzjiVUmGp+dLrolwO+/YPJWTHAmffh84JDBgya7n2fvNXF2uf4K
0JcLYmF8EjtnXflVFJ6N9l+42nQEvKoO7p/eMCaqAoI1y9RvPIqf7kJtvg5BV6TovtDqCLD2V1YR
m7EG5pml6AkwpLzOHZurDLKIy85NDeiGC+y/QlfQJYqWGOq5oRYAzcbN+UBoe6YDpJOQShKWBCbd
HHX8D/Vko6Cs2GtfEiJqthNOp4Ty7284uPpkqswCaCQxffUisVaJ/lgVua4wuWf9nRuL5DypQ8WI
rTLZW5c9QtV3N6habaxtHKNg2W8Q3u+kbge0vmhlvlWKg73LgkOqPuqFqHZpMMb8AgXdQkw06byV
9F7pBD7fLa/FllhCN/LgDD4mMF3GtfMZqszeBiR6lpwEUSgXHfzbbEtwtDWR9uGnAxXBEXKOify9
5hhGzJbGLBnAzXKvI0d4Z+ejeg8GraXcWxQlpPRtkWT2tWbZUOBt3CMRQU+lbDwUVIBpewIMS8+8
3/iGUWeMCevdUL20w+cO1oi91kktl4GCQ20TlLGlSzYy0aF14THBYxH8It0fWRs4SXZ8Ok0gAlOx
SfkE7H8EewOyh1L+66KqAPXkPFWuc+VEpvnDYeRt8j5YKoO4hqljHaVidYDyPWyEyQY5jfkAVrbJ
/b7BfoqV5fMNmgy1HKzWbwN/EH20Ogt1QI8ztSa8oxPoPBJ8tPxky+fFpfiKSQfl0DrKZrBiobJg
IksWRWNUgIT4dD01Mo8QH0sMneRoqF49usQ0kIY0SyF/QxI8cmr98d6ejjrEBPwWLl68I6EumfQW
qbSSNBMEnL+aLRJ3nNtXqtI0RJjnBZ81WiuTJnZVJE3ikBEzg60kI47/O6uEqrdHlQ+JRbAvHhbR
ZiUkT4Q6k7DLZ00gx3LolAqIZuOnso1BB7hLTR+hQvOmdCmGyP4DG+E3X+H7a3EZiOud1+64esF8
Ss6Du04jNOKEDM36AAbXmya4KRo5BAe2D7kikj2a5MJhKQABrSkXe5MLgXsBStGgjFEuyLNeh6Xt
eO1VCpj4r4GH8O5380HF2H3UjjBATfZ/ljROkpqd1HaziQGU0FdNxQDuPAJXT2II5+2qg09xAB66
IsXDRcTNirb0pAiM20K8ELwJeeKuLCsIktW+Vpe6/PdTucwTdaR914CTCRcRHtEZdy5YQEnXKB4x
rUzkgxb+mI5AeYD7QE5kIuROmCJnr6PThE+6+l318OFLYabFnJk7OW6yi54F2WuFI+zjrYWuj9OI
sYhZaWjnib1avmsBYFdwvJ0m6eR/k9s1Y6t9/EB5tK4kPu3GhV9pClKbJdWfFV+3QjN+eq4KaVXX
ai8Eq/QIbIVfKEeOveS4zUnz5KLNGudn0SxVpzobk8+wx86/5pzYVCuIywdxcEmRV4j2RlWCHEnn
UgkumzDtOIwA3EpfQdNlwjfBZnncSZ9yiFtG2W//uWeLpqcHfkxkQM/y+FwqClMmh8++W/mODUiK
pyW5aGmG/K7aucESJ2lYYuBdsOjK/+GRN/Owt5UdXkq6RNzU4dEVXRi5e7S7xzQwm57XxJIe0r97
h1S38VBqgzS+Gkjj7xIWAcbhdcp6uoiFNS9lzrYU/ri316dN+akDShRrxh2l7j+TocbNlsxSDInB
1Ky/j4wqZYUbLqrvef9HagPWInsv0A0+FcqGKfnQ1uSQgjQdybB6kMIrAPQxkIu+awKaSSby3oMF
Dm5/aL4i9k6vxmZzNuq+dicgc8HQKDzldRbMExCkUiby++aw2XHX3yRxr/deza3ungkXMMlMIn0X
H5eUC5lq1b1VOaiFLWDk4bIti+SYXaZsbqfH36epfLH8Q28+fRdK91oR4VktQ/LDNY4E40TxbCsK
1/xUrbpmAqdWu8ArIw1gjzIRlfUDTRqwUa1w0YSdhCbcKhOFqG1A0Hw3I9ivo7hOLLbbmQN4mMci
jlbOeTpBqP0LUmCX3ALup6c50YK9HFTyf2855HgAWynhDWCcTn6BkkI3JilV0eflP/Y/3dWsDgbP
GKmPOR8WgST8+gEgI8qh8QYlm7VomHPl1rExEzwJWxtxQFRM/mtWMOnLuPGzUgvdf1Enem96atvO
4QiTjfqtFs+VnIVBXkXXkmR/fBPuiE2X9VsDSIQx0NH0KEQWens/wpm274XcekL4Hw+/MlsNOMLz
QRgClFRuW1sXcRhPTGRL5nQQhKdjL31RNT082AgO4Uee1j/7TmxQnQ+3pL6+BuT7rK7PrrMTF3On
moo6HD79M0/ScIKOwBsz2iTcW8ErQ67dmgXTm4rbV1lBK8rSmUuVfFIGIAEAfqtrg+cxrwz/XOat
Cp5l2bQhhr4d5HDZM3UM+Um4TPTojN+ycULv2yHZfRRC1yhClt44+QAb7/B6WNjMM89GHcRmEqz1
NXfTigZOEOlqV9NIqzygqhf0HzRF9jVsNegWVGIXi5k/k1o4owuJJ6pyZia1k6A2GZNaOI8SkYRT
90Gqy/iQJupmsDlirkZhSUOwUYJ5lLOBu/MXoX/H774lUVvH1Nc26IIQ2QurwBOn5sWEsX2VaJ9l
yZauHy3x8/olg4mHxAg/cvdAbzIWhXOrxcp4Ziwo4lDJq8M9im4TP172ZnGs09My2elHE76BDqok
lmm7EB1blfeotAF3do8LSZxNN2zUnrf29gJAJxLjVjSt4S20+uXkRRtHRkc3yaKb0ElWAEU/uX5V
7431ROmX7BVjnJEz98WZvldn4fzegAT8Y/M6vl3wfKzeQrmEG7fkC/T7V2bl0hfAoZhjyuYyYJAs
Rj4R1aZvn4lDSsNWpQDDHXrN+4I2dcdHpJGvgXFhn8nZnjSaC2hgkJwxMGOw5+VbL1Hd1qAR4++P
0kJMD2CzPZtlkEg0UrFmWluttia0b+HQAC+UvvHgFoIbQC1ohrEazbvZ0lQlqbh5aC9TK9UTKRsN
v/KR89L5qfQhsWwu0BkAmBvwOWdTTGUNTOlt+gGhqq9LcI9CdBmeALGrCgLNb5qpJ/7NEqai61DO
PpV48SV+xYoBlyi+oiW6bGFFDpWRvaovoKs2h4xbALQIUVHHDohIc0ut7RBSOrXirKsNi3iP/Ria
4T/KYKDJlQT6YeCY0N3NDgEr6fYtZ3slTEOT2MjL2M3LgV96Hgof+nUVvUajEGsYLO/TOeLMF0oS
yQhBIXo7knxt9DaJthnM8+6m+hnIIsglgb7i/ZGs3rWkVfb+wIwIUfnJK+kcAhq1pD+LoO8QSdiS
vPFrM/GI8vII+kxp2ExiVxEPGTu+h0pcdPjpOtfMWFgGfpLk09fu5SkSMVgKkt6wVleAMied8dJt
zE1U8YqeKzMwmrAt1U5wRXIFVrrwHT0/oll1dJIqb1eIRtRpvMsgb97rdDL80J76TLtdDMgoMy25
gUbMY/coLox4qu908kkDbWmLmv4HtyareXtxMZuVgk/TWfmJwFxoV4JM9hFZQ0q60P4pIVZn9For
Fa1sYJkpB80/7+bVQXRNTr3isbaMmz0eCuN4ABFciNsK7gLEfeyncRZPkbY7NtA9lXJli+OI6md+
9OEwDAaectbQP0Zl4XRR/V7/NEqbVSK4JwmS4L3GsDBJsCxFOOdxzGiHdslPyTOaUkH+zkTZwr1S
9JKfLZtA0RFrTdquFnsnA2aebdGv+JIBo4KV3Bux/vbL9Rv7kLgf0QKk8krlifcUi6x6O62qVE88
1sCBuhFZ+KQLE+E+Cldp5wj0p1VEr0cSt3cy4SHm1GaPys4i7lW/2o8QTX6Cj7H/z4KjeOUroR5G
k8OHerp5oJXcNFRxN7KQI9lQm+YQD+fOpfHFg7wmQtkCHLjXzoBAXTKZseaD0UH1SV7GosBip0VK
ZqUNV3V6wfclAYflxmRGIrNYEllYjYERPFuHQeJSjgwzSBjbLDksaOCjzA19tpECpILwL3I0ltvR
P8tnW+MOgnWbH+LwVusMLlrKK1p01E3x5Tzf+QhDlpWfzLqGzrSRgfDoGKqs+2Jj+haoqY5Fg0yb
bHCyDWQnyXBw2tesOFpI9R2IdWrfknsIQDAdwAAthdrSSlKeOUGQkMLSqWTaarlIbtNn8OVEhkE4
YaGoXx8hEJISzuTPQTioyHPLZfbwbwj+8L/qwU9aMtYPyNoTcW6eMQ3wHpKKkY00yFkSF5A4BW0o
yn6yMkUxsqyBlgedq2Nwlk5cEHRBYHCoTVKcDXKrm/qUu9ahHXotwudzMclRNOkZoMJ+OAPFhoYN
DQWJWU66fmfs5auADeKKl9EZQ0xwD71EoNb40cXKMV6+BC3c5D+9lOOx9Y7+dNBWdGSIIlC6ArYH
Bpbl2McNd6ZRH3Mce/LoLBWkzc3238Na5SyUNNTMvkfOU5zrA2fcunikGRJs1JFEFGfPlWuznq/L
sHqLaGGF2wfyr4kHAnJtxcuG1S6qBzv1Ix0FXl7ipGTe62ZGoWkSTGLJ10Y72ayw7LWOWGYuVxyR
mGLAjVpa+VcrXiPIGvXy9qSzQzM4cMQU3nf24D8N3UbNFAegZAKUmS4ci0Md4LpE157oi75H56zs
imj90KxrwMINw8X2hIZqiEsID3CCmSwM+wIz9jhrlDkDuG5k/yRhSLkf0Gm3yKFe4l0y+KyZQ10I
V9DSNwoJIN7Yy+lgP5hQFFbjzBcV1MobFDjDkZn0viOAT6CW2sdmPVKPaO5AbdrYSOakPEFFuNAm
isrMDUrc7n/1dQlnaktEVFC025eazC2PRNcdqhgsR7HE7U0RCWDhEiBcfFAM4JWxU4AHmiJQErYL
ovuAmn0hYA50LcwBdpXzyqy3c/j9RJXDkYrI03eS2zx36cAoM4PuJory4G2bmUEnUe+k5u/9F5KM
KIjsIB2l+c3MVUEUtNPqyVwnSfbcJGoQ3jNnWVFrl5R5DOd9o5SCHklCCxKZ188bRJlMsDL6QRp6
WrZ6xJbdu2nGbCgf6OP9a9Kh++/1ne8Bcy9SUkeqdEtCcGpx7E90FdRgc5uu4K12/GceF47i10cB
VTjjw8EGyq/KMvLJjBUDq+INw5iaayFtla+MHzMY4/Atpp+XvPl1VOt3qV5OrCzxJ1k3ARLq71QM
Ozxr8nhmGhxe/dWcUveAUi9DUmbsL3WEAivCyCbWotopi6s0SJtUxkfx2gcsp/rk9xYcatc9mpPb
7YF5PAdb+4T73O5eAjU6zOgGKtIA2+zL1RmidR9uxPzRs2NvOjb1B14nTwNZ1Dz2jaAknUAypENc
9AJ0eC1FHwL4z2Ws2XNozW7BsSjlgKliIVRL+NYXWwLm129OpLKQvzTa1sDnaI6zSoyTmkdRfL91
z7S7BhI10LKAllEa7eT9343v8nub2nW81adVPbPLpjSwkFAxCvja8Q0EShf/ekJA1aqJS5XP+pr7
b75S8TKMTD83qCJQPqo2skna8HbgUwlv2Jf/rdvjGaiPifk9HwvDMeZL9qczByg32xhlKSufgACs
vDyllhxCMsiKbsMm4dx2sywn4NZ1BA49RFfwv1G8G00WkgkREUwRbnrkYsIx2VMl8q9HYuBkRDS9
dRRMD4P6OJPUQZd01pDwx8yJ4pvTJe7uowVUPvzHgHThlMEhAQYCACO+PMhm8GXvi409Pb0alml7
udoOpRyKXYmNVQe3IzfaRpVamc74eo5P5pt93Xo24C8K2yLUMWQ/81n1Rdhf/g+lQSxRCBGy548u
cZRlKSrwUJGH1BAjGMz+TiF2c8pdfMKLuKseT9gBMPyLzIFZQLbapB3wS04yhDvOjD5oN6HLLNLd
KBv2L5SP0Tbb7x8eC1YNJUvLXKT7S9y5ElSljSY/6utb7z7LZk0EmUq8MYuKO847Nq+IKIInS/W3
sYmbQvnwbkjPWK21qIS32ZWr6BktHv8LAAIxaEEyD4920oMPU6dqUyzwWg3YQgeW8d6iCOKYaKHP
4F9/IHaEF3EPPfehxgJa/Jtf3cBDJJhAb7svVGkD3yFHaLNE9I8OM5tl01dUFL988sJX4VppZOTL
vrkv8nBQCtVaGJLqH/PTPiAnIZPk2lXjJV6yIfKdbfldQw+mMNYyWWT3oy7a0rKPfr5kQJRXDbuB
hQL2jSErq5AzhyfXm9kSojmKkZ+XwRuHrC0y07hMIWOcMVF0fQ1Z6ilLGE2rzHCLIpH2SAJARH1D
YgiN2uVHcpNlikvgLQ/X8H5g1srUwQSdB2qOn7hJko6pffi3PrM9/lE1NH85LtHH7zMiTqDt70ea
AY4rMx4fQiskp5exNVET7f06zc8Jsa5fPUrmBAIsYE9+vXtUoZOS8csFcPqKO8r7X5TuDYFrdtt4
ujLIN2l39SgXctKMRAt05BobwzIDilC+PT0g6D7fjWh1fUXB09JqSIWsjVyI7pGX35bT7+bRVOGI
q5eHYYE7kaTS9YYVgJahPdfLym8hXUpreuQDpJByuydTNArhQLW8ghEMvJdp24+H2w4a352xPHEb
nT0r0/y73UWIT4wMlD+r1JbrWpkpKYrlYO+9myTjdXyOzf6m9LCkasmP8W4K4x+M4Fyi7PBFfc/2
DmnzJRly1WjQp8oIj7pmfHs+l6+KRh/DMzACd0c+V/pFXOL9JGc8KNbUXt9o4L7/TX+9Il8Sr1s4
dvAozerAC248U5nxl3aKUJdMO9qeyyZU5YIXpz3HAsR3AdWs1g6lI9ggqJqu15ZV1f/bmmK9dAPt
ukPc7JIH5RKqsG3ZKLCoH9HdeB3dDOWTWSlr/Ohw9TJriLljHPGSlVJFfUPw5Jx/1Fk4qNookn9l
96GQx6udQAVnKwd4ARI7flB014aWL4wc8bop6kbT6r5OJMQ+zQzkSASvGJ3xauNDzEJIqun5U05A
9DQ/LN5eVI4HRci4CaUeZfPWe9YaALR42MfPqDdvBMot0obpeMfrHr7ZZ7SbJD+4hjRwrn/2SgB8
ToBYVsaPINT+49SuYUYOm4kWOzVGRrltltQuZiI1u+7ai0Nesf3Fr5HGXSEKIKUjihvVS8eU7QAw
3w28purnQL+xreVuDLDKTaQscRmJEz9Gpy9Ysw2NrcqawAeI5ugJ3kzOmH1n6Rfx2FKsgRHuferJ
rcLRIvW3IAQNqssqc3LDfi6iMPsJtnm4uDshisibiBZeVTH8fS+8+630JhPfD5BhPJIyn5kAqnTs
O9ru5h53CFvmdjAnbKzGspMpAXkQS12Zee0ZXD0Yq/JGaxMJdkg95N62qdUfsw9jzdZATYl53z55
BOzG7oV2+RzemLd8zGG4EV//3uKeaC1glsyHkM2MoqtPrurcbmYDpsATR+8G31FErBTlAL8GKuKx
wQsmk3Qp31USY+oL7I2eWkMkV+6DlpeVgToQZk0MoP/+rqAXz/gbue1XbQcHTAHJw8H7X6N0mZOB
TglFEW78ZwLkt+FL+XAXIOn2/c6V17Ok7NzPDc4IQwGQGZ+RMlHfRJFyrZN22G4T3nbosg3B8FS0
HBCRSD/iTCAqY92YHlFakkChMLrgbt+ceGiVDw8gjfrnYX8FqbwwzZQeevG5998IrdOnJjpk8m5h
0ucuAQZRmA+ORkLiRdR7sDi9uRVFd6D5dGMEkbaHkuOZreeOBzhtj0jA4mdZci94QMwudTxbOrRH
/kPKTD++R9QRqg1NFiCj886DoK+XgEb67KL0yJPYapPBENBJ/RaP3G/scS3il4KZJrPUA0d74i1d
nC3v1kjFbnvYKV+aQVPbKEoyaOLJKWnH6qu+s2RLn69fhGa7+wuiW8/mzVetfI7dldgdSWaJ1Vmo
X+03Qcvi9ODkKaPHbehcIHCOjRP1Z8rNu64qBFALXHT/qkOZVVv0ZuLi7+7N5vaWBbyVzwNx31KV
j51cUM0cP6IUPCdnZrSNtdkVBDUNy7rIqfJY3wd01v+9WhPpcCiUwA5qQDVN9JfJ2NzsEbE/L8gm
FTL2BT8Jb+rTnLLlJ7ugo5l9KIQ9McGYjwKIvmEKigrqWtZxMSed3yFKImC0yYZkeYdBN6DhFmYu
p4GIfHVsQ7q/EmvpSnnb7E2SleO2/qt7+/OJ2A7x9fw8QKF5ETu/fWUaBVxWAhNrSvxPAerqIDZj
MxDhcJabQCoAOKT9EVvmYMoLuHVdOgz7uTokNAIfn0GNYeh+ROGGRhxWp7uqBxo/1/lJuT7JzfM0
8OiotbIeW6Z/AdpNwexByIxwAfSWEeXh91feAxsXRt+vhbGc/tJOsyLM/dLC/iS737jHqISBRDrC
gezkfsllIUcufIUqA/5kyyxNONm3bvduP4fW74uFpbr2gvw5Fz+y6UArPGd/QKVCOiCnZdIHRkBg
n695UfFXtQFLm8iAwOaZd9wmGAuYNWrrDXY8xTXQ2ZWo5FlkB2rb+Tw2wpaYG2nLSQRKTBfGrd63
EUiQRbTdnR1X4xmWoBQg82xwglLF3kn3b2oAwHsXWZjCmSfNkFvZe5AYsPU3UMfj0McDh45NBbic
R8pCY5PNdywqc9WgnYDlPRMhSOnltXA9MIW9+P6D8Lj4/wHzxByNvt8BTEwCmwaIAa1e7DiPOrpe
CUbqgjrWDIggOK7YrHqoR+6udJNaWHNsRhCVpDaS4qO17pEFWv/9GH8LzdrJnQKNQctRsu17Rxqx
O+aXMp3vn5HEkxVQEUA+mezF4ITKGnxdkqlgX9ZCvkabKi/EkadJHVwjY+eDhicsHRtoFGML3w2J
7UOAwrgS08yd3BLtqK9ZEAyVRJZ4hFqOPdGbwqQqgM66foX7k4RaxCaSI4Q0wVfRyyHLV430mQfA
BuSiOoheYiwVEgxNj6By0sRnfRKXZ4uKr4bFNnKTsYuWLnZs3dn77g0gn/dShAI4PKPDKYNzfVum
wBTsi09WATNoxiuPWbRTPbRj1xqmv28jOBcQtt6euv6Vxi+m9k383y6FaELro42LcrmyvsA5bjpf
U5zYcSQMrNdqINU2Xhjx2S0QCix9s0dpwSkVVsd6Cq/eSKNelv0/CFphHn0v/EYncUt05Yel1hqe
fwhbAK6xhMOXlMdtJyFsU4b2grqUS3qeZytTlC2WmIxKu4q13Zm1Tf05A6VrjMBjVUipTjuLMjFA
8xf4eROGiRV36FkGWSOtExkB71OW+Qthx3hFjc1fkztotDezko46GYpNklax7PpeKkppOAh8StG8
MLrTVN7j9iHGkj1LN+2gMi5FVqbEJXSW5M3WBN5DiovkPSq3OA1wEoYm6aXdsEcptQ0hRNYgkSH9
xOTnfkDu2yjrd/scxstEiCd9qdcH2CUBA/2kPXFk+zZ2REwccX+Hih6ua8PaIolc82bAdac7LXVg
hLnvRbUcWRtcIiTnn5zQ5V/t5XDGtXIRhrLwCXrN5F79dKRTZWSAWA98SET7FkuSra7LHOfr1bl0
D5MAdqSnnpoY3n5vZK7Ymw5ouVcuQ6q3Up//vbGXmPO1VMY0ztVXdoisvmr1SsRdaFD1ClMjrqv7
9W7DZfGhsUAAJ9f8hDp/UgjohUm0xaPZjf6zycufOhkkAgpDwzYWJ29YXgFjoopYFcQ6688S2OMw
/+EgU6e8Vob3D2sjix3+MDfeuZl9B5CnkUMfuzHIY+62r7a/DALk+a3B2xJtQOuErIdh7ykwL5wB
96XfhzHTZ4k/Ntm33L+nhxOkrQdSW4fGOgu/DalLWpElyKAEonEpm9axqBjffAF2oX9fUXQ+R0Lq
kT50UBnfF2sKA4q7O74Fg65nT9T1daa9XGE9rc80cJ4DND6BN0Kwi71wGq9fGyGOGv/n7gCoiljX
EYYx9dApTV3JKtSxyhfgdy3cgwB1Sl/5AWsf1iPXQJStXTGOHO3Ctudcqq08EuBIVhqcd6FutYS/
S7w6GMN/JYjo31XUVH6b/79lQJ3YLI6q77XjbOMUo7xA0ZwUQiyCuo4bSm4/IJ2cJLciLu8Hokyv
ar3OOjF1Y5X0mQKbFIjMp9+CeMLtV2uc3XddYZzEXtudbk1FoFtVyPdAnRfi1pyQOzNIgqyyJxfd
zbGj8sx/Sd2AunkfH4NEc/M7+DZKhJpe6DfL/7GspmgI9AEgVrd9jR+pmWOtOB9EP6pf7Dt4dloG
e+2lE5XCuk/ExXwEJxBKZvvte9jbSKmoRQlL99vyeOmB+vmqogluF2gXgQDHiX5xWWzBhxmJhTq3
ckJXmGNoOCpiYt9UtJsCX5TkUmqd1NCTk9AUBYOYCKX2+5px9Odd5VKA4l7z0g5lewWO24KBZZjh
ak0pUwCdhlYv6cQeF3Hd7g9FMobA1GKCw1r9o2tYNt7UK9/C2udGZyuzeImE6IivP3HbQTO9wTX0
eJXI+PnRKMvm7UAlpi5/ZzSpd0rbqoYpk9mbWVZf0yf8bxkNnk3GRhl/gPOeQlT0jEPpPcUATwdc
7RdkGT+VESX5z0ZBWS4FBmOSUDFcMwbC3Xle5UI9XqyUlDp1u35I7owXNm3kfF6OttwY7xPDgcWs
SHpdbEU8F5EjvFMMD9dcACN1+kF9bOc4LrrsqHor2713fBd+ml49LxtwakSLVqvPrMLqFR72CHX8
f0QOwJDVxgP/5INj2SGcZiQK08JS3iRB7SxD4AR7CMPOtJJuEU05mAsW/wzQ4DKOuCann3W9GI9c
4TqhdfK8V6QyM2Oc7X+r6Lh/UH7H1xoW50AFFX5zz1ghGmbiqcBaZVrZTtQ7uLf5/kPomaKN0pvC
Eyg75Gvp0vioLecSVvYp38L+p3IvwgnwPzW+w8K7t8Seq/hf5vAtHw9crm3h2A47+AClY5nT4YyM
jnAfz8m1YqfqIvMs5AtcvrL47efW2UtEVwBOQEmecH/ZJmHtErgsnzSaqltyla62DgtiKi307EMN
aTGaH7iSd5agvP4CSh3SHMPsCXP34Av6wbS1xhgJaQv/egrusAuBDE+wDaj9vqsf+pfRba5j6RIW
i/N2C+jcEzf7I52fZTcpbD5hXgRz1tFlu9ZIMhf+KrPqnr10JISQ30l+mgZ6HGRYr/fJqPsqjGab
Ie82rB+3HrrxpN9ZaIqSLIGQLcFGGWNFp0UYOg1oUEUVDGw/xy5kbL0gWUvpYN9PB+5FHldi/ED6
o+YZ4VeKOWXWpW/0Ltbbrlfm+5ERzg9qn2lt4Bl1E/s5NLaTHD2Rq++l1ZsYmfXEFaUpeERB320R
W4KH8kQdliKVK1Sv6UOE9lIIAFYelpqpFuOUdeOS6xtNZNzggRif3IxlkCTHMQsiZ8SO7GjEMTAB
S4CzjtGi7khBmiJOlijG94vkCAkqMjsLx6yIurZRfQWfjGmdeK59dRMEuOwnRq/5e3hicOPtFjUs
XGD4FwdmeeIUlWx5ENJ1YxUuCjuDmbFqr4eRFMg2S24VfMzSzwjD8Bfcsm38i10PtN/2vobu4xKk
A5/7QaVioKQC2Rn59oCFaZ5oxwE77NSwRfEhuPWnfaxz+qifY42gHgw5Tn8FfjXdtCQxvNa80eHp
jZYwz85zAwyhRjaXU9x/sEZxMeekwGk6Wrofnl6G2SMudoLa2JkMEd5hz2uxbQ6CXHgffHVRWFcu
F5aiNovPkYUbFTsJAKBL7hsN+0ih8uz+5St/IrDJurruBxeWnwqLoL3odHWBGfyvqYJBqaF5UZ5e
P4xlo+K/w1LMXQbAH4Xnjf0xkztd/b9nSPHsJpjGYYBjnmmnoP9TRNlRPvth7u8orPfOzAcbHcAA
GDwKetRDDGJ5QZIbyZd2dXd3rkOM+jJkAqb8+JdpSskYfYn1P0b7stbvQ/mfb3gaFu0wcpnkMzFL
A1zer+LzDBgRmu7frzvGGX0S0wyJ6AfWLJiO+ox3bYucWnTxYM3fNSGBO22tT9gmUOmCXoA6XBcV
ZUUOiossy/YGQzgNS8BQzY3OMPwdMgaWZF+4Uuku4e0jcN4hk74FCkjBdAIX+GgyF1t+WW4V2ymu
/ouY5ffEOWyKt1okoeQo/2n6SHIaIjohfVGA2fRdBZGB9PmaRugM/3AFwgehbEhsWHmLepyjmAel
NSuCvps605YssVCUvjrQfCA94viLWRVwJr0zSFaCJpUrXY0fwf76E2NGiX7dLSvW6HdE+OxH5cTk
/WX5YyP/uXg7QaRkn22pWlwG8MmW6Gn/tdvJO/I99Lb5BxE+tL6W5ma204jBs0god276yMlf7+mz
vOvwcXRvcR7aWiQgfppH9wg+aImtxfVAe+JVOQJE/UHLADKRWVqo1MszbCfjE1W9aA0+J02X9LzM
HDIUQjrPPokN/fnvutbP7uWPXCg9Yk/s0birr0Q7sOk2z95clo3CPiQTFH99L6Oi/+Tgyx5TALZy
Mzo3uSaC2IOImo4lY4ujQbi6hATup5w4SHn/d7RK9BwNkh8LYm0idk+PhdaCcO5TBlysqBBEXAzB
3xgsN7m5SWmzFRQ4au6J6KBNo/OBHLJ5kuQSF781sv4vziDqIZqbBhvaXqxM5ngigoEDKFHcCYK8
LqR+2I7Skhd7OzoqBKQ4MIoFIgyuRX6Hh3SHZ9zTZcsi67v2ctjC4GMfJJVwrEfkw9y07sC4Tn8D
tY9Cea/ZMWqqYrHvRbdiyn+Er/ghZ5DHA689KdwX5t+v6gFfSbMvWck1y/1U9uLlQABVrccqQzgk
mI3dQnMtOfxebOS07fVZjwf0hTflbFON6r+GBrgf9v+Xi4z41Loz6oEyUnv/9RglcGQNlh6PcOZc
hLoo+0HY8NUAVYxTPbDcDFgyLSqJ+I4BW+e5SB8WzlWv7j3fwflz77rdljIq0LkgTEgnVA2ePe6V
52f0W/7jRHb8doBYYM7pC+Yw4V5w4vqQ+n1y7FwmlPEkzjHMAU50gQ67+BQcjz444IfUmxLD33yZ
g9ya3UJrPWZZWIDTauEsQ1mWBlCfHxFoZhUBS8adpwqh90dGYd5FWok3Aq4d50dEyXN2Y+h5aiyp
un7Hhollq8USaXjKKcRJE2LOMlvZnq0OgLTTM/uMAZigCHZBzDt+AisNITfJeN0bwbA84C9AWEVW
1vma1FtaiZldBkxD5nFgNF12iVccnGrlaU5WG5Eyv7K+C7ClXu+3yYoU4n4yz9Ij2L2JxPhAIZDU
t1Fl0OiOy+P1AiPKeDBl/25qlI/vqodH8YT7HV7qPZv1feMbxwWW4fSiOR7MgSlhcm9J7c5vlfJZ
3+P9F0XuYJMuaYg6x2zTHj05BYHwnHWQL9HabGIus1zo/Ki5/M3csKb0FvlNJCgI9lTPw0O7Zmec
GaAjW7y6aAaWOz8GI1cZugswIRUFfJZpGCyp5flVcJCMTJ+R0P22YgJpzGZtfZ61HAZrel5aSDc1
81XPKomgdf6OrQ9HauTO4bWe/F4icAT5MK3ABic7z5yaAiBRrCHKlP0+1tDFBk3lh9GSN+XI/YUD
cAlp4M9zwvIFcrEtxVNeOurhwQV3T6MklSXPfB9FbLr4ojgbxbfrV7RXk+/InJ2LEb62WdJ/w9ac
BolgVB4o+CmEam363VCmEVmOMQUKhotcVRRgyzS+8qA0SBwOykEUHy3cFpQSrWTM6tbkqEmQkCdT
7BELCtG8KrPIumHUodyhRtSoY8QaXdYjvyhWLR+jvO94ugK+A39fA8agWbU5B/nkZhT9KqBzMJIX
QnuOvtdCSsgSfZCGgsnbyZhLBX1ISPyJuzi3wv5esOWNpZLe+h4VxLmal160xNwMSkjLf//MUn7D
3OqxnMVNEh0mR5V8TiW15ylHsuaiURs2MBo1r+zvxYy2YGvI/M1kpmRSaO5O2D06Kemh8l/UU0Rn
lc1A2CPZGjhk5pNAE+D8iJM/ESxFi+tts6amsujI9R0hArobrC9aOPj2ejJJ3dL8bGGmNFpZ3LpY
H4TzwMOYzzEVpsLrPfB4pvln3f2chvbgEh/nmHw3rhdyq880jhPecp1/AzJeDbuJ67x01N+CKNzc
0oJLQBMSwujrV8KwU40InBXX1ZROdIRXzmlv+PSB5GbjoMOoNjirbDDzE9vjnUoJt6iBnUfaYSNZ
4PBTlRRJhQwFTnTrfCGkHDi+rm7reM0p8K3ubNRRCpmBU2BauyeBstmSw1zRNMpXovYdxxYDJSRg
uYMtQNjG29TgfkTI4B23wbOL9GvCX7duW0DaC8s/5TAQ2dmN5krywoK1VKWQoux/KCv9mZlHMq+D
BZPzOEb+BPuYgGfri//UMMU4n18INNnbb2KFPuV16NPLFfJpqajRuWB9UqwFnGgvAozX3BhjTthI
Xv5AX0OLaurZO8fGv+zs6DRTniN4z6LeMNVY3c3IDJZFFy7PXCkV0EImjjOpoSix8t3IdapyBPgO
adbXi2bJiZt/eIifmBdfJqFxnVGnX1vVdVSfOHBE2KrOT/feB+kwJCetTLULslTvcvK6/QEVCO1W
OdR5oGId73y77H16H/Dnbx3VWzNK7Oh69MbaDoKcL6MVsy98xU7Mdpci761mnJdC8FLnRdwMXNVd
Yu1wXtzXI+zwt9KKY6zaM86c51nBtQXoSnVbcSgAP/t4v8LGr6BhBhajxZTF3p7JQBPJCgG9MCPl
9EdwNCd9N5fl+Xh042q0EgMSr81OiBiinRaBhEZtXZnr1yZ+MKaAEf+M+K6Wf8z4MmhoSCyEmZnw
A9koOGsPlYWlu695E9kLNzy4cs5JIxyCBU6KmdgwwtGb6VDlGnMM46e7V4ako5n/6PPVAhWrR3uK
ShPiWJZyz2J2BLKpGuR2kGpQyGPbGSlpWlMKdT88fseOKoNm213JCHRBDQComBn138+dTOgbQx3F
V1mFWmqp8nPU8RbkNcEFZIGaYInZXGSs1AkMV/RRvvopNWU57hocNHL5otUErGAwkQ7Mj3AcMm7g
hkuokj1+lbqIyMJ4WBvxrQhzEGt5vKB0EcUYosYspnOQr3e9kzMa0Y/Gu6Lnd9vSW4AFUrx61JMM
a+inzR5Oi+/03bd87VSVVziVFBdiJ6y66bQYtcIL5jyy1QJ23VXX7IGSusbZ0kO6Vi6+gluYKBbN
51gS4FWc6I4RDfvnq94MxQhYNOXf/KxHQXw1PR87OfaeHtRUO0LlpmgAq9MuqwUwHdhCSvKtyG+D
eQdhat1R9BmrvHWmPKsjS4CFueFh2hPLf8Igu1UxL+0RizTzRXJDcMtbIGD+THz/O0hu/OanWFBT
FqmbZwukbAmTBmUuCAw5fpTrpL7WY0gwnIIIvTFVdZvIrjSzkzXnLgn4nGBxzLRddvDpv73SbHZW
fBt/LSBj+XKoLXlCW/AuHx5veMp4QbJta5Jcq7wa5AdCPLaken5Wb7Wh+sHf6jt+JtKTSq/RH6Kz
00dke1AisUSIRi510wjsCF+uGwaJC/bMutBo+F/9p3Kzhjj1ht1iHkO2ZJf6yeTQY7/o4cKTJDXS
kIrUhoOwlyvQ3rv3JTP3okCuU3tIBFYZhxbc5Zmn4VkI/PSvEB1MD1yPwV7EJNVXKaiQgF5UUKUi
nCk/eLHp4RDeyoIkBdtHgwQcAzoFmRNTzQ1ZII2ItUWzQYxuxYoyXcAAoeoDjbntAKGGb7eCrpwi
vPdKkCSwK9fIQdrYJIycHsZtwNebbtdDpjyMJ+MfQvIM8tk8oOeybvk9DqxDqNu2alubl2PLIWmK
EgZNCDVmKithbkLYz+2Ijrpp97FAfVxaGcx0pBgLXe+j0tkhg74B4C57iTIfyhm6EG0QBWJOV21Q
xOgEk0VtznE4cJA6qxURJErJKC+mR9NXpcKaV1C5M2HCnVX+fP19JOBXXWW2r7bzyKM4Fkl50uQn
1LFUvRDiexYRIIzK8uqHiYzsWt4BFNYxqz7sitkHyDIqVRTP0Q/jpX8ECOvP6HsvVAw9tT42d1lm
hpjLtJq5ptdL8jZtcwSSGlzqAbgrtfMtTv7y5Wk50hLxVJKnj5gKivUz5PrOW0shv9vZLcLqNyTZ
i+hNinMeW504Xm6MOrx99n7LP4hBL43B6a8sYNAun4E6WtgajF0/01JQWztlO39eVXvnGQOfdeFY
rAodAWQxDumgrI/B6gichRK4MyI08KiID8g5R0ny+oZAk+XD5Z70vyusyDKGMHKpcPByDtOoF7Y4
W3/2wkMx7E75AxaPIifEmoyG8Cz2OwO0641pNaXgLWVtqV6kpJFsigI+k6X2VB5h0cvP3G9nddtz
LUPAta/OlHue4tlqYfaG7Yr0gOesZzHlpD9vVbPDfOgkM+TMNbvBKMaPu6b89Nx5Mjxss/gYfYwu
wJ1KBn7grumcErMhXYgr4fibChFgv8S3A+FN6K4apoqv/kZPkIwL1ZIz06X4hhn1c3Yeu/5HxgKE
QKYkvikfSClshqxDrSeel773zLlk5pTsytBJfBqfkpongS7LC41l7oJcG+kbVlYEhRd74JbzioxM
APaDG4DBtjkT5DM302N3dbLm734ViRJI2+O9kQoPpO49PSpS6wCXpofXI5aOkplFYh6Mat0Ajo3D
QtHj4Unt1WXwYWfZkbL944s/BDt9vXA9CgR6hbIHoEpVMiC4DOkoR0K3WSXfb/0LggCp4xFmQkR3
wp7s8giOdgBF6C9vm47nyEzNA6KWNKrsewxf3SLx4DXGd4tidgkY8wM6eSsWqgknssDSRkOjsl4S
pTSRI+PM5oKQ2EGZlmAs3+oIRwRvyF2JKSnywGSTmP/FmQrC/hB1fsPeyMaWfbTx2JOwyOvPdHoM
+brrv0IJQy4Z2Ma3+NDzQHEgPnEHcQzmdWSrWo7eDpyKmvrh8WasfNHZqNLJVzt+lhPtljHzj4Fr
vfYrnd8ntfjEvjh62PkTLqwtVLU8Eov74uJRN7rWqF1YRsccv3FQV+hMCirXuGfg77JFBWpwjtQH
cK4F07GTY/mLTdbFcKIZNdtVkkyLMP8Q1s5Na0aFZgOzzZjqB84XwpHCgx9VusL5Zxay9bbxsSH1
D8i7OVDHbTMVz+ihzxiTBEeWbDvY0hIczJu/YmmE7C0D+3ZibCvf8faNiiYyhm6wci4NZzKqC8Wa
cXMncvDcSMdiPgQPN1BGK6JsWz/rKVO7/A1NgIgeRmi3MjE6qWQ2OBVM+23Q03xUi3fViNvnla1q
zzeRHkpbjCz/pDdQTAwOzJFVnogv6zb8Vq2sBaylVoQvsfIuMo3BWaj94jbHvrFwLtAZuOuhxAuF
g0fqrSU9+JqzqpgnRiUi1o9Oqya6JRz6UfXpR0ZBN0VT2CcrLMJWccUAehMD/OskDlQX7GXWyCZJ
A6/jH+eu0Kh/q3NwLaNXkLx8b04q4fLn8iFTZEL7Z5jR6HjHCP9PR79K4Oer92/85013WPKg0qT7
kdAer2B3jDEfqD1UzZee0gtWOBm0F36v9fU7bOZHk5UgZa3JJAAaXiIdsVfDLYoyDLbiBnYuz8xV
vjl72BtkJ8HmeQrxMaHbhxh8giMuG7pE4fhFwmYoDFmQeKjdqcoyObfw8175rKLAhyuWn18ZbCOG
V5jDuYoaPu/TQSso0eBWeZzEloVnlnAxX1wu2krnt3nCmVhlj/vYLCc4gnJfoDwBz1m8D+ZuSp4I
fdq4RHDEYFJRGJAKFimgN3TbKSLpAuXZ0CiOJcEvCJihyBElDe9mM2QzDxDNJxTsxdXV9Q2rwtsP
HwmML+sw5akIcHMwk9YBxOqxtPttxOXQ0seoio+4V47NyI5fIDXbm6Sji9JEsuE5KqAxTUEPhwq8
XlGSaTcWIVrk+zSxwf1uBfyQeIDxfzbpRszL14RoD3tUrS4lf7RrcfN3+OzvJ1ImLF9F7icttfgd
/k5qtGZsGHq6eSG2XGgd5eWPWr7KjJvzqhIAPNGkLX/9MleA3z2gKJaYPJ0Zvc6jYejFZ+NjkVpw
A0qiYhNFa+W5sUVft2SjvT3EMZaguOS06j6ILrCp6WrGuNriamSEhRSzAYYWdEtggm6ml15hLxA2
9NA7PwXlyvzPpjJhj2B33T+sjxfHvsnH9eQADtJleMgoMFjgXJX3VfeyPZpzDEP0TvAtcZxMvrjc
rATEdYfJY1DhKBS8hWWmH5pnhWDpEG8CuOeb5wAERZ39dGzA3PyP4a4xiq4yOFqQ6CX0ZE8VQgMz
cdp5vj3BihSklUVyrg8+vMtEitvJM/ba0BN+tO/hyHoIt6maz4NJYnlMRWeqnmbZaEcd0lO6j/fu
OI4UfQA/oG3/ZHU0eLwefUrIDE6FwoGZVnZ/oBivfA1BIZEsYiB141ol6tLVtt6G2s4HyA5MFi8k
odJQta4p1FE+kQ06mvMatI3VqCSES8PqJYKIHqlcCzgalrQBnDy1VdwQfpRNup5G6p4aU2i930fj
nHvdQFvDoN5xcmqJ++PRRwnLy9DkrnuNW8FFE4GkJMyvf6vMa1GEm4sxSG48anOX59F5RwazYBnT
bRn0MxvtqMTrDxWaSWHzRydQOgTRseIekExzHQbV/4YZc1z3vkPM4VGu+YSC6mQIlgDtuzmWmns/
aPPUVS7LGNvj4Xhm21A548KlwVRn4MOSqrIBW/ptBF3ulRybfwPZpcr7sQ/4swel/0MIcNjcM3x8
Dm8ikI6hq66D0incpqgDwQGb6RClB2TBbiX9eEYpMeUQiQ9XYjaNHbNiGxGNVGcmYVb/d5Of2PqY
tE8wlnvowQ0237sVUogKAqIy8A7noNM/ub2b233BZd7d1KCJCl2ju/YVnA00ZJjOQwUh65k6wk7I
LkxdAIn28CGrCH87aDxTTsqd7AOwMRJkXXsq6VzgFOARziQlPJGL/cPBqAY/Tx852beEG/jARx/U
ZxvPTrHn4eMfetJ1ewtdeTsJa+bp6SO9cSe6gl2O7QrkcETtc7hS7iRBSzEQW0kh0L+VCoJH+55d
UWpOB789oX1UsKOUGSMkd43yzxPkkxPTsqcsgi377V3TS3UJc/B7WX0e5USGA4s8nPCytGTFZeF+
xyHH/lUfre5Xm4ucczLsSz6S+i+N7V5Jie/Emh/lkMo3vyiW9zmOIJBZdsenqiiskTXqKuvEtLgG
fCuM1+s78nIUwdxHljmQAy2vtkI6cfzCAj8dtC89MoZJ0Xv42niQBXKfRdiNpjwFj9OrzN2flidh
KwXJe4ijPLTy6hlflgSb22Dl6P4YzQbYF6qc+16ksVzXNUlJx9cxFVDecWzJHYWAMkNAPmuTzq3T
QvJs2T2UXDuJPeOkz5l15UGPvUfFmJsHg6JG8H0C65YghgqfgF2L7ApdIUvws7kciIJREpM2/68Z
XdXOELachdSOv0yq8mbktv2cbwPXaY03u7QWGQfwrW0J/gCwG3XonJi/lnQXdcFzAZDfw7FTG0E8
TvF7xUNjBwxj92QznKkDT+c167j7Ls9CMPAMiyDUjPCCV/b2CJGT/yNCIOcTSz6EpsnD3Ziohcd0
4VS29oIfO+sfhAZz2xlkTlvDL2zg/irg/PGvawwA6xLSIDu8tHaVpdKNjQ7vzDLcNU5726McCBfd
5EkuwHKJ3SsLlHFVCOq66KvwZOINNzCIpCby5AHyBI8FBxt03wEn+/WE8Q+myoQAvPDUaAK3L70L
1On5lI37QTpNk+QDIjNrnQn1eU5hlUuXpTqYBdcVFpPP1iiOnsFtZ7bKILEjcFiBztiPr8aR6//B
VnP4eqx7u/Und49LdCJrddY7FfzUbCFTpoZ5h2X2JHIvAwBBkf4eqS9ktlvhElWx4RwVnQxwBkaP
5f6bJRPNlSPpL7LshJs/oAYDImtC2bAfrVCNquITJlohhGdam3eXemB7SCJnKeMmxHZwcaUWDNDM
p8kw19oPOBd3zm6uKTqbpKSf9o0i1V1/TeoAx7fI6LSdQ/hIkU93ipTVHdVRy5XXx/qokUo5cC9w
7PkvP+Lg1vHqfulxPJEaX1M+dhXJbsBX3ZAQ8i3EgiWL/nvOeBqUGloCA7o+lL0vy56ulEYJ1B0K
2MG+HE5+Kbk4mQjhi1fOO2xAVMu+Y0cHOsUfGp+XRQ4KSSoKid30FPkQnEk7+Qv7PpVCMtlvnSpM
uo+Onmamdmz/oin1r3lzPDyC+1ipkNqfF7gPDpxV6iLBxBW0nC2TuEepFREWkxH9FcpyuskLFkPh
1/xTycwWAaECEvuiNwN+lEwSHy2oe/+UXdhV943rvvNQfTzQ3B3HE689934kSlUYgdQeviYIWezd
UrIFsq24MvNNRh47NJ8OZDpf+HJ4C4GwVqfdYFclP6b3qUtk8qMln5l7iekcWlgImjieBUxQCvJq
s7vPYcnxXPUQFGGtPiaj8S0A1+TsU/67DpYCucaozqGTwEyLLpvhKhIf4TwDNZPjvz5eqie6zrKy
XUAj8jnbJEv+gebAgtRbOXPZMfxFNpXYAEoxBSNes1yubiLkvQe92nTe0HbpA4kiCdGUY07VwJAD
v7tepAr2ZtK7eP8n0MojsaBmwChNnckfOZkS6/5fzL8HqCkhGzz4ivgLx5lKpqwikr850yZsy0SU
Fl0vCWs1Pr0PZXlDIOHOE0bSqQbzIsdh3omitaZ+swct4hdOWEbGUIsBYsPr84+G6Je1sl+fwLpU
Q20o80SSE3fIqKWmIjZVIoEzRa79skvRnraLx58BqEmzIME37ssYjv4bk0DMoEp/VzSlZTPZGNBE
poj56Z9KTlB/BJD0uVJLsJoFuXc6l4z6hq1vJBe0xoo3n9hEDA5HF6nhZNPpXjyZBV9KKVFbk43k
X/qd/PBgKM56+WDk711YejYA9epJHocklXE4ZfByOE8JVGnJgyRIDMNZYNEST2rqejL5H+gCTr4R
ONUULq/z1enhvt33A4B2TeGgiEcUCGswBB5QyY5vgRJ7BKDTcWuCttgz/7d7HXk3V4RE1a9NgpBi
SgxUdkBYafui7no1qF9hlrzklyOyALls7LxrMqZ3OuQ7KaJumqEVZi11BOahmr3kwSEnVn9XV98z
BTz56jijoPHPRFcvs58NCepfKjf3e0c/O7oNXqpbetRTSFd7XmHsoa568abGm5A2vA7FQTmpYuPi
ZmgtIDoVfd31F+8xeL1R0gSJdfYNfQZDRMoXqfqfskjatzF5UzGuwfWxfeZFcHO/kw+3jjSzzeL4
473ZNiA9vwLA/x2SHpd8o9TBb4Qrs453mbPjhEO+G+i6P2uoU7T5M3EavJoOzU8HzKVYakEevLzv
u9zj95oz61H6VkBOQPwAVd32viYp55q74yXabUXDfGPzfKU63OSZqmDy7qsduXJGHCdrh4yYI2RW
Z9MjZtNq7IE6VbBVbbBLZG6QKWI0U4se6bpDVG94YhupCDf2LeV6LXn0ANDmkPbtXbx51L4/zEuC
S/frxOGYq9yz38RVAUv2TVLJOwF20oWQMVLyTWTq4H6YVkRIcmGg20lRFdOQDyzJA6pz3VBZkHzw
cEsKKuFsGG7X55olxDUwRl9Z9w7BiZQlSqSfQTlXsI7qL4CoHJ/5nAXbg1TaHuq9GixMRQ9wnoG8
Yx1pzEfr7DXEhO2kPo/3e7NkgFw3IuevFq26xlQP2HrhW/kgoXr/aaOC+AtGeL9epOH3P3z0dLfJ
eXevtB+H7Q/jf88RkyfKJMvb+7ax94ddSMzNFNTp/JSwin775JeJatwOC7eCo+WkihoBNgffssxc
AU63Ycigx0LWbwchNQTsBLu7bNMURpGLAGkXNjw0hb4sWUzyWShGL3TBcJH9Zezi4tFry1v+6rKo
KewFJBAR5VQsaJMT22Ecakhw1F47R3usKeRc/f0yo01YjSqb9SukrzxdMvbqxGT3hWqveXFZifKR
ff87hxR6T/F5X1+AFuVf6qP83gOe8lIXcX4J4CtHe7z/I5OTMDHcDaglD4pyvkYxmn0Ed/yPg7+R
1g17Wko8QGdHm32WW99ZA1uLRMHEFMFGqVP+/MomMvqH//vfz5cpdRzgPd3wVgsi3JnUJ+li98mE
EuB0K+Dv5yPo/pdWnF9BvWlWeNfn1L5ka+lsujPxM8/yh1gadoQmFfx6rXtZB2lFl4lcgU259XDT
xhNRgHS17+X8b3MqEZp33N3R0RZ6YBu8H3KJo+Rz51Lv469Eokw4VX/ANqmYJJhUphUpYhGX+eTA
JgPApjwx2Z/uvj6AOYxggsC5P8+OcGj5hJDVX7hWLP5m9UrnTgpAS57Iy34ZwbE30J6SHAYIpe26
gUliO/D9uAgxJfZCMCo9ANMslBMAukpl2c/JKhX5ZEZAhk9bp0HsxMUEaP7QehZgUZ5TwiouPC20
mi/BWOikDDwKY3e2Sk0K9pO7cq59aSOr8dYGNzUsiGthaSTT1k9YVkUlj87nvGO/xx/WbPtGYe5O
zIx/Fazb4izP0lXNmdKaMyt8EtPsDTc1AIZtPGIHzBWfr9SHHBDy5Rf15Nttp/fhG8/hSRE6Uxlw
geYV34WL6s0QnRyUkKIRKXzTZqJIzf5xreW4aDdOLe2/WsWm0GrdBirC66tY1JOy1KoBKGaPAL/l
yRx3LnW2v/Iy2vnCmPSKSRrXoOuHeX9D8/MbaBthfX42VzR3siQVsF22Ux4xZcOIJGz9lrftpTZZ
zy3p4GzJd9LRSObKSWq8U5siiM0PWjj1gKt6QnO2WiouBQn3rqVEaFXJxRh+uboxOvJIMWjxKvPX
lPxzNQDi6rfMfgnJSADdRjhzHIU1r2rQhAAu8sfXjxuUfIp4sJzDVsy//vvBQFjclVIfe1NI8r9R
jBL2/MR9WEvYVib0fZgi8TZ8vrMvuFLJXCO2o02k/DQvGAz+qfH3fnoiTqHof0uvRyzpFYiIJvBd
aGEn6lEG0+svCR5d3HtDfg6nYonvQZ2XnKampszfMgmJkACWGbOuTSXo9TEYnowbeZcbQVnARz4W
CaP7q/b0suJSFBoT3rxwOiUVq4B6/Ruzl4PEPPMShkL9mn+SmUQlLEQKD6HMMYRo8qcySIo9WogP
xNeabG5HDpSDcckV6A4pJ3sh0xApV+0H692w/8AxH/Z+Y4/xMqfPqfQ4n3QPJk/9jK05I558y8xP
iHreI5Pv+igrH1Ik9sqtKtC4yyRKTAbGAL3G2dtk48VrvDMaW5mZXcfUuhMd2XfIac/7fyhGUjsF
Rb3z+mv+X6Amfr+AvIj9lVu9cAR0jzlFjYtPTzQFJxLQsc5YuKqA52b7seMkt6pzW5m9A3TeEkA9
iCkUKZYRA50aQhq6e7DsxfYPkGHkrH9gQf10gk8jLYsGQgVX+x+Mdk/ZtL8YuazkHK3PghrtrAKQ
b6UGURJ7wW0Rrw034mMmU7eM6nD+8TvJV2+SXkCok/wIus7U6FCkHM9gjTD7Hnrvi4wrxMLn8QSm
+ds0ukTsG5ghezIm1Pti3nM7hDIKbOC1i6YZO9rCxe8guJvLipfIyaL4diabfjCMwIgbbuJBpNA2
Pc4UpGYNgjumeT775MudYf9ozBPsn4CO18R65DpDYdCjn7vU0fgr9ySxjEOMfnksa5UrXV/wC2v2
MJVrT0dWNus7B/tJCXlmAkPLKKZlPRNAK04WcpliMYfV1Mj3Fb+Xnv5YKi/I70HbJ3sVwko0OrEN
AZJsi4rNXRahC9/qB4/d8/2MgjM3KYw0j3Ic8IlbKPdV11OnUBTSM47AiCR4D0H6/ATUest3gDHr
O6ifj89HG8LkBEzyDhvK7YZVyZ06AeqzQAop+egRG/5+xkcJ2y/yDLjhCdSv8JkjmxYpBmUHctkn
bsX0ItAJoDXtqpMc4ISODQDXyjGCbf0w54oGuxhOiQH7o/KWyD+tP20IprRhU/9RxGR+FoDL3cU1
iHxXhXYBE4kAHhnL5Ayu2/2iJobXnxHUssBDd/7LWJgwsyOMfm1uqrKNjYG/+2vtR9ZDgAmESPxo
A7FQVG7uksNP6besbfrNUP98XICp34c8pT4ddF2cXYfMxSNBdX1T50BAi8ARqnEGJqLjBBKQrmb+
DAbHcCVhMe3HED/36b+l4wReJ5nqxndsen2wArldO5/NA+KcmG8cNOzKjKLsXsx4zKtk9KQs2GiG
SRyjCzpUGr2WXkze6tlsedtMGZXFArfqVVGvo2QqSbhcA8KwrXB0MIB7T+xz9vyLoNZuqbE2WJ8q
Y8HQf782FQKIDOMWc9lRkuMyL9GSlh32GhVbkcwANNXt5Ojk5klqTau1euQY6k74FasIDY3f83lr
PMibMh73dFHdDRkfYPUoX8c660bq4ihbAFwsmB6kBNvpuphPV4vnc/k0ONduYyjXLhpJX+CCiYQ9
Ukw7rJWIks+HWKleXazSzDPJNCxpEYU1L2oBFFiwiKEuos3SNh9/CiqwB7BuDz7wTcK+ghD98sDj
ys2JFWAKCQvPCYoLcy50ZN2na5/4uqYzM1HcLJ72lhrO/V3IliY3eG42eufsFjjTObdae7AAsuVf
nvJnJQGO/dvhvVlHq+SMeygkYM7hRFVPtKIX0m77lkJyW9clzTQ6UgRY573ZBpFXbaWATs7hK11w
zEjIJ4HLe07k4bJTO+RS/mXTIDMuR9SnktR94Dm1q++XEEjrLC6xJuzHBAn5G4nV1AESsmFvrcOI
QJSrESgXlX0pY1FbQCGLFgoZBqD6OK0hhuFdZ6RTrK+H5WMV2BhJeg46fUC62nwD6pgQauu+qdZI
nPPd8AgxZWPTLLYTpOf82gmU4/v6x75+Nd6mt8PxFZC8o7LXTC5KCQ7LKY1/aWDzWRtq7mnfkV9r
/VmNkoUKL6t6/IziSabhcMwsAVHI6oQU3fopY2AWHRBVl6uRzqAyZ+BZKFr1GZWrD9o/+itnbq+w
6aqB0HBYXNayS5aPuW/XNVHCQD6JuPRAu02UBNGJzeSC2tmqCF4/qSUIhjB/Il+Y1YsI213kfhLO
rmncWvyiRNy+8Obp1kju99TQK3FRVEjlgydZ4QZ25ao0uLAZTSm1IhUHN0eYRqrmXGwYsuEq0DZL
LmMlgCGmuxW3/rMpKzMJAXypVH1GeKRhnh7qXHBfdoCEhgCC4KQk/lPgD2WiX2HpJQimzCwiLI6S
Pic0GpoJjt+x1lB4hDcwNQbfKtaszN0Py1L3kUpXz7IgwNe/NOXAwPyfVmbEoRtExVHjAjREkmam
3Glxd8OLf6R/7CjUdDmO5pX6k6FU5iMehpZektk9Ke/fckRIcm53rOW991Hw3QOAA6AhEpqDU1UU
CSte2g6cubgbvgQySmfwU1/GzNz/0n9qsgcil9sFEzwOzTIecQedGm3vBiVnTlrmJB8D0FLiRoyb
WnC91Yj4B4bpGAfebkjA56yYYqfGT78gF2HGI2+Wy4QiWzTNclnZeGQrSV0cOiiuEXvqXUsxm76O
lvMIZ0Y5uBms9RlLppq/H9UGakMIddcKZ1T7DRTiyJcvqjzRCRJS9177sjQxiTSFXlDmV92xYJds
CuKgRdY6E8uVHNnrdZtCLJhF5G8LVsYoAu9nZOkusnkTHBVU2ArQu7ZhUnNYf1RHHTJLWHP7BxL6
nyQwkPqKbON6ikv93p2EeU6FprEo+MAKEmnTOR1jY2Jzl+pQ7/vs8aQuukYHmLHMG0PtmOduiiEP
d7F1uJxxExihhsVYn/3RwP+ZN0i+3McJU2vfZwm58elbK0h7BW5+88N6iX10WRGzj7gcTL3czyDm
guhV/HB9MlWNey0NZMYtZvQ0W2FHIL5ldzOyh0/Qq2s+UeheHMJDj1IHbiE2o7JQ91O3ho0FZh70
Me6+eOz/E7a0vbxHEM51w9IOARgG14GaTeLDXArzpsb5WPel52320myhpCWTJFCpftRRQ/Bg6S+0
+24cZU28eSoNfpvjKj3peQWJWNoLeM5i/EVwGLhVUW59RYXBOebRzGgdbc1Hzk3JvDQ39gCBaQvz
xVspr2/jL+O5ajzY63ZTytx89YzOyYgKgfCk2U/8dCYQrQwvrm/wWdi99UFSxXaVXeDlvGIHZbAP
rOL0BxatCvhbgLR3yTHfn8HdVn6HQWmy9Iu11dNZWe/Z3584WX45kH40fGw2U/JcPcEIl5t1lBBv
WKYj2VRF1ve9XTuNGZMGzfKof90AkD5opzHtuhkMsP/hQ/Zcx1TnkkT9oOndsRMAQCyikbiZi+FD
mrXJVmRjxKtCqiJTmYIoqpDWKfAtCKYqtlCP/5dgadY0uRxnSkCOdOhjNfg6CDAthxqH3nzwLXLY
jRD0haUviWtVpiytkobFo6WhGG9RlN93OwGam0L+2BNr30UUzGWyh2TTK6RHJ0PDR/7PFUFdpVdR
UnhD56524Z0W5OaFA0a8whVV26AqXvYIaR2u9rrGw7ubcz3+x+BC/z983fS4UI0xQUnC8y6N7JZI
xdifNjVkf4n5IEDE6mvW0u5YRuY0u3Xx6Hv5f/sDjW1hNYvPvcozfsDtdcpTODbujvMkTqFlq4ms
I8eQMm3xvZ+JiAhkMZC98WP3d9F2PvcLrFdP+rtj9hPd8g8Dni+qgps6KFkLjEPHNSEzn7XvjehH
DTreDx3HBuIop0XMhHKkd+0K1mlSCWErTkOu6eL7cP5fmNsl0XKe3/LppdTyZ/H4K4FZLbJYnbaF
NxCxUHjWLNTuu0DhIpBDWyDMON8AcypmHtuB4ibiSfzuzAGnuPNFGnbNW3zz+v7Ze0db0k3eP4KF
zcUbHBkvMQylTkpXIX5NIYFdWjp2yE3SWeUqIlux3gBxyx1lBYhLqp0vEHpUn8zc+i9jNInM79Kh
4vNC1tT9TlftrhBs1ibX9HuGY3NWFDNWI2j5X2hyexCVw/+hGiGUKPO6ff3/UA8eCMD/PT+XU1n+
AOBcymAiKUEO1xxUQIlSeDpvVwlz1IuZ0wmxh4YMUSe8ApOZCxObg6tvumAnKFse95DSjMeBo0Be
zuVamZmV/uBd2/BOCRS6ACtjj0IeA3Fs0RbE1EVEPWa+0CKyWyFZkbuxvg1Sbu615pqcJsp1eeKF
TLeVTHNIdpE67ufDtOpAWxgppaYQtZSIo9v4Num3OT1AHtJdnyZDH/UC7eQYiF2oVHRjGJb7i4B9
ahV1TA4VPlVCRyXBuQa9mMahJNyUgZB/9Wkh1lb9V7tq3/+GiyBj6Ez1rCdk4vhaZuHbf9KLfC7K
vCHw/+GRSk5nOXMYzCuofHyp6Ppxa9x8yWqDeDK/KtX2qb2l7EIhohIQCygQeC/jrt2CYguYK/Q5
9Uy37gOj3W9GCtCkEB3ikwZvlx7x1FppcSV0gMJV3BlUdBnoamzlaYOxEXyNXzPKRPIhp4aMCVlc
1vVadTaQCO0dRQKhWzeggG0aX5RbXbXRdJtGzAd3yepBsyQ3tFxXBxLzUA/D4feLphYlDT5shr29
2oDYVr4MIiEpXh5BSKCq+Yqk+T1KVhyznuTiL6Bh7GBV2J+PQRpwv6F1ppDDYA2QPSNGubw2cz2K
vx6ARBO+cwjkLk9DSlR57Qe4DXcw0BGxI32obuYxG/GnFDKyVwQbLM99WLRXamueVqAVt5PZRL1x
Y+jCSgI/iA0fRE6ZtG0UEkXbO1D6BS1v3C7dCXCZ9QCr5I0+I8+0S0wv/lwyOg7grZLkkajx1y2D
CSIrdZHpx/MBsTQTkRZslEK+MESUDc4iUimgLIe2VdoZZXsutFt72LJM/whVWpQp0635N/m1xwe3
RYTCfoat6M5kyjDHihnjzAyzbflXhrrVPDc+JCXi4LPb7YLF7liDHhYYFAmYXj8FzehqgxAFuEQp
jjcBRNvgrJ9msETq95sC7bK2ZZDkgb9e7rf5n5aLTj9gvEFibwC2AFROkX3IxRJgRxaaES3mjcXs
MD5FzD3+NgONuHHhlo7kumCH3ITCjBYjpEA4cDUHu3zsauLMUySyYrYr0a3O9Moxyb4OH+JAIblR
HiArPPG+pdI6Mco/zFPbkSxlIqA2Pt374l9D0Ei0G7ndtZPJX6wu2LsCmowpMickKYuFhj0BfJj2
Dd46zJKkfA7LLH96kHJxbWAzaFDM3ILRuQvVIebHf+wQqYqx6yO0bGR2M1mtYEG4991SDYX1C8kn
+b7v0iW5H51wnm+pm+FjnrKpOwXp5+XeoWWIYwHThu0heN6eaWNIdDh59DA6iQF6DuBQfvNkkOCm
bfA6hZQycdaLz7UnTrcNQuCaSQyFpnfeFoodkoamS7Ju5H5w2I8h1PaVFrsvhYI4PzHrRaZXNtYb
rwYlw/hda8bizXG0h3YTq40u82X3kVI36uoOiYxtRnXmymXY4LYzkYEpfXmaYobOZFRa4aGjtG3D
mITZyzs5SMlfp9ltH6i/WvvXUq+N5R3N7lj9jTOlC9Vey3XFqOL5diWOvcDXl61VGhMfE8TIOJoH
TfuftEFktWGBNdqGXPcxnClENt7V27jmJO7/rZoKeRD+UgcdBbDcxgKVY38//Px08jo1fX1gOrDp
StPxLJ97TaIH7HjmkT9wkf0IhImS3AKFmiYdesCO4dl++S/zI8F/lCIk2ZR6EgkMzY2KhUdTwEY5
3cWv8rG3aqTIQl63waL1AIE7ftB9b4yFWY4RYxbZPBOVGtHbIhLHk1DMYlvCF/vuwN81clSFDfu/
PiqjPGt72s0ax7Nar8lcVI0v7XsmqAZ28ILjOIWTBZjvfHA+2PB7qVcFvtLx/R1jyZzt3QqdT4vQ
hIkVZgVx+ViEnJhJiXfVQW/ku89huGVHviO/knvxThd4mlgqI+hvKcUdLoxdMgIXyX46pX6xkDc/
nnHfWAGf/na6vr3Hbg0kP7mgxfXJ6Nf+AvzADahofRaHJDxO37zyfOkpNLhJoB8cOle9co2eIKFY
OPUXzr1pt9UYzjguUFsOR5jUWQyca+C5E/6MRFPiUEnPZVNZUrI2hxoRJfvEYjc2xEBO+B+b4sh6
N56dwfUHEeOB1eHi+73hhEtkCFXAoCVDvRZgMSCZD+Dr6RQWDxSyAQ5iMYhd8ZqSTYsAE/53kNES
u3CKxloWuaiRFlnlJ+pq4/k61nT3m/DBmVEKVT5zmMUFKpXabKBVD4NXLbB0XCna5qaj94KKejqw
dpV+cxLGLqi3JiPYWzBVYj93tYJI8IXxp8YnvDtStBeVhtarDPsnuLGXy4jGUp8PWUHXK3uBhHgm
WqLkeQ1+H4baV/ZWGGCauEvftO83sWu2s//18at4dfM/sLmoL4dxRtRyKeMYTVjmqYJuseccIq1O
GNsyJLn04UjNvciRrzK0t/uSMA0CVF2Zf/F8+TjVG/yl75tZWZ4GfEDSdOaXwJONO4cpemP8DsIk
EpBfdCgaNvsDeqMU6HOlUu0gGsMa/0GJbivKP22j+7KxZpwPx1FKHXeyBwmsnOmyycG4Wn738sKs
03h1Cwak1QZXVxM8ugCEMaS6GTSONwu5Jl+Xd2BGFD+1Rf5XnnFiElZqMcfVq2+MUDHgKKkSTSPF
D+0kfQe1vIIGrHuRD/VqX3HEWKoBfo8c18iij9BvnVzY7LpCiSYW/o7fpVhlCz/dukr0Td1yLcr9
Eddqa9L8Q7KOGZawGiDqGET5cDrzXveOzFgldYjDj4WJdwFbtqnama4ZGwi2/nAJqJxYqy99diJf
xYsoqfhTW9EPRQSDhSyBbzS//Potzn4etlGWhTXBY4ukRT/RwHgPoo3LjdSezU+lSzgom+22r4sT
tqs2sr2ZuL06Pb8iSq7KOJGj1afeN5q8rlUMgaFZMYrtbLaxETvUXbDUR7vG0OB7K0Su1d8nme+j
lSJERqLMIPQf3CgDBMRcLJWGyRo/hXJTEBqvft5AtEmOQY09gmmWS349435JaYcvOdWqHwKib1aM
eTi+2v38sEFx6sne0aZ6cpzoVXdXFB6xz2nLzsyU8iwbpGifN4u8Hu+4GphepvoDsYsrA7J7Abtx
DpAW74Cv10e614rTRcs8Cow+8zFfTc8dz8RdrbaHcbRASjfqG2iEQSecr3WaG2Lz7dMzF+OcD0h3
w8lrhBQNpNVXvmM4SU28mXV84tjbaAFx+3vYOGbl65i816IuI1ZgO4YS0/1rSNgtVLTcg8BabVwK
FilW8LdBsQWjWNz/Nrs7q3COEQ5yOWz7D3wIwRF5U1i8WOvUcBv2xz+ajls9kajrmxrm6XIX1v3H
5AozhQunbKoQvhwEugPEc1Ix+nfmJNeNufMF96jJMuI+T4F1p8c7TcezgdqtOewGbkhEgIepu8bm
az2OG8wa4m4J1jaJ/BasLNmFFFHhz0cQpnI8L4Jl8A5PPLAs9uaoSYmCTgKdlBbZKH8GhV7hTVPe
CfVdJOYv5eZjPC9bvtOO9WE6sD4h7YUFQ6UM7K/+RrlNutU2pT70BXGspAwXzqN0fx1dAzEHItlr
THb2h+Kna597FvUieOsrInx3hAVgT2FdoAzt/0ubYfz5XB6kfsmTmIE5b+eJ+NmM9UZfAN1GY0Ym
hPE9wlqKldqHUSLEOD6Nqfa03+i/R7KAbMgrtvXscVly4BtR+t/YRGFU3M6EsVW8bac3vJiWqjwR
J2fJk74pHs4WXevCNCGg/ZVVqscbkV00rG06+ueOPC7FNBl5GIBFiDqv2IsDH6eopSzsK/uc9sfz
TlJxYDZerphwBvZdKIAmmlp32PCx8WYquoKKEJMZsctuuWRPNdzAOzv1uKH2tVeIsxQOWVidXiQM
O4H5m9jabRHIn8Vt/uiBkpujBmLoKY/0dM8ztug14dlumu2MW7UlY89AH5PQxLGz4UCmslGmayKl
47SarhmMfbs2DWGViC8DyvSjUavrrpu5N/mOyokQ/IGIYCSrVLvW5iPUKvjBvtcArx7A+98EC9BA
KU4ZqnUcKccBpiwPq5LWGhwqmddYPu++9Hx9XDwnbs+Ji2ARi2XgDc/W/4z2XASExhBe1qrjb+1/
G+wtP+0cS/86lvD06JQT9H7XQM5PJEZc+a5Zp4PAWqGvXLigY2Rj9Rb42dWh6IB2CmSFDeShAeKh
N2KGXlESC7p5S8AgDwVMVyeAWbdumJDcnkSpGCGmpXR0unViIEfr4WyCjizRziZwMvz52KsxxnVM
1DZ5Nbfxhw1BS9EmNQRtgaTyQ0USxh4MCeO0KwLoDsSmXCx9omJKkZ2bhsEJMiT9/z7xqrngFybG
TaN1mqhZ+SDpp3VYOlXy588Xsepcmuw/O/28rLLHsIx7mlsm0HXaQBy2spxFeZz4DE6NDFBaapxk
79jQEs89YsjpoVEXpv1a8bCSFe7vKK16xDevDRFRq5hL44iBhS+FV/rBCZtJ0Fg4lEIzNxuk9Are
Bilzt+0a7t5qlxn6xRUWCoGzYi7GUpp7jjOhOAkeJsuXGKW6uN0PAQ5S8FxyGM05UksRJVpGln+k
u4wsEZ0zS5jNeej6QY/ByZcrVzPwriUtryO8OKP8//WXRp1UBsJAytxt4LdAgcbNUzNGQOnxxkrw
Th9x2iYe9sROnd8XJhu2bfH3sMw6kzW1RJtaxwGuMwAM8wqNI5709uxT5ZsC1uJLhEGGNzAzGBG6
T9DHzehGr3aUR+pE/NR6zbw1PNYOCQvTiA+v7bHqw8SujiA+YUE6zginhk3sJjXT/YrPG16slBoi
aA2u9zYj3nibju/wJRdia4+X1AfMvoTvnRp+Pj0M9E+iOuTajmm1GhecY+rN7CYl3hhKxwueJxvX
k/GGP4uKBoU17wz5NV2Vaku7meLel3in8DKvNvXmhtht034p2XvdL3+/A+xu/6GveSrOKGL6g8aE
O8zr8YnohMsG9iX2/JVmmA7C0NBBoQF42RwkDG8zz7WQj9hEJn97X65UiUB37chXVEx5EHj2E5QG
3jtS7HGAc/a672qb5WICerMJrR02dmwsGD+jpxHBq6jcC21l87YAdnACB0pioQjjwv0BzdoXhAyV
YJF3biOshuU0/KOWTWK6/ZBIhNVxlbsU9ved5+OLEydWmQ0uYR3ACyQj3gI6tkE8FC1o7JJDd8DA
o1IMzrFa5DNG47/3RsuZz8vScu+KXJztbXrcFkx7JyAbpvnsGAO6UJvjFupjuB043a3TaigiNhAL
u1FwmBpG+MHbGgGdAKTom9Y/eu67hVw07FsvUVOXKH1csHqSBsdqm+1yov04FfIJbOeA8vQOSu5/
bASRQWl7YTwM6Iu0fV+5sSKn2vGkA/tBTr6FLT4PYDQwZ+r2cLZEJe9tQSRix4jr7teQkwd4Rv2s
UIJLuPeib7S3bLyW0iutDbSEPHbwLo0GboJgUKihJESmDr7l/zqLLhoBdSqZYevolAXPNecvKEcG
l7y0g7a1Nd/QiDw51PbYXO1kIoOnvuMI2YTMPvTiYl7xIOTNUuzCEvSt3cqa3j9jL1m3rNPmicRu
2UrSOL30TiLQeIcqbYfMRfCty2Y5Bvg2ydXEz2aF0faho4YMHr2fZqoMe1UwwuY88CnNPynmBdF0
Te4wipsNEERLyprC4fhhRAOYPIboTfs9BOVsWintaEmfimzqyJL96koAH1q4Zr40Cw45cDD0q58m
H37iNDS9IOnWh0mcP9lpIRCbxHAyZ24U74yL3o4DTuyJk5r9GB0+GJtTSCxp+lwu/t+gEApkIez2
u6H96DI8b7ZWdheyQmXryyvX0+oUVmsIxWyZnkxaNShhFT/zeurUx6LHfhCHDNJ2iwC6SxGGAVni
t/0aJpDpxCT+657c6hOGoJYnFkbRZAI7ojTZFiMBvUw2QuHsIJfNOPhx+VuSmUI76GpfDGUy0Mp2
g+NEniUhdJMxJ22VKb6MiowlMBv5O4fviriqpiRd1SXMJKDmdLz7152vBmPKtyYOXCxz+4pwgn/y
fW4O08m9YehXlO37HSmJX6bHTqViFa7xI9+HTbv+wFGTsa8kF5MMtowbW9fkbpGY98qXt4SIcJ+B
Bj7wwBo9C3zhsDNvxBFhj0X4TP6Ar/Xq8iMMfy6BypO7CARFZkcAmL7NJ6XnFdWjnkn8bNpI/0Gx
LHzBdcFo2c7RqwQdiclI0xIb7zYc1zoPJE7bF6snT/zo6V12w4dcLqKrsIFasmcRrRm2VU1I5qf/
kdI1LksuwDvj2du0eYewRlFGNOOOhF6//Crp0T1z/jifJYFeg1ueyijEDqMwv5ToUCBdoLeb2Sff
bodLI496yOiRsA0J9eAQJETpQ4jkhqU7vQG6I0nJI3SDyAFKEizYL7rd8N4UXeZB+oZxYrsv9PHr
Ma67E96IOJ7x7SEDuGNOVvEHEI9cJ1hzPXh6zfIO4KoX17HXGrEipMpaPqoIBy8Q3042025JtmX4
6mAo94BEwZLGBV42IjxibpfE1+dAXF+yddihSNtxl6gowbmf9vLwCCXr22E72+MyaAujad/7TzOl
Jftw3fmsJwtN48uXp53YpRu+onj5cwLyu6cd/vaI0j0ThPQlOsGmqJXFThL739ufPRwqKjn7E1SF
XJCstvSvHGa5qg1Vrg7X6fXN46ghw3/2pKR8q5qqet7lKf3cSEDA27sI2wGdK8f2m8FFvC7phM2d
kIBbLdiO/KNyt2ImAB5qkBlITlZLsRfMdB1xo5d/1iJvIBnml61JQycODiwwEfrz3NC+ozEj3Op4
MopCw1oiq8XIXkUJsm2/O04df4gGjQ7MS0WBkbKYDnz4sirgA/jykXc0afSAmZ/WiLkaQ/4R6gKJ
S8pnSiK6STV5OUZKiHf4V+YqmuiIiJccMxqxEgCB/3sNHd6VZMcu78t0YUrZcEHEffDUTbluWX3t
Zw0XyfZPOUv92nVVuG2ir+7ZtcKJoVZsBUFkMypvwRCegDFBnc6EgvqEmyu26X9FGPfWXvwM7GXa
gir7o7kPwzkSMoEs6SSSsj1EdA9YBVlVjmBx+KYEnoE3unASXdPSVl7hRskv31dDoTAOkgNq1q8n
PLF7q0aJ0ggIxlVguzbAi/YBWD2H4z+l1B3uqqvvOvJSIbAQ4MuqNynn3gIN5yteGOnUpGOb/Ga7
JhZtnJ44ZgZZPAit3B0Hjb+7v00SKiCmx0slnzCFFOMl+hRR493XuVB4ICfLIvJbliW4cLqzScyg
gpot4tMvQspKUeZSFa2Bzg2qNuEi/C5OiEU7XZJ4t3Jvc5F6N5B9aqp8Ou/l7EzUmv7bGS+f0Fyl
zsZyodEzw6V78ypBe2sGrQNiuvRCyMMAA8Vk4+tS7WF7V7JTgcydM+VwgTFMgz9z6DcAmJKitZmf
4GeUjNQHChGxjkHezIRi0pBuMv9Lqd32djflt1hVW14mEE+RKwGjBpfWjm3Ajwev6c7G+xwEEtzI
UOMGroFlx1OnKo4rW1rKHlqKGYZSSTbpU+YlAYUlhjTpfFx9LM6+nQYsz3I21yqCT5qqBEH5eQ6q
Hs9s3v+PXZcGYdtQDOtjg9Ln7HUHxKjEbZSPIfTkX2xcD8/El8i56ZFn1/17GDgM4kq4ME2VEEPw
LrkO7okh0GxHDtPbUVv45qLJ8ooiJxBBiwrRpoQZZNHPWgnQTEV1boLJUR4fqXPkYEyaZdUXmgB7
HmXOAO65Ju/5fIFKPBP/cO8MhPAtMtK/Qe66vF61UhVH3Viawg7Hm1iKV2ppF0aowBmY13DnX0Cs
FRKWeB79SjijO8a/6gc6vLgIJwiJjsNq9w+EiRjnPZHP//c0r5EWk7qj5Yp59VmKXIw3+nCcZinW
Hphpy4aqkIjYeGWDeEPmdjfns6Rxh/TqcRpvMIXokFCeoKlaabHLPjDNqkI/AwonSWXIvrINp0E7
JNCpf4HVzanE9L10eu3ASB/0RWMhYi9blxFky0ANudpQUR9OwsXJbtWpXEgDuUFZ+BVmVQCY6Vx1
M3I8Kni7VsI7s2ZsUTf3YKiq+dGjxdfnsxmg229D124QhUzKY9wq0nJGgrGGODmpVwhz8bsIWBC9
4u5OsaGJOcICn1NkKRAcQsDAEPT2kV3XQBlXP8Gfn1Ejj8QkapmwmiLNxEXDv2pHYbjJ8II81fz/
gMPSW0EJNX5ggySAfStvo69c9cLz2aVPkZID71ORa6pbzLDKj8tOCLX75kWgChhvXeP9naCFgjGy
AJx1AVzozCw5KtziilD42OQZhcYivnLdbmuCFf35IBmfhfeUj9vMdNLaJKtL/1UyqeTdHJOecPAx
dzxT828dU5EWEcNWgv1RQVQr7ccX9PPknAQRHttAxxTX0/hIjb111qodFzNmWa1NNOTsSfsVh40q
x+Rcb4avbDxw1TF9N0XzWcfsujTEypazFjsF/q30G1EStNni4Rn8OahglhdOLXm96WuOyHvjNlau
L6fHQ0rcsmQS2kaOp9/B2xrMtdWgDU3sPzaiDAeUb5iTQmVCRDYUOFiVYX3TB6qM/28pQD+3Tt1T
8M52UtFjbx7pWqLPKIZb6IOv8L2WhmsBK1ufRU3pC2K/6C4oRpOA01hN8uBUhYsFdUJysL1uo8em
ohjlMUyXcpo9bB8nFzrAUE/p0RLYiRagARdhRUSmLrdpk+TZwjbZH2VyIvRchytC+xmlFb2Y1tDc
a+gxIEEWixnUKdXBhA8fQvpvWtUahC5nB8fhvgIy9xDIkIfiyZcUtgqiSNcxp0lVVu/ymVWnNNNm
TctsQDRIzddkxbl8KX/DF4TwkVOEpOZl+9r65YMTHUpP9rkDLQYkTqmZpg/KsCRguV/sUzEAwzxI
cE1aK00uBNkY0RoW9fwGLPQrRyVgJmoGWQD/c3d/wq5ALqnwzjlCGbyvsJLn7pHodhRs3pQ3BV5a
VSfsMmioOeRscwYOVGvuJNLYHnQxHd5G6Qlnci0NqpBiQLRMzZkpK168HYUKo+wzmU2ImF5ygFVI
MALIO5iLqvhN0/EoajZWz/3KOG2zxejwbz8CnJV6PEju3Qu0PnqTNAzrlqctouyJG0GUqB6vJotL
9+n9BQXFa1p/EmFiEkgpF7TNAtm0VEpB5XX6Hc1ZKVbSyT8E5RGPrZd0XNQlzULH4rhSNUFn0bB5
z+tu5hsN1AOBHs5RdphMPWW+ZIJr7V3XhqWqQnaL77P3rLz+8XggnufXzC90sT2vewvmgTAN3Hj3
vHPmBIR0Qa+U0irGlwVc3RLEVtYk3Xzjtd+9v4/SvpTmPcIUIgjokmZO2KlBrxnFf3LmozD9L7jt
gK+5rOhYId3TRi6AGF0WOvAUNaIMgEn3ZUMDbWuPr4U4zYZmv7vuTQLU0OPWaITsqLXRSzI5vQzN
6mhywGS46ed6ks0FL70UANCNR4unDbYDypUf86esPdwILpLyZWq2tYX7fE2tRtok13//Dy761p4R
ORjnVVWFy2PMw7BCW9Jqzi/vWmOlXeHeOwB90+V+0wIu0AerSsnBYVPhlWebS5Iy7631802k1Ogo
PC96e4PBwwtsqV607x0rFuezC89/CrxjvMG8BS7tUh62XSnqlUHlVqGbweaIfFBj9VHXyJlBgdut
5s/G16bhxt0yWMsjTWDmx6Yce9nfIuRJl3m4PkRQy3qwvqheNi+vbCIx9oa95lcZdAlyazMbqwyg
JNB9JU3rBDW6QJ2tVeXiWBlzi9I/nsUVKUsdDnTGH2461dDBDmO6Tg7cl8xf/vY/PBsO+2kYS68v
ehG8ri4i2YQXrPb8slPgOfBlINa3jU+P+1wIoRYc2Fk3cSicW1RVsoQgJKV40L2b7MHQidTCN+hH
vHCB8a42+xYcEI+CZ23r3cKTkFFV/U+uxaI6HHERHZUtd0a6tIW26EuBBS1IkSrLTcxrOiDUAuBS
mFoNifbuIXd0rhRDr1Vo/+oKC9pp1ZnfLRGABRDwWUg8SJR14d/PXcmho1YyeTSRjntLOUuNwXKc
0ED70kbKacOHuu0nnQWc51eeW3eM38GNIqnxdU0bySae1j+YGuhKfvO47jw27doV1VeWyijSaZnu
fbtFmMvlEJN4HYqWMj7kOK2H6XC2OLV6HB/jk4kMneyz03GpLwjb3I1NpZarjBrIrizp7CYtvk19
KkMRz2+tBuR0KzRHKsSTcUAeTaZAe3a6RGt37Si1Et1jZAOwV/joCI5y5YAgA7kzOptGzL1T52WG
EA3WeQ7+S3JJ4jrBSjJxum0X4RbyiE8qcC9eXnyGOicOLwtn0xr/oULpAjLG6gddDrmiy20wMyd2
Kxa9ZTAad+EuBxg3LSdN7H0xBfan0e/EKmhIyKE8Ovw5yJ18KDr8bYuzKIbKtOXUMuqgZakB9Ns/
1XMW1qRYsVL9P/lj0/fNoSisG9Y2QlSRCenz5Leo8/fB1nGLIJ03CjdZLQfWR4toLmJrqDHOXTP4
B8+/8QnEvljGxRrcIvhav8ya11LO/ZXVpHj2VpqOp1pvvKftmGPteMtI4FbpRZ+h2rVFfWVw2Gdi
u6m0VXJAb1EWgkZ/B/ds52FwIvYONjvpm47SxXKPhyA4VyX6JLsr50RYZT8ejz0xliXJOE4LqRp3
c4ZbGLCLwjuBvUSbLf6POfk1dTLt8v0DkX9T/xtqbhGaAAYGKJoiPo0B+YpzrEVE+/0xF3xfWCnE
Lh3QWS/7R2gBefY8irktrfY3cx3lTKqRgGjpKJHBpb5hHcEXoGJvBAIg0hhu/+1pOfd+jApWxcbP
0GaVVs7DodQS6zptnDzVfYEUc2DHgSfjHBn5UhOTcqNdcAmtQuwvZ0vyUfuwiemqOWHtJ/CKslTB
564S/WUq+g2C6Df1QMM+TTf0Cynv88M61iH8VHJDr/yUmDJmKvmHLlaZ4LboFqKlagyuO5lkkQw4
dDuyQwaxNO2LAqgeRuB21lLOXCdz965EazSeWNy3rnVLl9SW99y9gqzRPGSoKYjMuUWb2R5oyiFU
tcS0v9qaJZnj73Yc/D3Gm1OF1XudbNbaVI3D0b8puCHj7vB8ZTWL1JW4WnHRS6PPjQggOzLybvZg
VdCxPv/qh4fAlvLxi1cmjAhPeLMFMXMD85+rxvOpwDtMIzpSVwk0rmjb3Q/rKm47P4MXHxtl02iB
fJo1cSv80GndHqX4SHajoxM0ficF4JFcdMzmCQq3a3IXr9pKYL32MlYTM9VCIV8E/aipM8qoL4ZL
0O/5Q9qZLmmRq+MWFw+VjY+3M1+CfZ9V9fXujA6+g8DAbrclDsnVJ8t78YMfSx8c9OjhIHfrvyLK
ekfoL9Abb0YiyKf30KFvT1P7QM89Jkfc8dTFVVzK6KUba06J26VF2gpjKJJQ9hDlR+rMPUvKMkFm
X2PPmmoxbEXr4flR3/Yj2DQCQhhP4M2UUPmdnnjLKa0zLSCrUXZOOSMm3WAdt00mulBTSM6TAszD
WR3FBppiMKgZnxCOQPuwQGhndBfv/QBI4gCMxSqdSJiNF42FvbmT+cS1Ukrb+W1YgBREkNZaFIkR
2LMMeYX0EkGeRiILflJzjtJA8C+JL9UpaPDkve32A69PqCovSs94iClkmRP8hEM89TleUk5FHUVs
w942s5T6UP7VvZ0kBLXM0nmgdSbJmPEUiKg+5LQtUeauQrQk1yAbLI7jvrsNoh0Cq53m7f+EVLfY
vUxRprEkxvZygoAvmTaHVa6RYlNEeYCyc+9pp9d/xo0g+oNe+C4FsiUYjpEYJ+GkHe69NYpJAB9o
Ev8n0hUtrtQvyFoiTzOwGC95z3qaN5r0a6g9rcRrwoG2wmSw5/3ppGU9zy16kgX/E4JL3UDOR9U9
tJYLcv3kpDe8kLHNcdiD+nffz3KZU7KE81AzDnw1zsexk/7yyXu4MTAUpreBLaG7tKu+eaMITkBD
VCkjjW4GOyWqHjzux6NudkPKJ5da0WdlELz/OFJAZ/2myNC0O/ppihgeznr+UWJ263cAmba6dDBJ
t0bwUV88bEgWZ50Lfx7mZFUZ4UJ0usRYL+ahO/v+tmhi0SVdLqnC4H0A8jT5fcRVS2ewfsa9M4DD
JK53Ne0xULBiPlqYR7txs+u8p7SP7NHcBspn2Htqpw1xWVUpeakblf9jsAT1JXU+VqeAVevWadfE
cjT7zNVfGoJcl2VENpKGlNTF6YcPwuMUp+ZtXtigzwVsasgk6xlwGgQCOvZeooq6bN2b4LCdMCFt
nEEM5lLoZ2lt4ALUyBoGlLD630gTV0TS4AhpFCYsreKD6c1Gl4xSwsk2rbOmFN5e2/y03y+Ve1Xw
rNmvvBO2eXHY0gn+J8+2jjX5T98ujDfQ2TJ/IxJNfEFLqelcsdfdM/NLFxPhue0rJkYQFneldwa+
sHhNrFNIPAkbIN6PXn/qJehG93HjDpMYboMxxfwOtaDh1Vi0w1bppTVKJqFKP4nObq/JweFbcfQJ
8NK98roRIggNUP8iN8EfVZ7mRkH9qJcP5hNuhJRRX/vOqzC3z6DdT7hkPwdinBddlYxAGwopTFgH
EfiGmywlqrRQxTlio3twKEOOFSKeJVKSLfn4m+u5UIkGypjeevMSJk9GFRbzfqdVyPMjYdkNgTrJ
2tbJa9Sqk708goR/TO95MwmmdW/Z+ZFGM9KfJ7NzNGqakIz/0uedbtuReU+CRamtesGoBPXccYG4
h5J3hInvUHGnYu2I6Nm8ux4thP8FRUx/+widTDJ3a2LsB6SJKIyz7IAn5wuV5WxA3wPw8mKHXdkj
CrW9sBe+VAd2UVzcevX0e6Oo/+wUDcEou+I2B2EUUdty7Q7R/GSJQIj3Nrz4yrv+rkQ8a/4eKfrj
wNBgd55gBDZGGrGfyVUWSEhjzdDT1LT0PVQkHqHjjYkFtaLN7xcpGQnB61Lev318oQVF3gBDgPjc
MPAs3FOPEhRrR6fPXuU4cg0gwcO89FqDmt4aK0dTM/+dGHqXmTCk/L8hAxZvZZ/Y34HhEYQ+L/Fs
98+Xv+Xr8nl8fy/YcySoVif0COfF1XV//X8/TvlZ0OQEBKPXDZB+MYLEnkzmbHARfv2O5ovu/5Go
YyhsxCpo78lmVu4kBEF25hnLnV+2b6NMq6+ToyEQ/3Cdk1qYNJJSnb+kg75hnREHpso4OQ752NmY
xzTevUKU6MqGHov8JzCgAlBylZZPosI485ojyJ4gE20VUOua33+21M6uua22guh+R7VmGQmJV6vA
3XggY4xqStM7NtbFEgSmwZQarcUQn9OosOvq/uLg4v9nZXid6e1QzgErKTy2mZltBiNVRk2pLb/K
69+oxAdL+S/IhEyIZVlF7LJzMXl+MMyNjW0OuGyonjcdB558MjnxreeOLokKLJQ7QNg58CgiH9pP
EnJm2F7vWtOLav/qy0Qxs3xYa1agegXDW6c1sJ33e2nDb1IqTXXGzQ6AU3tUOzdyt+a0aP25W9/5
AAQ5vvfTIhEN5IWdSmU+wjqACbFNGq6b6+u9eKENL2Wra2ygyGhAFTParNrB16dcG/2xTWldK6bh
uZS2aEdp+JIoyGx2gUZzwaKS4oyYY4qiBiRe1FgjnldeBg5n9SP1ut9naMsOaVaVmV4BU4bYM6GX
BLbLVnBwut/Z+6VjuNMWeqxbI7cf6d8IFWAAlxTql4uIaXT8i1ToQOg+cmp++PkqkkkIRkpkXmgU
KZhtz5E+wHB/7kbf7S6GLVGi/iBa8xpZP9Nl0FCx4pTeQZsRAnUW3PwG1JVpAVPuddH2R/5N3W31
KENvzJ0UUCq2qMnUBTSMJTdgP/C8dv2uAZv4A/mPlOwCN1bbPEyXBilWk9Q4/LjnoMYmwiOMZw+s
cluCAlHZGqE7GpzSWhoKvdZGXaZobtt7gfIJooR/kH/i3cJo5FpiNUInSQ4XXPosTUpxK6ymMVUB
I95V+quMVqGaCNDmo+VpQaT/qPI9BzN7kwuJn/VbSJyyCOcTo/MsC04tJJoVWUoMW3jZykIh8TcL
VHn9JEa5yKP+A3fXhPW8rn8+yWAXycoQTaW4HEEsrcQ3qP0dGUcG+gToAAOY2Y4VZk/8dUyR8HuJ
VyqkZrC/SyapfJnBHV01i2t9lHtI7o2UOXgxSpHEG3MNzgFzqwB+bGZJObFe/ktGRxvVKK8GL7g0
efBr0ijnfs7t+NneIi/BNrvcNVv69BQe32mRRyiFkgq0ixFfSmSIYU6my5LY+5ZN78G3EyoRvWpl
+5NMOyDrxJyQvTijgIHCcufEQHImElFf41uL59H6IsnZlOle+X1FaQFd7NduXSgiP8ilnaiX0nnT
vKdrSSFeBYIsbXl67FtAfaZv6cEt62/74kqGKwhDAVU68i0igq8Qcn6I8PSiC0g3hJbUNVW0rtkW
1Xy1x+rHxQsHXk9cvPrbqmqbLAJOAuipNP9vibKHzh1+vHd9IfE9xkQTf9NT1wnGUtYiFUJ+j0Pe
Ucz6TlystI7sYyT7BJAa2vBON2xsp5o4dCECFUOYUW3hPGKcQrxefLguf0UBwU7HwKQyH8hpvNYA
Q+lOuSZrDlIPTe+ulcPOGhX8gJF0BFgiSRuWKARFCYaN77p4OLOfT1Wd9NvU9JjSLKAtL7gShBL3
Oi/r4iiOaUl0T8b5HpgMjF5o/DH3Ewxa9Gl/dJbuBPjLE6MbnOxTNaY5dM6M/DnnnudzX3GRr/cL
aATcTZvjbLbwk9I2EfC9Ws4qL+OR74ePUZpW8LCwXKVAbldknGtPk2N/qEu8r9a7ljemPDP4TW6a
wVR97T26JWY+Guh04NvhEHnzqBYpPHBjAOd7N/TzLEFiKRzILsbVgVFX9WrLoyNI3b2qVnkRtm9e
4nIwtDbCBwrNcN2PkRMA1hMNXDbmkwB4fKgZlvAAstq3Xa2MkftmItph1kVHpRbWdnCYgAs4QDek
NI5YAny57VcV9kSC7z/61VatcuuZo28VS2a/dZkVsdDs5Q2chLKsJdUrspFG9UbkpKvADXnRO0p6
fFUdMwcn4s4X70alw6/XvJtQx8RXSOONPDT1o3wPRXl828deHXp9+f8m3fK85yN3Iu2JzC4NtyZL
suko+AuaV6mNbi4g4M2BkW/L1kxfjNW3MqgJMeClQvQmOBbwftsY/LBPgnNPxmIjGW8BtZWBSkN7
WtVcNM8NvftfinbmC/MaNoYcwqH6UmfYYXeXkBHWawVURkPK6yBL63NVAuGXb0WFdfQaN+YHUAcf
BUdcVJNQqX8tdBuuxC++q5jM3+OHHdphhox8NQJHBqiaG/BPy3UCa8i0IpHnyrN06FST01DmQ0/r
RgC0BAOXT/Mb4Mn2706cZ8YcalLmnW0rPZsFH6xE7wbOgcPRS5z48Y5oFHiREflquYlQxBPvpQmP
uRauQAMvAoDJYxcrX9ppIjNkfx8+bSEsU2HzqKzdiElA3rXNUTmWRN4wsRAqBg3hrwk7EG/CfL3b
ewJ/n5CKTbVM81LPNgWzizrYx+jkQ/4q4EvINEoSBwiI8c6MkYE8RalQQguo5Mz7NvT3KH6Z2xUq
jByKVjgxiP7aSVmpSZj2AlVsnjmbM0PkvQrY8lJyGK/cZxOUkib4yPWDafHiEQl8EWMAys4V7J0P
JD72G8LtRP9rJY5eNfz2O8cXkSYkWee6FbuWB27sLjyvPLl0aHpz8/jirsBOKSJz6rfySPWuTJ4e
5NM9A2IUu6ISbdCy49vJpFOM3xeoNfoZ9JCVswVV7oN+eCK+1x3amW68qVGKBpTgKijb33bcSjqE
Pf26vN/aX9NvH56atMLtNNqDythCEsb2klxiwJx/GnzFOgEEG87A6K4q3Gzgf7tNJtp7TzBqPLl0
hfxNZh/9u559ggt/iqw1HlJcK+3WY+HmC+GRCAo8cCP42uzhKCStwrogEVOiy4rhp6YOFuV2ibOT
6A6dACvHogPzqcbBG9mogsNW5zw7f4MJvk7Fti99XGqxVgRLkBWOxh5NeZ02oQ38yp0MhrZA5Cze
yD2rfpFV0FE9THD9+LsvJQqAjRUG8qpHPF+Jtic1Y3RFAx5LoAD6dd8NhvuvvR5i4XhswoDgcvHh
hf9u0AAZA2AzaDnn7y0q9FhNGeZbajDFE1U7nthVeOxPSatP/zNJegogSfHb4jPQI5ccW/Q4ZNvl
9TxCYj1LEXp4s/5JghOvJFqhHI8pcI291QT19E1LhBOHWhOkjOtneGxB2DXVdDKGGmhmZ9mi+bfg
fwUx3X3MzbIuwxbsE/nHMperFrTtwAbWL3KNZ7qMYTgutfWuba5GPRPiBZkwbpM+00ypjygLJWdS
W5nmz2Rs+zxzJ5HHAwMxlPbNIN1+E7pMeuEpfoIEwZX4W21BppKT6sOJpuDZqFg9ktFMKmhniIGw
YF6BvsVKUn9gn3moVL2p6RClrz6E+oNW0HvQBTJQmH1WcPGUkHP11A1bNevSWFHLS1xtjoyri+RI
uXMZa9kOxEbZb+nXACdKTgsg/2apSWEuzYk2tmUYJdaqL0a6QUffiMI18zGblwOQk8bTNzNpB3Kh
CJQNLQEMWbyDNScvgB3qX+n2WD/xaz2Yh8G/kU3Y8wy7lXFckarMqbvpDRvOiYA9Zu7juHiQ5fFS
CwSQVUvmFF5yoGJ083gAE+sHBt61fByEXQVt4JGTZrZ2agI/UFHU+hqxizc1LkxSjcyOSlV1TZuj
6YZ33iul2YhsTfd//9rzSu87h4gcqt8Y+TwgR7Laa8DkFmBrIl17NDXzo1bjfvrfgMhVOZmqlhVi
UonqDzxR/nE6kdJ3Enxge3fJ7242LYG/MdE4shXb5TbW9ZlMkQtIJH9K0GOS/saZ3itHEwDrY5Bb
o4dkznGw3Wbdkz1btMWGEq1Eg9A0X4Yrf0N/EnQXxQpmmd8OwWZLWu1YIAeA2+Uxj8abyuGxbf44
ZhFYdONMQzYauQG5bCiQMHY2od8XUp7Ff3SSGsQDaW0huRZm4dc4M5l91BVv6Ipc/XgeQR2O7VIr
+LXXr0W2MG6u0F7Zzk8pOPXJ9eu/rRw8ug/NelimEsrcFTpBY8Z/JJRVqP3PVE3LpNdGRAV547OE
mi6X/hnzE4/aIZODCcx+284H+kTrUTV5fpjl+WebcTbMSJe//R6l2uhUYVH3B4shBfox5ifuj5Zi
KxlmaT1XEkOpmjftiAHsE2zG/zQ36oDRHfBgsvmgECEyTWdZmeYnHVWLl8KPBB85BTMxy9nxsN7q
KQb4G9djktyFe2ACjuE7rel0tY3l16xkyWEloJq3ITFcbBfPPmgqaDGrrbRpX02Q0XD4jORjDXXm
Sf0PJuOCC0L92xAKwt8qBn+jcrDABLanvY72c+uM5rUa7l+Bm8f0ZRxgZm8Fx1RsdrIUi8SH44yp
09szdBcce2f6/pabzTqx4pQwx95HQFp+2Q89fG5N3hLfaX0zef5z8j5UhFDSv5eXQLdwwFM7T2xw
JQbYPkiRsQTm4kJB0KpsxyzMu9OqDonR6TyoDXY4bhcO6PHpd5OoM5tGDSQUL9G5ENuUn5tQKyqG
PseY4Zzp20ZxOtCWls7wbgFQmQ8RDA9hiahpRo8kRjl3FRKW4vPTkcsRNS2SSO2z5kKYOT3t6MW7
e30j82rqmCtTqzAxcmG6P1d+cQy+qMma9ZQnA8z8WNgCUKcCcqsbCMLzEC/SCBTyEYD1V+SImU/r
yi0qxetGOj2dSAMIbMLKlgFE/EdZ5tHrOMXBS9Qbhe8Fui9JlKHHqnKWLsqYceg9WBc5CF6a4V47
tIud9aZy/Se5xc58vlhGea/WFHTIz/JmK/yvyPcd4uTN33k0V+sltkqhrKztfpDuodC2Ehano8Ni
xNizfXS0mQih/Rc3vB+y+htdCSZc5rN4oZZ6UXAcfcWy6Ynk0oK37qPu3OIH69cji7Slx1u/FhSn
QIcEpdgdV3llmrMM8oflMtIpjnqmvH24NMsSc68lfcOSv+m4P9zQt4QmONNF8yoGz1oZHR6Z5N71
QoIOOSEPYxb5364Wv4StnAZdjNYM5LSP1zCMVFulUKunpaOhO1wvouIMc+SUBvNFI07efc/SbKhh
G2V9IjWtjwDoPDgXRCOoBzrqOROGWdF9XCBRmxN1tykOUh4rIU2Y2qaoCMEv8GsJ2IZpSEDpsKhv
iHuPfVIb8Us1o/deZFZdaP3xmf5t0dw0zAKSoKoOqvHvatLmqu5oF2zTsKfI1x6r+cfbY/YQukrH
QO8gGd1An1ieceSr4ssRfbLrQKES/Hl2smxQa3MC42C6p7AXrPN4ykMPcfK1asHbcCkBlegbK6WP
5G8oN9lG/G+TFFIIvZsfKKP04RAyRDqFmhMyjl6DrYU6hNhJu4uKACakJeS/PLjuswGEUuVt5s8p
9AznNtczuMS00kLcUfw+AtWZ7tVm5pd/3jOM+YUjH12f/0akeafmpz+TmOTYIQXJ/g/umoPrCLvB
m9HFvP909N45trzCDcc2T2RMS8x46Mqph+DYAXCAkaMezz7adD/E7Q9s3aZGSfL7myejQCSc/0WJ
r1qhK/G4C2s1DexnnJPEVCC4EMigLl3H0D8wPD/F2UC3p7PhbMcqtBGXPXGTEcGjMESAkRX88KyX
+2R3INl/BPFb8OXqzYiAX5AY5/4GW+fOSSUHs5K3fFstXu7InwoHSrz331rDSmhnyom16vVz6324
xFcmimLv0+yWmD79s+JT5StkfBJy5bMxZ0Y/l7WX33RQna+NoJCWWP5lFN5ajadv1TndtZTCmijl
H1Wo4VU5L7znlIhmjz7ffu8XHMRcJVJ34sETCcrCPSvJjBYzVV9NXAqDdPmmpj+Xo7T6rQn6g5/m
WkizCflZLuklFZtaGJgyqGwJF08aGC27vVoULSsC8zwJoYf94VwDQVRDQYsez3QE1Rel+Uzej77g
kgOgJrmX7/RqlUyDbvTEINmEssHLZ3KP0a1NNpzmaAQkcHL9RYRqDUZu5L0SVsbD9KEsVQRR771b
K8X4/+6XIM7xQChEfsdjyf6Te9tPKt50BkBG9bC4CXukEzQCcp/Ny9+PlS+5mkopPAzc45PoQP5/
qXMl/4rR0OskwPl0GlnOSZ+UYl9BK/35wLIAFNYCvDUFWFcTAT/JgvIOiVyKQF5c6p9h4QvnUEz0
o/AtVJOQo8NTtf6iwVrOFlIbWWBhbmqJDa6xJPSZR3mxbKxeu/xuQ/RGfBuSHwssRjWnzATM2p+r
IjSAQ6A9N3ZQzBpm+Y/9VTqrYs2onJpFqI18JtXy5gzLjMXCe6ly9xKNz7pSikH2lMJGSzKYvoO3
0VuUt3CqT62RAaHgmHyZg+hadGHqRihdargYYhLIG0OrvgKQAA/3mgtenHYRDXg7ChuyQ1vxlhvp
0WLAMIBM/1PcwLa8LKzCnsGy2sDWGG5e1K504+qzcxwCNuHNdubspgnGuVw9hnUfGb781lfRTHfc
60FRXHAXyMONrNUl33TmV9blZSXFWK5B7/3u6FEXjlQ2up0iN/9/LAkJiuzwUK3jEjDBUc1SPIqH
KS7Txb0bBCt7F1moz0JFr01sIUMr+UjHncC8/OBM9WaL3prxZn2jRcF57mzgbOTCziUJDB1ZUeC/
pg1XVnDAA01V5Th557oM4TGzWSumKGsfU+9Roxy6NaKxT99iZl2F2REKjdKgs7018xVZx/Tv8G/D
s2tHzhiSLqjDFmyZLyz9lelUk63kutyu0j09YOudLlsBvTLRlGUkix60rdX1up/kmRn0CecHy4n5
4uQCWXgw3LaUKozHBl3i/vsPU6TCgdZiTp4mq58iHN138xy6JjF+JHds2Fsl5DMxPtvl/S138wuq
tn8I7hty4t8ky1hNuXtkDXGR1uXmeJ6Pzi0jjOkoo8Eb8tqM3qeIhAOqnFVMf64f92TyuC3nUO1m
P6wzU3xq1+zgrpZrl4xft1oI75rWpd4vPmSA/y8tKhBV1O9am3Oe3Sn8yxRL0d5nhSGPjug9q0xl
0JBAnQAWVuK1hBQSAVdnR43GQoWlMKMWd+TLG0DIwsc0LWiKQihApF6UiTNnzGpLxS6jLGRzsN0O
32C7ChOv6g6YnBxm2HW7FwMniMdIxK/v49GHaa+ORFYYThGvgNApgTPaO5p6SZ73utN3k+8WZEe+
GlLrAHv+XecZIDzSESyg0fLvIgw7SSrXs8j5J0KO37oM0EP29Q1qSW4TRBoJ96PB9TYfdRPTq14z
zs0iV8lJ6l8QLpqhIyuMjSgz5WOJ0s/MOxOZinlaNjKM5/YYRfwXgMfn38p2dTCikY8qC6oQBTDR
pEQqX/QdzdxXIlRJfqObye6iHqJ+jgJyBBgAZCFrgsLMkfkfmBX6w4obJzfj6zKcNL0lZEMXkQR9
yXL92/hc6RU+HdYNHdsrI5sr89eVzlpB0xQ7L18RbxP6QsffedTek/FtEwN9W0M876+bHST4JSm1
BUTr82WUonY4KnzjPYjwia2RE1gXzHJF6QTfePMYu/MaLf2vxtXshQunkxFH4avrH5TC2hre+72R
UrBUQdFHID/Q/+v1YPrLrdrULpO4wGDzYfg3cmBMbVKbflx7xZgRD4bnNvYbRM4AIVcpumwNSMOB
gVqTkfoSn3kDxBxIR6PtnqIvqMkGRoPFDRXcCsxu7vehbsdE047bp6HEhb4stSjfbJaUVkgCFx4a
LD6RXr1ipWo8OphV9SkJU03oZh7tuEgB7Af8xVJQoJeJ/qEDm89I+lQFDdtB3jkW1jgQomePppLt
KzWH1nTyPIPDNwxlu2cxMmKJzfxVdOZNw3KMjmYf56P1DmtUkL8iroAo+ETTlPDocd2irSZAek3T
kvrgRY9F4u9Kv8uWL9dsd+20V3RcNJRYoJPY5NvfjK+Pyov0MPtFnrfZvQbHRprrSBWbnn1HxuGb
nY8UhrQa3RfG7wJx+Ifan7RBnlhApAgpMipRUNi3q9EKWS7waFXLF6clp0VooTJ789T6rUws2yNw
V3CtzV9RUQSom0WnlqIBf4j5CygPTdHGBzqf7KUHW7XPGrR7H3K16aG3/0nLKOGGN7mgpKqbh1o6
b1x3RqmDDhYLxv+LtVBJLnzCA0goqCWhM5J/8Z9scbvkD3uE4GPItqK7Y1hPM79AbYwJPmy9xnmJ
IrgXqVa964E6NZgTsf3NMPvJTIk3L5ZVeRLcOMzSr5f57hHSmrZyGYBCZ1HcIAGVp+FXvMBXp90X
y2rd4xECnWjx1hm6mgYsjcskfzRlzhJzaUu+fDHKToAVLMUb2GnIH+4630oZEWE/rcbY3NQ/frI2
5s7rYvgG/earBIl88ZvV1H2KPlDszwOFXpQ338xWV0fbrYYABFQGiyBcFkWMcjMWyBctsRDKpcVg
yhUt1nSo28wv5SiWm8EnKgbPuGjQWCBA1cnJK49Cl87p3emJ5x7bguLQtOhdEzAaSZCxzPNVhXMe
b5079tvZm7LJRj9IOvmpHjV9YtOa66f9QpFSsFEIxLFfWiCP6izTqVq/aIQ+CGNPJmwVweiKNEFE
BOXu4kxEHD+iR8SrmnB86n3XXwHe6O2zJB3kY8zl04SIhtXNsfHv8W0SC5egTORUWvwXrYzVYi5H
haJ+tU8v2O6OOV7j+xUqm16NYNY+icSTnj6ttxGxISLn9CTiHUOjpFxFaCg7PPGaqqhDlUxGkYMC
ObVDM6LJ5XbPnSuvpbEjF9YOAVKSLXhltghQ4OiR8MyfkFjhad2l4WzlpNj1kem4ne1hUWG5x/Xr
hDvFKaJMEFb1JC7Bkgr4kEDuHe3nhyIwBDdQpRZSbUb9T8pKxypJhAnmn/QFyjW3pDTgZm95PfvF
kELAzvoQzVEBv7oRh+Higol+yzq2rxdbwtz5nPONOET26lBwtUBa0yrsWAQNtw/9/CWXsoIC3XtR
tgfjOIyxenSHGVa5DqxpX+xP7Cr6Ghp17VsfBJU/+EizjpDtaW/e6aQhKbero0/Zomb/eJBVFhql
eZ9iVBpEo/dOTtavvxwSajhBNuUt2C9ViabO/KQHNoGF21IgJS9nN5zwQLdD7g2jckxDLeaH8hU3
xnXSOXWPmryIpg2/a6T8LZNgVzQAeBwDKAfhElh+eDy/feUl/AcQ8px/SlNv1GkMJB/Zdf0yoW+Y
9cWIkC0hJC4t6857aMYsbpaFJzk/R/K2VnOmAJZWbCaWg8HsAeX5twJDJY8MZbLl+eDCPsAoWss5
zTVPTCHZDf5WZ/quDJBgj27CnCBM29tmRIyu20+HlIG+4Mf9BRVbFy+g+fFeSdARfVMqrj0NVwyc
+YDp7Dq8itQxnYqACZr2HaZ3bJHVMcVfcP+9iA7nXNV/AQD6PAjjpYtfiLKZoVCzh0b9o3OpX8LE
iGGSsZQLBh0PROEka0in4XeLY1GWNw9nJubx9E7Lo/OAzQhcN8rNUHvGaBbM73RHUOF+0Dm44heS
WFqbclMuGF7fSK77E1ExYIoWFU8WEtS3YiBktADfvBj5KoeNMa+YtYU45n2tQQolBBQ8WwXhW2Wt
TffrbmCblwoOH7D6RnAftwMJsqihjJMJyie+abFhM3nS2XlrDJNjVKH6Svfgqi9CRxFQhM/sUkQx
6CzsdQdOVpRmL1ahEt7KtG06pErlXl2X8S0McRdv+XdxnPaxmpUZ9TFLOpFJsaGRkXALkR3c9nIh
izij6uV/lY+JumnYkhm2BxKu5K6DsWxnm+sn4Eo6GSThZ6hRslZa3RHZs4OenEcYnCu7FgQI14r9
G3WxSb88Cn+yh+n1PDdY97VGkZHGGo88/nw2KfhIWVilsE7JnMyQ7mQJP8P3LIvEv4+uG/5ovCSB
qGvIR9edwu2yMPrcGzQSRMCeSePK3gCs4Z+cb2p+nhJmrec9zLQHgkDc0jPx5VRYNaXNqdQDFNXJ
SrJcDd37qU5sY+tT6YUjT97+gpkTheIY6jhHLYzloBEzWTDyjdu5xwsgM2ZJIBVQGeBRDBsLGur3
NMiZH2PQ/wafGc7ikt9l/tAf4iEqfIt+3Qi5L5WSHtjO+eZdk3fQmLwPV7W0d7qpnwKE2fIBfYZO
ptkj2LJUxGdZ8joR9vrXaMVsxbM3+thpCS3W3FrVekwI9DiW/DN0qYGVAcYMWzv7LvBb8EFcYMLr
fTdtFfd053fjIVpyHaMzMvWwZO+/uGzyw924GxIEmGKxwE0uqzLwT6/F0QS2aYnnP+Rc9iGtPMCf
S1MfbBLYQpp83OP8niXXrorDa/GhFxp707QTTlORqdbw1Vv5yKATBO2H0oG0MVcrdSTfoCZSm/SV
8ZoOrCddalef2mX+12dmfBG9hBC+IQ3hsDpbPGV1UJ9DkFf4uoiAeHVbUTKxVfD4VFGDbURbC0OM
bZamfrp11lmOehBb8p8ncUKM1eeDrw0Dj2Tyrr3PJFdja/0jzEJbq0RdOB255ceFOd11Kl3nyrc3
J/DLEtnm3DA3jzBZYvq3T81CyDrgTvtdQBvYHC1E2c0HDroRf025s6Qs1l47sqjfKuoctz8t1xC7
XCfxMSnCDUPQsSOtmqbBjVowVFn+RyT3e+3KghZxV5rpchtLx5DIxhN7NPjpWlm4AzjXOU3ARAW4
LxSGAF9zSIm51A+KJE8xp95TpzC0lM1xcNw7XEtO2a3r8P3mULHE7sTc67NUox1htIQI8W33rDEy
R+BFnK7xKX/8oASX/HLkYr3Ys6ylgpAEnXpu9qbJWLCD5DoZE5RJNRQ1xdhBrNYhIEEzEg86222O
3h5Zv2smSd6pysZK1xfDaUCnRBeTbyJPG/zfbE8tYn0ZMPzqQfNXzEqFMIC+wXCWYui6gwyhLXr2
rYCtkIM8jmRD8wNPvk394Y5wPFZtzEpq376HGg3iTJs/1H787sYseEeP9gqk/QObUAo0fkBCJjeN
oLJ+QRQz5uo17wS3cySdk7pXDkDUPdmKJ31fWsRm6x03sj1a6EeyEqyJgJjAYcRTepS3Ggot5nVh
fyh5OesEGWqjAB9PuhhUiyBBDtdmK6C9db7x5/LRQ7pkT5h5l84N1QhsH2AOtRFl6lZApImJqHLL
gul2C7WXwq9EGEAkD9ozS0ydcpj1v4z78la1IY/jYgFkq3PbS7QONzt0zYHUHLSmej41TmvWY8tL
GqTP7iFD+8x1BkM8SZDGtpDG7bweTq1jKaj3fzlIZAjT5tA8owJRAc0t2plT3U8TCTG3qvNlIE0o
hfoURsNq72fCMUWa2gTiX+QRX65Y8rVOYmAflYQCSxDfpJoTmJwPCkRGE6J3DXaL1bSXuw1BOlgn
M4KI987ANUFNxY8KdyS8rTpKH8fIG9PdEx+5uK5yk5qR+e3YSXH+zchFGtaOx0O8JiSU/9AF+Sjo
aC5rHQa9d6nsOyWv6nJqi9JP6Ed4fPzXVdgGivWsu7mWD7cyjH2zzd/fzBrnPa3INx58lP2CaYDG
3fqwnobSSm75/OHoN5RZS6XUUOxhHCrSfQqWIV3C3+YeLfKWtoXYn+qAiC/tIEGPPg/inOt6zVdT
Zpj6QTzGe6vjsNNL3Ae9O2tbYQPcwwuybkDH3SMtS1apVihLBnKeZm1FowEsC5U0+uPEHlj9vUTv
eoyF6FUlbkJEnjAPpIyQwAww8ZJAtbe7RjZa1mkDp0NClZLJ6DrqqaS+T4VVVdTBzyuTePEMFKHh
z7AHONuLIVGpOEie4pMxN5WIwZP66Nvp4fbWLg6UmAqDpH0SglsL+heXAvyqKb4a0aVFC6C+ZdUm
gDIvb8HWbcUxT/Fbx9B2uXXjnQdecdCTa0KguiVg6ow9EiLiXXj9ZwlbIFpyCPhg0QD5+SYxrgei
241lI5IOqFPUezt8kuu8WF8romDRTicoEO7saB21ajTS4kvJfBUkXKqb6QKwxdRP9PcW0BpOt0GW
PNwxInqSYnwPyft1LdoaKGFumrcBs3GNdVtdJguklHj8lVz69MrVBvgCFUVS74vQv7VLD8r1aNR9
4BVpXkSUJ1X08rIVcBauxuR+DQyYhV3KglywOBJcYb9cQIqwSYaW/EnECYIntzG2EAcyI2Sk72hj
Ww3z/zN5+7u8ajeTJ7C5RkqBoqRdbUgTZL2kbntzoFkw9f/hlCHXvMjuFu+szPft4cfCTQrzdM6o
09EjxfCajzZ3O2r7RRccGhxcWxJJBpocqsmQy3o7oJIumvuUAFofLlivhR+NfsNmxtck1svAodmd
Arm7jywRWF/JKz7bTl78iKlBsfVEyKwMURbEwgxyeztdLyWSaMo0xgR6HZ5tvXAu2RBJLSi2CqBg
6Jgrx0DbUXlSoGeQnYCKrxW+vGH4hOzdXoWokcZ6CKOa4fnwkDh6ik+nqfnWHgcOsgnWKryTtAFQ
3Tzeti+y2QMRjcMAJTgWptQyCY3N4H0ADDRCguKgLLBogLeKL/2c4K3GaWHGWKqqNMzxsfZt7PLX
WEH3AFuXHpRQi2W28NksH/SbX1p1zm/HLFbLqDWElMKM8yPGOHm0uvEyAcqRKYE3D3D5HSkppKZs
LLSAYHFmR9uKNLbVd8X6SwXiMjHLgZcM7sJ/HAMz5DqMHSLrIvrAl7u4d+GJ6Oi20xHQQXJgMOGE
iHe+oiufPZQUTOmilrg6j2/gwf98hoTS4S6Avs7+BPyvORAz6guZ2qpGDzT1dt+EtcuEm/qLfs+O
qyoMCGHu12UdRpLwignLEfB7W4DhVdGo/Tc+AGlmUNDesznsKZGYu0QsP2EVz/JDJ9H+YUtENxfx
rzm2fbhV51lSYjLRl03vazwQa0RqjO9mUUwYyQaZTVvhG/EB5Wu3mwna3vpUSUFkX2Ody9O9ALXX
rST+UHV/B0iO22nqOrUMqfS+CajFFoGuXCp93K7m4pDv2/watN+JHAnafY5orP0p0ecgHVMrRA9h
/o9xfCQAX9C45uXg6xqvvZEIG908zIdilxx7ci5AYtMm6Po/zvAMjTzPlHhlDUPbx10qUpooCG3T
AGaD4A9rbdq6w7tuYEmoEq5Xkkaztq5Z/YGv1WQITmIeQo2GSimHUSmqPFq7hJUH2OfTF3Lrkstu
Jj1oZi+V8LU1VQ+r92hkRq8HS0zn9RT3nYOxk8GdcuOyGHcx7arQ17ic/BZWFL/ZWRN6qmm+AseZ
rsYMzz1ZGghsoxsagCVlqEvsBJhAd8qn6x61Zg+pzMKU/bRtbFRydoUTHheZJ6rrkfCZ4jyj023Y
b4X1s5wPmtt8N8Gkk9SB9B8QZse2bI//h5h8NV6KXANg7xqb7S1n0BdwevStyHkmyzr+tHMFmE8H
yOVcmsq6KRVreB6+QXJYzo6EZRdVxK0ELhl9/w5u59IDSlO7MQ/4jHnjno5bsdmQsMegycwBF+vT
8U7YhcgbSPx/1HbSVoQj45taiOEJHCrbzOGtBhbhp6MmPKQXCtOhlA24CFIySHsaaHPzEAJ/T0/y
OTDcjaIlIwjtqRTI7vuzzYfwIedCmhgJgUOE0fvekMLNODbUAXItNGTbGKkOZjrDIf8P6JrNI2rN
EYEi7d/KbwjVLhJPHbrLNIYnfmEJc/Ge6M0PtDAmVVtrg3wKnkiDEy5jrBheumylbxKRe8RkS81W
mOSDeM9tYnItVVGYK4ax2OQFFmOxF+kfwFpdRfaPXCkWAES01jXXuI8QmRHL+iYwd5w8wO6xH+aF
9Lzr43+In5Ca2L9BKeDFJJJUvkgptK4Obm5B54R/CPtbvmUg74buJxnnkh555wkYIC5TlEx4W/w1
yKnuuATkkixWT8aar7R2yvzT+6XUOc89f4kRiwiHpO8ptTfQZWfoVf627gPoozPUaf4wRrYyAweK
ayAJMnwR1w5yy8tHTkokeD3kE7c9ob0D2ZmWIpTPfL4Tby0Jnpr5yeJ5WCNg35fJMtxMgkqeTvsn
QsT7mxdumeo5DiZGcU2TyFcb6DJ/ER5Q3HNs/rYg+0P3AD9a/rMZK7athlbbkay/CyANWolBGC1r
NoJAZWyWweubjHqTTiL37nifwJRuE7XuMOzD28phU6iTdL/kaWLX+lMXkf1rgrUIfzP9226sZJ5x
CfAhh8RSCyNBeW62so68ogzdAmKwSCLWGbFY3ows9n7yG3M+qte514SgrquC0sRVvPS8wkujXw1m
A2Z16quz0CLZhqW9vHBrODjXFiO1LVEK3dkGcbT86raOF+YVNSIKUxQjILzVVygfsC1wBVCvZ6Zt
ttABDomXreOkdTNt/jp0FhDtVzm5Km9Vn5EkFZmFAYtgrCQK0OUOGucaDo4xL44yPBVxb8UEUBFL
xpCIy/2r5qlWA/vm1hXnsiHj2LTN1JooebbgPdFule/Raj0hPUBunSNtvFwgTQ+uNAnQPay1mB1t
6eFXOcZV+ciDafo8kFp/VJrLHa46wzBAS4mwjW0MD8vA5L2HJeDqY1A4Uw7Ck3inxt4jGqeAqKqv
BUo2BKdEjPcfe2/NBjegcGU+3mJAJ3h/b6FLw9b+2Rv7kAmlna7cqhG8ha8Hv48PCZuHBgjI98yp
jBBqOdbGLNcRB9gj7vz58cnCp2FbbPmbHUoOEhWf/VjeSouqGVggZg8ghA+Gg/L46OslO6lp0Qs2
1jYIvt2kPQSNHkICtu7ItvFo9fg8eeRWLh9shvZ/iRngKu0FV3ZcuW52eD3PdC4FN+N5JzzwenI1
LJoU7eK6IDo9rzscAuYg3wKwgcodZmEQkHQHfmcAxVDBN9gBbDpbbixgXm90kYhMTBF01sifkbls
IoM3Rs6WHR3E2BqbFrUS7bmiEsvScOCcif4bwURMe/fmC8ZXvRKnAJVX8zwBqsLBtDsGSNThzxTz
vIoExWS9T9PdnpaW0po6iM/6TI1dW542EWsh+E3RkaQ+Fkr0yxz4Xhh++/EwUKeboir/ejMaO0dy
xYMDafN7S282q8WgEx6T+/939i498cBMNTRq6AVDe9hVtYctUmm5HppN+Jx71XYsSSN6D6c4I9Nm
zMDSam3KtD60xuDKqkXEMyKk4M0twciJasNqyqRx5NDTOKz8wauhCff3UWFnZVsvHpGVYuebYsqc
WbNAJg/w9zDou47mJNsMekbSYVi6dUe2cXja7whTg87UN0IWWK3dY/Zm4+tlhpsyQoXZZUo/svR5
i8JmW/U3eFj4qOCz4NafodEbnq1CyZPTcoy94Op1LJKaktcTF/ei71ApZfT8ALSrnG7+9VJNqBrx
YdXmdgkgROq0bnwAeDrbC6I7P0tJfAt+bG2UC6P87yGtAIzLVrSidQKyHzp+4zNC3LTNNX4lyVKX
BCmjZ319Zl6cUZ/1khUGJqpgxY6HjaQBqjpQzhGOvgQZXtHbF7oTGvkJcz9iW7XWrgUAZFk8dURM
37Q3KzWh/aAN8udGd8hcIwFG8HAZgHGmlDcsDRW7vJ4uYessVfNsxGlUF0C3hBEWuLqQGrUqWb4K
L99CTTsSeawgWG4cwP1cFqbEJY+d6PpRugtR7xLVwsVbI7GSvkhcXt2JKI2qNDNc/y8iGs3HIYDB
erH5FocgHlgQpzWdSvcF5JiebAn9m72wDLTco55jedTqv3dJnHAGsf/2z6gOO8XMhxObzo6FG6FC
1/0HLc4TwaIJEQow3R068RLLu/bDBUETKO4YdOj3Y3Bz4EcI8Dtu3mvt8oSlLIvCtupK/XfIIQ6L
uRZtvPBSxZlN0o5SSJvDLCxEFKS1jBNi81gsHNAkO6zMHtoFxd7VKko1SW5c+EQYDZ3d0zNqqX8C
/xYzw5eiqiR7lgoHBXas/yhUi3sf9M+M3tgsraI2KwcjkzR+srd6qDN8lLAfJ9Z8VGP9gf1tikVO
+UKtfPoALQ/GYp0eP5xLNCegB25/mvUGGCALzUi7GgDkV9+GpLttf6qMGcrTrsvolrUHDyLT61xF
tNDUhtGxQhSx7mTIhbjGSH4SPZTSU8Ych0jXjEpgCEmm67SOEP5QjqBgBLdeTC1Z82c1cZxEufXn
TsyIMnGqC2kE9xqc4YPfs8ZCu5rq3HEpmjZyF/NxwN9jZ54mfTP7gfBY328I4IZ5elwg/dTe/yem
Dzrn7RuNIAR8RXmm7k8UIyfXVBw27hPlsaeG3JYFFN0yaF95/59A0NWpF50WlnTjbvCn01/8Y296
7dEsA92Lc+Eq/ZONECq47Eg5Uk177zNrP40i/dM6c+Yb8wFS8sVjtbIkAmmVswMa2/2aImUCBdjC
ByrsY1cTntCmRs15iOxBi9hBLgN0EwHNCVZOZvXvqOVdyDCQLypW7iNqGZXoi0A5U+iicuMm0Myy
8M2xDYuIV2OOaVAQ5OFweCIyRKkTBrbuRB1TfV934teAGV05mqL/bWbXf5avdra2zLnztJkNcyDz
X+7aCYDRpO+lVPjI7+xgAA/V+juJ432u/RSced+uPnvtZol4ffOzJoqGk9YfW6Rq1RTd7t11xHT/
7Rf7gYLTCU6m2FhGnGvA9ybXkio1Y4WbOjaZWa+TdYP4I8eXjV9sKdQzfJdjmIZJdEZFwOxVuAIu
viY0I352jYysoP/1f157/VJUr4m4vkgGfRpnwz/Ojy7hu0hyEpz4AF78iR4zcILQicLGLgcP22yS
TveA7vMcDRBbu50iLzZZQvccAI/71NU6wlHu/24WaflMSIDGXTIO8YVzhJbdLyd/IAV0TY9iCQl4
TWPBW7fBaoWcrQoi96jEuUCeJ5b6T11cbjsKu7jv1MTEL7YH9gc4d/fP8dWXC/kym9tb9B6JctwK
Iv6OIQffIt+Zcd9gQglOrnt0r57aVFlTplbX4pJDpp3wCtRpLAHEPtAlwbrAFEANnu7xZzWwJC9O
IQGn/9a3HayR7AtTbWeCQcZROrlyeaNPKdR6exXctXgZNC0YMMNsebqCkpl2orJDv9iL6gl219sU
4R65W34NP3mvCFwohYAdaZAozRjOLjk7YkWr4qz6LeNeHWyddn9zxj/iLUaNHsWs7EiPen7Cd6B0
7DnxfACI9dHBHLCgnA5EN8il/g3pjca2ozzLcmT8RI54N0T2rnI2AnO/0di6ZfkonihIm6wEsutN
P1/KAzz3P3uM6gX7BZddNC/ecBDblNx5stq+Gzm0z0wwq+jCip2mdxmR9pHZJpRSRNn107q8XuIe
C+lqs6UI7dIP8z4dAZ5K3t+j5LJmj4OgJmT7pRqUmbtx6hy1SWDinyRke1htxPxlpb0ZOFThNy3E
+C8aZgJVrzcyicSU+mvyvyn1DoRLUffB1uHDWrVs6x6m1YmVtgK78AnMszlplY8P5oFQAgXkjVTP
nxLmlVAS6c2XRYjkaplH7m0IjqUS2Wi+EwwleQQvudU6DDP3ZMPV0tKjm8cvOhzkoROLLQ7+LK7A
ysPi3S01i16HEQaQFi/J31jWYeazhA1LVaCg7FAbgifOXUdtsCNkV123sYnbdS6TqDocISglZ13X
QJjmYreVPEmRYeNHrTg1px8Zrk5Ivcb6Ey2SVHA3pHMhS4cQhtlFJ4msePeQjvdbna8IdowvwGIm
t5aEYGToGrlCEGy/29liDGmAml98p2p5ekyMiKpaNv5XhFAI+H1kaPW+YvTYiGfLik07DUUjgzKg
aJq/3PKvtj5bb4c4/5iQfi/VUVBlUg/OzWBTq7tuTdmB+2vnKd2TusFmW6TDOBvw5Cbj9WBHqtM5
p/lX7G2Z0XTSAH2UadAlXuquhmE30Us9Mr60M56eYS9ULIn1rUdhyZOCz0qzyq7Pue6vHt79rb8K
Jjy1rOZNR/iylHE4QpvLC8YHC+sPcoUDapEWEbh3j4j8QUkptKCX1uK6z9c84Rjp+4ICis2YCx/E
pnfr2Dk7yGAPI0PvXy5O22ypCkEnHqMtU0MW6GYiYoguhy61t3gF/zymRNfXksO+vf/ogWYYLnOw
FrbBLE3yertmHAzcmI48t9uUgEtk0bxucCM3APJloMP5ueRjJ0Bp2715RaWpwLGbTJVtpMGEqV1P
HzYYgW7fbx9lMMpbRS3IbprSQ9qixYWqxWFUlRNjwrfEpC+Mby9JD6o0oInbO4YxcpyKEupRWIrs
Zk5xHOHstsnxTFnaFiD4RfJqJvpWM0Ltau8QuBAQhpNOZurpu83Pm4/3QKcdH1XP48Ay9oBiWRw+
A6yzRJUAIazukf7ElItg291SEQHzUTHrls5dNaBKZzGW1UP6SZtirneCRSm9dRza6xMmh8Mm2ilN
B4ts12w4tUnvveTz8eIj9DpmngGgsXONXpVY4pQbV0jO+LNnqnnjGfO0+oaHdoBw8tc2TzIeqGEs
+PTgChD1LKRN76SztiVDtolQRKInptfNvIYw3+LEzdzriHZmijELTnRVS/DTD6x/Zo4Y3JdgymSp
/M84rwSF6U3K6L7MjPzQ6NOyDGixG4gQ71C5f+rIf2gYdQ8XAmM1LljTjgHsHF3TF9Y5zy2j+Olp
Cy7YyRDHFem30fmrh4MCTwOAn6Vct+v5puZty74wigty2xIA1UZ942M2WwbkeuMUV40wJgmQrCv8
vYxb9qC3TzsI6K+zMKUBXBr8i6JQjp8Jshmb6SiYN1TGxw9O3qOMElnQY3VGRnMssW8iUsxmqUFi
dyJPoZBwnhsCzYCzrQM0KK/upeSY7Q51dvv4XjM/mhOpkXDdPOLN3CPHlRNOxNJABCcCuTPogW+F
f5pW9gGwapzy6EKsfmjNJksMksF5DCQtmqkezkIAe+MZ5qJWVUZouK90P8GHDk7eDltblmakvir4
+OrdgOftsZWIDeI0zEFOKRnGnZWC93j0kVnakKc5ik0AXVHi5ED1pDWlQr92aAj08AFYHdo4CgaH
qWiMrqu3QPfs4nNN6CkfOjLPQh/ABsoY0uW7oHFHUPxyACGJVLiPxbc7be2XmqjsuJzhoK8yyOm1
/QplKoUmB/C8l+MEXvXa1KLwFN3Dfkoh/iQ46hDCZyHZDOXKQA5Vz0h+6t5bMXfCEq15ISaK34j+
WSVffhE3ewEC/e5hrN5Gevi00Gmcl6yk8biORrqC+Q82U4IQ1nNxnU6kGxuF8C2+dspnpBZk9cs6
9LtU2C8sBKOGari0etrezD5p620Z3pRUih+hiTi+P9T8i9eBgV91UV9p+5yQCPQSLoiFlzaG4Lm6
6Zzaf1cXs4aEksz74HlQOarrRPOg+okwdtvXtTU21Y3NSFYP/FQ/x9fOvEV1G/rDsOzUFw1EZKxB
ZyHQn+x+2PhUmlNrcCZQnnlX6lKoOePI/D53itr3Cy6pTWz+eD0EyoDbxCmAMOf7wd4gnj2G/aDm
ToMjaRtruCPpXoIy6A0BcB0GB6d32jpQvP07YNJPaqyFqZ0rIMvQR34elE3lLx4n3mMSUdHGapEN
kYt/xZCTGDh/garFfom75lkZCEEEp7ndREvieSpCv0SoPd7c5JYWfjZFGh+Qgq+lHq+AD5CGJYZX
6vtBECjlFSIvWzzisHZ8PzUHirKOp/XpShT9LsJs3Vysfbi1bXv8xJ3SQeCDiVlbbyyMFeTHycxK
96+hzDxx5rBLS+TS5Sb++FtFKyv6kfjr8r7CTmhQ4rJT7zuOu4S+Al+zDCEYEVEKFTpXSb+JN+8s
iuSctKR8Y7eKzHan1P8LN7f2bBhpollgsqzgQDG1MWe4TNTh4wGeeVEqfNL7p13vxMsKktUYhx9G
dVBMz4wJfMaYbAfKW1HgQE7I6Y7gd6I7uDG3P74XMVB/C2ivgAoHJCWhd8geIsHGucUrJaUW6zDf
jEOhSIs7nASnDuXXHOwr5lhX28dY/kPhCV0NfwyIinJ9VOIPfBoSaokrDUBPW2k0tQknLQ4pYygb
zyjG8KUzqbVcP5RNnB2AxXFDOz0F9FGgXYSXRoZ6AT/Dx52dsQQ1ba/KB1u5xu7IUhtwDWMm5ysL
51P010mRIamTdN4rUaHR6PmVn80rdg2MJz7LYMHw4Cc8QD3sZyi1CmNBLHgWERypHtpotNvea3Xl
uaaFPIuYWh4TM2WMOtVjzjESVz3eEzCyyEhKYs06+oGRISzGZg0jidQmYXEBVMeS9Q5QQUN0T64Y
9rP3frf7n9jYbx70HSOITzyE9lLB7hvUdtGerWoZjasksmXGes7vKTS10SEfbAGk3O8EIQfe4Rdh
slRCbkLAjvMr6ToECYkpA00Qp5/JO3nmG6E8SqWaWmqJbVBxtCwa9XMsxj3HT57J/EfzxN1uvzmt
FMfhqiDPVrhY0RFoz2S5qfBo1HmO61+j6NCA6W0EitDma9B1V6cDWYC9pcWjdHs73/y8+XXLL2I3
JII8b14xARPcAm81HCXVMRCeQ9lL91TK8N+PDDqx29jMQi1QIMb3oibSptKKexghTmMqIwqSANpE
E8MP8MaEh0WMnvS0TMGPgCCoa7VXlzbX4pUU3whArCx2kMF0UqlDvgYtNG7P2NQr4FVuEozShDFM
nnx+1Sp7lTct3MZSfY/+po8fwZvmlBZ30x3gy3Sey4ijZMBTk4lHkEfhVl2wIW32P3lsaerkBbn9
ZFXD7SSjUbpw+TJGMdaPTzhTvi6qRB9e5tRO5NEw/Xju4c/689IUhyc6DA9Nx8dkyC7s1lrB2eK7
xc+PbkXbwZ+hCz3Kg1MX2h+/A5CTe9bd8IaOJceO8NllsuW8gLXxDjhrmY5QrfzckR5eSBGAGlBx
0OMNd7zWW36fJQErxeNhkJB6Hb0AdpDhKKPnkoKB/6qR6jz4TBdjN5vxMbzPAGVGGJ2goI6kTtyd
Jk4K2yRrwm9QGHbeGJgrzrh5QPQtKJIRq/+LD3hq82sHTkCEVY2edtg6gIsiBZ7gvlmFGZLsXrC7
k/F+7kEztmINQKsZcumCBpyrD5l9fYPI5v0SGIs/f9fpSiWJDnj3MT5OXotfQ3M+I3qKzSToi7RH
v/HWesY/f3QiDVmwb2eZIWLrMC9re7pHFNcJrNCiDtn7t2mvKoIm4hs78aQprzVs1KQZt/WnZCst
aQb8/ozWUxD7ofS6jsMEaaSwTka5FORyUiM1qQh/omlcyK4ZcAnpuIy+X7GEKj5mUYApeoh+iXQb
FhcjAApsAfGoOoSUUxSzv6E7sw13gDoN30xsjK+9g1BwBvd8Q23etn5oE+qzexocBRz2X9N2v+vt
TAbzPMq9v2lnTOjR/evhNZhQyX/xpOsd4symiP9bCGDUkrx1ndHintzQxH7zJHtqbfeFhHE+Q+6J
UwGTLiw5DYNyEYX1DN9oyr+jXvb7zEl+05dn+YZ9aFBqjpRSShvVG/+pM5Tqtme4MyZGLliHHhaC
XOVxs33T+bQdMYTw9jZ1UZtj93DAWSucHT7Brdicp9ziwwMuSzgIJdlz/uE8qsQvEY2tCAGUzh2L
2UcHjP5V4JUC597Bm/b2guh7gJ3t8odAE78ZcOqVn29UR6v6RKlMJkQ4pRJNv5aCuFXGeZ49q1k6
beByIOni5JXN8ED0oG1dM9Lc7dqij4O9Ia8+E+7DULJqRlWXvvEhU2P9QmVhkam5lEwAhklors68
LzUhJSGbyW5VV/2k+0gHYu26DjAMplERfS6EXdFcwcHacFhbeshWKa1D4vVK/tOuHjkf0xpyXZ0E
GuQoY81cZgdWROaDvZ0jb2DQ1yeN/ikvIBNzgegxefNYDFghb+8arHHdn8RNq9VTNUw22i5+HTTw
nYrC0mMDvhm+1+jgT0J+4O5ueSOPTSfzQCfvFzerN8u15QxbNbOHK1ePy/Wv3MCFsWyOwgYx9CL+
cb3//ViyDKX3lbnRj6qF5h2pI0e76v7h2HMcfXC+krto495eSOTujZFSb1M+kYVm1bZU6rru7k05
xAaZg1YNguNMS9VC87d7+x8hi/qkQpCv89oc+TiPjOaj6h3DuVUHjF2ybBlL80WsuZsrNbgFDvVG
QyEaxamSfji1PtQgLnATY/i8uNN5VM5wtSCD+4XSE0nxM2hWjI548ZL4bopy5hsOqhGLNxaC06D1
vTdlCCZVMGC8GwlJX5CHME0CfDBp3MByPMIYwqvvgYQYJhBV+ZCx77EuK5jiaiA08H19GTQ36HBS
vqazCb2P+HAwE70IZoh51W5thT8KCTAcAfjUi4qlvqZwqJpDXKlYwpFc1pq6yuypFXJjO8OfwErE
isb+/HIQl4TFaA3NLmK8tVhS2Khyn9Oa8XDVXaxvc6aNBi39kX+zDcDlWMzf7AkGXkAxuPtNj9og
9TqhjU9msMPlojYJu7iu8C/63mS8letkRcb9Q/jRx3X/JdF73V81dn+GK7gWO3gRhrSBFTrbgnfe
V01J9K8I//oPKqwjwISLATBupKhZvYQGFHJkuW94ke0dQr7ns4YLRAfG2pL8xP5zIvnOuI1Tnt2z
uHaqf9V6IoFskxyDhN3J80qcTig+DkGvir3zRD4a6hV3jekb5fJTANkTbT2uvHc2libi+u0Li15W
V0nFOL0CZsIQ0luzySyX8IJo4baK3m0oWc3wfVLlTBkBdXC+EF5fdg4ymWVaVumIor5Gua67l4r3
9xCyGzg7wNvsDbTvqt3GrLVGC1NzkhpYZHPgQ6ToeeKWExA/+aCIsBbZYbmbUWPN4GJrOCgQi9KI
JGmZdte1O6WQ0T/ztt+WD44uipgDAfNF+PQyJwAyc9AJH98lqmmDTd9VoWJ9fFj96kyXuUYn9Z0h
+45d2+N6SwjaELgXXGrWoCvb2F78NluDHYPnL/u/st6Z87YfqNi/Vqyj4U41P4YC0Kyya/jfoNoU
io2gr4xbfxAftI9AYSPKnskItKfwN7J0/u0jQIAS9TTYqkfXoAZQEidleAFbqmVOFWNgTlgBJIhN
AXpPMXuFdpPf629hWYcMEJO4MbhFYSBetV6E4zaFtgmkY9+7/BCDW/f6KX/GbetbfshjYuH1XkRS
1RYl0IZ1AIBJ2ynkXGnJZgUdxxV6OTz44eaijiCazxri/2OUNHMBDgZKkI1LQkYgp6oNmpndyBlP
7bj/xxaCwJDX1XNOW+uGdt1mfWxneuGPS/Z89qGjv14tBoPu/tuLVW1zVYH1uM9wLisgMM89zYh2
wcUgYrr73F3C/U7UGeVRzfLz1W06TxJGDuZF6ukqpp8HjUW9eocJ3HJmUKbuoEOkUppMc2uV+TSm
WPn+H/2YDx6+MfHgI0ey4BgRBr6GpelycxdcKibk4V3UNjjo1n/lRYu96tTNoASZ143kYB5BydDA
KpJEsU8ldwV8jwDd3Qf0ZFTMRVOLQVJbztzgWQ0fFKrnoiy3LmOuV8scNdI3LRKKCE1LaEMLB+mA
EKvo34hBabBERFuvAFPD9BPgeRXvlQqxfzMS+ty3YhdBguLMRf/5BSlkogmXZTvxafL7exhbtxkm
1I2DumTyEfl/1hIxASW4q7b7wfBvuQ+cNjziykaS+/WN8iOUhTjJfhqZ9jjtECBhwatxRZU+JZii
WorW0WswJ6xUbUANQECMx2CtRZa99WgepWYJe051L1V0iIwbbGSWtctmZOHgQhaY8Y5KExhtLldj
fSVDweLDFHN2znUKIvPZlmOra5M3SgwqC7wcL82pX0m0t3mAefo+Q3TSEOd1EfYqMnyZkFUKt6uO
dHjutj4VFoEssK8mcyXCmUYZ/wL2p8RrUQh3F4kJyiANjTBsHTsMhtOhLLwwqPWRGqytaVN3Tluf
tbPEBwlbL54eXR1Z4UpCiLxKqIk0NT9px27DjPfONi045BGwG9qFFU5PAeJ/AKgdPSUzdeq1pZIs
PnVS/CVSVrf9UzhRFvVJI5Vf6JrtWN7I8yXpprxkRgROQ5lbgVjkpibzOQG63GCfAYS/PIunTF01
v7/KE9bDek+NVd31QLMco/UUtY8fq9lq5OqZol2nlWoxRs3sIKbXbbZQ2rdFQmyqAYausvbvxHm2
YUklQzsOljtCGabcf2rAHHGNuldi7a2UgPm3xwqHHv8Q4SbfEh3X6fa1BxrKXOJhpHh1PkYHqQgk
At8aPewA63REqu+dENcr78svD8tcGFXax6bSm2mzpLQTbYdOw6aGQmitcmfz7s0mBw+pQH+TcRAK
od/cu9HloUwdZevo6BREdUIFUWGTGlYCmgT7I9bwP4mVI898bxuJWrp86J6F84EGUUdFxKdLFxch
ls5TNpTEUArccl8W9R6rIT9VqN4TcwPH0ZRRA+xM7AbUqqYt7VVd7du1iIzZS0ZuujLZQQLgq9im
4+16GvK7hDmRpNb5YGuOP1L/fBbuT73GnQmTzfBGyzPp9G0KLonr6lWyI5BHcZMRBpFfeHo1c+SM
JMa5GOZrRPYjhfuSg9cJUw6Rp2ryHpo/1MCk63NLBOiwWasAv5Ta9+fzr4FtpOXMim2eVsGBQPkB
DxmoXINxSB9ieYN5DM3ETeBNsdTwRjl52L7Se+zx+BziB4sj2BSySV/oL5Wc46CX1yK8o7JwNFgl
6A2nVNRyhRIp5dDDhFIBLNd+ZKuavua6xg1E8oiE4czfSvYsXTv6w7hkfIx7GMrB729LB1A/a1t8
xtkDqegWL6LDXNpZ+Iqexfe3hPulxXFctZiCuNQgRZJFoQuuVvjN0w5gMMlkrcwCnV1Z4/OZW0qB
qV+qLukh2fRtvjCMLvJ0e73hS61PsWa0zbv+WoXKFS9unN9GLAwuA+T+lml0ZbVHJws6GJefcLv8
AosikPUReSPQKg5w/6iE2EBk2SSIg/NpO7sKO/etrwZB+7VDAVfrvEoe7bHYbIAQFSQGBZytt2vd
y3b37EyIsnAlFkbFi9HZk956+wFEGWkje4+Xlav40vyjHlHLFhRH5SqYXYk3FTwySWwK5D2+M2xL
dR7AGSnNd4noP4qbe+0dvWyjK9zDibBLmfJibkjNqoITOLMm8oqk0rOKNCI7gPKkw+pNNa5HkqSC
9uMxGYb6PX/8s5oJeJXQm2kpoeIt01mcK+PooKpyYFvBHpi3CMP721GL4Y5Ko69FvE3q69UbREeI
e1vW59vfQO9cFExwLRaOkey0MbUr1QCPa7pcSAtM/wvM1thbYMzS+zD+5XaKBLddxzxMNxh+OQBX
uzpJek5rjIeHsnUC7PA7yuVRvFu/ymDo3nfh5tCztWEYIwiSx89Ur+LjOKZQRR7WKiAqcvQcpfjE
5iRr3pXZlH81yw7y0oYZmcUe5vwHxv6AIbRzqeweDj0SGBaYiRzKYmrGa91oc9vjtZLMq4KeyJyW
ESicVc7Lk7L/2PVH8AwznwYntNHG/hcsrf288bs2hlQ2gc/b2DmjnMGmXlPlIiXPNK6Rd42BVt3C
B+WhmpbrkjxugTDnoJC4r9sNYQEjTrJgsdjfz/d/Tyx67d4jiTfxxvbhiCySk2nzh1DTgxs1KSLO
ClOcRan9BNtWvv0qIjSbkoZuq/4296j2isTPUf5ZlFvcIk8bf/8Z6D91PGXm42CFZnrSLI4QzdHp
XJdlcbMlI0BxiMqZXCD8UATo1jcEW45a3KsEge6YxpYhEwCcS7p1Smw+wkm0lwYWkyhy8JtuPSfI
wsFj/mkpVLczDgiSARKjLlPlCG1cMcNiHCeBX0qZYVIHgEw1kVzBdEsFqzB2UJ2ySxG8ot76rvT8
dtT9Wj6lDqvpUTu7RrSspURohQyKqtgnk6Vb+nPBhBk6oZypATRYI3nMefR/XTanT1s7lWqoYOaN
ZTWg/e8FgAGzHLLd9Tywhe2BraqXH2SqHbm2zPR4nOHqtyZJgFaZZ0eXhiWFPKR6G3D6ucIozyfv
mSgq881/1hDVBA8WmMGVbs5FMG10bw8M0RCPWuEI4lGjeqhulos7Nwe37e+uy+9bszqyQbH+7yps
gKUgeQnFLx16RDuhDsdOgzPgm1ow45Cn/4/zE6+n/T7606suPZTP6UodCoOoKyuEXNURRYDKx0Ca
Cq7PRj4z0SHyczq0JzsP6LjgQaej54xDC9HW0pOfUQHDgxYyY3Aw4ONu2xWXC9MaC7hiJw/61IeE
Bh2o1yCe4S603ousahzfbBB6q1pXcupEVk1tvJlmHZDP/N7NnZEcD1Uiw30LPEDD/sRKUxasIJo7
5L5pvyVK8g5im79vyrixq2EqPE87GaZEinap8jiFfRvixfpZTwZ16kho0sSAx/8EUpLyV+nWEqDw
Ekxk+o/g3IHTgldcptNxNyRelt4oYESRGj19pkdlGVzV4O8dLFtWqfShdYwtTBOpA/9gHdrPRJyI
mpQCUfEpZkpT07NGGvIaazGbUCPtu+Mm3dQWZywt+mMHMJ0yIDDmPvCqndZPm76gdlu47biaYm3K
RjAyPjtpC7k2qxz9sTlwYswXqFasUFP562ML7oC8Tvf3xENnq1EiOTEgzzfjiXXwUqRS88+1Ig4s
tnAsV4cI/twhaU6O63Yf9HLG1gY854c6YqkVj1Sd5utNg5Hrii9U0syv1fPcZpwtVPWinggMjvUY
0T4pvP9xy2jKtHB69W5N+4zZqUVAWEMK6tWZODagJ/1iHvS8dL6UNbmK90+BRkES2R5wN/dGwnAp
1M6xnQ+Bp3Edba3l43zAFFySD0k3LNRH7Ze1EiPosy5yONbOjeg6paNwQyArSdFErSW/HxiiiXhW
CCraReAQ6C41fmsqGPs1SYpUS+/57bjbdGTTMCgIO02SGNx1UI1IV0jwZJZN3d0qn10DhdzIFM7K
LzfLXCJw1GXlhOVDTaoy9XwhHw1tjqqjemNfACCYeZmi2WGdywWRE8rdfd2ir2/y4KqHfBYYuI0s
3/LuQKmctv5FyVo3/gYzedVB8Blxor7MB3zY77bsiNzII4uTySKSBJWF0Ui7sytjrl6qqecPmVcv
eHSltLVUH4Nq7Wlk3WfBpzuaEJi3Ktv56xIfJFJXaZIU4Y6qt26Z3McIaEkJCFimqOQRtb+6SCBz
wWe8e8MKTz5BAq8I5L92wVeXLV2qJym78OJsdKCeyZ7pCVfFi9C5mPpWmgszKbHsEPcvGpAlmh/k
2wrOD/7d/FtZ9TJbwaVzQu2+KEjmiNeJ8LKzbV76md15pFiwHZC5OrQukf1FMW+rVFX0AGYNDs/C
mtGIHInqOhsVA5Kr+dxjcAXMDFn2S/uJkddFUkO97NKujS8rBYoJZuWwDrUwtNzCFMQtfSKpJ9PF
P8X5IPDtbYypG8JQE6FehoChb/QmAGg0k+WtyqZtqSAZYbHLx8bcc9FoadwB10AjxO8Ep6iscxcj
b2bKY0M5fB2HZAE9sd6XOsUGpzgfqyWNsKYqo0IbZEyeOlmPOHbkcJu01eM+APQ8VUEM79LqJ/+G
VOAaSdK7do2ITE8klv33Lqe6kN2ZLresLhECWX8rCEhtu9430nnfOqThPGLuQASDL0LDO8mbtHI3
unKGhZ1zsQpW9rRhlX9R2o/VlTyRqoQur5wgk4hcFFJtZC3OPxkc+5xfFHfXbunUskqKY1xIHJbf
61y+PLLlen3dpNZZbyguRubmPCiUqkAvP+YC3YukzyW7KYfBbnUHBaGNUriqitwpnWa36gEk8YJY
En8Hjkn5AjWCrqqgvtnDxmjujUZ87iaZDy3pfNCgdJmm5P4yqGILIk9QFNPDJwYZuUN1WywgrnVR
/dc1ymuXvdd31tMnHXu8ND62mDSXs9CSSomjY0weZuE3eXoOFxQosSnc6WoCS6zIVchfna2LWpOf
nfYTt45DPKEzG0htISREAwJKmrOzCUELGMiAdc5Yc+CxXn37QtVcnrAgflSNXSLbaxWhIsNhenHf
OomiQswO8LbuLvB417i1WbLGoBDIGE9lktnGcZo86i0Wsf/k8Gz09BdoQ4oNBQrnyIUstgvV88sZ
EaglRNprX/LyIgyhMK9n9IsX0Eof/QZoCUQkgw2RpxLJ2co7uGMvkov7mLC/x8dwAAOLBBXU8mk+
onj1hJ6SeNIrkBbDx5sT9ALyfO6u/7iA+1zr/me3CXl1K+5erpRsP0hJT//x7cR0aLC3mcxl7Bn3
esfECN6Ee2XVkKRwz+o4TWA/MPDMWR4aQq0BIlOEMMDaalNH1QDCegYrxsZbz2aikkrnlSpLlAZG
nY5ZAEip6fSciu+uzcku+ytjk8KSJIFtJuk3Vbo9lFsV5tyzO52Zi1xjUzA6X/u44Dg7+Kx/BBj1
gKdiQHxHK6BlL8qeTtkztPvVVA7OAuQbM7Vysf+mGi4ouG0X7iz5lDhY5uuwAtkyxFpXJCQzFqp0
3eKpspVpl+5P6ZEhkuYFpx57CPnFDsOCs4ZUD2ubdr/NbfTTfL7NVlu6ngplkzDF6kfQlA6p0TY3
0JwB7hrGSTXQxKSXdFFxNQ4Bk3BzqOk7WriU289BmeD7Wxeh8muhrJF06j8d9jh+i5A53ErjV8Hg
rIGFXsOZUzEe07rgP65fM+AWfoqKz8Zsi82T8NbOFUR/GMjei1gaTVBp6VBACYSq/db0VRbLzk24
Kd3K2BmMZqkkThYYXhTrg31Y4CWRRdyGTgd7ggOMxz92wkewrSHZBdF3kizaGKxc3DNyLwVi6F95
Bitwp5CAYK0ZHXI+FvsHdQDryEXnsdxBRk/V/Cy31fl1haBLpAlUzwVHXGetCFal3PfhkokMC+MU
e23bGUnRPWgHZefIKyhagbNHjMCnjCSKWLOYYAKcvoIatEVICMe8/K7bYzioVe6cS3td9vdhgR82
tgD5SCr4qCaG2lO4Mcnz3xIGZAkAnqaYcGRXpss3dK6i/VSvefEw02t+zeaLdPRaOW2xYRWyO0Q6
WV9XaQ46qf1Q61GYD9KFeSqze2BWDYbbnyS41jPL4uFW29BOjnifTxw8TqIsoyWj06bic5ZDR4yH
bEvov0NpLwGrbdWquPEk7wZW8ddAPFvMSFurLbfu3MmVQ4wb2uE5+1PNlMWp56sYkwe8lwuAG50u
1ZNO+1l7Dwf7iRkm5D1KGYQZTW5VNZCBXWSDE9eNcEAUwHTN9RzJUA4iY5sdXhV12uSrQUgbEgAi
xxjYZMvomT3TvdTwi50+L6KbG0VlB8ozusxBy+lWiUxEYwWZae4hW771ulQdm9R+tHsj1LAZ5zAJ
6ztIJJgdeAgn8DKSQz6oRQDu0L5pwl9qWVFlUg3TGUTH+q2tiYsfkYq3rqUCzEy2bhaWwshMjNd/
ulsQ8rPN4OUjCiOk72UcyjCBHLJPNNgfGxn7r/yCHVBzChdP+PArcMSjUW788I8+DR/ieqVGafu/
ucHWq9N6M1ewvL3RTBlMyS1aHgS1QY0C7j8FDs0nu/f/q0bB67LEV9D+azKB3+fW4aB/+smT+x+F
cw+cDfZBDATTEG3SkCk3Gwu+ViTvOnlKnlgkzyxFTWLfZAUoSkk8k67kxbon5sAU59cccM+u6WZu
lncW9/gRdICAVr/Ukvp7YsZG9hSvaZcBbIcoXE7CuB6ebHEFFZb7GTgGRugBYkW6yyHd7Ro1NugK
6Z+8HNPxgMOKOq4c52VPyX9bb9H1wTUp1h6YNmMAyv/rdUXq0j6/hzybx2vue5fl2H50tLYczMZK
craIx9vlaC5uFBmE4cXCxd1G8lvjpu+Y7M1ZVi892r4LwAPRdjTEHibVx8HeyDTzmlTn5bifLu4g
FRavIgqTzzyDvE6PvRUljsYghCNjV8hJhjuLvlLA+HMn8ELklpGDfcUU8AxhMcX4jWYdlxgGu4qK
sUtmJNUdcNFgOXYYhPKhxmik228XzXbR755ankna4+15lqD3aoq7HQ0Aj9mnHlLxg+hvW/4Y8wJL
nS8/xf0DWkon2ddaGAMBr67ozyA4B53uZNoAouhpTxtaOi9FpShlfauoxXP2gNx7/db4RRtkWcAY
lycQifulkHkWOToZm3cLdWo/cCPXi1MkPkkmY7C9UVRuKNoaLstuNKTGRBOdXAzsYhSgYmj9O99z
dPt5ETp/DBqX61j4T0d1JjY9Fd09R+lUDZPJLAWxnLHB0kXpzckmMONi7VSsbWWvxEhDCVNbhScz
hbxtYC5/+gOA/6WkfAOXqYRpbWgbD4a5PO/5nfGB3Ksdrc47CDYy48pmF0nJFJ8G2T3Avryg/A73
223HU3kKxB4XoPAIpqGSiYaIKcbzyIylT2quxWJxefuAH01fPclvXs/tJJ2o0tZNv5N6PxyGsmPQ
CuV47Q/J2PAr6CWY0SfTW3wULCCUUCheBz4D3+7MfCn6roVGwIAYgdQtEvAOvx2QAIDTGRWrJ8g5
p22pnLCEni8DgOsRCqHDTsu0RBmqstW9VjrIlCU06OhosJoTcbcV1ph3WkpSs98BYpWtEoyyrjTk
vlGTsJDXBWjn2ZP3u8z0D2aGaHBAzqp5x6Y7MhjMgVCB3DbV9QP6nKoYUuDNX07LftQA7/+wHSAX
P/T1ywS2qAB75OahAZhtw4XvS7p/y0JwBZmNCZR8wq7ujO9PmcmJO1vq7qwrE9NBaWDaj1vIiKv3
fFulaiI0BGkFCEUCox5lks93Hly2HbZT064eXEYaGXXFdgj6vo00HDknsaEq19Q4j/DFCJVyGYI9
fF5/gedbKUfCmbSoTdUYA3SWs5gFp+8ZpCwOfL+BaP6v0xg+u6tIHo6y+yLsdqkTna6d9dxEjxiD
sIqbZrHp/S+XrACINPGxI25pqcymVwYmOjhwiAb63J44Yr0D1oG3583kpJLrJBCMY1rb0zLoJLXs
VYd9EeJLvF1YUiGsxqpZPE0nIIKKnfyhXW/wPDKcRxgDQS7qnWCD7S5ZK0/oPG5VFNaU64JKn/R9
fY9RTa1ZVXuN8gqnwdfHKX91qRHsDcVUnmdAojlko/lzzyO7Or9cjA3U9TFq3NMEgda9aUbdDq4Y
vcONpRGG63z15dL0Xdk6SMCezqyuZKn8ygyQRHV7qptvvMZx8208Tv452ucFgCoWvuT2I/OzMizN
GVfO5qdieeHxYE8zlrR8hOJVHi/5PzGByr295IEdMOtsW/cEF72RxAyJy+h9iCV7V7WjfDdamt6C
DsLzoIpKqWrnn1Eqkw7rkqlpGKlurUEnhwdO4RpfXRmLsK38YHYr5CxgMU8FW45vJOdGvx1a5SwR
ATRJrb5cmqcfozmT7z+FgElZub06Py7YSh+xNSA+huBJ9WM40gwxdJJFiuSlk0m60bkpXM9DGRkk
9ZtEvpmk3+sc3K+W7yTYdi5iYkhdpsh3nHkx5wD/RlIzVFvzen7/8kZoP3RuXPyWxm93RF1CW83J
PXyxcu9OcaQ2BzxmSFtZsKkDNkxMWIJwwf9utl6Caa8Y7hOv5A8D1rUk9T5K+al1JvCc2rRa/OHZ
mXM/TKL4j0mJj+HqsSk141lW2CbWXI9sN3R0Y87bKbtndc4DidtEglMsCjZLrGtVfimkr5oGgfUE
t+c3f9wb8vw5CMR8U77OGKrn0S83+vDvVZ5OPnaXjU1HutwQuIYOqPijPnaWHLzvTW1hpamATdv/
hoexfj9RDNm4tvt+fEGNvUbaxuBF/yy4oymaX2Lr4hQvLYmx1jWDV/IgmYKJzN4XxVA7dqaRvEPG
Fx+gKXD2KKKxVKDNNpZ0jrcqSpEbU/btu9NDN+SDJvOLManbXAWbneaCetOipuvYshg71xFXguXS
7xpjfh+GYrQWKLldt38sZ6ry2H3I7F2A8HngVTKeQQAmDXRH+MUNnX9H1xt0L+fi4Jd04CLJPs2B
0rdkdZ7p/BPIw3RWXlmyODX2nNigx1hl0xDLoQqY4M+AKf3guPrzw4YaygXdzgpsozf+k1p6LyVL
Yo7kynlUUaZqGdLlbfsZF8hBcnvC+mDHgOeUIlCNy7GS1Gy8ukKHTQYyOZpcK9eBU9szb5jCKoPe
+zHekItGaEUCYnlBMwmZM6ydA21pbdr38f4qgPRGaswniNKI39bc1s2Dm5o345lUzWnBCEMX1ItY
/mm9V+ioDNImF+U6BzZFpqWOK9tvFQUfcDRL5VoamsrmVYzgIhZG1ol7/Oaza8KZsgrdAV34qYUW
Y8nHkBBvljqCnw9be7K3rBuw9EQEoeFNh6NKwMdc0S68z7SdekpKR8XM3zIJx31FUXfHMUykWFfl
A10W6hCmwGRHjz9NFTJXTBMQdCZcioRxm/9ss2vJmleo3BYDgiyf76gGvF6J5tsPPB/m13q8sshC
Ji+TY7/QRczhqWJCKaQykxk3+0QpZ5Q1hlOyc2O0RVcQqcXcfbfCV/D4RsehO81Plrqn5jO1S8l2
K+lRE1B+mzwQHjFmiFe7yi+ZW4AMq946gcoKwlFS8Y2FHkRLcbMf3hul5LVASemQ0RfkmsBjsTzI
sjvX9KKoTekgacG5Qdhutknb+/EZpFBcV6NyFaKgAjJe4k0ggBOZXmUQvYLWFExtVr0khM4mes4w
bAMruZOUmuFx7omBLfsMtk/roTySo2M/33lOBYlu/793tXPHgmfUi2V+JhSYeK6vSPMXhzk2hu0t
1Z2uDDEm2a2EJ0CyerjqYVHVxfTzFNawz9Xiw+ElhQrrwRmoVlcrgh4u9rFGZARqtztUU+neAd5I
CWnQqRD+k/Hjt3n8naZNxL0NI4yn1zVVSp/ry5Drp9KmyYX8YQEeIUagPKFi9X7chbuUfGWpom/G
+be5db0GDbJP+ntrjGFIQTmWjRi9rW2FMFcMICyh6Zc68j3pqZXmaqT3C3sSTKcXvNtjzXkRju7X
9PVRROQ/kFFRcMEsGX+DEeFNQUK9SFcUKZhFbMc9xr+k0+HLCEv/uIf2szz/lN71X4eT+GkBjoem
hcXDBbraKHNW9USDDH84zHOcwGEkT0jgu3G2/qN6sVVF6YZIR+JJmfm7bApG68QWqf8VDZJ2cyAR
iV3Ral5JUr6oXOP0iVPiM7JIaoE7d1PbQR4JoUSe/f5nAkbBCFn8pwz2hpkzmUiru98qTZ/GjjOh
daNwx7V9AFQ2jI3b7APhBs9DWRP1ZK2848ZuvhOqp8OxpzXcVWwa9iRCUGwRDMQNSwZR3Ojb6tdl
pZKF2b14LLhczvqbmlQzgMoVIr2YqMi/8DHHoZ8fS79qmmfEXGyMRp37C2+nVWYt1duDoKIXYXTL
ZI/TnCkRLBy27GvsYcNcJASB+lEmbfDq9JzdKELSp7Y7cQZnWf8uLVCZaislGdpcWaWNozQZetni
ZrCPUmT1AS0IQ+VkHUliPR6pAOYcDxIW5O9AxdN/qNYz0UQgwlHE7ZbmDslHyWvi1Mq1QbWT6EXJ
GLzVsJjGplKfIzc95xk/FTTbBaHEvJQ7hHDfaS7NmCtiOevqZo9wQMpj6R2aM/QBza5Jo2EWZR0W
9fa0XF3uOo478JNxAqwjJzybk3tme2H8qKN5l5kiqwtcctLp/dm+Q3+fH8k5kEGsDrMohI31TivC
/yYLuIvBMCOF4YdeEPjIFMpAQSfuvbQrtaAJw253s1qcO34osXFuCw3DiXqIghW0xBMMACTp8Oxs
diCBE1nLuuZNEt/ys9S5eGpQg1NkN7x8x10jJcWGDC3v+6BncDTXetBEP99ALgB5QTh3uzgFZX6Y
gMZVa3BpFKJ8OTTKgiZwWiaNpHnoiCPAuAw1pdEpHjTng2+BRJObKh5339ECKa6pihnB9b2ApPLp
TYoILXEkMFXv3iZptDFkwpyczR4ohWAnJdBu4hoTLY7Az5dC4+xN+M/rGHAup7Ql/KliWGDKXPzW
Akk/YSzMdTskgFYoXZ4RC7pPd/aE8R3JkaLZLvNajCKfkm6dd29DSwbgxJTaTHkuXY/XB3z7nrtv
XMe3olaDLUHDX1Dh5nwbhEIzyqpF4WmvqAf69PWqZIgAtLsRQM6OUancjuTaR7fwJ/fT8IyTmKlh
lWVpFyLSUeg8EtSczw7FzKfl3kjVDwPxPK11CxDDJgLDag+oqYZFY9BbX6pfCu/0atOq+SGQquGx
69sJ3dy+a+TMlMt4bhAxf6oRVJ6Bxyzz2IlC2sDE70k69JVD425/YZU+yglP/v1Ox3c6RAfTWkwo
/1gv1GmxshIY8Wu2/teCag/xMmm+zAzm1dxcmXKg7VZs8i8A42EH8IjHQRgnplZ7Hpfb1ZHyvyrB
fWCZ4PDoxmyIl+moeLH87bEaofqSCVq/yvWEu0oMg7WzKpslRpZxXfKvi0BjfnLuJbJmB1hRyr1C
hMLlo/5b2924k9HvyEH1tiJ7c88KlEavCuQ5J26s7/hxH2nhPQUzq9otzhdVcXcmazCljQs0yyii
UcvvrE8yCvIMKK5Q2jiHlHECSkDI2KOpZfkwuJaLg3pLutqUhzcAq/mnL52nuz7/0LIxzGwkOm+8
Y3cAeCv8LqgU5W0i8/wFT6c6f70DjIv2jCrUdZHP/okXN5sH8UuXuIcNtDcMI/8giOucJilT7q1V
Wj6zWJvg3gtESKWx6oyc9xAkx7LY9mPCDoGijzHnMoLNjn2aO0y6bM6G/nLaKFhZxTt6oKCdEaqg
1rc/BczXRAF9CpNJDnJweQ+kW8e4redK239BZ93KP2qr0I6qiyR7I8ldiCo3N7Vdy9O6fTKKISSe
7n+Z0WaZVGtZHBaawvxaNg84G8/GKJgED50JPt0CQscGeMzatKUdgeJUT20tCHEQubCf8Vxlr9rJ
FXgUPHUM7WYlg6w23lcM3WqFZ3KsCjaq/adQfyYVu3YXEg0nlfoZfU/vQraeN2Cm2RxHieudH2eF
B/d5JfRiSa9mutlpsbxhtCEPp1BHq7OZ7cssg02qYawDt7Bbd7ngOVUdlckjgNgJbErUzMaNPCkw
EQ4P+FLk1EnWPnOt/WG99ddepdo/+dtuYg/EIhQzr6nQk0gY7NZg1h3IURCFtJiA6A/zyJbh9E5r
mvVz/wVvMjRgFJsIFWOg6YxiaN+1p/Cd/sN32CwWMWks3PsAev1ELpC87a1AcStymHXWMkOMPCW2
OFEqM5qM/nQjxjp1gqvgaOYKNCi+8G9Wi/aQne1RTj2s9uqjdguYK5WN/IvODt2+35hrhGQJgptH
znA1hWicEIuhhN5p2M67QEqryn2q+b75hZCHGNB9fiFFPm2tHpAVoAUHUWJ//CIJ5Lp/Mm0tqkUq
IjiO7dVRgXHXNSZ5gJpyuDFPlOdIYw1w7ReueQ9xH3lDVFahFewK+6mQHsVJySIyu59A3YTi+scM
cx90ZhAAqAn0F/rsNBb4naRBFZuiXOaIqChQSW7P+Vzy6TprDFaKXDX29nJiLP68B42+yJC+fP2A
G0CLR+oj2TU5GMWtZGBsKrrRYUi7nO2YJvaiFx2PIO00jiM0ikoBP1VD8G4dmpdIJ8GIXHR0l81V
Gancue0BwfmjARU3S4gCkR3PVAM7S8IsPLrTy0w9lbgZ5inCbeWtZ9Kk+wwt3f2AUhLt+JOH7HAH
RxDMS1s9ZV/uArIhgOqVoJJeFCU7dpmOB+YnRIUMxY/3LLfR/MfGS+PhWW0S5Iizlnbx9JGd7Dqg
lQofwerldcqDrtN+c1EEtU4gmyFsmY85Hwf3poZmEwkzjb6eFnCQzJAV97BXbW6RL54ob+jVwnQP
7uWv8Y9sp11TR4n1RITPcKNZdrd03em9MP6kChYX+i4zrjW20lvp76wdjiO1y0aja4MXJDB9frkc
T0rADcExtJ5YJEoUd8/m5S89jExX/gveupAn3FQaZOZ79l28e3hNMsRRk1NkAGQVHgb+4ErcQogk
AJaXxj2SUlM7exhXDzv48MJblDuP2jhP9LP36zs431Ol3i0pRHKpMrBBQ2V7mH4dqmqOkTm2qhUm
WKnqCkSkLDzv9MQodaxbc125uNNuzsXMxJEfbBf69+iY4X/wckFo3wFNobt2i+tZuFvJPMgyTlPi
KCrNDUnBYMACazsClWUWLy89UDinhwOWqXUku/8/k9RSBEAEvAEYo7h3TP5UN/6DCv31PZIWvuxq
lyDMNnfbU1+zpojdRTWaDNBYgIVFTiVfQLFcVFLu6cfo7UdlPjiFgxHk/oac+481aZTNzLtdekuS
wzJSdTsaCLGIiAB1ZDgTQE6SHDrMrAVSTuejPwu8ipkFM2jQByJcN3/h8dAL8LJ7DnXEuUJD55iS
4LgDQ6f4yK60mk8ydaizGTdaDlDI71fBtFMDcM58KhrQwFqooXA2cNK3CgeAAfNArRL6Pj+A613d
lteEjPKj/LyNbHOOsdcNFvPJ7q19CnnkNrtKvflooxLGHaIAdaTtt+Rjg5td93z89Z2hqcy3vkyY
95txapQnMMubrt+DRa/ZL2GdyY+gNXNF4Y7Ti+e19mpnf37whiUbQ9ysDJlpppXoiAgPmTy8miAH
sX/el6Zn2gqD6BllE1PynYnq05VbGVkBqu1ln+TTfNww0/Qyx9t1pp2Jm7RkwJzlqL9+kuyyXHch
s0p+tniWxrZh0VfNBMtoHdr6h9yPN3taDRkqKZkECkXaQxY+I/yJdE2tXMujXyZDdfUYLFvYZ3WH
XNgldhKREXjG7GQX2lJHZTzdtoqy4iLLGtHLBIMKqk/L9MGCteb0G5nGK+xRrSCiY8MrVPoUVU0z
iyjWD1j69d62QUeX60ygOHztUd6TnriOQ4OOFzH3LqIfYpKt0At1yrALI8fObGIlsrmP1GpL4WZ6
ZWoEfB2vT+NR5Vs6R1DVH08IO6WVWI0exImTJbAgnUY+6iMXetItaCATO5jR+mvJpQb424HPJDdv
Ffa2jm7owx4Yi+pbg4PLX9MhwYBxxAJPUUsD+Et/S/pLrzK/8fJuiYEPqtFlt7FIf1hZdS6H35ID
68L4j8sXQY87WLUfK1JPqQoXC9DPHboWldr/yVYVALvJSgQLfcee8W3tcWP2kf8Ng6MiCHKCg6TI
6GTxGtMm0pJ8MMMtL2JVghHwnttF4+1mGNzCELJHXsF94V4BMClwuHeCNslHxXRdkDK+90kM3YTm
9kW7cSr0eyepRA7iYxKhhpW7zqvyFlTzpHES9sdFbVLLPC5rZcOko6VwvraLxHgMF2m+UWlbLQ5c
/XgLFh0kAEwtSOz0URDC+JQ24sheyqJyRRgTvlL0bMck2ONX67K1/VGHKrvPhtoCqdhqad11erx6
jCcFMu8oIr/JYrKBRwYPL9m1iuH7wLwPlNY0TJX37HW/KVG2aWnXuf62M3d6Z6VAa8UnaOb+DqdR
xWhZcicCoeRB+/hD7W/o3d44ZKBHF5YT+y6zyrIlnE9wz6/r5G1cPtSkPInOg7xGsFVY4nXk5nzf
G0auGIk8yBNG5WHgjmKuDKocJgWPxfPZOn6oqOl4igKsRX4rKo9piBLViPlaWXWt5YRBT7hPMWfL
WmYVfnhp38AR+F6ATysbcKMjOEHXhCfHtdlLm8dc4WFhTi0nQq2xziWcMufEQOqsgv9DYZ/Y+0u6
O1UMcprmdOPZP2XH7zs4e2GX2pSXouC8oQBn8bSrot35ONyW2KJIu0EdhScLl8D7cz8fWKgkjpAn
1P0Xx67KPfWy9T3LmSH7EvR9zAN3RrfQLFfQltgY4fOqCJQPeQJvBc/be5wUL4637WyBfiMo9YpK
TLUb7sASl43JWgUKb72XRm53rSvUiNbAnw2Q2UZPAHpzQLbu3w42cqvNAdo6r+9ED6cdC+h7pQfv
w/qxwDzhj+sVop1tZMRR6f5KlGIxgTHmbb+VxC3kZH29WujzmAjFq3LvzK9xADoi2JA1ucElZz6x
1N5LnHhuHozDt0ahYlTNLuYTrogVEOlZ88kzOjbIIDEIkYZtvAkV9R8M1IzjeHyjRiSm0mO5vMEy
wqe2NoRvBY0EY2+hb+joZBph295GhHuy0wH1n/XiElZZ6Dk8L5WpFOUeW+l5Y+zOHH71ldpo7p78
7/LKsfC0mw3zEHSamhi5hnzPISS1VC9OQTzca6kAvFNsHLvXG8Dch2pFHQMqeG9/CCkmkgJARsUq
hZOmNiCH+dXIcFJkpEFJch9+9O16pGS7fwddNKEUXIHZTdftleAso903p/gm+xWB5XVsUUORs6fr
0f3KJfvhevIlwtCHNquSxPbtphgkowckfFieaYUrm5KxMwlh4Q9DWxJY+vCFXIwRon+gieRvw3S8
cMmyET+Dp5A0xChQLlGzsoM0dXTDo5KDKOCmjfbJDzLLv312ERikW7ds29Fe8xyVrAILzgoe6ZTT
mIMZ0g/FH9cP54F/rkpGp7JiBN0c8MiRbQCMAkm6kHSMkqPMxP+hiUbJ2o5H4YSJoNh/FgNkNUdc
8HLDkLjSAlACOi8CMceuEZnrPKG7qJIynU46AYCQIyQlqzTu69k+SXgtACktIXm9NUrgw4BQj9IE
Sa7jUrJwXGp+FZaRWtK+A5GhSQOsjgkAM5EWBLhWmuujk8nYX8okry1TLWKqoufxab9jUTILs6f+
GdhTd2LJwMbEIvhxNLRvoPNUeH/2ka2bG6/+dNpBeOvJcZ83U9W2jEUHR9KEscqFAt8JEVtJbCX2
WFd3WyXGkO3X3g1fxz/B+CeZXZGb6XuGRJvHIC10OT7Q9TjRMHwhhH2uqaJPGcKH95wWn8FmWFci
JMYZcc8jQL+Rb13sv15b8w32mWvJWxK3VjS8WvbhHCNecAnkl6mCe+LQsOPo36sVGBzFeGFOI/j8
LqA+iDKsbDziDoRL7ySPkN6T5kTeXjO17GofLON0mP0j7g228z9S8TzoYQOjRKXfcb4vNEYcWUgA
tBRve5lBlCjZD08wVls81tSzHPDgORWdu20AxbjO7GTKU3m4PMQ+4pKaEu+cBtJCW1zRetvNy/Ac
LP0Fs9CaUWSwpgyvKFcqsZjxIUtkqcSVD1RWHnN/dL++sfHdf9nHocrmPPLmx7I62EOzC8RpTK83
FqAdiplOilOWHUYkFKKtETAIUmS5VX7H89zxtyz1x7NiZNlKXiwu5CCSmuzTFx54fDcOSj4+FbZH
bPROlEvpP4O6JYQwIA6RIEY735aBKU0paUYxczK/JjlPiPmOrulKcrdpnlQUtpqd3jM+BEOvW20e
+S4G/hVKTBl+rmaMOw5Po3209UkuYWzQruT3TAVosSK1Dwj3QKbLgwpfi5ej0PI6s6VSBfSqNJoV
/uv5esnaxDaesTHpXjV7ZeoXG21awwFuGMnzSjjLDUa+AWxHGA3R8J+qioOpdulxCaFOmvEvFGbH
Ha03kxrqyP3CBdwkJOoBWoJ06nBdmudyG1S7iqUqMR2DYYhru2UBAZ4Up3jKrOvdPSFKF3SaC87V
HRvAZ55uE91IAyh7RclUe4VTT5srhuOfxNd2TtgqLJ3vYdxSs9kaeVSmrNkcg+n24NfaMHim7ZZA
2SnABlAR2tc1CaLXp0WyaRFgKsrYVtjwf/rAEXZa0WyGXJ056huiJy6avBdpNXba5dsjKABaILWL
oxLO878d6nh6oeDaKdZj88Ia3/JtOm0FrB7tP1aDvuXbGMIaM9eCr6vMVSm5qXVQpR8MUadWSrMd
V9aABexThXmvBezxV2m6AqQFdI/m7dXWvVvUa/OZ5KiEJvYmsv9wBOtK/TecKGbiGgxGxmNPccNX
auZ5SFidL1NtX/UK1fwx/oAPBW6QXveRVnH8MiibpOay/I/ck9jqqZf76D3J1LFOCifjTHbr9DJg
yxyItvZ0NNaBT1/9W7MeNm9JuLEGizHtXlMeMtId/n2oEevHOMH+28lLmN9uYU/VTEq66b+PQ2Pm
tokcS0P0KVak7OqNCZud+czTZ0umLKg/9plLsr0CKQuZg76Ktat3vvqRmxW9qkHgiDKfjokulOEq
/9PlgMw7Fl2DMeE1/hl/vw0xWzTo1HIzOgToB3bBXTiMBc54yTWDK/+cHEWtFSDkOpypQ25/8dRs
BYoXTSoqqcOEGJ+zrRZLM35lPs3OIbNQ3cbHvi2eCIqxbUnaPLjAJjbSdF4yioAN/q2BZTVKQimY
sKqWjUeQ0jnf4NAHiIE97pLfUE6S9JtGwZVwtzzTWXWfb3TAFfifQGZy/FHkoLQFl7U20NBQDM3C
hL6TogITbG/xASXeZcXavK85vyqcUIK4buONhAaeA0djopmBXJFVKKm/snNf4VcLUJuzCLfEQ6Ru
lDEypClofMfXIMzIJe9OgPZRWRCLZGpXVFJslL/klG+x5RvK8W60pPH00sLW5LhkI5Q9s6R6N0iS
NJUI3NZT4UDKKFBx/bK03bbrVwUjuOuA3idJtEKcATbNi2owp8iUuZY4+u+1sc4doIc+c4NGHdx+
iEPI6WuTcaQCkLBQ/+TwhF+9J7uwK3JY2aGr9IryBPgxIEvF9pdOUUKrflkadhy3aCjYZbiGyRQe
9T+Xqy0znnEfti4b53Dnl6e0jMYsZk+lLXz/4KaIR3Yi5CC4Z9gWat7SDkyK5xVteBT/X1ax8+LA
Kk8/G/CkkiN2FZfsuX8ov8kD/Q7c40XtGyZln552daKPo4V2Ud3KTmANnZRuhyZgZbyguUjJRSR4
1um2uW23R3tIt4rIe10yFpRWvQIR36CUHgK/jZJXpd8Nnhe5eAyjMtDo5UX+7Hg66iQMQUUvmoFZ
Q+J3DMVpFMGoP+gk3dH7ac2j7Gj57KIXiCjsDqO2B6bJtVXK74AhNE2QVhGI1uoK/Q7e8iiyhpcL
hRV4hz4XHIpKroeho2C7vDNsX61ZW+ijJiR4cyC7k1IJXkwQyc4u6ZfN68POYWj2iS6FpmfdC97o
m+7CwsDq+c4tpFjOz+qCaNZZ0/zZhoNXDE8f6N9mql3b10TR4Eg6KCsS85Xr8hcf1K0XIyUP840i
/EDlpX+sd36RMXvuDZy+oOBqv6YNHWxox4HQtVL2zFdCBHM7VMIzuQAn8Ot6CxVWHDuzUqQytz7P
BO4g/lHWx3GmZO46rvpIf5lU65d9ivJ7GpFIkpamaq/zJ76Z96/c5CD1YgdeAq1G1puqXIvQ6Qpk
/u4iQzyc2JvzVKCnYzlR2BWW8kMKaua/EfgJ9IAcsDJFcRpKYFyeM+QIaXowct7wd10GIaej3JAJ
3tvN95EQQ3gh4sRq5AnmW5vOM7Qkj/1zwLBWYFQ1av1LJRWzCytffq3gWZ1Q3JyfJdEaK0uGJ45U
Riw+Y+CAepPGbIFq0B4V1KwFy4d6s87fYWtTPfmL1VVgBql4sLUvLOP803HiF0h87EoB1TSTdfKn
ZeOhfCboQIIL38VdH/64SVTv69NvjsbQvYPzA4KHKUJx2vDXaskkr9RoA0le9f8Ayuj2h+psos2y
4LpCMm6j+pHpm6Dk3r2kxCCVviNzcIo5But8iB9LtYtpFVY1uzYUhOdMvSi0uq93BTyT7IEJ/4iC
nI0oSlWsX2ncSHf+2hrsia98fwApjMBJ0BaiNLzKWjTL2QDgRyTV+jkzIe6I3Z6BcXBZifhyoUIP
mm/w7bpvFDEAFlHClzZsuNb6rk0SkF1c5CsE7leBh6vYRg34f6sdmSEd0Ywj0A/3pVk9WEg2AQho
oL+FE5PHAUpg9NnIRQ2VhkJt5Cfx3EeNqNOlurqpQrhFTv8m+HraLII8zXIWY7QBzwAf2PMhBynf
QY0SBdyusR8eZfCNorWmqVQJHgO5sa3Co+vJd1mCCRRD0UAEW80ovbdusU5ftJjYlYK/4jA8WONa
jf8SPVMRRegtCeLuHYe0BDj1n9OyPqHPh7QntDSbK+cm8deDXUVTPyG5l1UIQEDulRIH8Wl42AtQ
X8ybx9BHBiLRCqr/I2YslgrOHJDG7Aey48SNvWnSI6BLrVdbLaWyDzpwAMgiw4QK4OaYMawGCfIm
JU2MUZkzBjpkJs0lOYv55XAHcp3O38m6r0LnkvcWux2dY8pb7poED6ov6tpWPJ6oiQz5vaGZldAW
2bYmOqm74n0dlUuU26Zi2B/ttUoNS2i0QDv6IisCke87YrThBgzhEoVNB+a4My/JEI14BK2Vj/3C
5SnFlK2qn5QNk5lAVe9DbXVCZvp2/rUr77f11WM2n/YkXCjriSmc2mlZl4lxThioXedi0NbwRIMm
jdinweMBtUId0oocVNfys04k/GNp8XewkiJ2IicWZ+vQiNQWw4FFVa6UqiMyEZTzGA09GqO0VBNq
nBwGnkxcYmVMUhj8C+VbkNXMky3SvL0FpXBJo/NPd8qt8EATd+kGqBhucGWh41M7f/WmHo7O1w13
SHPywAbwiMuRAHxgfET3GkaLTT1CSkNac6/xqxA+saaPJYnv3Au55Tbw9z+57JAoxtD4QbEi1wTS
pELKj8tGjLcdZTaOYjCTS298+YyYhCyYv+wCjDi/psi8MMrvMTtX2FMboPa37paOpDTn//SEh4iR
zTaIVNJu3CIlL1O9KVxAW+/Y5yIgpXySvKrQJaJH0Inqkkabx9TQkI83MWjYt3rRlUDbgoVGt7Dy
HvQ/gP+ZuAK/Af5IKievwYAAZ3aF5nXM/BEVNetgPDY509Mpu40NiS8wc27j9vqpj6sOUtYA2yb9
NDbZFWU2gA0+SQA5bKXnvpNi3KjZVZARXUShsup+ETjctFDeI/+Oi9vfSzPibdp9hxa4KHOie+8x
8MRIi2dhVz0GNefr4Fwl54wCwl2yxqQYiyBPu46DVSybreAOjIMs2YjA9RMnUMg4t0iWYrwXKcSN
iguD96feuVe1F3k2mChZoZTwjWMRefF7H/R346BGUZ8Rg9tSnYb6FAkT2jN9lGvHvfvObSuV7QpS
0LH4VKP2CRm3O1MPUmB+OH01tuWYoq05uKH5o01aBXBLar+zymCH6TDWrWVPXHVxZ3NnTNXWCeeS
cqPyQuPtm4p3QlQbUUOmEycQ1TU8CfER+98ydwsDASwA5RKiD6T3DOG0QRQh1gAuFrXueqaKR4FI
sJqrD+Sj7lfjmbYGrLjVHDy+XNMGdNgCWxLT5B2hqQgOSGZwEqdJNmGV2UnMFEc6fOAm6TLbNSIQ
6bkBLLaSctDLIUpYBCfofqFwrT/yNkhLzRjYOS1RxH4C5qavk4o1OP5XI6hglZfVkoB8/blWfE7M
CnBi9Ea3DsucfAc6guh2uCZEMNzM2x3Q6sgdcTRxLs9VkZ1E/5foR5w/8XN3ZjwwfM+sbv6VVmvQ
fQDHx48ipVcD+iajoXHTOdNxR4WMwiKh33bB4EeQ0SaXjL33WRNZxd4AUhTvebintKhamTHLDBMa
HzUATdw32hXCPUWVsi13RoLQf/Df/byJQbvSRAAYUsyD8jhZ8NqFHmCZi1M78X6XT8ToihsQjJZH
5pGUqVCsoNRD/x4JyF4IThMwpD5/pa3pPqbJQ2Zcf8Bfpqbgqnup3gj4Rb2NWNhwcTo+DWWDfHw3
aSywRjpyg0LT+AeaXorJ3Dc+K1nvHtiIcFD4RCdIpd7lxB6wCuMsR1n9aQvegZCEsAPyfuwAWTVn
bVSlhzkZBZu3gLFgsfVURY4QdTklWi2vEBYgoTHDy44rPojPMJUjJmHo+1TNa8EQwbt0O25BjuGX
xo6RsUGtmQqhTT+I3o1NuTFNqjDL6u4fJaFG17aBlGZOBohMx0Yyj+lSnfZTh6n9oUCRrMf6KpwS
ypOCcxUD+/EW4TM4YI87SUta6fyIXiCtVkACd19uUP7KOknf2NBsgAIo6W2H2rH32At1i69HPqvA
soNsQrD4Rt+sruIu/kwAi/9QAUt7416yaH1STP+omVyJ0Z+XF5+N2awJKUgaxQrrA5GyBbH7MzWG
g/qBRxZxVm3ka/zxWmav0zPbGtzjqEvUNMPoUQ56xmql+JW2hcBJ2cFDP48a/TbGenfzUmMsRUEM
STrPUPmQ9BUVHjFd+plhKItibF2GDRNvkS0sbygtj5eEMJEWqOSqQxxZWn8FGL0DRcn3an+lw/Q0
GK82O/N4jzaGAFHiXgf5+MitWwCca7QyC0U0IrJ72g7FOeRUbhJPm8nhS2TxdmN3r48CJO8+tXUr
CktS8Y3hdee+nS/z3T5o5bYgvmH5fA/gY79M8PjLRM+SxT54H2CVZN6yH6ws7FZTwaAch4XVY2bA
RciUhW7gnQIrkbJwGRuHaFPoHuuXHXgEfG+jp4K3aabcUC2pwE+jBDS68zQxlrMDE5nOnqxE/uQ7
wyhaGdCAc1y+0ShVNkRNi6AVM25D5sD3eETKIrexNqqs31dLFMs/msdkr5XuLoQpcZS6jfQf5cQG
BlB5dEuuV6HPq81+nuPOR+SlEpGcmvnVXUB1/m4oUhtGfSUppO+4wdTj799mwnIyOeXdyYHgIGiT
vIWzr01dl4fzWsyRicv2ZX+zRI3IPVpAXqrRUTRuLxsp0Au6o8e+kkuVATYPO5aNWdyrFnEPOtOY
ITkUbV/qpKNSt4XsB7Xp5f/x3LnBVYCDy61Bzjw+9AkOnMaDGPwCWEFvP40SgX4BrgJ3wUQ6uL5x
myGoeYzTdxlM8YBCn0tRYdPI0415E5e2jS+ty3eOz8FyLnaiomnNyP5KTA5PxlBlotMCMs4qI8lB
yt/9b1QxPnImrLDVcfh4nIFUTklLjwas3q4j0HUgGFsuI4migyQs8nfo3zhqGlUNOXHZZE2n8hyb
P05zUHuDO9FfSI/fEEgIyE1B1ERDoUbjoOYll8AZbYg+k9tCGZP413+POs+JhcLodt4/T84PhA+V
HmbQ8pi23Y32571o8cZ2wppSsSUZMK59cSZeN37xWPP3PnOh7SQhjFoNmL/xmMKv7dkh55mi+R2b
pbJzt1lNF1nVbhV+JP0AZdjbjeigmXxogAERLQQSLY7TaCrmLuJfLBq4VZS9NMBgyB47d8qsUzOs
PjUuTMjPHKmmVj8yxAVRB3PDZnqtrHE7ahn5iIkS105uMWch8o4k5+C10gGTqddGv1xSGj+3N9wz
0Y+KYASs0j8IBwtDL55lHNn7tqFUWtx7nAL+EKjJAA77YKEgifOPakfFy6c1CT/PBdLB55VGFVA0
jMZ5J3UELHh/0UgGP3LOXctRAAcGYXW5j/nxrc8FndWoAU5lo43RUt3WEvEI+M2a2J84q514vBm2
/Ej/mxwm3ERKoxt30gV7blstCtNnBlKT5DkyzW4n6gUZ56DXiuk06YjpqsC6knDcSiXmzrg1xxkw
mpvhMYri7JdiNIlVE10vVHVw8Hq4r12ab11Mla+2uqpcVJc8d3dauUQRl668b4BxCpvEbp5wsK0p
BhzqQDEqXI5Iw07l2SorxERrXGH+0muv9WKcJ7Z7mxEX30HiGC30b24Zll7gOQbjOmB3Ji0Xu5Ij
oHosSOnQ+Ze4uVQ0Bg7chYttOrt9ZbRJdMP9FsrVCal00e/DxNnlOv512TtpEYhbD0jOKgTFUY2h
w+6Vxck40Xxm+0NLSQqp+1sXm0qRiMvgbOrPnsufxr2qYzH4CJtapNzZXt4C9fbHNazKSm10v+aW
pL+6NlTKreW/e18MjsK1Otbw5TWqxR2XnDWDMxhvbsV2ZY+IJ8p6cmQGcvVCy8NczbWNTz1T5GzO
J2M+ZCGOOF9XCg0ghcKb2c9vG9TsWVwUdD3baCz2oy2kopkVEt9qDotzyF0W89S4rUPeyxpB/YX8
bEmPe3aNFtLLt4No7PRIhGjBUpUeUJsU0neYJNzUlpYI4OBu2f9b0OrJpP4f9RC7r9p4cukcsghU
+YkaUahMTLfNdLTtHiwwMgA26B44y8c10NvTUbL0whYYgFNKoZgZ7I0r0W/qVzqwV/UBwmcjK4Fj
xBq6s+q3uVLozbowQPP6WT3et7hyA0xGvAUh/uJKCcDzVNoEItzNBuEUviM+kVjQQEZm7vmlhJq3
DSnCSEbzdhYUXM33OmrKC911H9wjpwSqtUaGg1YOVnRlKGuKdX5c1emKSXHWnaewN+fuL304EIBM
HyZSHVW11PhijbHjfig0GNKd/1B+choZ3dEFFEwed9QcLD/W94HMsz/Ex6cVntpeWcJoW2RzLjBw
O7d+vbYg+M3lXoDHX6FHQ1KYRL41062xFg0ktBzVKSP3m/0yE0e3oymdan2O0acW6O2UQmcUJq6B
zZjnyfN1lsoAdB4GgKXn8vTRzH/l+D5QX962bj4MMNU3d5iWwgB7H4hErlTTUky/JCe9KPWFHMFb
2LalOCHb521fZHltLIAECNWh50Px/tr/LCt+BYy1GcJ805DWMwxy4JcjF7YIEwKQzyN/NFMwg3HF
pJwKH/HvG9FE3mwlacJLHja+28aKFDDXUgFaCS4Sl4VncqAJMRt+zJAcXwD92nGOk8ofwba7sVgy
dMKmge38RxSr5WiLLJ3o1wqlgYPRFUgQoLq6DExteXIM2pGVvvA3Bnf5d1piNGXpkQulL+1WanoP
XBumhJAnfHloFdwfidtkzPTUVHsWwkjFneIlc3iTSB+gZ7xJxO+9rB4BgA47Cijly83HQyHZw5OM
Nn0fVUxR1DGDFan/ZkmTtOnZQsWzVRXUH6mqsHJvZdstDPCLPhdKCbAkbMYrm7xSvBnMX/Osxaoh
Y7sPdh1JWroABRWawJ9qzKXagEGTeucQHGkL1HUUvWE5NkXLgbb0VQ8Jyx5nJ/VAB2CaC1/l+Wev
lpcIZ68xxkVk0VgYgY+BAhAt0Ur1ZWIuHj9hwa2BM02HQEmv0kFF7q8gWizxNpY8QKUqINgML/9Z
d9yOE82H3MIZ5CMdNSLP5eJuo/UkGEDPWZHd1MBupw/HUkshbIJlyenfZgQFAiydjYYDxD3JyJBz
pUPHlJG2Il6sFSKiC3JH5JNPA/9hEXaNouqtoOKMIMNxsTqNAk4cqoZPvmD6NxDOShaL6KUh9F9o
F+BtCCaH9uxGjwSwkmp8HM2xYGY9dffkxh7zIM3EUvWRy7MqE/Bbx3WsAgpPAXj6zGQbohIaXLnr
CnsM43V46fsauTg48yynxTRyBEjn8yiwa5uB6xFUNZK2W+YCa2Cc+u2PuDLMFif9/iHbUcocSsHZ
iZNt0e/NRmd/5/zfVnI9QUv+b/BizFYl7yfc7oUlegfLox6JpTlGO8fHASC7ewGMf89oYy1Xu0cM
m2ds5DGvxIvt1RTtM3E/mAm3pw2Fc965PcY1kQpdIgQ1npy6wRyAC13YQ2N8oVRmnobVz7ttEUXM
Uum/FDHoJZH2vXE6u9CJ2cecRYv1eh3SscGD9r30cxsE/tHNT8xQIDX4fJSGpBfaoo04Aa0GanRm
ffATd6DtUfX/MIvK50nFbLsJeBHIJ8WqiZJo2igtgZk7J/hw/cZtazgn+F6ZUNZjuOrIqF9svY5k
Zt7zeV/7UZSSs9QCpx5Zi8PWmYKwoiqB1DcypBeKNWwG9xzQ9BKA1WHMOmsNbcXJWOom3ReX+F9F
AY51fTbpuuBdx+7WF0zLXzVGiWpOU0C+9JVNMBASl/hLXkcCwrZdypB6aZ0n5S0qxbQtu7SSOd0Q
W/E+NzpWaHfFmK9vmQuQdR0YBVNFQFAlQuIVI5uKPcf+uLqezb3VCvVrLK4IDLo0hXZ8JARCKH5r
Y6Kk440IEu/yjhRUOoDEB5TtJVVd/RDwjT4BBLqxkxbjmc2h+ou9mHDJBs5BJ1ZhFr6jlEoGzRY+
yl1VdrWO65XSrMJBs87+XyHnRd+K6HQwXm5LeR2O7cs7R6a3HFVrXYhSnnS352Q3lo7F2g9OR66H
mKzaawWvPNtoNgcVvLRuk7Uj//Y7/SauHGlYSM09zoCNT879K9BcbHMg4R3N2KInP0YYeW1aWOkN
VTR2pJLi/ZYw9URPfqPMypotHT/ifEGzSizK34zf3Vq+tCpPfaaeYOrc+pv6QekT1QvESDkMyCA7
rUK1D3sztclrwoxNywWLzw+mnseGeWlChwOea7s1diyRW6wy9oI0ACHOqsNPqGQDbZy0vUVvS+84
kIN8Jt1Ro8/SQJiFZ2iz7qI7QFIJjvpAm29V8mGqAybNp/MDPRiCl/JkSGniYE6VkpE39Nj0859V
bBL+NUR/hCpvt+iHkbG5YqRh4+h+YPHBLirFG3mba+iJy5S1cc3ru8/Zg0MLK8M0eDwkK4XCxx2E
BJouXTMvXiKQ+Qe5GeNgHK0pZNN7pGtO6y04g/DKRnvnicbafP+G6tGipmrax8OUfAsrWtgnRyfh
NZrObyOCNhEaIQehw7CZrPVSXeAqNaLRyfPITahjZvDUEBN0KtSzNgemLyJ3wknApSPmglEx+nTB
BaAgiKhpXX4XJE68AQVC0nonocTH1evrUimUok7akOos7l9k+phUy3+Wu/gD80/fUZdMJbfdQNDD
V/IxQSV4iihTq1cAgnR7jOOKGZUe9RG/7y991ub1lvn/6oVdzjIsbd+EvSC9TqlOyJV9LS/S28uz
0yHsMSu2yu2h2dOEGueQgmwx/bwBEpJHVUUU8F962+Wf40kMbgUUuvaXip3LxmtoaRFfrb13D2HG
uDQjR7/ooDSrXY9zMCpGTBc3JOmdFevvbSR7+AYnL6NRoFS3gJjYOW7zyO/zUGCixbsMtNRE6qFt
Ce557ZSMdQII76M/Kt9T4oyzIQi5mzHFxfJlXk3kj9BqOh7g5lHUdcJi5UUamiXCWe0j/oyJz67c
lgb0vbzxpkjY7U/E5LiUYP2cHqVUsPuD9wO8VH37wh/dtt+GvyxGegvoINAsFgtkunOUMopEJZap
ALku0LRRTEUBT89Arv4KHFh2x8qwP4scSXBEOkQYHydKyzTPs7ZnlUnopsZ1lUFpRcAid9pmtpXa
CPMpToC3I494kCnBNfwJjQJNnAO32UPvYkbDchginkJiF7NCseJoQo0xv/5tvOoYJV10047W90K+
18oxvWYsd2iUtlRnpYxJbFGUCRki9na2OrWrMVvQfnUfsgJdYYoKDsYqFeFJ3u0Y08lHo/x3sRUF
oteStN25gpymgcpYpna7W5yeBpmC52R7oH+eSTYLI7PX3TDp42E5DDy1PWx2Djm8/ADNm/e0Q/Xi
my0lUPRDSkN7+9ampydpEVqwaQSRHRr5g7S4ojaAS55Dhmm3k/jd1VD5mVRVbhTbRsVU9Oc54ipJ
ygWCOVMnAjN2S3ucUOfgTkWIYQLebcxe30l6fARfVYM9q/xURGnVZcQRxU5yLeZDdWtCtA1jDl1j
lh8gclj1YwtjErmWI1wuJaimJM4/bF4fqK3IDaKMBhPRda1UZkAZ9e8YVVZipfZVTBszLgOdqN4y
CPk4s9QE6qMZsqUlu/g+qU8EJ6aEc45BgapQQFoOSVtyj+kkEFOAs9Y3GbW3aG1sbseq5+sBTeAp
5XQ9OFbZwTk7CY2MPTlgY+RaQylkGnEhBHzQyLQWP41/Jr4d/T1k/EPQq5yPWOhZtXT8JhyRcbF6
XYVN+vlclG+5pG+NPr4L/vg5rkLM0BVc1OJfy49mA+/jzWug2yZ/2zdLelhz5FrECy5yxjXTl7BG
vDvKlSG3jF5w3Q2pGEoFMMwJgLgWElx8N++uUTCTB8Yn1Dp/kelPeww/F7oQBlwUh39HTHUTCnxG
/1zG41oifJjNtJVq0M254RFaFkJ4EpHCWuHqTnZVdPDO3zwP5RxA9uS3sW6gRAQLdqaxbzFm32t7
ey3ONOJlw/ks9UHhIv4GUJac4b8DTcxfX0cnPKD8R8tHVTQTGzZDyKwarPbzLzPvP9gbaroaDxKT
X22xLWH5BQ7bzq6EhbVS2W4h3DvmDu439Adp+B82+VOSNz5EUblpD6OqY4+bBy9D9C8y63HFoYTZ
ELi9CW8By0YSwNMAJc73c3Z8m4tum7FPaahoChPC8B/ypf/ThuQEjOsHyx4979NW2B+iGVsK0FTY
kdee7e0JUOjCXfQouxsv5uamdh0ixs6jTvau4zRphRCmWae+i5RTovH9YRVxg6kHw00j5IRnuBah
4jTUl0SWlMomcdP+18n6Y3OdCVfRy5bN3Y+FG2Zj9yMpF4Izd4WSnxHl32Px/GcR+fX5oh6TUVz3
cdamYjB7RAEGYETB29SppA7y0KXx9oWObTJX6NgIBSiwT4pGo/S+Tj/Qu/t3/46S0DP0QMM30+nj
4tV5JrQFFVL95KRfx/Ytar2bPZZDhBOYsdZb+Asy0XcaWFwZ+bZYxIP5r3OcDFE8v0UxauBagANV
5jRiLoVz5OL7U234itcOy+i4N0sCHadXUfM44khopRpZRCWH8xfoSzzOmM3Vjge+EJl6VVeoXoou
ojeCDu7g1nUJi33Inm5C03fAJOaekpPYTcwQ9oqEnaHQ0U9VHX8DI6AY8NEahtVI20JSVE8xa1a2
YSIRLL53Ueza1iOTZuew4nW9hE37NfCSnyv1/wSkK4OMA46WD32hlvephGPvYYFMhTBH74yokGqs
TLdXpSgw9M9mWjyxBTHklcy1q+fQ6yy0P9OVVMclrnZ0Bdf3B28qRyOya+J9Gp9rQUIBjFc4tYMM
tSCsAGp/C7n8d9gExc31ZDMD9MTfrFiEQAx/FBaiPxSJxWfa+aX9Zvok78md0OQqRtsfDPpP/de6
37omj5ZlmgyexI8muvR2hCU+6Pa7xMPURJzWDC73u6KEtY8KaHVtb1NIFHyDi3Tx+sdST34GzzCf
aTmutaOOg7gJVrJHlDCVUPo6pBsR+gLk3KnzW7NoYQ3K0M8g3b0ppEsaxYcmKLCDgDmnVOBAag7B
YaXMv5hwW1B6JpJI8CvnTPinPT/5mGtDt26uL17pAFf1eLI0Y6CQ0cxozT0Nfg4D0TB+azpK81mV
FO1487wz80ZGHDVWhy+FT9oNH+fo8LhfqbA1FyzkkB7qBCpDlcIYJEKXi38BWrtqLAm+zP8KI+Qn
XZrYo0xae222tZeMURCzFe2TqJ4IiufAtfWtOJDPbsNwoXxfSnc4emJesxh2uluMQXj4T9VtqB5X
akE3bkxsUvjSiNTD+8EDrriMsyOLGRoMsARoS2e0hm4GYzZHDcf0UsCflmAG7I3hmCxi3wyDXkpK
abyd02OVfdPg875pGStsLVYPBe/0HrcTF2JVRt2K4PLzJGhgp2xJMRuyKazYrAVJr6bJkHsaGdYr
0P1tlfooiJzzdG0XTI/LY+LARV6ui0y4+rZY8UO+s0l/nlDlaGWInTHFK++rzH/ZcvvvbY3l0Q4p
3Jp1IClnKe4dGqyfUi3+dpHMTINCMJowt+oG/rtK6PmUYrg/l2RAs2ZbgbML5wcMgM4WV0+IIXiw
DrhhwZPP02yAaFGrXPqndsydw1ovw7Tbx8fISWWHP9gVbXUk7yjaqJndttEg0cQRo8WmThhVZ0sE
dc2DdPwTmZrmV4eTDRDhWoBfY4+knfe+LyNd+Qa9jxEseZgSI9usTVRgvvfMEQCrkAABd8W0CUCh
Pui2WTlpOyPnmXz0ymtJSFQetpMSZsHHNxtqDfitj/YVhR9xpVCOrBJNUcPVjFeSIBaPYlYNtuIu
n4IOChMq2VMQxsriKC36J4jJDptw5G2/8QV1/XbrpxDfqklL3JWRlLx9tWOqDOuIPJcx760buoCA
mWcgXLY2xcNbOoNqrb+ykjlzg9hWAMCv6d9eYfb9Oh8a08+2jATLlfY+oNfViQ57g+xpPPtNcvAR
iZZ0FCwKvSNrLxI8gbjoUkockJsRXphhm4KjDDfBCtvCKoMBiUCwOINCCPXPanI90nxz3ytkB5x0
A4e0uyXl0sRMCm7KJ75iieXhcUMtH58r8Eh1B9dG0F7wi+jmeEr48oxdYaI+ymbUn2+u3MbOS5uB
IMrQusBh3mmnkzSIBC2E5LQvmGclGY7RciTFc16rq4vsRqWq9MrPeESdqfDP/SbKb97whBCB3VvU
7D4u38ICJomoBUvzdR13LtOwV+vL80TMkXtskrt8t6QMOu+FCjNeA5SP5zDS+yyBGYxYj/9J/K3J
9uHHgM65sHiTLk562dLjJcdqbTzTjKPmrZ3RHE0mDC0odi1YK6EiFr20MUFwjwdWF13PthqL9pj7
mrOpvt4XjIrkcduX3GswFvMAxtAgMtWwvajYvuqZcNgQAZZE9ZwPGZk17OKYMTeLkgpuOwCJMUra
UDuqqNFUye+iZFpJE2hYetKcwa3APykoeQ/dYUc+4AYp3j/DpVhtzNU33CpmC34A58qsHPWzcn0u
smlvKm7aMNlJsL0cXAviH5JLbqguoeIVRL0JEUrS9WzYnUR8dAprYL+Z7Wf/5ekzipVt8DItgLk8
a3lp9sAfTeA79T2dlKfFoaczsu316EYJ6t5W6Hewe29hcx8GX5nxcg7UfYxYtrHqPtFaTxAOY402
S0uyC2xFbYOgFiB8oNgg9fZz6FqrbroHn1u28fnWpYjnMYGgJVtRx08HI0iH4uA6QyTWdf5VoHGz
aVJQt3F36F9202dUYGoBnMukEnaN+TTiPvHKbz9g/tjDD9aalgI7AkQRzDTBBbQh6myKIuBU6T/G
tCUG2Jj3hJEHdIDn7wRMhPMaamfnOGVYvy2q76MjqmopvEy5ycL5MAhdUTr7RoKskNXX5izM3WeK
DmL+eNX+H2kVcZz+9gZQDRhgQbtNonVlDgjuc4CwLsfpL/r3ZF2AfZLKdwheQtaHrWehr6njOUQc
7nf6A7JaM6jCbrYtymw3oixqw90TPLNB1VnTY6UuX7F0IQC9D3ks83ocpYZi31m08Lhi4/lWaO3J
MsyyArQc7xN4M/9Y3vhTuhwo6JZsYUkjUBYA02MASTVlJChfClSv81kEtI5kvQq46POq+qWlTwce
jeljpFyLgLd+ELD5VMwWwCXzi0tvw0EDdlvdOttxsaWtN0sQyORyMHJmtvju40ABOZPcyFQsOXZp
Zyk7qZjatWA0+R8cBQz4CJeKqDMnQR3T4TnSJOtCtZju8UXgXajfRtsvlXqvzmER/zI9gefv2QdN
ybSe5ZDoAaZzWYkS7Tl12uIvE/4QO2+Npds5flhZ9KaWyIkf7j3ls0gMETu6cakHSw4vUronh7o3
VdNEk1oR8Kq+wPFetSCZX7QtbT/Sc1uHJkLvsLBZsLfHEewWHN43Orv4tsg8qJYch4e9ECN+ctkB
XqtUQz518fmhna1Kw7nVYZZSt3toGMnSLTIR7SSVmvLfaYWekdIDLKas8B/3R9MsjOFDeYNwltvp
6j2cn13hTyilWFxy5riGKCZA75Nw1jNzJHWVOCV/ClDNLQO/yC6W3NlecexHsPpNEs6VpxcYEhgM
aQnv/IjPuR7pDXWZjydCOjhfnrUAGLf8rS7ZCwTcBlB/TzWjBIreEUb/5arwQHiMlCkENW5s5vud
4dULDqficTjc2nuT9dQa/SS3I6Q2nH6wI03GYJ4mNN5UqYKdRvC5uJH3D0EFku7BEXHPMtQZesjU
250TkZSLzQNj7Vw0G83PZTJaHU4smdCMSyvmnuRAYCmHOlzet9wkuau+ASonsAdItzL3hRHiWAet
WWzHbkDig0ZT31gtkznLqeE0oASr9DhNd52ePJiDw1gBrjegzMaMEr7Pob7kkN3GGITxkDahrzXx
UzXEzswqpWHcVy2JZTDm3kjg62k81gtUhW80I7ZjBsz/Nm0XC/OUdNwtUlcD6EQPqpSnJsqHZgJO
2MhqDVKVtMoWfC7AfLbQ74LFS2AzYHSxGgpabjJHMmdfkDXPGH5H4bs6v1qR5D9YmelBTWbS0w2o
38zVIY0xyAmZB63AB14EBWfXkKEQCkGSA4upf2jSUmb4sR99U8GAsSHCc61SuGTHs2zPoBeeppXt
ILYBP6GWpm0vrTcYeVaz3FmkI/nDg4eXKDdJKwVkrbvc+MqCels6LI5lPc4PTJdtL76HIk6GZpmg
YLjZz3enBcfz7MDuqwZNwrkWfB0fd9EYKKR82gpi4gDnnGhZkYVB+/zVDBjFTmLaDL7Mxm8Ltgxl
chVK8t5WxjpAVeyQhMSvJOW6k1yPHmlaNnChwimsaKfxJMDAiHJeuyykhOQ7OUMRv1BMZ62WHNP2
uSOLSu6WohCg1TRYr+TPETq2cSzRdqRduQJg/1TR42KSaZHENUTDHeEv6VdNvjhZogVwhiXi+cPY
JDu0YnNySyNVUs8bBocn+UpwyBrbYXMea/eZy6aXx71CLg3q8l3uf/wdN2PiFgH7Q9OAcEdmweNt
TKduhJLqoucOXH0lYev3P0tQyegvWP1Qzt3Absb7398AAx00ivTLOSH9gzRRhWrlxMeKelibYpG5
CN1rrMjoxtD19zeFk6W8bXeRoGwueglZjyjG0TwKYoyI3cz0Z7gy3tioWBqR6tJ9a92JtDIb/cik
x2zv+d5bErsd1qFsQ57chNaoOl5H/fdUE58aB1i2Z9IXWvmNJELNEU8JhNc+v0MhQ6HuVRb2Mzy4
Vh+4qBHA0vMLxQBZYBAf1G+fj2qeKSf5ruTivcaizHtFuhcgS4gUFJVyg8/5zHS2V/APttYqLKz+
/XYM9ul8gMuSWqdWnevkRBLQ1FEnXBfYNLGTADQe8ew1H/BdJcpdrK/USHzKvDM0btaepunEDdvX
NNv5bap1Fr6axepron7kyRRk215csph6wyySxguh4yZ9fAx4RtVmN/lpjM+9xGjSmK1q3CNP92yH
czG2zOnppLD8mA3ZRyyRHt1QVAWkkXYmMLvbZwMygtU0H/iXUtx0RLJ9r0PeKPfn5fZvagoSE9mQ
71pzHQpWMkFt8KFHnrXDGYscN+MGN8l83SMosJ9pbJkRm7XMQs6A0VvKtb6Pcmsdl9KikNG2pqXP
rmCZ9m23X57tpQ72bLqms5MV1cukgw0mfotbYj/KGQD5UbAzA91zsP7iJwD/23NQOKdX1ovDSeFl
T3M/iRdBodskH5RMhQuvz1OOyScRaYfzudxns/KRc9n9JpyOuvdMItycynfltoUb7wxRw/fj2p23
GCcMbYcmAVZLwIm3yZ4ESUk8NLttEYTTM8LgOy7kFpNFAd3gV4i3DURsibxgOz2j0B0B/rkPTlxJ
h+LkLUmzInwEx78gjgq8x2LWkmXeQvpv2lQkXPdtTFFxPdeGM6uRMM64T8Un1zhcw9WPhvxC5Pwd
PrRh7Vv0astmx4iLFg4/Fmy3gBHnN1N11HDrW5hwznC4DE1OmU3YY5aFpUWZCej1FGxz7hS3THUS
vB0muj+6TQEaAeDSUXM2lpLzjvR/urRnP3csito3O5c3+3JTuO2702B+KIE383AmHwKcle2nShVn
7WBYmxNUCqMWBM9lS9uDYWAJxBNmOVKhUD/iiBAlw9ImaYWgZxkZbGwp5ZN2YCTzexfzxaXQq913
AdynBgSq2zL61Qy68FUVcTsGKfDG27+1teaWz2PCj1S4EF5Yf18GgKDCfQ9cGw0mVLvmjcOosrEj
VHjNgVoYcV6KYrU1lPKxqRrj9nZ8ZTulW1qSwbhL3AYW/5hU6vaISDZppZ3Se/ccnl+YeyufglJF
4Iuhps7YmkC2d1FYKVKMIWzDI6koyYNYdlk5/ngBeUEsh6uN3sptZnq1hDPeq8ErJf8q81v5ugkt
wbUstzIRbmGiF8drnbVZiyKLbsOp6i/lpWcP+RInlVff3ijOUqzWeSih40PmYS8oIznwWOMHx3Lw
i3mAJcakYEcLkKUZ0WW0cb+Gq3rEOMvzLawBNFBbxorHVQLBRRJzzSuw60645DPkoilrG0gkcsua
HQ2uI3oQhtECB5QtXAHY26B2AdDFD32tbuCkT4eN3amZnk/qX+Apn/gpGzU9RtucxaQfi3/j39Ze
n2HrVuFFVSeI8pVun4Eba9LOSiT5tMKA/caHJfR0z6FaoYl27/7wzX3+y2Bnq4ZoRjLGrbHiMwPS
B3nug05Rfvo5sknpBXsr94ncm0zS+WIaXoCq0da5QAPFmZLcWjHi9O0x1RpaN+bTnYxnasIUumHt
M6BAImj9J81XPKm9DCSBaHHNSefkRzsrMOd0OPBHJt/8TZOp5TTL7f3Tf07X6F5H5GBYqEvSZY6D
icDPkR7RMoD5BmFCsoN9cwOq+rp9cZE3AeIqWiC1qO4QIVx+8Nx+jXAeCDSi9mOKo7dtG7zz2PbX
z8ZJ7i3YEke+j1HgFgaT4E1SHzd7s65F+MTGgbYPjE10h4LgHmiDHb7kXEhm0dwwxdZEircrlro7
iC334YGAUKrQtbN0wryKDV+4r+F7zcQDXl46ufSBn5bWIOgeSAMcWpHj7EBF0/va4elP9B3WImnE
8OxjpJ0mX5U1rZ4h0RfDql5wo26SEXgld/x4AZJEUeIf1aym1WQ1YUwTBWG2MMty5Ve8u/G3uyx2
5ME8Eadso48w6atn5yQ6IpK7FMx5xaUOB7YMD5CoGNp+6BsubSZdeo3WwzThhHIFMTgli5Gn7G2y
HNe4Dxi5QwZk6T5OYtFdL21R+KYMnNqGhOKTD5Cgg3bLdP7MD2EES+Tq0tYfMjqhmaO8tJyP8uRJ
Xo6hYqYiMBpL9B4SiGEo7CK9SOpljMCMj7PMvWTQmANsJbkwRLYemI7uskgnLITIbdtuYtSgtcYA
b6LBhDMdUcZTrqtIHqqmLe4hkV2XuPPANjp8fhiZydRquSJXi/I0g9Wk7iOKjwteWbtbk/czwmcD
5fT7txhY1yGP6caEZk71FNh0OytH+/NhKFBay/sN6/TQwM2QyQhK1/H/QLl13Mg07Bhb8LE3p0k6
vVBVMmhLnzYPCg4YJwwjh3PmFKZmIovOP8nbarsrcW9fzEXQVZwlUPIDDjaxRUPl1RBc4pI1RI4E
vbsSkdv5vE4JVs0GmsuV4IUwCF7p3GcgpuV/9rLoioJFVe2JESeJcb4T05ZIyfxelQwHcP1bB4QD
EK0iOvZhT7lIpCRdnDh8kP7MhzOtN6ckktXXvQb7qNZ1XEThqKKiVQOalzAS3cVwZkYown+91NKq
B+dQ9/LrA6wdKyKJWTcZKbq78cS4EYO3Gd4jPb73VlOFm9bv3rgbwJB+Zri9zbeIBT7bMyTtsGwU
T7oV5OLkxwNw5OkzWGpsaqXXLsm++aZbtuy5B2e3pBfoV2YfhkvbspncXyTb1uADij4zkxkKDBIH
bskX/EGpOrYxDdl6wkN40e7akeIEGaFf3QqF7j9z+HlUxWsWot2xfLM+2OuXZBQH6C3AaORCuQkG
DJqtp5fZaduvEHLQJXTsgRUyJ2HVmZexc9WZIHulP4GzA6OT8pUmJj5uG9M9yA9+mWxoHlG8CGYU
Q4t/MKjFucYwoC3qSWtepl91NJGOQVwqEUazAjE4Pb79VCmDebPOyvvfoXO40xKZ0JEa/YN1viYo
Yf/S8+2gSJ8Kq1I6TvUuCp3h/lGsHxW77QwkxbWBp/jKZD+bdfCO2tHPlMzjSJPR+36WCKTmC5Bs
MSngG8qAu6EoFZ/AHsxwKnw8UfbLWoZnq7zZayoFjfl52YYt5yGKVEE18/U49U0Gror7f65Mhtsu
VbH8fpKwkPnmTxnX/6IcmNbB04hptyAQ5UhmQR4cL8HiF1aqZgxv38WmhJpJYGXlAhfVQ60YgR1h
UwDqCs4qAB80rResyjFh0eTXlGtCUlSihOiZLGMrk7LswMrecYX6oA8ayePTHKr1w7zW1/WWnBNx
u+teDsaUpqOUW8nKVnAlxPyhWN19zFioujQUd0ZqBlyhjgfY6fHlFC+4hjwpH0M/2MAqq4RiB/Xa
rwG4jDknavLoZezujeEjtEOZX1BQIfSPQX6yXHHyL1++SN4qsqujMHtCp3y26zlANUQNkrz2ixmk
QlfotVnD8uwl7WVxLWPH0wfOTjFbl/uuevX6b5RGn7v+9iC5RZmZ5kJAaENnV9teVhvknLKvoOqC
OxtunWA1Fp5V02e4J2myJ7uOOuVG9jMw3Rx6QOIAS+JgmozL/rREC2LUwzIsVMlpcIS5E+PBysgE
JVykDYiQC/ucJ4dJsCGL3/QmUxDyblKHOmsOT8IksNEK/fcKM8R4oQKjGxKcG4jIeUNCy1W1mtRN
7XkXAXJ3mgIYgQ9Z5X8CvcEl/Ht4UDUT23LjZnJ/ToFTOrFV1pTfLF+3RTwQss+OYGUnnv7wxlhI
C9kyAPALZvE0OjZhOYmq//+AegFv7UbpjhNtRl5nsfpvUZbbb1vUJcSm+AZ0+yT8+ZT7OL/5R+Ib
J+3Zz5gCHfk9GG6gjHa5cXJqiCP9Cxv9iAjSo0oMOHvW7AbYlBbrYIq59ZvpWbYl29OW2B9axJPH
pQUN4KwOEnnQEyBH0lM8PtmT1OmQk+6knScdn7aWkbFbxhg2adlqdOA/LxZEHxtXFJQU1JpljKP+
y1Qb/aiK4QuJL856vn2TwT32ty4oDvYYYduBl5NdiaSbPUlnowexyYvoxFCEm7QZ5xuhfF+kdgku
IUi04fvO10wAF1ESjpiHRVLB3iemIdKREYzK91lch8NBMoerI7qfD5v75DveY8531jhSwr5qqlDG
gCNT1DWWJuOAlUFPvwhswB3SOiBnN8TB4sOb9sucqpLqHujEAkNJ/tLnJuYvfphlzHoigXKdSmpC
3fR+62xof7FsUev7VBGfh9SiYFJWRuFYTVVuEKn9W2YS5kUQ7yYrCt0KqU2PhckMYWOalNlvS7kj
RlddzUQIY1MgX9rTw3IADdcNokDASxLcOq0nW6X19ADUaU/1Am0t/jFyc2fkcdD+1m+7PQqN1UPw
++n3g1EP7IX7C0RUljLGpkkGXAN5rjVNytq7PyJ5u+PBlP0wlqYrGne/RFMBA40BKv6E7RG24dF9
mkd/rtHjAhkw0gpkeEzC0ivdxfP8DecCWHtvF5gU9OPx4cZyhaC36D0b476lYEnBJfqYQIGJhXe4
ctMSuNRTzO8iuVn7ygE6hIi2OXhg6buKPcYlSZ1CibZJIQCeSvCgsAWi49Mb7n+VyBBqcMSWTOqm
aOLSq5ciZRrPWcZ2LnylHbyg8mP5BnlmJ2OMyCSvTWonGk3qTZZRFr9cZcv3c5nhN812PryL0cMi
+qHuT/2nbmxEOzUV0z7ixHr16oH5sHK4Pvg9eLNZz2vmI1N1nV4F3/DnxeXB4+WMfOrZJ00tsSVj
qpzbkzvssbRyxAT4zaXje0jST8n05A0IdB5tVAnAiLuHBgbUXqm5UeQXLDlHm1PzvaMdnTUcvqIW
XKE2zlct2HDSREYHnC2RNDkhTe5TBU1g9QoNkGqJ+OxXk/xdvV+H/GUqh8q6RioJujKpJI+lqQYk
6m/1qjV3wNYbqGNxytlG+sqKECgfckKVt/Ved9OLzHiuKG5x+jSF4B/6Zqsc+iB0CIq1FuuErUxT
n8bKzauElTwJ8NICilW59SM9sxzZwiCy/6ryQ8xVrdsgzzVhCZphzUHvFKpF/f9PaTy88uOmjEJG
PxPuanoPLoUikdrcmWLUC0SM/ZaKnpjUIh0NabYUsGfI8ZYa29mjpV1pN0WFB5AiJDrewT21yE37
TJQ+hp/y42aVP2KRXpkJj28wWs4ccId2m94OfU0A/9fHUiaY6bdvtMkMZs7OP96cYqG6uAz9ac0a
79HPJ0q57QpYyDDT+Ccs8vtCN3Y08kVDNQrC+HNwEXA6XpJYHuc7maT9wFByQ8yTeblWlMG6/fbu
FIAdUGw5WS7WANB1uTNC9MeOb/Zc4cmB5KL2sc9rLQw1A9obi5ax+PUI2+V8iq4sM5N/8ejCxB/R
Lie7IwAXcWAIVKJjWQLY2S1RM2mRVQsiBt/Q/Vuj87YQ7+NL3I0FsjsUFiqRkEpo5J+GPl6tOuAw
QF0cWGh5z1TimMR4ZmJSz2TB4BcRb+K4IRSYgGJNk8S0gDTZlU6yxu9bMKEqhccQO3OmsxVAPxBG
s3mZzwrWgQOYL6/UKajG6cV7fgymDdYmOtUP1bH9ia209W7XtXBUotVPf8k+tzp3hVUU3XqBOZjO
QwMv62FHuD3J9Md+bSRtE01NhkXmKmuooNZ8HVMZxsMiNkD+TUL93wc73s6E0iH3AvFlaJRwf43n
hWnu3F1d80lkKpnUfctiJwWKpyyLCwXgF0vGTpCg0FQc3/vWcRA2m4uFyGVs63hByKC0On88a8hx
Uim6MpIoiQAH7gMGNu414hHIhZuinsPUAv56P18FrjTu0F9zYObaZlj8XvCNp65f+HCN8wM8otyQ
FsVSPrsQHJeDbXioc9HbLY6S4WhSWh2Y+Gj8EbcPekBRgHMehZQm/v2DW8fU3Xdl+SH7XnGV2928
VGgCKVlTieQA7SB2bL6dk3Dcl20eMGYvmFSRBOnW3HhcJHgKmhZLECzI0Zx7oKeqzNAub1HCLVAp
Wa8H9vi1fKxRWOUS5wsYg9LLDE7O7//conxg30IzyGRq8IEquY9WL+YJuyDmyCZ4dfM1oywYu0OT
natkzCLOLls2hHAjOEIZq6b+axjO1JN+kyd7Eyn7xLxLvl/ik7h7+ZxmyWkmDSlsgoIbiPAbMScm
STawQHakL1oNSnUNcH8MblrF9QBFs2gjuqEVaB5qvyxsKfVIIY2813CmDPEePib2kwiPNpqYv1N8
xZfhjMXT4TuG0Y5D6pfnXZxFeUW1V4eB52A78akg4xu6S7dKJh9q+8U1bS15YCzstczZPLlQAQ5w
MjQyTymAcX79xt1nspo22pB1ywDleB21yCKmBjNjtgptU6YPivwqc+5mSV0rSNpsPA0ejF5ABWHD
wwlj7AlK6OeWEm1RLNS/hAO+29X0aSgQh/TcIRGcu2A/V0xMN8L+wnFebZUc3xghIbUxffc+mGCH
nHTEZxNuRidYl4QtK4VZXzx/QEQTvzX9LbkhXSCO+k5Fd9K5LwoFchEoPIyfzHBEHMJhSCz9YtJt
nM2ttXI15z+XJddrA3ZMzpJRbjHhV8trspoR/YOZnUKaIEBggw/YeC5sJcRhtBnCDdnOomDoPam6
SwSU8ES9PhbZ/LkFY4ab7HNSZwxO0yi80IDtXys7Psz7/vvmdG/SdT84QHdE9ue93vuEX4Ar5jo3
g1kmHL7X+SB6HXl1c/i7bnZyAlUGBqF4vEhcOGoeFiJxeGdsAm7YWCh23ydJc3RadaQ9rrsLL6X1
kgkV3lROLfdQw3tvUGhHhmV08fabaL2ybBd952VGO2NA7cpX2eyKn0LbKJlHUJssA8PN+HnggHNL
3M0gByEuxszE5SEG8qV2oOUCke2WGitMlLVzG1hV0P8u64IPFMqZppEceZMGd2vDGh0phVA+ngFv
vJolUiMjpl2fHm2oOYCe0rNKIJN4fkoyTXoXotLsD3TiHBO+Ak7rDO8alWdS+/r8QRU3ttqe3osm
5HlKTh+3RWX57cFPYlApieYDdkdEhvn34Cw1xR8J5QLRTHMXkGW8SERa7QGk1MUt5TYfAdGoSiPR
+So7pcQfM50uMjV/KFMIcq5WwfLBHTXxoVEf0daVuGkEygG1sd+QkwuvMBu2j6kbGwTJg27NTtMJ
yadX7hlV1gE4J61IFnOcD55U75uIXDxdztgls8zvWSMB5aE9ugwel9vHEeFvnmmef+LFnxtlfvui
s9B/Tbu2yWjjwMkkH+d8Nr8ijQXH7Pah/dvoOAJ3enVRvmabmi5PqsrpejjplRLZ61uvGzynneyb
bv4tXlMTRi/Isq5rDvlTxOJ1WeqYz8DHLnU5xcCExKX4hqRU5SFlAGOyNMaDKTHRyaU5Ydgv3jHs
FFjhd7OjfN+agetkXq6rpTP7ikwH/hsUs6wii6CfjSF1mSqoMNq85/qx4+O22f05CpyAFoVHVyLD
/MttESNGiFIBdowPT6mTcTLQfIjmEahyZJ8pqOxrOp/T9w6SugRU++CHYM4rTxHjzrJ3y/M5YIEN
pySM/4ymECVY/VXx3Vo+gqbhhVjmyJHwbncbrl3YlD1mJzDpmtYv81LunX6IuKLQ35HPW+mxvtTi
BUfPLT+npa+URbJhzS8DP8KTu2OYqRiFkDRhKE5yQs7HQh7VeIaCo0914AzkTwD6ElNh6BkKYsZo
uE6L8dU3yBd2p/VJg7rpbFCR1qNmyOzd0eJeivHWDaq2EmLDurZTzhgrOrZ1qRYmxvVvv6Q6PQRq
dq3Fb1VKjXJ2ebvoQjyiuD2X+8emW0jexOQtrRsfZaFyxupa2ngs9JvWB24S6m4D2gGO2JKr+YIM
hLRf6bvujkRpBCYWr9qjOB5NJJDrEQAVy1pDBbUD8ECfxRRp7j76UoR4kAKLdmaKj6Pxnnn7oOHl
Qu8sEAOla43uxv7FQHOm2DK1s+aUvfX2QDMdfEvctDn5AhkfYRU8kr7aAD0Avqd5eQzItqFwXjy5
Hx5L+TnM/q0/EdKgTGoIYTSWwi4rr00M7Ltcx7UfSkoDoVyNGe0oV4KAX6iVRQugcDHwbHHsx7m1
KjSHYbodBZbGcLvf6j6Il+eggHpNh7kH1KipLdzo1PCSgziCeHkenx8x03Mfn/Kryz48KOGrNAXu
gLInaWa4FCmNlJYr70mFOpp08kQbbwdtorqkuYnDy6dqmumHMnXO9WyteHCF+/BceKn1+1BtL9I3
3E1bfdbghFV6SkoddtMW2nmDV5l6dZbzvBB4l8hdNRkzlXePkYnTezlKfwRkfIDD4A/2X9o126Mi
1l4FxktNLW+5JpWbhVDhRhVzqrsqmrAY4L81cNz9xXFZndUzXoEtKNsCwArBosVlo4e6Bjh+2t1N
FACDmB7Zri1EfGttwXRpxGXbGMYuxhxldyHK67nsL5uITPzF5rTwe9ayF8loclJFE954N6Qanolh
T2KK1WKz/3rquU/qnQ8WkGI0LtoJkmWJR/bQusE+Blx0C6Pz+Q3+zSfM9+z5Ld1rNwBUg/wCBmcL
2V1IwLtRuO7Z0oYZQJirbgkfev25fF3YO8nxisbmGJVjdKt0uf91Wc4B/9BENJ+Abs7oxsvxHDNf
lzQHNb6Xl0Zm+vF688RF4RAGzqESQp3+rPkRyiifns2G+C69sTp8lKHJ1cOizzTjqkMAu9j4/b+W
kYb4e2Z3Zn+mKbUlUYjVom4X9j92KOLDKX3Hrft6A4CBicSap74fIzGDTN97+LYCKOTMXuXM50bL
acwE3PB4e9BgCDerdu0uPbivMIsfrSnp4IDTbH+IGA6isgYVlnk7KzJuoUoUaSsUzlaZSgF3ErZZ
9aKCTwuhRQQyFYL3UM5iWpr4nwB+GCrETt/+uf30X5lexZn9Vqdbwmr16p7uRW31Dx98XtS5blAp
gDzFv/DgwWlgcv485tfqcXgrp6o2n7P6MvIU5U0daS9oznAing20Wyroa7+YBjGKl0ONWED4R6zg
dG1cAMy+e6771TMFJFD6c4slmEPOhuCif+TMEPLhSN8ER0eqKbfqI/h2xn2NNYVO/ncLMllDna7T
QTxKelA4hZWNV75sIsyzOyVK/6vM8hu6oj9BS5woQdEkg1YuPA6oUPhhL11ot0KHCqH2tMHv88aj
e6XHoWwogG3evNn1C3j0ey9gUkGP8rGzSIw8MDp5Zs2E6epT12dsWPKyXj1qWdus5Fn72b3Xje7E
x/OwIPGYQb1JqCKarzmbKZh0GGAqH44hdsFiH9PcPRZFHbFHPGrM9OYmBCimbHBnW6bSlCZ2iYHf
0qvUAFT5kcBS8jnyCQTBDLJAI3eVnnD6kzf1jdUa8bH58hnJLewqHqZCyo2emZedDKwB9DB6/zA9
nfLRtPWTEhA0apuzdWIlNnpYe/Iba3JszoQsFgPc7k1Jlr+fN0xit6f1F7GYn52DuzS67ks1Ptgr
BKoRhdG01Q0quqZXrG+WqarQ9oNBuZhaJw80QceDh1ZaQ+iSi9SJ9ZIiCzfcfOlLphrVJS6NMGvS
SD6fBVmrkPxcl1BzkAJSrw8GGO7CIwvieEXPdlcNoISn0szWXHgm/F897EnUWdrqkkrHclo9mPUt
WERR3JLZTlrx2uVc7eaQoTGoNii1m7v6Hob0jQN5R1w9AhIUWuk/1HCsB5FuWyxtwUKta/h98z8m
5OklEZWw3eoZUJsZ5YK4rE6W0+aBxK8fKiN8oHNP0a+guG3ThSqY3lq9ObeePvyCMapb5gNtu01h
wUeznxMukSCmXfkYpX37jI6rv1Nezb5YB3imbbKlPQhuw9/MlHHCr9Oc7tR9IHbGSA0rHCnH2hWs
Wr8TvFR4vOqQ4MMQz2NKXDUi0EAxFLHHNAaxaN/7DltZQLO7XdbKO727ijUW/av5Gd5Ynyx7R+t+
U1cvyDrGKD1xr+6Aw0rncrwhv/r0cmp24Yqe4GxqJT5GHTaMbzl2vM+eAQuZlUwOgBe53DAnVwmc
80Wya7bWV3xILw/VAJDpZ05FdYLagaF4L35zIaSof421r7pZkEht3wDzARKJcfIDX2GrrA/V2SNu
LeYyesr3KFcnd+IcKXHLO6t2R8mKU3TTTobPc/fCnE9VPVx0qs8StqoBmC60h1D7SBqvHsXkFbj4
1C2QuT/iS1T4Ut+aZkSCT2o0/nnXeCylq6OhHLQBU2eXOxj9+n/ffAMQGgRI/AiKTL46laK+jXnC
i8j031kpTv1NbLOCWg1HumRyrTlJYS4A1xAmZO+rCfDrjrW6V4tIajJsRPA3g6NRLZ95XeuwE/VP
YvursiLxGOQXJSqTBEA6szeUd3S0la/tHGJrSmPvjsIEK9KHQ2ur1235FNJv7DBP37quehzUWAC5
CMHw2xbTCNvvSkQpUevn39brY2h3MIy9Ax6hAffej6PrJvvfRCLlAPoEYzZCoq/c7HyjcJgoX9v/
9Kf9axEcJsOVpOhZOMb0ZlnlKoq72Dhe53xRPT29bMaRiMsgMnLFl0mhT4z5rCpVjSY5fCitQMxn
f/9JJelPpc0TGIAC49aY5AIqVIvG98f7Zw9HTw7husvgMKBe5Chwpg3t5q01uClieY12IMs24/sz
pEtIWTjrKmUwA5cEGb3tG0EL2KIpx49Pf3giD8vCqKUUi2Ci98VOKlJ8c2AlYwBPAUe2MQMtgdmT
rg0pxaMhcCN8wt+V8aLfKag/qhsVamrYWq4wlzVbnFConw3CpgfBBuXD1UV52WPXgQqolLiTPehw
Hzm2BXhE2xUmPgfl683sY34NNiG2ji80x4aaBxORDcnAljy3EAkGGhlM1ovMoM060oF13q1jfoOG
yH2JJnnFZnBmz66z5zpQZUjlErTLxNsfqDbYBZMfvsOsRpnV+UckZ1z59U2YgLstEGOiYL73ph93
eb8CmFImeJCfDYdA72JMoZ84k4lYtn1ERO0/z1MOEGXZTjdS/OTj6L91XTPIqbZhUuq3p7uDsIQR
Q1cOBG1VPbrdWFWj+tXm9+Xex1cheWjIKl/NFVEsQzgknalSxAHXMWtTe4fzzjaIQThk1YYa/GjH
MFd+Q1aDqi/XyvKd5I+pw+aKJrf93nRVvhMekSFTD0jwGjLdEit0kxEl2AzEecOjBffEMSenkYgS
/HcRzKzuANhbjd5k9D7f8T0FsDr3eoioMc2Z28s4UXCAVOgOgIjIpKzAj6kpYP63iq4VVDumvHSD
3p9Rwzfgd1pAYbvEid0csmHQz4ptakNntqgz3LBiHzdnS6QHhjmfygehknL7rj5SXyfR9gv0LNzj
tXhwCzWudAfkwjjwKx6Y1BbD8koVpFk04ByTwCfpco2kDSZuppAPK46n0bL4oer3e//bBg1qKc7i
oskAstO+R0kpri2j0bTgI09orbu4lBlR4RzwJZLRNIX6QFKtvQ1mUs+Mlf3/Ja8LD6twvGX1NDAN
zAaXCOTGdUaPWrLS/mo3TZIa6jVSodDneB4g0QIkcYkMG3yatiASbSZmtO3P4uQi4Fmlc/XLSkK+
jhfJYPBM7JS75CMh3DSkdL4tyoqESbgZhYjzSkgafJKMqzANn+ulhBmk9Tzow0pwMyGQNBpCyjGZ
bSzsB8jeUUQicAnYTon+VZyPtieXWzMdFMKiZtE2YIuNvrRmPUqg/7O7yIEONl4QPFvWTBgOOI21
2LykZuZQ2PSS6QtnlMVbayIEB9UIj2fL13W82NzAfkbGEseoto/7MAUhit9AXhq8WQ3XVskPeGsL
SezcbqqTnKOW8SMMEB+ivyOUB+ZzIEJ19bzDDA2IQE4kczo2YIIt/KY8ebbb5efC83vsYJWz+ulw
mTApEuslyQ7Dnw+OmBGeBqYrOq9wvBpQlQRX5AB4mlLF8FmQZZXiFEnkfZZKcXSDhr2mPahzwVdB
7C2wWo+mDRsR3VHCHe/V3xa+IVhd3VUMyB/9l7E6HhzSh5E16ht52b0EbErkR+pwVgCFP4VKfBTl
/o8gw04q0we6FBNbEYORv1SbxPfyMP6aQne016vyAeePYDCpiidG02RFdJ1P0CxnYkcPatM/z29s
E9N2H19rorpVHPSXB4cO3PKZIqqJmpgafhVIYT6DL3zdK8UEDfVDzyHAU+Rk6MndqV8mlqQnzsnR
ZFuSYw9lE9bNc2YMtdlBXaZoJ/Vxzf2ikrRMjl6iN9YTFEKsvWVyGV1F4kS9ABF+dY7HHZ7FsC6x
gJIVrY8gwYVeFxujBe+kx0UzFQGDPhXJnUJytDZN2MOB+/cDA41NqYt4Z0mO7iFXmGYEItxCteE7
scUYfYFtqItX6JXfYkFmOj2ry79Fnf3u8B1KEoOBxzGaZlisSySWUjtW85R9QPPq5lqXsgNmeImt
VR+cRtoE8X1mLh/k7Aiz776sYh6GwaXP9CSSkM34smq5vYxM0bxdtUz4+WvB289rWw5ViqL4VW7J
M5C4sWB6JDlIuriwkavkrJRBzrf3mtasd6cKrFgRrBtZxQ63EPDJ9ReIRNQhO4wvbRrufNnXcIPK
QTC0EtC4o3VQ1X7bTDvJxeZc2QdZ01VWpOcB+AmCRzI9octDMiYoBFABFugxSCYe+zunfeZyEtop
87/8Bh8ociRIs/AVv97vmGkesfwFRE6P00RdDTV0vYBou2xxkege0az+kJQPb9TKD5UPpgi4bhz4
RKXefnLdHjmiIoshSBqiK0KdC/PtnfpRE9Y6oiSmtywfqEr8CmHtjMD2Je920R/w6J4SjMx7aZgL
rU9/cIuNVSdDO0yoXmoX2e2XPj6k8Rmrnf+mCMawO9rxt/d+BJ1F6UzxevHqt43TkLKFkXG6KZMJ
zHtrp0JthFtAumga74SkEgJfSflkNar9SkfYaU1VGk6nDY/hfBJDFTzhBrP/bGa5ILs4mKNIOlhp
gT5VtiZKG4csHK+96/F7qiJQV74fIvpP/Ithpz0Ht5aCppDttJ0XQgsgDsnO8B37sRluZwbgFM0P
62IYEHR0z+khJwlup9ApDomkcI4EoRaHce00Bk7Mwssbjt2JsGNAl9FQnMvh8WYROA6OwgZJBbU8
Db7Jbyd+Fs/7GHinxZzm0LwidKyHOfN48shzambgFXXyEvKCg3/i1dzqrBz5h2QEXpjdEubML0YZ
jXBXJtth3I5Py0uKaVEatgUqoX1PyEH+II/aI52ne0/PiHjcchLWae/mX2Uom9pqoEIRxD6xBbln
0zrXkos1jVOmcra1dxBs7FiPIxtv2EVkW5ISUoMaG5jk8zcN/MIdV43SvoYuakFcd6QaxAtkKztw
r4ef5GN7rMUGqvSZbjIy3UT2y/xObj+IkDRA2LYUPomtxyd0A8L3UqPqnmDMLPGZn9QrDz2cdm+Z
Bl2MQU0o7JTnHS7LG0ZEeSKaYuQXOyUUr4LxgXhNBp0odcRET8xS82ZhT+L03L0KsCR7JeypkdPM
yjcX5fPd9MgTH9tyzxqSdMjIDzLamL/QONedgCZQthLfTNDMyX0x5vFsAWATgfMBByfLbCrh9DuI
iTAeU8u6SIwqdtCv+05AZHmZG0VMZcT5h1XaD8UowBCfpWXaeXmyPdvMuea/Bbxwpl4UszXv7im4
w1xEpFGSl/+DX0/MJNVhnMICacVnJvOHVHOLH8q49p5M9hqtu92g3EylhhbqiM3zJdezhypR7/Oc
JHvlmKV3Cu4d1lfwQ3T07FLw9vH7KmaS9Jc9g+yo/4316yKm5wAdhOJtRj9dZ9maoX4nKasJx031
nilY901+ngRj5INz5YpvTksxj926FavDy/y8bp9LgOjxPYXJ1hBExJf9YyNiMTgpLa/RsgzJpYeE
V8uUO8CABQsfXRu6nGgj/9TDFrnzU8pkxY71FA1RtXRVr1i5scoAGSxapn5enxdtDfimYqvx2LX+
NuOrxDEQJs69CTTEnEepBunn0UJ6990BhpMVagC0Mq+yktDDtlZaXjV+6ms5eNrWNDkiKjnBWnVF
JPMUsAT2QTbIstba+XBz3r+NUDTACWmnRfhoJtWh+hAg7FkeJJIgl+AiCIf0NClosNMkPnWV5A3+
mVk1B9TwlYsGnBa1Cq6ho8OQLyxjgCDVPzjjIXQ5L9O5hClG5+gypDwJN2tMavua8VNHLdrAzGZq
Kwf5/jaXzuLKqRaaCfQ3KTAmKyIO4e+M+vHdH/0fCewH2DS8VEpJ4cq0xZ486QHKV9s5OzkdhJdC
tvkjcY9G5+FyEFMUbVs1EwV9oELsKJ27RL7gea23TKX8Tc/yn+jv3w2FlIR83AK7XWhBld2/+5va
sNIakOgmRddWwySlSMZAXd+/S+xZw2TiJ27v43aiDPEzVV5ZwVgau3/Oiw9zEV+A312LePtJfWEI
ylZ7bZZguXI3gNw0g+ByYdSQKrHuNtRDvqdD1EtQ5SBQzBfO6LTkzj2JvehGxyb4HmVd6Tg12l0b
8IjZzS+SEe9FBvJMtGtJzmtTuMDNZp4gQSKy5FxTKlREzqUiQ+bPEzSoNoA7ky3Gr0S2i8CzxOn5
mJhl4S0FeUmBTVLE+LNCpSZp2PcDn3pDZWGHdF1c9wLibxrD29UdjGlfbyDQSnAJy0TBkgYYDJVq
3L/fvbPs0mm/24g8HPUqv6yx9lVuiqLTr+Uo1BZCjdReT41u4huHs7xqE4ZJH2Y3vorL6oHWiCVs
AKHp1xcZn/7Q3JCzDWeo3PPmCZc5GJHlYP9EL4X4iY0d7QB+kYWz7hVWqvFyNtV78MQbovXg9kkv
yv9jVxgLXqI09lBj/n37L11ARYQrjiBBAYi84uTGolObrDfkPtSjBtqJ1BcM6C6StWFK+DSJyzKV
Z0FRviFpq9ABeEaRbIB/35xsuHXlQpku4SxbOrtuVBSgPytkfw1wnUEFVsspYBfIYBwnE6MkXh6e
IdPlt6NyjDMC63CS3FBvHij0GYrvk2N/kx37EYZCKDK4qPSCS5tHm3uVp+7rlaQTAsfB6VRlycVd
A9WaHArc5AtcvG3tIwGf1RQzcEu4tCc3GTjkcJco5t9vCp4yBW9MB4OEqxREwUX1vbBM1jiQSiM2
SywE4jC5G3Ju/xsgOVDfTT9uozYto5B4Rdi9xJYuNFoP4cIKoSBYsWA6xWyq96WNTiwM7EgjhX9b
a1QXCYbOdtOT9iiLeThMoFVGsMh0GorZTTix1w4ffzGxAhG87KGjR/CCpvCJ0sFbOJw9dE9z/Bc9
tTb911+dk5zB4qhB/Pahnm2PLfaoz/XBgmxsW+3CF7uSxsKftADoNNTeI3p6i0TNfCgPiUV8Iumy
29OFYCzfjRNc5vCFKLSGGG0N+a1s57nhwwn86zN8y+YPO3ewFF4o2FUtM5CaxMJW2vqs5NThGGnQ
JBfSeUw9IKReXyLdZX50u4uuFghdlIva5tQb6yNrKD77iq4YyksVzxTs7FyGar859gu/AMC7VEb7
wm1YAHmZXL2ZLMqDLEs29fvAGxJZpieqf11Ag9PjU8suRjtiYU9KDoFdAV7WRX27eNEOcJ7Hs6OG
y2RjQd6owrvtXAaVLEze688GRxvJfUw9JIxSA0dEjiU74Nb0+ErjFSYa4Hs8wq7RTmDoqLFRpKeR
IGy0uRNP4fSPlQID1QXf19GFRbbMTvb1aWJnhk/GUwoTeYq1KIyv0c/oIqVni93H7PA+i8Atowzu
pBo+aA/4+HAKqJ3DulS3K3i0jwvGbi+wCnsb0cAf/p/lmv39IkYhTmTSMzGG4WNMkek0n1/bs+mE
QxmG7IQLgUH6uGY3veidd5Th9hoMzxZiq0elb5uvzlC8KV0n7Im7Vx/DIfGSqbcqRDr6YFlu0/x2
/W7qfRF9JU2ZgGgjshdfXq2JMGQ2yN2WLoFaUmJAlp6VIn2GOUqx4vZME0Pn839abeuPVrPvyAeB
MrYgcEdrLoz6PGZeN4RvRWozh3xQu34eICSPOpcvFhNIzcEInZp/ELty666Ay3JwmStN/PjscJ9I
H28miXx3F+/c/NtHLGzrKIGUT6vpj1a+XM6iTrw5UCcZ25eteJef1PBF8ZdTU3iIXdJHBfSCAakm
7eEx026/knNRJhRwVdIGHH+OvOBsta8RVd9d1JhgKJI7isD+g1yKPTO7WekBUlXr4cbbVlMR9buE
LxGTbqPeaN1XSdAEoy9jFLPx7XoSBaCs9Ei/FSrR9Zawx9DOnoUeZEQKDhzhXooOE1m5VWjJz8D0
Sie81uoELShVZ3PKNYPFVne1yDXSJv55PDW08bC5T2sxV1s0vUB3e1je/JVgUzyuL9yYZ/0wDB1M
UoCbSfCvFzPJGTUgN/JEvZoGyMCSBtf9g/jRh03CPFBISXedXdgzmj/0PYJlC9w2BAxOoVXD4naa
G8b++Ter8g0tLFxQtD6/3PRwCbcXYTiy3ZvKxtmstfDAyLq2Mva4NIqOZGPbqU2w1YZ5rBXZ1ttQ
eEG5UxeumyQ63qrEhHH7xoWCDfnWQKIhk8QF9THjNvOJV6q6waNlMPMW+6jJamjZ17dbZDGzy40+
Ha8WvJQdSryiqWMRd4TSOXb9t1hDPIufj3Nxk6Fv0dLkAwf7zW/eu8kDVkcpAsPlTHItwVch9s5d
QAKQeW/ehc90e5HBgZiVVcK6KvM4IJ11tneCDcsoEUZK35hkKmChNIiRnvk2sgHMz9MTsM5g2BRB
789h7qPE84hx7vR+pNoGLvpRoW++sSmSvKcO7j5jCOePzdFmDTDwnJSlIEJAAsRkcpWRr4987pHV
MxYQhAK5Z4O4fs+KkP8EOQHHi4WP3Aa4pmS7k1tlDsU93ZqtfwmXZCCd2cEuM4hgVAUu7yHXZFVe
ERs9GxlBoGaStvaJzNb5gAFfG3KxYp4Ixnqcyg8Ciho/Z9usWYNd+vA4YN7OlKoWTEGN89bCt5g+
6voiKIj9OYuCc/0eVqKTn10mPIxh1p0dRSk3pyeb/HcabZy7RKEHtzIeO1ShrE4YA8xxxqjX4Rlo
fNKJisa+9G7xGBA5eztO6nZHl9yqZxoEdl+8sijsJ8lbygezd1P9hGd64njO0yNA/IXBkYAhH99S
C+Tt48s9EnR+PsbpIto0CcTB1P4Grs5Bvkg8Iu8k0526mg/mXTAbLOL0QpTeDXgf0uvCx1SzM1UI
gRALD97uoTxClrEjsblqd8yJ/vluBorpSwlavTRgY6NODgpWDypaZ10D64ID5DxLsQAH7JpWKuBs
BZ+05FPJGRBSXtEGC0RYSnTgH/jhw5cFgQLi6eVMUXHWpqaBBXBfy+dWhvWaCrQEUwRFLXCtUfQT
t3RXiFDctY4h2XWIzm8n/75TP1iwiu9V7v70+p3HFA/bN7evIAmTxKwiJu8ir3am7pRr41punNjT
T0EW8vsdLQS8DCc8JaVdRXuYpG/ly+01AcvGwbqkj471I8+fHbGlAwr6spX0KidYSfd9GOoHsCYg
yvgixMZ7f5lO1CJGvYWj+5k1s9YA4lkD9JA+etGyWoNVBeI0AI0vC6ZxPEV5XDNUadO6V8GYFW6y
h4n4b0TZaYygf++CgA5XFb6mwVhAv6aQOFXvfDZ6lmCn7xnYZHnaubD3lXdgQQscESqS48dfiq5m
HhVR7K/Xv1MUJs7fNxL85gMlvOJdH5eLNVQLqLhq8Xd3iuKKWSIC+7nOhEcg8sgMZSQVdnpw6sOx
+1hqpylO9AzGm2wFYNakcQpJPqqJVcFmeYGu+dA0G75FToLFdhkv5DC1Dbs7ooBaqzgP72qumZTm
mmSH+yXJTgXRQw7KUMAeqTC2gjRulUtlKbxvbCeaWmbHRQyPXh0d0RFnCPc+w4nir0JMP9XaAcx/
IPOZeZJGxfGCvsOGuwwl2Y+kC+ubMejAwroUb80alHBJ86DKBgq9OvOV4tJPGNmgIXg0X+fdCQJb
ZDlg8f7VQ9hqLxir9WC/V2MSSe7B/+FLpF4+6DNabp4Q0rclECmI4VCpZYZ1WWJ0qceCIPzzRUAW
5aoufr1/6OftH7cWXhsUcXTDnq+61qv6CdiLSW1JGidlJj9gynB7sDr6HNkqmLk4S0+HMC/7H+Sm
07AKixJ1CGFdrJtP7MIn+dfSpeNiDDmTJsqoJDDJhmd+Hx+jeNr1/7EkH5KUf4NMjuwk/GKG9Fb4
1M8adazq1v3GJZfk610TkrOrKtZVBnMvdNVNqyRmWEh+6dykjYctzjYgZArGZTwdyZ8RIrwt4c3n
g3Fda/ODUgQmU/l7KS1zopGLM9Izw7kGElOug7C4lfbeP1eMD9sNkgMlfDdHs/OE2X/ne+lQm6rF
vpFF7C8SxpUkDZqvcMHON+3U0XZo/E5uOdNzSxRI1k5PjWD7u3cHnrQVko6KBkHvmYUrqe8JREye
tf/mR2nYwq2BQIelOzk/TV3BPVXJy/mVJ5CkiIrtCXLawE9llu1ltj28HBJUk1/YyX9UgxR0Yfcb
hEP2RT86IFamfokOr2pkOnT6wf9wvcNDjkqBzSsWSdGhYDXigl+knlJ5oM3r9xEyJLHJseWvaHO9
Wwb8M8+yGiQBBtubo0w8P37/Iz7MUMZR2zNqJqyE5u65bb2vXzIfGwvHm8t4+E+yWlc8m5jCkTBa
vWMl2lApC1K29CHl2VpNiLTRNSo/MZTYfibDY1eqTt4ucTL0s9kTX3X0WeX1kSscL601iGcPuJ5/
iIv1wiqcISgEC1oME4HcHGEviZmjiyXsdzZHVrFfw41X+4IOY7TU8yOT25h94tg616foawSQSOSV
d+TTdYXatvbU8n8yOwnpAmMjpN2wi1OAcp/iHqAT9B0SPm2JqeJr5i3ltJtD21Z0tfIg4wzwLW1w
b8fuXGAN2VgNRs8255jHlwV6ZYFsITY3tZ6VqD8j/wZ1KVh5o5Mr3moKSsBksgGodB5DMZ4INypB
Dwl7PIyonwczhGmKK3GLR4o/g5vKaJkgAV5dWImuaen3WgseT66I4pa6bSOhaavwoYwY3XjfMayS
7FaWTfQ2PDcGBfZqgRmjPYiph69ohdh2jOtgAFm+U3UksLUo8s0EIvqI75rZsQ91hqK9SyQzAYv0
V30PS1IksTj6weOp9qZjWNeiV2/+JAOeL3Tg62orXgM2QJRhuv5acPhFN1a7flEx4I72+8BPKikd
CPOaT8C+sNyxHTjvU9D8bBdCptERZgqx9tW4T+13ZM0b5UdDacUsJnomxwV/45J6EMmHBMzSHLWc
Mb5nZc/QLLG/UApb/dDy6hpRtfmS7XI3WC/1lqxNKxc7+EkVS9OaogqJgqGaiftVODbcd5k+Nyz2
plb8oxPsEHu0EWfNtH/elA+w+AaVkgl0sf/ktEvPLExM6ZH51pxeod3dz+aplYmucsh8RZQDcqTw
etT5I55qBPOyuqvB4cfcXGOskbI0ORS3ObkIR+y1T2gSKSxSOAd4WU8t2kZ56J59xuLpRtKDNCEB
10IEDcJ5fjaj8ktSmTDd4b5UOVjShX3TAnTarueIJImMfWvNDmWLxN6BlVXfc/Pf3enIbrHbDK5m
WaQpcjgZDZaQfTUrJmNFYcYLXGARFeZ2BVuJYt1Xqr5u46PwiD8/NspXweKqzWP5CgUDNogemqXP
VwPp+8UOSX0mX8ZBhmh9gGN+KLdX4OIeGS14ebzs+1h6yk0oWm3WUJYSZcUy9hhBRFmiquLWPJPZ
grU8560I/MKmtKhm8/713lHk4wY770NhtbcjNN3iScr1b8FMCUg9iwrIaplxC2Yka98T8oB8a7Tm
7NohwgKIbHIOoO2NHAnDlnkpLJxsyi4XhgM/znh8Q8kIz0kRidGxQn4Gv+0VzFUbk/k3sjuHGHYT
6UArJZwEqLDsCclqRUfrfOCj8dgKr2qWQL7EIY2mSMIRw1E11Dva51H6Yfb8lblvEv7eA94eT8go
P54zPc8CsQrFF+En1gmzJ0/1hKo+LrqfO5MWc4DOXuNBKrVNNTNPrv4uUDis1pFsbAw90P6gYKYE
X5dBlpssKDe1M+LR1I9EBOk+xg6KcNOV6Y8yUHXllTB4IEAoLphi5GLt1v6nzH1E0AAshYfH66H/
3IeCAy6lkstAUxSw+76jLHBvEOC6TpUw34RfSd58Up9HHvI3XPC6Qrm+dlifAaQejRqYPBF2LxGy
ZjzZjk6+n/MKGI7cySnmFOYfCs5/88wKjDr2/RKurxmXRhGOG22O9tRB2GWUzzVuHelVe2cljfWD
Me2iixaoiWERdHGrPozfUs+OpI1+4jsLMHXdc3m7ASKiOtQtcyO3vDEtO74+BwQOgizCSVV6NDbu
Vtmb/X+W0j0Hc1sweqF/Jqe9TyFglDmFMn6tv8rySjrr3qtwlIJeruzP056K50j8TUedpzhhUxrE
Ip8yrlfwDheXR4MsBqd4TeU/2erC+u/TgLWCln/ApNrZJ/vgPFx2Dr8VUK+H9mEbwYU3FkMXSXsQ
YYSo72/W6IPYozn0/05ww6eVqLkqksfDkLXM+Rq8NkG6cQsDwdLqiUk1rbjCMTheSX05d+B/Ikl8
AifVee+RYrbod4VCcBCce+cLUL8y7+toNGqRe/7vONkFyhRkZeTIliu0KOYyQAp56Okv9hay7hId
iOkE4uFQzgQ5HWyyMkaXyOPf+HYS0OuGbs6/FmgRdcmRlPND+CxI7g7P/ORtFCkQclzv+M18jcbt
Oc977yFykyOkoiXE8ZVXQN5x6E7O0DgGuDXBO1VBySKQPEh52kEo1Bp6VrZtjXj3bKNS+jGE0Jc3
yGcCO5ME9pGycUdUyhOYJ0cDHRouVKAnYAkMVpgG1DGUuO1eVkftcj6EjMJpDIZSjLAeRkMMne3f
G+FA+wsCygSa+ZaVqN/O+lcgkkdv5SvgM7BbBDbpmWGGZ0tSC7XnADtJ4Oi7ONNyqj0f7p92gJ8u
PwMa67h7gQMGetQFTe6+QSmKM/ot2O2MgdnYKPOHNIcjQW7gvYrrUT8QTi6ICjh+QvsCa/lj30rC
CE0UaaPSIdUssGD4b2PdAnapTluPlGC0d1A5M4Jp8VTo/1K9noyYZRlFvxHhtK1WZkeN3rqtXSBt
JQcd/6QmKHU+R/QkhFIdDcXnzM3azEZsngwsygfzygKoyqZda+Tjp0kgGHKpx4HC+nqOTn2XrTWo
TYzk6rBZOK1R7X7+dWAEA1okcuaRRqSCBMx7+TjrP2bXUs3k3TaOrZxLAyCI7tFVIsDTu+KhLHIl
h1otO+JoWg5teKuld7YDRd44r0xe1GHhCOt72r1I3Mf67ktMj/jqXctJkEQ2O8n0/cF7jdJy32I8
YNaBizBXO3ZAtq0QE1rtUaQAz9pOxPIXIMG6q0IjW1TRjvs5Cjtfm3NpL+0rYCT+t9Um5WFyUfe/
qw671JRg2WPGFtfPqwzyh3RUKdgdFldDgFQZMm6MQcjZ9PQcKSmRkzcvCEUUdldCx3P/csn8nUv2
qtXHh/jLwPhl+zVmEDd0hLA3zy2m9BLVuWc0bufUtsMvk1t4xo1qQYw9F8eLetg7+qVL+qIxkrbp
I6CFPyqHCfWO0jtYaX71OI1wYSZRC8bWLPpeatSOUTVVFhOoT7GvRSgCLkCZIKC/6HfGQmdN15Ag
ct1hYPVZD50AG4mk2P7r9z02gOo2bCg/Do7RdlyA8i8lyyoXSCanShCPYv6Q67bZxZL6BrnfK4L3
gQVPj3LRpXrp3LjUd08agYsLCi43vQ+PJ/eiApNQnc4kaFgNiXTfoyLsavt5obYOYeWeihJ+fhpq
nm9IT9by6PMwQCNlPT45/WCtNYXKXVxnAQ8qHqkVH+cFupY/66hzjx0hy2O2EnmAiiYnqAcgb2nR
VTb300VV1vnR1NRXilTl8u5Cih/IvefnsRhY31RTyCJjTuzEOzzBhTrp5ethtypLiIJK3TL641fz
T7QCFw1rMfZTWBnHQKzL4FbWvGpMn+Cjylguu0joAuafNzaQrzB6YyKDyG44CApK5XmKy/ie6UVU
ZUXM9DJBXubQzyRhQ6mK8pWS+Ifc0WS4llbycLZfgdGesSdWAQ4Swnl3DDtQDf/3VJiY9Jha4eB6
y7HMNEKuWZpcuS3Uf6DImLkmBpHNa2Fvg2nO6oj53b4cxzof4psv8Qkvlr6Hrq6EifE3uC3fUB+m
id5m4yQIRCYeKYcp71srJP6gICH5o08D0Tqvih9gymDzlz+ejjVUMqOGR91d2nj9LU+8mQOGB0bj
tNySLqVOTv8oU+ykhLlkAbxSsUPyWBNTBs+BPjH7OmdleEb8WRlZ8vuYe2LeZTRCB/Bt85wKoaVO
PA5rN8qlRXzANgcyGpI+ycAFCHayU+hYobSG4+Pu1z10jc9Fza+23yEOg/P0qGEKowekMYudv/re
Vu9FCLTu/zhMXdlwPqCl1j2+xgi4fU+Xxp7rIUFk8w6a5lC6R9LqHlHctawNc2+p5t5zSiWVvEA2
DZKr09hl3P6yFWJgwOXZN7VOguUuZ9CRlPt+Yd+ce3gBzD7vrktAgqZVRfVzoqMTLk4CE1AhgJyG
z+1Df35WjMvIs44j1hunBIucU9KWRz1RBmHyjsYbyukyui9sI41iZT2dzpV6mGvNX0m2y49POgB/
i8FSWAK4gA+RlnagOKv21/U2YDS063+pPEMTvQe2wfVUsndVQkRwvkDMZpp5rWZHPR/CLkJQDKJr
bc/jw2ItpnL/JGb9mXJKlhcgd282hDZK1zGyfcRWnfyXEJ2xMKLyyet38quMmLW7VhDMYFJzHpeX
YYQ6ZjrAMV/yd9g3uy/qL/jXze1F0WcBzHIHSHRSrN0Uxjfe7x1Ls5QidG1UPTvDLaMih4AeXkEL
/yeAmDTkEs+kHvFkL6gO/b0Q8tdKhE8uaPUL3SPL0ff3iDPXSz09A0IJJCAUw+mysZaQGxQNTOM/
27dpjP/j1KS0vQKqSbWAyO2I67yePoaDl38OBiOivAZLmsnllfj0GfN0caDEpWqWua2t6u0CcKVY
S+rATwqEYPWav2XKvG78R2NYyfhhVMadHlEptf2oxaG/SQtPd9JUuraZxPqvU5jDc+LmT7uQjF7p
b0SokMGLuv1XYzWPeMQZPMkAevlBIzwrslPURDOKkSIYM4GlXKbFZsOya14TURGJ4NtiEMg2r6cg
rlLYLjk+sbdId/10ekUSBwnDMfGSKEu2i986P5mwo8VgdusdN+dwYsw1vcvYwSjjlwXPKQ8qmsws
aYBsEovHFr56iUl9wYYqM+vszCk+gQ0QZ7vYH+ZSTqaqxvSY6rY4XAc/yeY0UWbhOj3EkIC4zTeK
wkHqf53Pp9vPgti8hWbeV8yGAo20Bo6/2RqEdUSuzmhwK9d6t6YmTBzejF1fGAmw/Z2jyKN/B7lG
iovZdhAhfqednrFLbhMnXRaQW2l5HuR9WMhqlqzP+RarBv0C2iU6mZbn8OuKnPN8EVvkyj6wZ25x
2kvLqTIGAJtISK1rdQ2tSP8o1hLrvOfznivZoIkao0MquMEjLeyk89cdQyAd51LoxocGSVVl+FEY
ehkjP4E2phk9Y+txEcSqzCzPuI66wzALAYfjTl14Tkx4KhGvjMK8hZKAzqYdfHscQ6U7pvp0cUIu
wNnH0MYNoSYZyEIld1Cpqix5z7t9xJUNjco160FIqcuKf544a2dZwkULI3ZqKiP863rS4HMHC5SX
QidomJpX64z9HQFb94bPZft/OeabAddEfRpjbTnXhcqfxHf136H3Vo3JxjmcxxNmfx+vK3Aq+20c
xneWL2Phtn3j9dsTrFVWoEdfHysb/dhqT2hhgEvh8kNc93dlnphK8fEoYREnF0OYEqpS0U+CwT85
pFQBpKMNh4vE7GO0pyFJN2oGIutHOkSgZ+8U2VMkd3hMvylFGhriEPJ8tm1XK+e0EVyHR5A65OkL
TizUcToio9edqYWVJj3AlEfXLKZlv75llayyGbnv4cP6opZDe03LkFooup+NudQ/+ckbBD7+EbbP
QCv5BLM/6d8zts6FvdblwHhHYHP/1+xZOxUW3kXAHFFz1Ho9E+ufypOswT1LSHbgMs1qlpsw9eEc
yRSqYEjGcAJRPuQJsXIs6ZG+Jw4sXK7RWFH9V9MTkMf4NupAgFfotoSyvC10RsHuiYLZJm1hBX6G
pQ8xzJXYuF5Ee0059lhM5JMxzCfW2UMxVmSJoPyJCrNEBI3HYoevtroWk92bKK9g91qZ6djJHbp6
1T9y39xptVHL/g5KbYJ0fYiFRqxp4e6tx99KdT9ZTfXjua1ez48ivFCMB++d6C0gIwhBMqwk8qVM
zZVjA4eGaeGiSefTTgtK54aHswqtt/v+dKWC8LdGdY7UYjxWllMfFZhCo1La5PORigySAEMQ3+r7
fWbtFh1+DRPlNJsF008O/vqCkB6WTnxcb+RvGNpQ/KtL0ZcP9VXDoUAm6G/wcKdNKagtyUGeY0UL
V3o7FZ7NYe+JrXJZ4GmVZP+4tyzV/h4pW0zyHHFXYUXIj0Pb7+Lf+As0pw9Ctxu6SqozA8u3X+8s
4XnayntpqAhjZDyO4aWxbHP3hwPQ48PQbufc5T6Bfi3EnSDC2fXvL8iNNDrSmVvgnKtbrwsAhgeX
3NuLImLo/tuxpNJJ7nHLDmfnT60Odz8OU1K4f5Poih90eYyjyCojP4E/phq/lnN6aBT0qDAyCWOr
3gA1Nq0m2SseYbMy3/Vzz/7XeAeGDWzTthmOqpA4epG1Z6CCV7DNhXPY/LQtUwLvBNBJEs29mUtA
y2uJlr3hCD3jqlBHKKoJkkj8QnWNel5ClL0SuuoGFXai2nKYd9Aw4k19uRt5J0O2xqdW0oJuR2Us
5+i0k8CkStJiceAjB2/KKUMHwbtZaDKfk8hSPuazbnG4W8YoLF0Q52s76s1QRlY6PKHKkNutr6Z1
+h2WWUS8pRxjFNHJbpWhpB8lHYA/XA9a3HDu66ioXT+bZp9Fmdo9ashVzcLVDRHx2+qvlZxnbqpr
LO4ta0nNf0ft7ZXiLESQVp7u16uYyKc+LwdhhDJ618KIX+IRIxN/uAfBP21tdDOhkz3fu+Ih5eK9
Ti1Q+tn81mPDoNqsMEXGLwpSsLGQwViPh+nl8so/8Szhi6U1natzygbi1x7S2jLx7qq6Vi+i+/am
APWZsrErfSCCX69Flh476xyKMVZKOzpJ3C0+Iuc30DeG9YK+Ez+ZI87tJXPpurkbhx89K0dKR//h
4bEfPxP6R2owVKEWgxLDQO9ZWbpWTfeQ1riK6gUyPMDl3mseoWzLpzljnHgjmWRDJY5jNDYI9zLR
4ZVA9g2Y3UZg2eYlSXdTRQ9ZLTGLti0hhm84i8fY4VpFHr+lIaynfWIhqX0A5nKiHoWW5fd1OYpx
RtS+lk1Shy3/PxVJCWa8PDApgTCNnamo4PBOP+a79CMNRkZ+00X65dV7XFEPF0XSNhXM/WJR2vTS
IjkSfmJT1Q4s9BP5nSplsEAhnn3AyZj7b3m7qoz0D5lMunRaa7VfWx9+0f76010ev4DvPaxBi9hu
Deqcd2E4legdn1xpAQv6ieAZUtZ4wZhzM/p60vJBDyCnTCFJAxN6oKyCiX9x9WZcIEiOyAQhr2VH
3Ym5akQBNjb/WU6cao7ObFxIhcI7DxqAG6x3Ho7sWKcqqdfTEhKIJ6JX84enimnJbPCHcSRrg941
Zp/gYPPB0O8YCEfdwBvRRtFES4Ub4bzOi9vHqQKDlrFBYTKMjzvcZgeRqIYwbmsSPRLAD1NqMCBI
brVRnomi4HqcRHOZKk2Q250qdW1Ljtut2i/OvodhSOMd0cwbE71M0TSOgE07eXM1bjPE1eMpTGuq
CGT5Be3cAeWajVxeBzWZBAYIHSCLsNEjfnYRmgUuWUUDVFnHCTMtQB6wOS1yOKVBFNnKWBxQv5I8
VjEAVjYxnROS1g+hLGr0vffRPTyItkE1bSyxfyQns9D0yxl0aO1qUVHpG8HUskCpGhv1K9h7cCx8
B+ZfOqSUi0I0WGbY/46Fgz7ZDtdQ+MmF4okkn5Skqf1zhq8Hqg5w4hPCartrnslx+4DcgmsNn+YV
PndNDq0u9+4siFyaMYEpKahDURyHtKtGHMQ7VMWL8mknvzWq9q5IagzRYp79vB2T5WORGfZsHinq
LGv4ECaHnIlMbcK1T2sqdPdkPscJa6uwRCAg2xsUaw37YUM71AVsKaZ8kVuBZbtogOy1saIU1h2q
b4BHXOo7ZM1CagucanDqSWTHfDZF/1Er01/r7bDk/pzVeyUZ0F4OB8j4grKF1X4Ue5moBKgYVp+b
H4+kWJTuqU326zUiq4yyJEmt7Jh4ZBqFP+Nfn7wyrHbILte42p/fb4zNu3+KhhS4t6x0XUk0b77V
wyiP9KOfh3Grz1m84sbGW8oL4qrPmx4JH6PjwQkybGDiDWptty44AKFxhGjAEkC2LEKQADOgUOeL
D2yhp8RvUu3PhUS08qpkBldkTYtSY323jHzyPvsY5rEAJDae1OgYw4GeFcVvZcOtOjSQGBUH0aMm
gIrMyQzvc0GrMd4hgOi6Um/KMwHyHdWgVVh6lyH++Od0+rssz6aMwH1YUpLgnW/TPSU1e2KHXgBe
sYeKYgO7g2mUBv0V8OSR06WLiO2Z1wfqZiunQ+1wJDpjnN6UrBeILcgGNV3ceGnw5KCSrEA6eR8u
SnETydDpOldCdOmtxF0YRoIajWYu7quU0IIWUBVR1hpPbr6OUVr+i3Wo++pby74UN8jDfPi5U2xb
h1NShIzchSARn2bQZruEINUQugFVL85rb6atwiH0yUBKB0FWPFoOfnArchQWh35lkhFOgkrtcRrx
WgCIQgyBSBczeMw5P5PlqhqYqdDqxc5mZm4a9Y3Am3xGDA6DHX+zpZB3kZavt9e1aW14gO7wiAf6
SJBsdWPBu/adbZK1bTxn6ta7MmztFfIXksYgKWhXc2rLRmDQCEhZc50I6L/XlScIKHyb55vrk0Po
WFTqfM7ldUW5rmm11RvgxzS0QQpxJmzn/4/YyIJBFjyY5JMO+LSAr0kOaWqrzyX4LrIUnW4Bsceu
Nr3ktj+gulbcBdMCxZJX3dVqMv9EYhSbKODyUtsgF61y6G/QLUgw5NLr0NoqgzPiCEk+H58Z5QiW
OkCKuLFtDPPvh4n87TF1dOp2bGy8AP0+CfG8bjzondNayVwyNrXkGW42+ObYL3eBv+EljMYJyleG
5zJcZBohf4INmTEx+aXFsBRKgMt1CSf6RpjeSU7ooY8oNSqn3XlzlSCBSmtVvYQiUxk3msMSPcYu
4gQyFHjclbFNYUvGJM6nBarXgdYgki5CW2A6/xX/Yty4jaCyl1NFlArihkkEHmOnTgYSXJBKzG/K
SrTirtosTjUY5IEn2TcrudzocH3tFHsQsgqjoln/zUVOyFzLmAzHjd3eg1UcVYtSAfEZVLDpclUk
ZxLJMap5iZd49LJOyMZf5U7qUMStDV59LVN0TXg9tXnwjS6hG7Wl67pXYdrL77CTY6BTexcwPFl+
bW+bxrZP7KQctBKQkqBwDrcwpzcSkzUor5ttl56b5FFajYNxv98jlRxixR1D9i+hnbSAszVxibrP
1JTpdtFxzqjaYQ4OwUTs6Zy7RinwlSxGakpS0OnICCIN6FgCLNTutZR/OJLPcqMDTErPszsTRMe7
zN2xVHvsTU5bPEKmCKu5pwMnkqRBKk1F9tHpqKvySoLgysVHCJGQeV1jHd0P9lzmn0Y/AD45I6k3
kJGkCjzSiJJ7ITCzhenzDeKBSKLj+sTlXAVS3gxDAP2VYtQCkD0jD+cL6azLLpBHKJ0vaNoFL953
lOvP7k3Wn80P8Y/orKUf1uB1Zk55tyGgID67BEg+m3wtDxCr7A7r8gdG0YEPRH9Gy4Dlfy9AfKIj
nDAs4gZ0tcDjXuC7lT7YeleNjVaKgLmb2fL2/rWiO9i/d6Sok0fxvurxfbUZqRjG49MEBepMs/NN
udkLYsAlS4jU+8Dhd17yKkatnDiQFBzmFZR7lPa0U48JzrnefhZBYRm6Ij28vzcgE544413IWvJH
2Y6r1nf18/WRHhkRCHXmZ1krg3jXCBtQBU6hp3+RsUypO5sDGQUZJx1bTkgskCy25P5dB9JzS/JU
bw1MpbrKsX+oXeDf845Ow+fm+l7Nv+9VARQgbsBBvpUUGOkwiLg408jiOvPXXVMhIyLHJHIdzJLL
OcoX+pjQR39caBP33GLzNUb1B5mg4oVGnvDp1L5fFn2mq6WesTL4GT1nogacvMKgBs0eWkGZaM7C
uxTdFsVqXIwVNRGQVrIiNG/VY8KjSmc3UsCdZHxtPyScIM+f9O+iWIocMobZ1VhZjnG/B7MsMS2V
hxKvPe63GtUYsIpkCSzPWmS5HA+CHmiDIHyMcjE9RZJNq0rdl2F2sHUHQGEE+XWsuYdIAKNSm/aM
9WGgcgtQeJ2s8edKyMHm/GZ59zsyMZmW/4mv94HYaKQoRnv46JBSsO0C17QpB+ttC+hbRMHqw12T
TrhORVwtvLa79cWDT9AImtuPLnWPWRWoi3KkILg0r6gyymLIfN9FZVnY8G4KT41fJeYsEVY+Luu+
LthNxEp0JfKLC1s+Sem8QYrrEQ13cJaeXRzbudYbl9nLnXhDM7HkwXCPpVMtOgfowoYazcc7kTYH
0vQbshkdxPv+38Bi+ysxOHAA55B9LVvzQzRb+LgrLjtuv2CQ6rSWcyVXBJMeGpUuF263ZiQAZkBc
R/5i8x+dQhzW5fZWlti+jNW+l1LHKD+0nwbs2cr7JRsFbeFuJwR09Rpw98dB0ynl9UHITs0vPxYw
Yl9pKcE2Rxr4kDUq+AvBaSyJQbfYlda7SO9J8tKqmkDeADP1RQQGwAnykDOgQKMihVTRpkr+q7in
BnQYzT80oqaAML9rGR4jFqSItkavKujnPqniLMBJKKmXwxCOwPy2k3ATxL+3eeZSnmqiE7XL7RFq
iEc+axXOiFFu5M6+iFyKy8+DeQHKBRJMUvDu7gbrxG8LEndnwyqhqSL7Nda0ueF/MZxBwe6nkuNU
2TLYCR4b58wuwbw69roYph5xd0ZKgdUotLAWJ1rlt2t56wS0pPLvYsf3H8icWMYG5zgvNaKxDsIV
I0M7dgAHLvAzs6EvhgxewZiBCy3k66/vyiSOJJUOTYZdj6NXNJ/8uliKBXPq1NT0AtWX14tfak9X
Ll326HKDoQabjHIkEXigDxQnoc0P21gKVqutEsd0HKRI13+6D1nSrabcD6Rq4ePRkvjvnXxWnLEY
1Lte5GbQ5nUud55K+oxzEKCRyoEWY6k8GBoHb+rmk/q8PW/NgH/uyooOIBqHBN6ln4Cqyrh5aQNj
LJPzxpBOcsVoqwVs7KYyztnCfVCcGkwUcd8/0owdjEr4KvL6NyZOT5rDnXNZM7oUQ6RB5ZZDAFDH
e4ed8SPdp51k7EQvxd8AKXdpBHF2fTSFXmS6YTijoKmjKXqpzRtJNegEDyYlom8RmmDZSxT2Yu10
WVHXC0LWg3nwOLo5xQVJMhp8/KTKWFMZdarHabOo042zl5hUdQ8qN6lVyGYM2dQm40zU0HLPmlEf
78e+zqk6jWqPk6kQLhmathLpcJI+Rp48OKMQo8LLj07Vk4hKuI3PqUyP9Cm9gYnK1xcnyK2PY1L+
RL5ebiXg1EAdU6ZtE++tqAEznVMuVdCPWgUxwKYUAMkCnNFu0LDYhk6APnXTTyyDhCarrIPyGYE4
ktvQxljZ0MuJUzeab0SteWwzCO8Nr4CTd7mzWwM20emkQHrnc8/BsJVAssOj33S6N5R7Kh72pjyv
mOEAK23K08doahoiiIte3EqZKU9xnQ+TsKylH96R2uJw8M7Ed4oLEi3PYwdV9lkQMe5G+gmDMu5I
67hmPXAiq82bD7lpLCEIGIQY+b58ZYtDrZUM9UCUio4EhUCzU6dxoFy3qDENfMzfHruTgfErgpGB
dlkeSFZX4mIEWB9LYKoUpfKIucRoaLdxEPl1qPMMnOr+4aRfr/63gxGWKU+2/tjk6h4QJGV+/ZZ2
WBco+DlHYIarD9CDt16qZ8rw41VeUUlCrOVpNXZv+/+6k1cioc+oyJGRAM0hdBQRAfMIiRLiEoow
G3gXoIesClmDs3RHOpohUdYAYg7bmWwrOlQHUWJlLWc8OniAjJfNzJ5ittxT09ieo1IscdNbSVad
kt3MJsuAyg24dK/iceKXiSWG+52yCigQZYbUmUGJ8cbSOB5BB3K5MgoUikQkHRGN9Gj75PM3EJCQ
+sITisk1ZqM9guvuGnL+J1rfs4Jc1bnCcQEyieAp82WxZK5i7H6p2KHCzmdg7W9+Ff9EhEjkDu3V
Y1ZRAaGepc0gwcs8j3GEUPcPDU/uMS/NvoHt4/k2KMooA55lt3bYuQcWzEM4xVdfsRuvsTbp3S2+
K5EJWMtpf1wcixaGqh8psQXdtDPdMJWSEgCzzclY3eoRgnwXvLbTGyIKxDS1p8nVABRX3em6v9Ht
5Lx7JB+KNTR2tY2hRkzkBvE+xhr3KuZZe9rvJ5hbFpNybFZBJkPqWv5UCkn1PDif80aF+LUgaKCJ
tRdLXz+aipgUK5pxeBKN/1nBdIen3PfFaLFI6A/VoSFoYSVUHyvBnzCsS7M4TAc0RSmwewhfbwgH
0EX/j9PRoE03+4gzkEUqUehZraoAL1BL/X6NnSSYIDqBbiG8494WO+B+Jdf4vOnlJBhqQHlWTpwh
nbtH2JoWz2SXk2jpwDvcwhtYT/ie4RMo+RmOubX6Y1AYdtanX1OnVAhz7ih7qSitkQfmlRXkMukm
8ZUuPqjEr7/u1TTd5ObOuZTjf5ptNK9eg+lR1bS8jdnD29hnLDVeQ0+Rili043x3jItUTRN9UlQT
T9m8kiBz3/MgtIL+dlPenT04yvKFv5f14Iab7HluRrXP9T9XagYdinXxIycJe7Z/zUpoTSGiVtvN
aaMTct4v3tBZqq7pfgPIzpi6gcm5CsPZiAVqp9d3eHzyFz6OunJicdvFnOb3Moyr4y8xAxNReFeR
sY/2Ho34t203/6S+KbO1wiirdk6ZV8ySYG/gFDgSu+E4QhCjZYd2pF8Kii5DOE9nmagtSk1vVNX5
azO5uS3RxGqSKULOrLeJRn+uLIca3kgXATcf58VPS3d7VtCvRXXA7FdmWEBZ7HyToe5jaCQW04pF
g1Or+BYlknFzbaX1Y/vDhQqMvomFXOpO1/tCfYLTx0OqR/VoHC3zpoFCne5f8RNLZL2NyzqVT44q
hlxTRK31IzNtRYTO8zzBlojTI6N5UPqMg/sDWYT8RP8K69gfsI1SExrLP45Wc0HxBTQhTf4M/P2r
WRHA5Jg9ljuiAdp5nHBa4qjpejkV+LY1tOhJE1gseHudV0XSf+1WEcO7Au3UswtoT4RyQ8KM368h
VzfxW7rBRRwlIOJOCNKCvSczcUTyDk1id9YbtfrT4zRNWc4Lru9atsMhADOJhxM+ngxOalWowPgZ
UrnomrHYArJvd+H9CIdvlvqzHff2QRTJSDqfO9T+XQNZCHRfdSVT6SikKN84nt+nzLwHwcnpq7nF
nlFH0AbgTUmk2b7z+NndcHJLP1YvO700oNQ8S+INzay9qWyx97amZFj1mDbTuN0m47y7p6p2hrvP
g75RIsECvDTdShfzRbNtgzvtGghyubbOwUEW9Bk9mNBCcJ2GpP9epaqYwh4JCRiTz1XY63LMGAQp
vVe0Z7DkJYGVRxttpGTq8gjcIoMnhFF4h4cUcPvKmCGfyjZRmuBT8LNLeTAbab2BN0w1GPdYDgVf
/WFsbp5T2BJD4vCE2xNMinLPiBWABWRl16nyfn9Lql6Att9leYtL/qR7RdZzPvfRQCPFSmAs9VjT
1NjcoOEqtgCNStVUNMiLh4rSb/a77L3rYypjR8u20Lp5gcDbKf0f97meH8O3mIBtlWBTOTCDE37A
n7vIj99mifEoFrDjcE+94qr604NNDvC/UZ4RdZTxPq4GgyrwJ7mY62Yfo3JLklStJgq9I3U3NrtY
URSp6c1u1AtL5dPcT6c48K7lP0EuL9gIG7x0/ouHhUYjsbyuMt0jzapmh9XNhkxo52fvcSrzc5sh
eBZJi8QrIsdD96diVWrp4ctMwV1/oHHzSFVjp7khORM3A+KTLw9oEuEi4Xc8S/6UPkED8Atw+7NM
/l2Tsbuqjk8LtXznk9jttCJRnt+vm9/QSZxZmHV5UufKJuXAdhlJsY2iSe2M5eOvd8D/PQ4qdvgH
RK0UIjvdm5ZWwy7oPcJr3bKRJe7Kd2T0hNY/sqr60W5ag19F1nZ6k1tyNgmmyVh5lx5lY7V5xfeF
e6HFuBju29+o1FYTnF9+U4nzlc9AI2XpGrdcu9pTnoeuKXuOIccMpQhvDUVdiFfo844jXqfY+ayz
b637vRFt4zWw3vMLj3BWCGCw6H0gDBemhDOD+NyI/NByZxRmfmYPNJrTPJq/VgVqtl+mOhmNTzMX
S4RB39AxE4mMh6EuravJIm/2xyNa9oCwmkxKWnIYkUs6YvQf/HRO587zjp1ZNyRlZEJXnzgOm1x1
caa2KwG9IN7J3JPSy3tdJA0OAqwq+VySt/Sbg97NsUvorG+eA7alsb/w5gjACwU+eW0wnSQtEbOl
w1/qlRd6gamx2PxQuqwFrd/B37wFtXQsqgf8Z7FS2nqANKVoUDoYHa6JP5a6SgDXMdCmLRMqFGgJ
TZEDgzPSl4Y86d3L9kyUTEQ1mVoFb9MpJYUXjmjWMfq+/MzFabXwW0gl0HYy/mWV6l3KwkQhU/sb
ow1DdvxxqI0XpsRG7eouIHG2w02/YTN9hEkHn5p0ZaxYc42Gx1kYQFb3E90nw22fncNowIfBIiuJ
p6N7Nlz4zLJDZtpevWp+93bp9okSRfEyzZ3yci1MUEeV50qvPsV0Vyj98WyNZh0JyFCm6ouu9IbO
ld8rToISsGfA3E86T9a7+ngeZn4JODUZmfUzUxyciM4V+tkrOzkwlvHX+qsAB6hDHgkmj0aRPJZX
Dy1PVj4adIhtXTCTLiHo5LVvq8H4C75ZkWqeJ21rV/E3TlZEdeGzIQ6erLZtYCN3ktfDU7JzvJMj
xiEbwoA7iHUqiGww+1zCsE37xGJ4bCEqG4iwZLIwXnBjmvPKmRGQTqkFLFPXhxtPW4UND7kjBC9h
RBVuksx1lIfPro1IXyC2lFtg87v5Jm2u4oW3ZNuJ4TdGy0/QQqUokbIFLM11XSCpyN9FbWwBrFu3
xQQSpz89zirSzF7QBmOFjMZfVHaqztumgyxC1qb0XN2BscqJBdVb5BuCFc4jG56JoZntQVvi05sB
bbE72LcxP6jKwTk9m6EugCLZB41Oo61P3sbLFMYttxyepp95ssgBggK+gu+3aApZqcq3dy0jSrga
yJuLrey95qgM/Dc/l7DI4eRxhPJxqzoHkrrwGjOrdVQJ5sha1oWSPkHpzjhlGApc858acEXOobJH
KkBHKwOX+ZAPxYc4l2mzefLTlP/d+4GKVFeW/l/pZlrUE/k22u+2mVCL5b72B1ylj/22NTN8osG7
u8sdjc5UKrpYHaGeqfbh3UVOdz7F7yIZdU6+tiOYfIs+saSjySyAE3EmPRzJj33sr3eXgv7aXi/u
tOXEbrULkBZ7+aWRjteOKZF3D/PjArKQIJdOoNjJx5DJyUyhg60Af09S3xoTl87Vl6Q92Bw7GlhN
i6inAV4iztM7ZiOSsgNav/Hbz4b9YLGDNFifn3LqixUF+dlJBe3wREEA8Ry+Ps6jVpyIo1gqUW5b
mXmCCLwAbjLnc/sBjFSbq7xuojY+Yj0IKm8sZa/dgaltao4N2MjRX9elVSHKLiLKz37ajpD2VlFk
COnbn5x7ivJ+BCQ92xVokU+vSStd5Qff5G51LFvF06w2mxWtdwB3CvYTc0rLJwKulj+LmNPqTyjK
Ts3FIYSMfu0NwJddpHTlK7QewXp6o1xqOjHehn7ldw9jMmbl+c6sUdX6ikkuubfff+UwmJGv/6P4
wnzzUd6I/9Gv2LGzddk+3WI5cGXrw0oIxQc/mAEjcTd0D3bc9Rd5wFZKUtYPq6RZErfpID6kZIrp
DKqBKZRD9ywomCw6F52BKsBRY1EXRoog466v6VZn7NhtIfTZNHyipVxIQQlOL3tT01FnCRG1CI/K
M+DR6w/CPqloojraEwwGPZCnKYAnWSQlZgRyJj79H3ExNPHhXU7OhuJ12ZgO2+dRwxh8wg4h/dPO
+SpVjNTE08eW5tkJt85tOwqoEsyfbJohL1K6fSnDQLhLZ+fI3Dhp0ORoJog7MrVGL8RbBFBLYzFa
gG2StOKNxL1HhpdFh3uIdnsGVBKpQ/9AICMurQcy/mVTLskM2mYDhGl1qtuGLJ9vLerBY2ouTVBn
i2NPpVBcJKOt0AFbsbHuX+1xKfzF0GXZ2qk8rCVXn5i3TmQzg6+NDLqyVmtVz7MYzTSFGWUUE3+f
USXtArbV3Vv5i352ASz1WWm/J7j8zp4IfWj2pbe1x6NbBuHRo2OymvC0Hpp6GurppN1wNk/WgPIJ
yvGOUCS4D6P03z91AuCqHt/mVzAvieGQIRhGG1ThkBJZ9oHKkzsNO75Rsbs5ZrS2SILpGd1Q9igC
dHJJgcNxArOg1+ItmE5qOharJ3b7sANUyWQjmjNtP2vpmVYN66pjdkmrEv6BlJEo4zp1SzytWPnA
wGe5I0sv7MFGDwhpCMmUVDEEzXCgb9tcb1FVVD6xZcKsThPEmLFBmTf8Zjk88f0per5EkW+KIPx1
g7/taNLtnPRMOhWxhYUn5B7hSXfVUXBkNWrIRWSPpy8NyrOZRpx5gEItIn0vx5eZfXQxKOjWecN0
JUnjAHWn6gIOgFBlpaDwIjijr/hKlLAWsjyrvt8aKho3XbHB8vOTsRzNQpnqjmkFQvlOiAIa4I5d
gYWlUdL4QiNzAB/ftKBempn9C4LTacc/VjHY5RaqkyVaM6E1yLW0J2wcxKgduf1zCT/b75hF4QBf
rSIvhmne4+oen+YzMDLhP3Vbpeqo+4BolyePMEBtiKWBExfFzt0qr0Kk2nbgStglBChKfpK6aqfu
QaxuwJSVdKK5R1Z4H1ekn3xY8U7qNmzeZhNzCSGXA8oy66XCwBYg6HcAIuP1L0z4EiTb+DLsMQ8J
HSN+m4PKok64srEl7uAbTpgo3t5Q9Nz8lQIBOPi4L2U41zUehatXw178DRMVzHGFyv26qaQg7qbp
rICtPfmY5+SDEWTVM7HXss3UAHK5KP8ZRj4mOgynS8JvwX4OD2o0NbbcCt+pSGLwFa6Y7+5xDa9J
0pcIpD4jvgR2utUn4hMQhMrg3uT1TZH0/3Qw/Ai+WgxSS0q145eU8O5tmlBrKxv87u+/Za/O9Vpn
1qfZZwlIjWPixmNURR2lThMjfbjdXdv90TatxLMMV/5hR7WO3qRJMM1d1B992CEO8gqPeepWWCqE
gZQgc74E7gALs88fEOcOlcXH8B5eIs+igeW3w3v54TCDGPiAF3rG4uN4UW8K93fRJbvWZgzQH7h6
mAkjy00TwM+W4OCxj9EjZYSqXbxzFOxTAVtR+c3QhCv8y44QPFgysjhsQpx1O7fx3U90kko8Q2SW
m527cFIfcdJXaEcU1olj/ZFqmKHur5oCnj4xS3/NcKPdjiRMW8/16v7i5XDTMRW9NqGjuWvHMi48
T/C7RbHdb9IbOJXkeh5uNJuoqrYWLyQZnouXohZBj1UYViGPSK+nOjNpz3Ztk4rMXTD7kG5nFcQY
tqHbZwNfg0TkgfbCzbE8dw5meWIYLs8AAKt3Lf8nGDUGn6Pzjba5i+OdfyIXUqg1vYT+YMaPEykq
b7NXPg87qQ0q6eE8ddGX6EEJnpFXGfAN7iDZ8dM06R9s2xXV4HuXLnXb8b6UNBu8+3rb3Zy7WrW0
GNoSh3ticO160JkePAYIerdZR9eBkMHdIt+YEm7ma+BGac/D2O5e4anN4KPJZ033yfq00aTFfbzc
kUV+R0hWcHSOKu4stXvCcF4b64uCRiaXw7G4a5sM+IOVjqVS4dM7xGT8bBud0I1wrAnhwbm+R04p
NFI9WB8byO8cqr9fcsAZ2gw3YciKyYERdlKB8qqg64vUuJulAIRtcs5ukiEU8nl6wTIfVZagOkGF
Ow7mdsOiGF+G5ztpt551NUj+MSCA5v1+uX1P05MCrXtwwjT51hHU/zrswE1TARuxAu23F7zIlqfr
qN/LgXp/W3WyY20YDJa31uDnZiUWwCurMOcP0ahG6YSZv4TsHEElHx0dTsA7twTaGUMHi6rT3uuy
fX99PFuJeEHgEj2Y9+j0lrVn47jICInPuGbz1ERZbdFeit5xuQ/OWNynjrFs/0awk6KD3/VO11zC
0NuKdLeL5nl0WIPgOlHLf8GLkkfpYMUl7jVoKjWDHsSfik4I/c9WvE17Rpnrv9VePLaJVjGbdaCi
DU8CigLxDWB9wtgTvjOog/p9ovFJYWwipMhDSUq8tD6b+4XePK+YMjeL5dDMLTHna05TSeudDq1g
R6yBNdXCnl/Td8h3QIWsDgAUJt8JofZvOItcumoerHBjOGj3P7nSZ+pmvNYFTFLxAQVidO21JGDd
2NGddiPkcqCA+837E+umJFp0TqyVJEkyA8wbmtfVtrx6oGcglwY8uFm36NJwg7gRlQcnNKUXiec6
fo5JwWOYAjFR+3Ro7rk29sONPgFBvgDB9Paf2KFpBPi3CbQuaJcPdm0kh3rH3JZHvx9GyC5zHIPg
81dN2EV+nzuqB2/Chn2m5igF3qTJ1LkuMPXIPPijaA15DDj0AuTq4XGevptO1z8efXiSA1ix/4IN
dcCGyaYy+YxjoObEG97fN8mpMj8aHTqoWMu9lk0kJoABKM7XiH2r1MVG6g/1xK+NZY3bkpQlkxIK
ZNlClWS8UiyT6mCcc9E+9ZEmNPif1X78E95o2wVWtCzj3I1XPL7y3D4HqnAsavY1lJMfCEuuW88f
ChydhlQgXdwaMmXPqLIk81JQRR0rm8FyxuMVYEITtVr7fNSfNe+gmjylmrZNPC2KX8PpUi4LPArV
oR7UsMwBL0fEcji3aavGwYdShwCJlOEW/6bQqSscOE+OX1AKlBGLuDJQnHh7EevMNqADjUKpQz8g
2KRoIMOrjN06hUXTdKdfShTeUKAygx2bYF/pSDU1Amf7dXfaxtgsPkNPekSIodzYE2odFMuOvXMG
ZfRgrI+S2A0MhRrwG6jyGMlKN8xpFL9yg4e4LbDZb7oYr0kZVir/ILnvlekL0N/N1QwTrnokZ3t4
ozpKiGEVZ5z5ySa3fpBe5YL1I4+9+9Xfta6Xpa47hHk2A8t4FXGy1a3L2mQKbcO2LTrmCqXJ4fkI
dFP3bi29Cb/P4w/qPp3eOgo6o3ygTZFU31eJtUcuOULqjjj8Ww/7Er4VBBGmpI88zfaSCxpqGNLE
wEAiOZfgiZp7zecATPkcu7SBNmmus8fdtcywCbiOU6pmeIA3tkihiCdTa9R6+QTDIjyP9JL/UF5f
MEspqZlFGmq8FxkwQVlfsvY6lBYu7WVDDMZdKRpGu8z+30UUb+WKfmMe5HP26SON+OpeN15NzY0r
IfChAJkcOI3euvvFzQ6dy8N46awBhufkFt1U49bO2Rr5rWAveM5Ie3h0SN9rd8F0g5UAKkJV/lrH
zoDry9O/2EC93rAnXNTA/Kfdsvk0MPUfa9TPmjD7t+Ujw2QzWSOI3BTj2N1Dd6dR3uIatkycj+Am
t7R3KB3+3ML++6r5qKbYyENzIyx/lmwAMmK3gzvrvP1e2zqL7Bn2lFeN2Uf/18LwDe4Dpd3P1Q24
fjjRxfVxmK3xiH8FBacM470TGkJ2RK9E11KgiwwNFoxzseVcOkF3i0SfLzYEFWEbaBYPviGfpmNH
qWRbiI8jCxMSy7F853wqXx0kDDJcrqSvW8fhY4pj5N04S6m2bItMrbDuJR78SULGFxVloC/V/PYp
+FSaiNRHY0cR6XUPNSZGiQXSOA9/QDsWO+6ixoEAGkUPYhPJXIvnijyXLC+taaVJxpjpKKcuWAAY
vhUIX2bXpE62Ojz7KmxMQQ+B2Kexq0jm+u3hYDvrSEQ6V/zSYI31rWJHka29WKhaFAHKkcWaOKfY
7g+JR8VdJGUxFKx/TaHt3hto9dPbCEWijamZ2h4vMz13Y7jVWA1eN2q46uYgemeJATrxOVuLHK8y
2PWtpEPAP5YLYFf2lbnaHxu/8xh00tvYN+0I8n9zK0NXhaQO5lz0mWzclepmBJbbXR5as3XMXgi+
zYIjUiTJgb1coFnsTB7h69er2PAXCVDfBV1P0vLqSVqEyWp7tYcFHwwFqclnMNyrQFOJ54Wso2/2
6resyuksyA0OXWhKOx8rS+1jgdjVgWJEcP1dr0/gDa7kAbY/JkOM6Zu7fCzhnJnnUecNw5kzIm5T
Ptw0OwYiSA71suDkpb0pQs/EYdnqyBO06hEFKdItlIRGffPrzf2NZZOOzRECN87g53I5siM9vZ1C
HfiaW2XvhbJ6TQ3T8rFM6ZIuWDHZIRI3JNLI36DG8b55eG8j/7DBYpkWzJ4IbWp+1Hg6fwf4QAr2
oyoN/E5D+JD+ZbLcgn0io62QirPA2s52e45p3F/uMlctnf8QfJ8qjxll1i3R0bK5ca3prX5OQHe3
kpRUH0Qs+pxttMhzUZRkAGoD/IiEagvwbbdN6LYjDQDWhIQg0vsJNpEmrMQoz9gYLnbLyGnxdmC2
TbUfiB4fsAxt5tfDEjdE2bIFnuz5dEcYr0LiDVqVRAbeP5/NybV6+k9lmJBafKHF6zyMBkT6CVnh
8F44QGYPe+slQJFDv/j2roaDnvW/OuMlD6wy8PzWpzRT9AM4xpcnQNIf80OImgHk3fWSkJfM44po
klCxwfbRLyhr6Op7eBz2LyGQCSpuYR460pbiQpv4Ezydmkv0ShNlXYxF6pb9yVhNKi+PBJ6Ynosn
VOtVnZYTz17aYxd6bAfzpI+faysdp56C3OpVxb3jv7bAivQBWkXsHK62SjkPGNfl9yeRLPPMcjOC
ZZ0fagXrtp9XK309jGZ5v0Y7T3MRkOk6Mygvd5mfM4spsAXuWEftMAyNA/KK06m5eluDbSwWxaTk
+qDwoYJbsp3QHBC43rIbRKtUNIpYtpLtdRRsp9wVmsEmOsfWl0q7YZBn7ilOlvDo1byiopS9Vva9
FXA17SqRio5qKTdJzpSt2LaKESQsMTd3uQBTFF3xw7tHM4ZHFQC3zHJMO8XWru3Xba1Qd/9CV755
VJyQIp/jRykoPwqnp3Mv6pbGjUN6n784Jz985iAxcKu6jGKKuAcfvgS4DoH4CDJDO7zivLpKqSKg
JDxziScfxA3FwF4YB8VQUrlDA19RTCOngCBhFuMKWSuRWeniwD3WGc9JRVuDAOtWpQgzlfFhpPfE
7wliAbhEoSsyFZDMHEhyDrZWoW51a+lz1ZakyGpAYJn+LYs8G2d9MOvjT4TnVvdiE1OmpsA+ZqkQ
dy4L5iIbfWL+Gbxgxhypfn3p5VFVz1RCziyZkCMnhsI+3MFNNjD/+nN99adZ7v6zr2v8b1/jUqcp
ClSCUnhqhG4nWJqVn/ONGXluzCi8sxOioPhJROzu5qzdGD09Z6D+fgHb0hj5bqbsTk0MXMI6YtJA
5actl8GGNK3hIDztz5jG6rnZ4spxj9F+0l1Ad2TE2e1rdfklGzdd/JJunq20Md/X/1z2SJGF4VyQ
LOH3F0tRObOmSaMDYmvF/CDlFzbfty5H/x3RtgoV+ud8Vl4fxHRur0ZfYfo8ESmnnrs6wjz9Kw15
3C1YtSjwoJVy9jM2B8otUa4sz832OJzhEiVbh/cNqv4IQP+Ujy5zkw9lobdoJh3ezgyDGazdFmEv
nfIw5KX1djLJAKRwou/AExK0T6L7xZ4wueCw1WPorqd2/PDH+KF4tQLMEsnQ8YtdZsqHOPHTc+rw
+Fp3mIRqDxWIV7RWNVTLcYgJ3u1mi9K669AJSacOZYB0FV1IW0+wYSX2ErU8QYMybGz1PahOQHq/
FMn4j8Uj6xhHa0z4k3lwYXFQTwhqTDmzW2Dm1gSa/vJLAk0EEqQ9yC6EHAEM3uVcZrCPlDpIE9zX
LlybvfmrF72Jfr5QDPJk25szorbh89HwcrG/ocqR+xnOUipXBmkopVj5vKgPY11eSBUIYYzddg7S
pdAcawgUM6bHdeTAr3gpdYXwDSjD61agDLgW1pvm40aZpBuzOA+QpKTXSXVihii26VyuX6unezlN
X5aLmQ2i/RHC3LvIzdlNghdH1m3POL/KIyBvR1OgmwF8RmqegFSJGdx+PGZNtU29MyK2Q7wjcItA
3oozVbA6CUM9W8kDJjl0/y1gPP9q/tViMHUxt5rmIvgk9mnl6ReUwDi0K0SBG1o47s2b24AvLG2e
nFqLuKeCMdSvmAM62UiU1q6vXF+PVAT/1C+2gdWBvCOhRn8omsFs7apz7lEy67ePZAWBjvoAy7Vg
fm3qsgrnUUw+5eR9m81n1I/fIVkPwywstj9aDuSE+jvvBh2amy1L2CwRMQsbzj7Jra3b6ROEuB1M
d2t1+EjDoVN2HgmwovrHQv+ym8N6YZRV2prPKLhLCWHOMvzJwpoXUdnrE0+Fv7ILjVgGNyd3bXJi
/CR/5+RL3Oy9vfvz2hvJxBw9FXHZ2LBX/j3wQgqzeMUOStz3vZts+1VhMurVh/9nEc3M2RXz9oeC
C7FifRSo047mEeAxv6oDg/AfVzqV0S01ub6/hBMKrhYRLABZfmKa++R/3tugTDHE/GjG7qNesmD9
nAURXYY2GTu9XQ3eG/QkUrn/aVMHA+YhDseR3ePu7kc72KdagT9JtGw6982IcU2MumnDgV5Rm2EP
X1QfSGYDtbXnaXkFmn+yvmGsXLgWcDxV5hvly5PQ44k3EZkHFxt/K8XSEHZnXc3FHcag/+FeCeRu
y713Oul5WRPwcDKxAl/CF63Sr2LfVbhiSsj21iEXlt7ejjWduw3psNEjdIr5ipNbqzeF9YntK2tk
1STDd+B/xG2sfikpZZeORiFSRpKhyZZ4541G1ASj5PnzeYrucmhd9kCQNMPxF9+Smg4Wj8NfdsIO
WqHWSZeX+AKKRSPqvLghI48SM8675hpbCK59Xuy4oGz9K031bYpRprVcZ8tFtEWnYkuhu1sWyHKZ
7GfwHX6cO+rFylSEurrjLaFUbDw+RS9wHTkbGKjTL+Piqh5NBj2j8qvZrHexAeHhFTjm7s8EsFGz
1fqLIYNS2IUackPuac57bGoJWItKNlp0WuzviCl0P04Jmnnzo05dGVi/+ERvn2pSzJ+AX2AHvMmN
3yRBs8DlyCNkzUSLkY5N/pPHIP3rvgdiuWEg7GBB+xaS+nuy1TW3EWeYi8m/IRZq4c2wydLsg3Ov
2UUcijFpV8lyfZOrlPfRHj59bFz0TDg6+dm4aWxaQhPFYljStDiaGTdt+GqjB2sU4pmGGkAJ7T9s
kE3QLowbLWczALYB1HmtP9kuXo56Pt2xiyqKPyyZXoKQukGx/ZiF+tzJli9Mz2yg2EgZ/vruWSLW
hpW0UjBagsrQpf/75c4lKPY50reLlEYtNTxGflWnAlP5g2tYhKVrsGd/6VteTQ8aQKeq+ltGvYVH
b4RUQc2u/rb4eIg7gJ4gfRPcjTmyCmsbIbUxRmzhknC7J+ceip/j5OJHSPmpQt2eUotW5AZUvV3Q
GpZTohVQfyZP+G1jygXwLV+NQfTWEOoMntob2xklFtKQZf1NvuwSimjc28FQfzkv8wElDbkigwER
BNl65J9XE8TfeLIDTTE/uPv52J21ipIR/A8Yj2sHvCg0RPn4GiEpw5mw/gRbV8Pk4kEZtAG2rBfc
sK9gZ8JAQtJNEovDWX6sxMeh0sGSYR80TcRUhB3GUcfkwNRb9k27Ga4swLvtYISwXDkUrgy9409Y
4snsr/uz2S9kKPKqj9IKt0JeDuYzVT6BZpbNoQYvlQHfnuwemnakxCcB21c6rYNGdmZVyfTWbqu4
g7D6UNojk/5nIOh+LxYZn0FOpPVQGUl6haBO+Dy5RIFKZEL71/He3yqn6QFeXbrMXnRlCgWHmdcl
7iHtAJ9r1eyEKKx0PrJS42qNN+r+3rFQga5W7E1qXCY5cVIdYFxwNqRD38g6/PZmBAxu83qPWl58
jbIvKdgK7tLNqwtAGbsEsaedVzbbqX5exHNwqYcwdlYr9SkdLalew/N79M+GDA+nFVpRxckf0ppS
D/7B777pGiXZ1Zk8gPpPp9N55X4XypP2j0w24q9Pggz0bRhQG8UEmUSODtMrH4PUhkN9uF0rJMl/
qbmIrPNRsEy4QOAN/IOQRtSkcpb7NE9JZqe5ZedPgd0ZYRELHSAdPwyvS0qRVX6OZZxtMSyIDE90
lTO1h494Zoe/2SQ2c8CPFl8VpnkzkrbveLo5xkEFEaeXI/y/gsqlu4WXa6GP0dV0wZJoQXanXeYM
6NLmwqAZ+UC3KS8OXUIdTPmSEICX6dYDpboElLCBAhbVDtjZV+MawJjDKqQyBI+DUMJqLnhHHRov
jtXSlepo2hXJM0sljkLvul32xko5lzOSNoOfWECXhg3/73ArVcLdyQATVfHPjM1UhjagRf9LRKih
d1uYJQB7vWXzl5JsFxxsNaiPHNRRJt7a7jamtbFL661HAEh0CjeC/EWxteuE3G5y1jERn764QOKU
9W1cAuTkPXA+Erw5oD2qmbCHRVgQ5ePcVaGhJ6eMWv2ZEfNnXit8+thb7DJTkt2opa+6Q8A1U12D
OIOvPlEqEabsQQEIuOIU+504d31U9VJBPMtOQ3FiIrIjvwiG9Q2RYjXHLA67xiXtTuQzpU1LgvIE
E1v60sdt4PNV6Q/BP54RjPNZSyn/yn3+gdmp6Jeg1GNmQKbaB3N/yFIyLBvyIkX2NhiWetNN3p/H
tro/88WW6rJ7TEj7aQKsdd2BMmdat/OH4mqCzwJ6sk5Uouh3bQi3/gXbA6XYaYpeO1Jlyf+CObpf
dxvIkm8PZT+LOu39+IX7LhuLa1DCYOQzRkRPqtmAn2xajzShyfOxrN7R2bvj/7RIWJiUIAZypve8
ggDW5bcdEBQHXgU3ps+Xaz8pC+ctygN3h4XlqU5DqSbxR4YekL28JbqD6cDJuuCDBsrwj162e5+K
eS7yt2nMJSYUlvLxQWJxcZaDW4yvGYjXFRoJhWcErh0RFG+PUC5nGghn7LIeEvLb9gNR9FY3oegT
lFbuwb3hiEmkjCYtFQoM6PKW5fWjQKPKoWDX9UUlro5yDJQUXpttXIGSWoGk6r3notQ/AyQw/bpS
Of+rMZM1quY7j632K3ohfu+lkEeKKliQBHmYYuounHyp5rkk0Fiv3TUP7/TXi468VfepunZ/rtMx
BTKa095pRvYpqqTxbvK7UUD35rDauMBczpF2dHYfBhOnRyn6aRNURkeIILC9fnYwqPMiCP2ra39f
ZD4M19efmlZW1phoZ8DieGIhkGKg62K+XoUCHxrV0PgmbU/r7ZD1XMh+vBofySBsTmH5Io+HKDLc
ADghCN8bOn/CyEwDWDYswTPfQkRhPnaCWUcPoOEqgS6z17fe++WQ1RlHNP8sLUpwQsOJlo7AETFs
FIIorDH+A2eJ9VV4WGmUdGoRlX5oJyLW146DFTvX+CxkjtBsTg2bpI06dpYTAiEqaqLYr4xtbf/2
M/A4ZYVpm/yEn2lyGzMefD3wdJdr7xMgDyE8+DVt5N4zS2YUE3JnwnGa8eLyM+vlP6twaNOJw9nu
YfMH359qmyXzJaG7Fr/+r9Am7//jwsDnMCgSctQwR+pLTJ/XWExd9yrdxyiLsm/Cyy/MT0mAtEFy
S7BWUeG6BnJyv7bIELCAYdRxKxIOi7z9O+sQpxuOXKN9RqKasCw91ipqtGQrko5lAzgN/K703AXT
ulr7EdxZ9PE1GxIuLBYft3ALG35yBQ90tJd/ST654H/ZomUI0fPff8eGCiBHkiEgFPTKZLfJ7XPv
Ipp/E0EPQEeuNqL4YzdxYkwCwfsQEutMGvk2NE66A6DPU9lm0T6GmXf4rGPlOPpFf5T2PBrzp8xJ
ce/WuFzAi3nw5TjSaRpv7UxHgR7veKAY7akQ4WhM5tsBXSH1w+zHEj/ypVDYAU+9dz7veGpcRB74
GB1cvNITuUbgNtG2ptb94LudDxBb9gFJYU+OAAmu3VqqWZXYx7Sn5WUZoPwSUXrX45PqsXqzy5JR
MMh/nKTYVviCF3dIQebWh1SbQHkwsoMqElpIBMmLn3bFCjj1u6Buu7fsd/hLI/3PmKg9fzG/lZQM
PlVMv53sIOGTRxFMGg4bTyc0zdtGygiKBgZeiMnSWcg3eS6bpMUqRjjZNB1VGnBmHnEOrxdasDVU
tOrTjP4Zlcvb5o0ttwj7uMhs7dDD3YaGxWzg0QtiKn4BeUVIDZDTvfXROkem4TV1EA4dCDXglp8H
bCoBLvzkf43CZVfY6x2wIHKl7opBwZi17lyo+B+9mXZvFdmVv74NtOBzGRUZ8P6OTzMxiIu5aJsj
yAiGm1RaRPsnAp7IZLfl/aW/gRDvZ63Xer+sul9q9jrWInxBh4vW2MR1C+yOx2qhymLOHbyy3smE
e6dWB3PcwywqsJtdlHJJeD0QJ+iZfKJZ8fklB2Yeh/KVDhb+8mu62QEAqLk+LDBv6nUou+GrRDIe
CP8vZ0R+BfgT8elyVmqBOho+CpUOvzwoFr45DK4JsYFR7fwlo/IL7VnELX6Tn2NWeKRrZpC7X0Sh
q7eEGVG6sv8O5oWHBA30GzoO1dCBGG6zNkIGcCu+nCJDYXQLtXuwC/dKKftTZEshxiR5vz64rP5x
AMGTZgaipB2BYDb2dWhmpMtMf0n4wSt7cFY1VKAqRdQm9dUefniMqWhhhyouopxdzbGxOYf2+eUF
gDfXv/1MNnYHG1E5RR63fJB1hD3b/Bgmhya3mBWVGnuNEuOehM7nA6IiPuc7h+0KOXdYrxsxVqAM
S0IotK2Z0/t/+7kziDtoapCLQBcA8HWZNVHjOCQrbxyga3G8S2oRN+aGdoA0wsWWxj+RQbmHqzcJ
nxesf7MTHbeDtVCabDsTgCYzZaYN3N9gcDMhBPRlzPXPsetvLsqDKCQsWl5Clm0Wz5ddlvxgDB1i
yxTr02fK8pocyHkPYbR4YfsC1xR1LUaSfKq6qNTOp6fBMPUp523OtaIS8lfyNpsBLmh8fJwfxyta
5oAKrOeqreZeHGhqEMqV+6o1W5KCUYoFJHbTCVN8bVDnjBo41IPJwcAB389DVRJteC6V7Z+O5Ith
6QOSa0hLDoU95EeMamwyvivDd1DR2/rwSlury+S2uivUFwPeNJ7afOMETVsA9r+7Nn8a1VWyZgVw
j2nuMDjITYQD95nQK4QQYDbuNdBQi9Qoa/ZvUHMszFEpvvD4GbZKzc8JoSJ7OKXmc8WpquKX67Z3
sD+TSKT4358HnK8nwYUJwiOj3GZ0VV1XWQw077bePv1PYN6jw7aaACTgCZUnS1cJrhMD61HmZAtz
8ZJr6iGkx2wKj/seMrrLqUv2MQLkqU9/m58BkGItz/aDrOO3DQDUwynY9ARyOrtPpManWqFGUs9q
dJudaZcSA17GNeMa4F0m1HB+1LOyNLn3VGiAyMIGbquOuUvCSWgQWo9ZH53roQ1HfmU78feuFUCL
MIowU4Us1wm1W5H4QGcqKHknyE8oVdwzBYi83WVyeNN4BQKNMHMtdGEUmEoBphvuFXW3FBsD5jII
TJsRaWjBBLfmwYHbiK4fVR+viFbUrywJTnIqCYFby1q7dBRWrp1Gzu/hTuLHPxSUPdLK0eiNRcVh
+d8h1xTvkgaaUEAVqIueJE3m//oMtMEpGdqBrBFKceCXoXHiAuR8me0y6+px+piqWrYFdnIFheQl
Bu1rnDDXZnUT50I0fGgmHcar9HBCqm+PARa5hnLi1pukGsGCNPFgYM3G7Kmy+5EXCb3z7YeXT0FS
i5hl/PiGfuqjPJ28rL2Z0Wli3SNfY/ZRftA+eaS4YdJV/P3nqt5QXRwbIxZtJz+mCk8sHRFLl6UV
WruKh1kw78oK3hh0M6SjcWwL7ErHoLb9atiukck6qaXLTcPvI9gN+b4FyJ0aHXEjrK8m+WBFmItD
o2bxsI3gH1jioRzv0c9ErxXJEBEEOs0aD8b/h8gFyfn9S5tr3d5h/W9zWaAEKVJMwBeLrPBPn5Se
uztQfCslkBXys6NinpWZwoJas6XOCkIw4g1diK6Hv/FivvzSavlKY+x8YYkQn+QNVprBZv5BzNmE
pVggldeIKxwdgDKiiSjP2n+Je6P7qI+mh/nQi3RdlWh180m2L2nTI3GTi8ADp+M9DA5wuvA3BLwq
B0FR9rwppmHOuI78HBBwJ6BIfHciBZfqjNsiz9A+tt+PugTlqWq9A3Qebd2muXKp7ltjtayCscdb
IxWOLqM8iPpVfW80f9Gqg+JpQQPNAthsaXyNU2BLFidt/xgM5tMZddMm639lxnoTO4kHGlTvTwU5
9CW4W/acBR1SBbfGTk03Kw7/XK7VOF72B7v1ft5H3XVzQCWHtcIDjC7dM1y3ZyeAg9U5yZuVcpKf
gv9undwTCmAsMS+0ielIadwfHNzpumy/NnAYktqpbnm4yXxT6N3ZasR1fau85dTzWG65MhBSWckl
V11NrfMVS0RrjzyNQIKPRch6RWJyvS2FBXbXsOnOZdmy4ST4aHbAVMLWOwIWPZKZZ3yajm/q/8PU
K/K+uEexa09iKB3jH6CAi0ixhVp+vmU1iWtt9QwtOVmddwETyQmTj55L5X+wKS5dvz5oZIJh0fvh
DZRazemGpkzOU9EJ4W58YIxcPzI/bxnXXLBldc11fR8wWcFRRilty1mZp3ZUOyQm93/sycOFacgX
SfvepUOnHZTuUpp9H60Za21NnjsnjJHj8q/vcTELYXS1pKdVjh1K2N5yAuEqWF0mpIxDl/DskIIm
o4Lkfnf95yA7utY/liw3JeIecISAEdSML8WksVptJWKcPo1IXRqEayTWVOlp1f5PrxWpNx7B797+
o/0rWpeMPPoAXIRtyxxrcMUwVqNW0Cvrh+VxC3kJPTi/tN/wEAxbIHimCzINkqoibyD34mVezW/L
yJl0SJSUW6OS1gwiwxhqDS7SFNLW2BzOI5fqRgu61vE9YGOyNC2OPVVS5mLXf0fc/O5BergCL/AG
+D28RBzoVch6LGj2soPfH4U4eV0NQ8vtRR21JGlM1pVUBaxeBOkcKznQvTxqAPVfu/qdM/nFeJxp
6uXdIGqyxefxv/a7IVbfrWn0dvWXmClfK86rRcaqQwI7d4RE5OSoZcUsEjtqzoH19M/keKID1q9l
QXaiPQWhac8Bo5JKRJHR1WBF9iI8MrTWiVuRrqnJdovk1K1LfzFlytls9OGZHmaX6yVH+sGkf5QL
MF1M/5D8v2P8Gzm7Je0b0Y127rxk1qH9XDVrF2YVi2uwoCzCDclQEERcW/dbX4Vd3HK7bgxfF00y
jMzyLD22mBJiG9h373beqNFkFHMzn1eAY9B6rLzlahnoTSe6qdOJVd4sbgSeZq2tk4g+z4UbwW+g
zJGcyMh4DO3dVbBUPTNXPWjbj9HZH2cq5IS44Q6ZwdQBEEZkyva343U6IvqxjqHRz0Vi3/Z0ZI23
lh+2BD3T7W7X+uzfzX0FxsJ9y5zFzoZSzjGo46GCmCpVIGMq069uuknFQnT4x6dE4yA1lKe1p/LG
V8RfOYmNrGBmpRK/B2Bh4HzzSnnN582HSpN2gpFXf/HIoez9z9ktBtJLmWvHsJEzvn433HkN4fs4
QUFlBz+rPiMsxuCsE9MM0Trv5dXnQJAoPvwMfeQ5GRxYvtk2qFqcsLSfRL7vVOs4Cf/TC80MCB5M
Onwm7KH0vt9ZPPqiaG06MtMYDy7M9ohwaKE7+egoHDGiZ6uStPiFZyXtjhFHf+xfhb/hc7PSUydg
970WU1NUnTbBpYucXoyuCC5JbMs0Ep1OZnNs+LBI9f4onn60XWaREO8wKJyJ6fOugcWlJbRxUHYe
QadEkkNp+6TzgWTVFZgUOkp3KY3zuuli4ERXVfo8SRldOXFrD5zgjfNn3tGrWKvpwpkdKHLseeqp
MrkFgBEoUmOWxepaGvrg1ruhUaOqDRKO6qWgR65PBrKBbYIpqbzZqP6gpvEYMgPQ2FzzG7O9bGpN
4GunMvpkn4FR7+UckleVOALuL2t91MOdWcavFF0pod9skDerrS1TMgfDpF06KCr2ok1Re6Jkzaa3
jZaa2AmHBYY+97Io/BoDNvEnwY7cfO91HDYj34dTaOlZdstyS0Cl8Xr/BaezQfxydx++TRVj25uB
wKuoUIiWOTHdolZ+AHRdRWgK0/cBrO16ACmSBjw6gkh8n9S6wVJETBdnE9lTa5LN644YSffSsl2K
aJIe9M38ijymq///LlA4sqJ5Y6EQIW7dRXLh5WUEzuCUonG++RUWcgy0uYOYRG/T9ENP1YcSDs9J
IKi276VuBuGVXdzVBNP8DDvDq+3eU3X6yDBTAH0rMN8CtbumKE1u3fAWdl+ssNsI5UlQ2qzCKyYY
/0nVpQsWImL3BcQHggh9nh5IfzHTkb2BcEMWFcozqEsYyqqe9QFc/hlvK9dv/GDPyaQUp2G2MTHb
/1PK+IdIjW8s8UAzrYecFrW3IHkWo/WUV0+IyNKsf9LqZqihWePgaWHxBTEpbper4qkOwai/QwvE
gzbSssPePgAFjKjFtXGIMcS5zuVcBDk7QS1dhE6d5M7P1PXGGrLpas950/vys8a7VH/Pvex7PjtG
bzFREJ9+cYylXbRrK/qulE2LYbtVOSPd+/KOx2WfoCUrQSpkL/B9+106eqtcjHxtRpV12buXdmPJ
luINFoHKKLl1WncvK4RHwv229/OiJwygx5jP4A1OOivbXHzG5NAKZ1UF9HjR2gHhFGlAX0sAgaZ8
HONKh9ZVwxVivhTnCT+bmbNU1+7vJBoCVOsAE3jr2fWJTkC7bj2vTbamVmBy6cAj/M8iyhUEaO/+
rqVCZd8v7G9z7+EL15jATyLjPvcFGO2YIi3o4xWPjGNvcgqaYVbXMDtygQWxS9Pn3cwShXRz1Dyk
SEbi3BM8gEJbIN+O52QKC5KvItZzdjed5/k89lPtxC864Sk996jXSGTe9TYEWDHB/N/n90DvvZEt
rLTVqqbkDBZATW5uc8i/ey6G6qLfYtyQx9PtdMYgHZiIfJuzuO5ZcCr/4Y7CL6XtGhvJgHqxXM6l
FGNFr/C8xQzRdcbcKzgxE2fFv1EJCE1p+ClgXFmHdyUZC5wIdmgWwyz2xNnln+bwgaSKeB3CsIPr
tCS2MuK3BfZsnDvSUtDa0gBZFNTbkcP0+iWYGYbDXpV2i6k0oEWieAHGQRqKFhQI600LwLDf81Fz
z2sQnR/Kqde5BuG4vWC25hZZixR8plBWyYK+2B2sOh1rnseSA7Bfp7On1Mj41TC2DnfSaYhGAjT+
92BsKriXiUC9286TtKxsbtMeKJKf8B4axsPrkDkX72riTK8ajIiDYv3PaDNN9PKbdK/qW0Svq7Jt
nG20nG2qm/cj6yP+e1qzDUQ0RgIJ+WHb/Ix3EOgNtxrVZJOu5Q+0jb+HGNPVylWI7jQ+4pSF0uAR
VLs2JP97gIxBpvuyJrZDPN+U+h+QmgfPDywdjmo5Nr+avlaF65rnPUqEDe1vbWeUtI+vv3BYDtc/
4kSCz+uSQ8CaxqgAJe/jJmQU4Jazymavk62ccx9SIh5NHAXOTbWjuvV9kGUDOoisLOtoy2xEhK6e
zM0RRSZyfTOoM/1BTLde8sjAU/3S7MCmsA126xM8Kv1ypEElfqE4MQgjSpIpGyPGTZfNsO/5l4VW
2VleI+X3zXudgOLm4C34KFie2QH6rzTRra+K7phZ2BPl+8GnL7tOthuBx/nw2HUDtaEMmOTusPzE
X0HgAQrU8CQFx0nx3wYx0cHM8aIzmre/8PtulSqNBAn5tUlIM6JQX36UVyQ4Yxvnlhc18xfBf652
Qxl3JQoaOrCs010sNWJp7bxadznKIY4ncUUxpeLjWvS39t0BDH9v6XN6f2gAlkuVlsfpHL31Cu/f
9kdZHZ097hj61eJLsB7dYHBnI/yCyUYfny1qbUwJ7dkpQnnN4khwN8+t+O/XyQAu0jR60OzWMZKm
bcZQqIeYPlJoOdu2bWUWX9u3AJyqSMtAjCpJ9YMpUONEAD+40dFl3u3/nbd0h59S8YOn4mR5roY6
auIWHFZynBAcyL1jzMH+mERJWHEOHTdTkyJIQZRPv8LAllYgvJwjCMNAsslsLm3mJ4w5fnNiQo3w
WA109PPXVLrUt4pDBehEmX9Rz6J0WrD08a2a+jHBILZItUP5XLyBFqQIAOQGKGI3+5oKGsXwPEFm
Yy5mapN2sV0dUAr2ygUax/q+BS6wr7cwPuClny4HwX59WWXxYW5/Cl7BAMTr2UMxRW7j0pxEk7/x
8Y/44bwMEYEMubm07toMo9ANZjJ/GdcTDH/f6UwdyjYhQIs5jLlTZXOiq56tDLpvN9GfQHxhIBLN
sy3jOkVysmy+NHUyc5lELnnCIZMh7+EubgWUeBUHsmCu3QB8PhEqKWv+718eSgPjY73d8KQIREEV
CeLZJVjyMEIHGL/v5cx8F+xPq6z54nEGlzHHC09YM3JiMeNXZ9SwuKXWz3zW7VB4d3JTyKUToAnY
PgxUqU+r6Cm+4dFasKF1Ul87jGWMcHm9H8lFs3bZeTc35gmzk7K/n+Vn/vCuYwjUYQpTyHAGaFJJ
FoY8vCfYRSy3wSr6ppV7/PaxYXcPCYBIhLqhF8QyI2PdPUyn7ADUGgJNkMd26itgT0bTA1F0ANWW
3T24gC96h2DF91LksnZVkkraSvGOlhXx57Hvi6Z+Xt/RSkZhcyxRLe5cfEymWI1vAdIKUTQFFvLL
yq9/tun9gAk9OJi0ze0xcI71Q2OWwHxQ/y/91lR/wF8Fs5GkfXWhRZ/ASzWFrRGQWe2CQWPVnTJG
/iNkUdVpGCywr0XnGRSnrHy0/ltqXYkwOSV0gaa9dO5l8cKovuewLzAK2d3A3BIGClZGw2Hwxo2e
p7XG7fmpAovOEfr+wwmDYsvUpkb9IUq0jrOil+ojeW+Y8uFrmcSrdlCLRnQ73Mn0zVlwkK84A+mY
NjUumVZsDJQo6/gCMUTuYTdMil80SMOKWUvr3N/IatbmmvYTNsxB0bmqmrEKNZJupc08K7leieZc
rFn6V4aBbauNlzC5RvWP+tHXms85WsupK1M+IHKiF//jhQh4RB77IaGF1CL8tph44ETaVGjpq6Qt
78YKC4U0sQCjOWczNCGticYPYQ6krADFAphdv34oAa5/JJ85h2WQcvhryRYLKokgK5nDyhGN/Ufl
UYHDd7mEQIGvG/ZfzTtsnjikbEfK3EU62xSqrEI0tpmMlMnK8sSq2D/DVehifmRZNvGoJQbu/64b
WMJKdFNQunYSBJdirRiCFWMTpykW1GJqWuzLKetPWp4xH9TUsXu13bu077XTGJFMbTyfJcZ+Rqc8
KLnjqe2X4DrUMl+YL/5y3ZTbCKl1J2r//OILKyqFM1ArRFEP4b/YtRmIT48tsEMOUYQC9oCuxnek
fhGlwYfu19rjnCtudA8QFRzEG7ACa9fhWTV7PxZGDMDA9Qv1Qs5+N7x9U4Cwhv1/z7OurZ0p4YBD
HuxhCDCQzI9OAQqYfJ3QH2DG7Kcgex7y4tM1H2fukln1giDP++Jq8vitslGx+IafZPiu7YMXdOmG
xeFu6JGVIEVTtu/cvzNcMiycU+eAAHjwmd3ZPbo0innr8MSwyWVwwIZlNEo2GYsfU8NcYw6T5sxy
EQ9phdQ/ITu8qYv1PGAY4KgMAE5F5b/Fi4TNP7t9RJ92gSIbAW0oXO0T9SxYhqDGULJM/KNgNa12
RLF+BCL1wZOdfE/IESXL9ymAlUadgvZWgSeMMBhneq1bWWMAycIy7qXCFjZiJUhGrIye6rTTTPnf
4L8VVCDEWkQA3Jvk2a+gauHHO5Qt9rgzvb1jhHJeo0q5E7R8m3aipwm/aEiaEl7Ps5Z1TGVlajqg
kEHWnoqGJ4wanhMmfToTyJHcOgwKt8sYAFpMOvNq/tZJi2eaMCOq70oXMLp6gSTB6bX/Bn+FzTx2
xAm6fH4wW4Ysl5s7EZzJF7FoqI8dMGH0p2LNCpu3jYY8qLd3gcHfmF78bOo4BaOnTtegx+T67F4O
XLwD1QIFbAcgddZGngnj/Z9ptQaMHaoes0SWYH65hQDjCh38rhzj3jrKj6hLzaSQGpiGcnLbZj7b
iTyqWEZx2bOXi3gQletzFWrfLP/i/XQDAFhB/xWa1Y+h1M06t2f50iy9bnaSZ+LiEM/86KkWL9nN
YG2JhhZ3/LXbsjx7OZPXeFA1oH0+CTWVWkQ+sC9MJNnhWMK8eEAk6BnsXakiEXWGsms80XOD5gLU
vj4aL14ELbtQ2X+CVDsFoM/7o98WaZ8xbXADNOQepe1tyx/M+1yeXf+YyQ+fMTHRTaljRcUPnFjU
R/OE0iuL0yTknxjY0VSqrBpzPAf1iWkByNCUxzNw5cnx3YixOGb+7JSkJUemRN2vx94sSqNTe1zN
IyzOdOnnlMmN2qt9gP5OgGeZeWGOEm+o7bpl49gzK09K79QUuqDgt/Xlk24O3FdQbC10d6wDfyFM
0Mjr82lJrwTCgrZMtEjTMgfhPA562OmXcLODkB02kccqZexYX9sSySCFM+4zJwPqQ82OQP7sTtBu
UDoLtjJxkx1M9LkI9wpzQ4pQX/zxU0E+QUHP5+BiweChVnd4xVIMkVica5Jtpg9lgsMVIRC+X7V2
wjm4wTJQOfRDggU4gXM/j/RdGQ4JYnBF5elzSEhsTMvznPsSqTup1f89uSfW1O/EaOyrVm0rqB7v
yeI7JATZWr4fagJK/oncKlIGgHxuE5HhbQPejEKTMhkL5QTr5s8AawsCdyebjOniUZ1+8vxtQ4Wh
PCwy1cwpNfj708Dio2f8NdpzhdohoU4Q56HxThCsJr+8/Pp+nxiyhklG37HGEA3ZAUmTmI5AfrAJ
g1Z9ebmb92eq2y88l7uA57C5Xxn0Pl28kR6OQeXopEqCb2Yof5g3ua51JnMJQoh9ZzyLEoQLS/R0
lFhbhx6/D/ABRIi5A3NoUchq1/gCLV6yEN7AyUcXMv/ydgU+YJ2tJh3ZbWE6MwqWeVASky0Dbyr5
OCyCj3mZippNVcCBckF6Dmif3Tr0sBxZgCAH0c0J024Gjg4ZvPLgWT51C3MFDM31t42grYXwlu5G
lNY97P8ZW/FHWHrD0uISw1wVpMOXxj/sWfwV6W4porRDJlt2IyfU+Hv/r+D699ng06T441w6WtOw
9mhsQojzu2Nt3VydJzgte/24J0xh3Dt82yRFV0pbFX8gjxYfnPM3+l2cnpH9WQ37XRZuoi9vsU8M
ByEcV5j10l5Ceap1YSe5kveqkVb79zkeZvNU0ocoL1o/IJB9aszfdBAfDM5ZlHLq8FVQ2f6azKiC
iuVlG+TphLjPbbm8dEU61Ux3Qs/kSQmIeAsGoMl3fJ8rt6C2bQqlq4s8uacM5bd2KqlbRJ1RrCCc
cmSwXgnjj4rOkoHCa/Zxcah0ovQJA3Hregp7v4SVy3wsYGH7ezkJ7atq5lRopVi5N+HnN9qm3XiI
YiqYq4/7Y6wqSGE2oOYquMmjNNSBlUtXXhT/IVizE1Jiznns9RLLKd6PIwriNWzupOFPE2UnotBm
wbb2v6Ak9x3PO/KsBWuz1x89lQ/CNzSlApGadvsSG1Q8r5lPrnx3lLNma5tL51ejk+QeG8jfIti4
2X/bcjTBMM+kWsEeIga570XU0kdtg1ND3vlo/Y6/+xpO6KkRrZtx2rcmiHzhkchxVJSHrSXuCpl7
zMjEh7egK2/xXlE49uTNqT4zG47NXJspMF8rzb4TPoDVwRksvTXQl9e7wrz8UHi0mDDm6iCw7cE1
YS/er7yUdFtiyKFROgAYlSqOEPsij1mXC8PfH5Gl1ZQMSb+s/71WLaglbiIePNWgfOTiT7vo/+T4
YrOBSTdCip11RUHwK8CadDqdrM8ynaMdnhhn9qRqZ26yA/ZYRQgkXE5ySEMGYSQxNieyvuP+fm8S
l5R7OFwf/is87++3hqwhl7nktWP7tXBWI+wEeo1Vtj3cKdY+bVFY2t4ZSMt7bE+TdyAHUgtvnrPz
XjhBiGzAecfk6rkw7QFqWynEC5xBRbx8yTD2gOKjERYqhsLiTFcPjtHkUx8QA+CCdoaZ31/brt2l
GvSB1WFC7Fr6bdF64ci41kLeq2mCtUOwLW0CaPEpPNGtIjZxdbPV5uGI2diWQG7vEPGBDOLKykfP
CB828cl02/v7+i9WPGQ/i0AA9f6SYqTHZAa3gnUv3tINp/l5iDHyCw0Acp4LmDMa3Kyi5Nfi9bzh
TezZfV2Z6yDJZ+f74I0Lf8+1823OZHD3b0LS5/TwObq72kmyT4K9KRRi8QXvR7Er/qUAdG4Rn7Hx
IylPXd+qCdMWM4FAukq8K6f7CBWgtr0B++v2r5oNeXkN6M6lU4ugRNpHj1FEafu+UAsDZzEtSgRW
rIzL1902eGliba7dw//axPvIlcLjOYxvTSr4K2BZXTMUv+j2NGVtymyTPVYAJM766WHrndYEFqRv
Zkr9QSmhQMJhmB91u9I/Xp2h9jEd9P1Z19WCyJ/ppd9GAN69kOq9teYYWubjGZk2m/7MH+bu55A3
v6P2s9Xrb1lOeHZIrXYP/EtrZ69vthPK3GF4fR2ygzWQcW3HxY4xc5/JKz33ScfW0XXXaCrFWOR4
2fD/go9NvZ6HUr/vPkKQQ3f6ftpelRwXg6NGx0N15KxcEz2eqIG7wFu8NgXjoczhWCfd656nKLCu
qd1kgwMcGGvYnd5cgCV4pQR1QoF2aMWlJ/PEcy9Hh7u+WlIsP2UmqZgz9uhIHvKcfTAdEGjD01iO
BglxUFCqe8SDIwyes4/4XUjzk6vLsHpji02EG+4sLLlHxPtMQEW/7eSjZMP5Sqa8awT/zHj9W7Tx
9OOJqPffy0sdSZICM+GFHIC6UdbozK/6OX7E4Dj3UkyUoFzKObiz49fqA3H66WTG7iYrjFMsTY5K
JzFG7JcIZgWrB11J1MWbbQN4ajT4t0x7xvUs7leRQ7KZmXwQpnIvlCSJdz1KTG4FF8sSS2JGa/Jo
8t4cF3V6h4ehqiY0BLssII52GHWdej10029APqnZZ3WB+tuIMUB/XXV9711S5GLzbWMcsjG4bo5v
e/vNEiod1eD6TxMK/e+saDBflah5nlq+Vgov6kAmxSVoqxFL/wOWyx9wcPxXTZi5js/aqK+d+gpV
fD6iwuHor3K1dk0QuJWMdmxErB3DHH8vj3skS4KmVUScrVlZfUVFxWq/cBvVGW4v92NwMtE+WBi1
qm8fQEulKkKdhlrcGAz56/JcCwXZr1ZkXOTLn5MT6KBcixsbqUbVl7XLzV5J42gEdnwo7ErGfIH/
5VpKyb0S/anf9OH9XTXK2BSasOFIKuIsajkkXxX4lFKpGRcuHfcrWTWhqhRigUuVivRZmecpXkC5
WPmaGYnQSoLyZPQs5cVP03R4DWE9GTQ02tQlBz+IBpLSKMmql5ox/fNq9uVOeH/nMvrRqwikh19Y
jKKYz6h5C08YDgVXh4zEbHNxbX6qoMIjhWJ0KULh6Udegn/wDv4N3FUBoRHXPXRCRasPUFSAkrJ4
wNC/aW5wNQa5tjh0PnnvatWUJkSEQ02yEWQbIbeR0HuUS8m1uQ3WhmzsWSwe58+LVRNPD/f1GXpS
BG5K2GwnRFKtYfiGPbrcsQXQSseovoy4HRMpqVCgV8X0a1Y1VnjKvMInlbR2Y/9cpIsi2V309Ai7
dJCC6hQg+1aSDUEzeV6urKi3wI9lxd+s06tmig5WsRLLUj0TuEx2vmnTQD535figHBKqP8ukWtRm
vX6GGp9E1vITo2b+S23ZCKYs18pj2SRe/qE6w575/aM1DU9O1E8k1zHytF1xByAyFkSJNWeLVU6G
9dWsqJMkHMT44aJH6DEoCz6dUk70J/5uax5IJ7qJRwfwo843OLZOgMduCcOu8vQEBoMY586c9L6m
to42/pdTzM8D2aiefcn3sJmGxv6aX3mdzbXzCFV56NLTp96dK2XlDEhCxeyhW7ACTENAjGvU/5f/
IRkfCXWxvQRUDYVJD/Qn3Z61mOU9fwOn/V5HD95+q6x7peb4TBdO9vya8qPgD38xIA92jDexHLon
3xn/dy9v69qiWTiazUvgTvKvOUNio5T2GL8cH7elznRGnTRZeFoN41dB6A/a/fJdsBt8W5TAAlJ3
fAKZlb9ghMsJgdwR4w1CvZunycUHMFf5WJE9N+lzI2oihBsSCOW1NBBxDJvh7MlKcmzbmzl++wuU
vEo/UjuELsllgFKnvRc5YVB7H/eQkU40ZZ6t2HYMxfWeUyv9whKfEw9yKSg4C91hwmztx43UFV3b
d7A7knbnw9QN+PXfQEGlF6nP96KotxrABmpGyfUrFw4qtvvDSoVby+u66Zv6vQyD8YR1ZtrYwXtt
CWYSsYB2/sT/TIANEyuSvWUeEX95yVc1X36FcXd/+hFG381XRpYTaZ9BjkbenavWsDIW3MROyo/a
u9j+8n07cYVVTTfQqRM5xiTzP0IxI+wykjUXjgQqhk9YC5iDxHbo2kYYBBOTg42rAfPbUdcySYDT
G7NzbWl0Ojtr2IdJaFaM5bD8vPwDSjHKGOf08Z9w9hC7gdg5kf9iU/HDl79/DJyhGAC+rf6BbTSO
6t5ZCbbaGzB4GgFLrq3EKykPI4Od89bVAParIVLGwBBCJC0hcPrnV7nrdLJixdohUNQ+AAH1onaa
dygbgBTVCe2jKqpSegmoYuCpmxFsgUEsHzu2OhQc8ypwPf5ct+W8yZN21LqvYu90sj0g/IFg/bnh
duKP/NuBRdF4i28SbB8OJhkJXzWKFRmm9sRAJrsPJb8awGLIPGngN+cR6rSEM320VvWzHtQr5/P6
haCuvKnfeHexrT0Z8DqqmXUiWSRUqIPYMAXpAU0rvCQpuPRvhnwXatXcSyMVvqg3wcShWIzt5ckD
cVS1+qddTsTCF1qDBm5568rc0WfRlCeFdieuWNnILE0foU49lkb2GA6iv+0pVus2hU4gGHYvpPZb
7+dTZE2Ok3x9JFnWXt7CUxccdbEOrPTMsiJ8EkqM84GN+oZ6iyEacwg0iOMkiYiC2jB/go+zzSqu
8G3k7vNSmwJMIxzMXfOUdjN+PeP81RKRbM2GDkSCipX69lQF2b1MgnWWdjiZLpF4i7yvjhysnV40
OyNn+otDUSV53wAFQeNp8oL1OaZyqitH9ImOdvLAReHQu4B/OjUbx1nuoijcpNjXjE99YO19w+q3
LFur57BlpuQNX2/U7ekA6g6SYxODl+clo/bmU1b2ROm2RVkJIlC0VS2GwJIrImkIuxBHKcp8OVuC
OUaQZmSBbVBn9zdHoTVSJnrMac2wjeya8PWbo6xLIIuQu2UobvcmLnovITty3F1gBuCCEyv6LAx3
kHWqsBQSdNQbLpE43cYxkctGTJJxC/g2QqmF20Ex9L44S8yA3YjqFXRmm23WIO/zQsiIsJdYZV3L
iM8ipMhCLa22xk5aI7QQyCOsBDS2p5BnQYyWmpYYjuwkPn9xOdxdKcg167qR+XSk8ntRqrT2/BG0
LwaFcCXkqGtn+VIwUR2FU86/9ZI3n7PfHbwEytVj6Y74QBJEqQpzW70e3UUtr4nxM9Apcyc/2zcZ
lfve7tv7SFuFlFkZbtLYCAbfVsV73UGgos31IktzfwFIqlT1lrWCyyMZgKNYKIIB2a+9nUz5tIgS
1IpCDPdXT4DTpMjkF09IFxYseA1PZGryoHVuR3CgQ8bfBNY0fjeh8Z/uqJ6Fk0r0J0QCsXjC86xm
x2XkJkGNsycWLq/G4Kpmob6qH8Lpt9598g4zenkSAvKj1R270MRgh1SQQe1BOcZ5HWZLR5imwSi9
Z02yBE2+zfFYgMw/xkfsy8AFURNwwrC08nAO4qH7fuBP493pXsKWFa1hMlSPBfHOiPqvx1W8fLZz
yLOD4qF2FbANMOTIplMluqjoeSiIx7lOpGY89SLCRB54ruWxMMkRL3bwC+96mzMvEUJCK3YtZunD
KYubvJXNPbjluSPFR+QCLElWVOeRUEbQmyughsAbQJNzQGjbJye3xVI2RC125fxh6jc2pt7NhdpX
SVNzvaVSFnZxDv1Q1ZyCwrhxpkAYUB3ljIX3X/2ubJN/WzTxfcbf796AnkkPMYPPPYl6pYITIPGT
wKHOrPqgyVLtZKu6uC22SoHd73VuezQOip35FvoeoQVoX6kFcnXje/Zh88aYghMK/iM2y/g4VcBf
dfsmkSnZy/hWr4t35me/MRSWCRxk0MuH3sVOQKbupB50tarQI3eoLkhJBVlGfSUT+zu7dI+4bh+s
/PCX+xdOwsO2D3capcotYzaw81ghD/lt8Be5YVOZYopHf49CUtmrgMZcaJS4TLnE9CqlZLGaXoMK
bZ28RYiqhuD5KLqqUsg4Ecdi63boMeqUprP3wm/P4JZ63xUPGGw2ypwjxtru97HJn/DcmTSoF1da
Sw+o899zsgVvjmQAGhST+KMwFvhimP4cI5f+TBvAvpycRW+TFfYM4QDdY0RoPLF8qazFrGq9mlr1
bABf6MS8WDcNwS7o3eIcq1AbvAs2eTbKfJxrJbZ8z6WnQle9BE3qhviqvdCijwxGTaHIBuNK75Qz
QK/24oBL30+6c+Oi8ejU4yxDgY0qZRMagC8HC5a2Dm24KJBW0v3qJImR0mRPDydU9gwvEySRKuAT
0Ve1PikSlckrq06z2Xm0CVtQBsBM2zEOpP2ziCOugYQyYe7syoOFzu12gQ63/S0F+9uQhCPsYzzO
kg2Abay6K0/Wkm7yoxTBtWwohdXuYNvb3cg6T5xfjPXuH0ZJBT/Pif0Jr2LouaaW9jvKd7Bb7ZZd
Noj1y8m/DctoWlx/vtZ77vxpuaVffyfZfLIMC1QTaOXEeMR4s9On6w9zL2JPCsFhHZcTBMQSeJIE
p0FfjVz1em9MZ0SdbSDZTHJomXoB30T/5CzmUVDNzOtq7BE9XZSGuGDPpG4ZuaEAS/ROvQ32QEwS
gxQfM99VgO0+nZVYpjTMJUiqvsKeOn+WUdFywualEj7p03PY+EbcEXmMaPZr6kXOFUjdzMq0qrw4
WO2Fe9w3m0GU/zasX+U0FXA7SJIBYY67+8O+y7X3xj+CkJ1/p32n2HWMZ+7VBeg/hfR6fxnf4+EK
MNUFe1nP4sJ4J8AsGl/rjakFoakHr0kNO/rPTGieha9lokwwQYkUWn/J8RiwxxrvYIQMH6xXPkp/
te2JTNiJTDDgS3yQkJ9xcc2dOd6OgYXPdzZM0tEl8knpVR4vwCP1NvOD7ES80IK9/3Yw4ltbe7Y2
kI10zC8r2mr02wTaSjSg8Itck/T1SzerxNbBqcDX2QAPYBXPH6ueOAPXZhn6iYiuUfqpFDB3fLmW
DXF6fVAKXSBR+RVbTiJzFe4o1GnHhlHHhCRv37+eWpogWwMuEYIsd09ZVIxYu0agDaU7MWyQfnIY
3ZbYeTyE4vjwr+K7xJJ4E+TE0Au5Lyugfp9BAmHylkodNbJA2tvqlFfdS1TUo7Ufe8znj3KIMOLN
wWlLDQS7m2BeZeHUhKppUGwwXjCA7TnWmlbnPbyTur80NlDZ1KRNwGce90l3EzbVEaITDB/kXJYP
rT40Sued1qBlyGBj7AjIuq6XNZym3CVILSNknq6VdHoShfOs4lmhdnzGGhthkBZAQPMjtRakJ9sV
L6+9q8cb63p5f80NyKdYyJ9MACWYxcDJJEt+C5xYQaqggyTbE6+a41yxnq4snDKpsKGKUxCDYu4w
4SBoQj64LpLyahaSuaEooXtGvz9d605VZS33HfKujEg1WTyY27vYHedEy2u7RkrSp0lnt4UkQC93
mYWmt4xhhm++9cNK9kffUi74kFwuCPL5rVmUBXxFF1SkVLABEgypAl73w5VGflVCm0W/2xw3WqI8
SvvMQAyvpVTTqu2KXsbRQQNFKiaHSV4jgTziLX7QGRIs79rIFEtSAWabEvOmsCypOK9LjlZe3C9u
UjixjCG3uQs1QWFrY9bX8uzoHSKSCsxABFCRn5NfEZVViKCOl/RKS2euUL22ziKnGbNAjGvqs3W1
ur/6+QDVbot/0AW2Og0o3i8mG3NZ649GNkb7wLsMBbA3olgFRmHEKkLUzxvvi02H2q0FS5EDJQIh
uv7zsMDtuDXnI273JZkqRUVQ57ZXEwEF1JZReX2xwtp2qIDJXPwCOiGtYJsAEoCJjYwGVkXY4VWd
ceIN9kkgz7Rgu4P5T6/uSf9Mllhj1+62dw8nZ+gNlu1SNIIxBe2+r1W3/ULmr64nyBAIa/btfXfK
oaybrgnTOidKzwvTAGgcdR/84tcW1ak2SC70FpiWs15+liMoXyHuDsSFSwuMkgYUDqMMS92Eoixe
NUYrXRPkfQq2EJBVPcT3muJ6HYv771k3hKKRJtmX2X31npek9yQTfejebgEBzZ4In+bqWINp/PsZ
/A3Ub8MatpwcbnoJgxLz1vXAUKi255SXrNGuPOUjatL/vcDELDUlZhK6sITEsfdWD4TdyDDGw+eB
QXoskeOfE88uY08VNKFBJecxVsdoHAxN4/rY+X01GVsazhjcsdFsQOYWnuuC9w7fD3AFeuhL604V
faV2s8spQKUxODQ4BBj7ssCTOhd0O+3bcTCWWDt2UPfPri4Z3T7ISwwaJU0jgmqpcFTKRIU8eUY5
wU5jllwDfJj2N7G55Jk1OJbwM+LqqjKS/iPeNoUZkfLEqG22l5H0kbr2FGAFc9XYL99T9HXBhELa
7D9y5+7OrAP+D66E/8q8+BO0OAV6C4+dDY605scHhiDrLEue5o9Zk0KVHpabbLXYHTFEdQABcS09
1Bha2p3e00ZvIvik3gFbX2xrolie81Vq4FuRZqFd2aYEm3lCI6yzqejQIIo46nLwAV9jeOVQAY0j
n3Xd62C50RsG05DVdc6kGqsgbqF8PpVRGRD7A/6sTN7B7g7DShhrv9QQE9ra5I3PbR92xip9d5zy
nJ+R5BBAjep7hPoKYmNzVZEShWQ1pltrRFbN4eJeaUVbA7QbVu1sejAxJU8nhmK3D4sat+mrJPZr
af06GnwLG1I+tbjMPbaCmuboEiWwn0JiG/Vbe1Ip35l4jVYzcOegb5otAKfLCaNLVBpFB4bPYer2
nIAN5HPT5PFe1AbEFLcf0sJ1d42gcFNlDH1SUErvqxPjDkMOdqlDArA9qbHyrVRzU/snofgPV6Uv
GZwswpSPpdIhrJcoZrF1tBRL0Hz0NPIup+LA1v9S2Gs9XSVILe0dEQNnO06woFVdgNEWcIGU9uGe
gYXMkgNcyb1cZ34L/XLCFJLZwa6ahZqbA/M7blMQPKJ5ONKhW69+WHVr+wl8hZyZwv6Wm41TSsl4
wiCIyeqp92fPQkjx1q948S2WUL7JnzUxqPl2xdJes+nPJ6lJ7a1N1f55MbpNcca6jtsJ8d0avbwx
ZtY/e6VNwsEe3LAsxf7Y/CQ0zXGsJFiRCtKuYsrRG+OmqGot3KtzCaFQsvRlL6fphLFEZ53h48q/
qJiQ19P/kC81IufG8jBUsdwkzgRARWetIfWm8JmdJ4zmhCgeGTKRoSs5IPBByBxxiEg4hcFa5eUU
a2MTme3oiW0lcIX0BPPOJgT7cdXC5kxDOKaHFmFjRJXWH+HwBNTyV/ti64NVdcCY5SYitHoSXqxq
d4vb2MqVnAL2hYQEBqwgccrXLTzijzF0bmrbJMLt/MW79kQ/Rgm0P3Y28VM8bYVK+0b2JXHDYNl4
tmTzi+UhhDLWYaE3/yu19e6nerOvgW7+RpD3yHmhEkb6aYfozVIk/m92E8S5EEp19VHcHzR70HfI
m7xcvNbT6stdLaLdQfc66gj8+NVg68bAA5TlU84T9ewTyVfo8aNqMHpsX942VA81GWO88j8MVLF5
+9wrt7zxV4QANug1EnzTF/OK8rkvzktXa7qdEkNwR70/ig0UVzbSMZ9aBDER4Eg61SCWLhMSJleI
K/sz48zJN8u9S14owoqCrQ6XvZbpORxph4GM2k+K2AfmEnAtFSgcs0VwD7fOKIYx8q0VgVuAfyQB
HF+VtNCIpxzB5X2HcVInGu/yU/L5djhGpZoq5g5uthkKSuoYTYT9Ye1zKrMnv303URFo5wkLr0UA
Sr3kfGG0SN7mpgf8zdnfUPmzXLxxDFq6XRJlG0ri/3dwHmhsEEZty7796ve0LynH//U1F4QUTwuP
NXx0T+o9KVYzThH442C0UWeP7fi1w0TNP50b63LFoHaIYMjgwrI15v+il9AZVfV7G/MV90R0uqnM
JhrdOiZORnrK5DAJvKw0BqINPm1nZiLYoVKU0F0B/NvwOxDpqHjM3f+5MPl6c/cvLv/5L/RP5TSH
9oVkgDeJdWJuukwCqI70HcyTo7CJeqWB1niyZjqVPE41YhwrZcqIz0Ht95zstbEJsMU3qJ9W4taf
QPxOmkYwIbSjAuGNyItfjKSoPrhEacH7y5Ah0TpODoSjMjqiuAfUoTxxOqWjFwwJOfVlD2q1TmLH
OHiunOjmBQUxHj6vE3ZfgDko60ZoZ/Mm1j1eeh5SP783cU21Rp0mNU+hkxYkBPsl1Ey1PCdR6PBm
oZtonSBz0JnCYJCDaOjP+KnsjYqIJzyK3k/rEDqTIf3HtNL1GG/atHAJekhtCfK2XtispQPZO5WV
kCHHCc/CasyEvwfXMy7OCqwlrGuxAcBkmK1WbJqPLwrrwRpzQR6kxhWw1RbV60a+io4FBkrnptTg
lmeOxrdMw2fYnqIRZXPY+inoQeikPH9qOH6jub4jFsku9dqSu5FgHKx0TCFUKEZ0dcD+gs/yN/BV
OGWYcxTxYOkHXFUGJHPiO53yzbIckXxIrvh6/m8BosHf9sdcZue0nsny16Q+U4bRV84K7RMtPc63
E0F02IRP4V28TXggvye6Pwzw0E+bZDAQjBRIi/am0AemfH7V0aWu7gmmm02mwTkU3G25eZJqE4Sx
TLvRzHCSYlyvwoRnSnxN8nZodiGGQsqRnkh+hRKwAB7WGqfwfsE9UyrH+rwczZpdpc2nitV0TWJj
jXFui1KimekiO89wrCAhzbqyQUF4PH4HVbjC7gDKFP9AYmG5KhxKgbt/+OdKprqFgYGyTgJNHLGj
hrNtMvxY2vzops/onFqAduWPPpvENE/A6TBmMCrLbmdJcUSjRvnMzvVKJq3IsOdiEDd1cOGQJ3Ge
80MI17LEW8dWpn6lTsUHaumUJudOLVopWFtvokthAaKun+WAfCKKYhY3DbgcqzLLbNAGYlVkXlcr
2x6CNrPwyzuZnkwiVbz2/dAxkVu0Zt2PrBkrrjg4NBCuwAVsRnaasdAljCx0WDsIMukHSRMHr/05
K1PYp2IxTZ+s/1XUeDwDsYYal9amixFszfmrONP0jdH5UGsuEWRa3SFHuFFF7+euTE2fMH+dQoDQ
gYmQ57KdPZFyREUDSP/gfG7j1OsFmLzLEMf30kVFmrV+55aJUgeC5M2BwpVSmSlMUMme+9xLZC3D
+coAZAdQBun3HJaHZToQ15XwCcnxh8j1lq71X/tl6j5xKi6QFP6Scwnm+P5iGIyfTOH7eL+9kN4W
iOpalcv0bt/pI3jwNoHm3CEgUmT4yUnhhOlkzgU3NfMCv59fxsKtX6crnawdr5kKwdBRRNGtN02c
JvwxP2xT9oRyK2bQ9TCHX3mcwM4+l6OxFWXGzBxCx6OGOBfK0frGQFMCInYnOqW6cTXmFfHiw/dg
1rITAJKJrCRbOFV7ghislW5kBfQUojTmB1ah+s/pnRkO2R+x6UnXG/8BKVGYZ4MCUnzUy4NJfsfH
AdBUMOnOD/6Oq7sbNz1VAieLsSNbuVX+4RUinnWRZKOgTzXamCTe0pvB+iAtDMzx5OB+UQ27z5lX
DaEVFq7VtNUgHGAlEizf53UAJTqz0FaOtWhD6sOU1mSfhDTeNdGTy7keQcNh3CIcaWvcYlMzhkeG
RGHSimW+NDwa61QjxgTnJoBxeQwklThPstLraWYCf/czra+efc2OhrdtInpzu0TbYul1tZOHg31W
8vVtQOwbJtEoTnqQeTB04E+HnAENUcYawfsrNT0AAjCule8G+QRHz7kulTpuc3BDNeu1VMUx9HWV
wrpjid/O8lz62wOb6xaH1Ajwy1M5HXsJjyRUXfWIHmmsWu7ljgSQgBRUaXEj71V6kwLYPTAxBapr
m+AHJy7bdcAIR4HXq/X5js6ET4LPRduDH/eW3QQW78aYMqbSp6btZvupPSbGbAzAggVCBRmKzYQE
LhdURMQ9vyNQuxPslsuaYMHDEUjsrxjLloiSJ0dEGYDfr/HAshZBAc1rQnV38sIqJ9+BhmVLpGrb
Z54Iwyy3PTWSeMMJPnCfEuulKdKrU945RsVL1iWcaAehRagoYCpottpiIH3MkA6eOeQRjBFXtaGe
YbnISYQ1eh0pftoKdCE5PaTAAPI3zUimgP3BEGDNJ5/moYuic0wEB+LkruzCeo9qH6cV2KZ8aR1T
0eVAAsYes+GjnOdW1PdMADdXnt3PASTdNnBgTcTHxwbhcDu/tbKTwIiGpFc+STfz1uZcGmVILMBQ
R3mGDS/m978ucPcsFCUe1vqzrQuYomQoIDexwF2g07wkK2K/edFFn0D6232odqQ0whLarX+VD7sq
gHPspOD0hnzdIjBz2RKEcPhLnGk5L7A9lWUz9vNPvieI5fQBstBxWsVgCYaBUttK/YTLk9lCVD3t
jSlNSbwwCuDZN3bxC8JNLTy69L76KNEWmVo/RSZfPX6+Ej5s0WYJPneJmEP21++sNenmvpVRUAFB
51EUICt4U/v/3jEhH4ldrzw9yi4h2GMBbUKRFZZuwv/e+QLptDiY902apY+hPVSJJoHIhisJMPuf
E5Llxcg7nXt3iT6QsBjd75TMnakqKqHqF5U6VsdjUSjTkDdI1mYDT9d0XsqlFSeDIuGDg3sntSA6
xHaw7KuK25WoC9bZ96Fh9G00ydNCZe6LLE9++gOFzXrTYxZhh/TpAg88bSGpYPo9bjwT1LA/gY6u
gdP5kITEBHf9fMV+5YKTmAkj5IWWmw0llm/4G8qxJ3M2mqihu7p2sZb+aPh3/u9kN86DXnfUMkrO
sYIoJCmfDIg9CAfLIqpGc+hSuIbvnxFyTUg69O/DHqPq2spipFmkwdY/scwevRl+fyq663HSBIa9
dDDbX3EPJu3qKANfZV+6E3TgzZ2c8xhHjJtHX/ECPGGjE0VHi5dSXV2sjUOm9QfHJZwyUyaYPW2g
lE+Y+kr36TQysnmImEH/CGsVxVTSE7InSNrzda2upTXi2aI06ru+g3YtAAWOqbJMYmWPCucf8Bk3
/fLj5H7r7Gwm0ht5F0Ufqui4X550aE65oxuSYUhrxFAN720bWgX0c09vuSW3r8T3svoctUtnCmL+
Q69IbDzlyQMypUIG3vjuc5Yz4VqHmKFJ/PmMjyC6qGxlQ2yc0tqxgMtMQnQdp3VWl+adQxVBUvFD
mWRYY2pE3tlFMA/HjD7I5heKTfgPpTnM+/CsuwhJ/GqNokIpt33qYmaZVkwpX+jl/R9lrsq1WlfC
gnOalhiLtMU/UyBGtp5SzgggrIdktfiPwAbL5AdskHvo6GB+jntMqsnaozwhsFpVloaaGj7i1SMI
2DzkiRx09rXHYjUfPNF0BRUmU6s7JyX8WF9/a8UFOX2LDbmWqNTkVhO8wTtTL6ATfE281fmEatgK
KAgoouTl/yktuSgbdm9MkE+dEBpHqo2DhSxbFAi+KReuYFJ5TbQAKgsPBq1r7/Fzv06fCHACUlU3
dP9oMT+MGpeDMNEISzlhXjs3rA58naXqbXDdQ8nCEvvsaggtMGNV9r0ZTyRhXnZUgGHnqKgiXu+J
7iqwe42JKkBHoIdqEF1WPA8eMBIrRnBsqfDPhoSadRV/bwtpYRO6owGUkqzntQnGOczQErtIMUz0
x7oaTWFNjZ33Q54DQfV24OSAMkKNVLxN7Neex48GHuuV3Zq9ZBk4hjV8Nup0KHbGOwZNQm8Lz+3k
EIGUsU0GnMGiR5Ipt1Qyx8+D+9KXHaQ/KiJJPCg+R714+qNtIXiXQRN/tj6ywDRqBXHUqo+vExqs
4iPTSFZmzLHjE4n7tPJSBzBBY2NCBYCcKQhW1guNmVkw845ZgT/1tas6uzoTxXsrtRwFl2khvGfM
LcjkCm/ahHupgULa2fRd+l9hDfD0qxG1zmFrKBtepxCXtjQzkV22P2nnSjoIhw6Z6WY7WrTJtPHg
zSfXCo9HNKva/Rlm5inA8k1rIhaZIhdweI5mOKgwrZgkeOAOG8mpxnE42Ul/E8nsMeRpzUoc9yaP
FZAhc1jwkQLkzILNp6KegBnFMAydps63Pl+jw7UEJzK9G+ljT2vvR1Jcc+t5FNY30jZ8xAQt47j+
pF3HvHtcV+GDUf+p6YNKlXMvfUXvPsutbWbjVa7imogt2/yYtFsN01CYWjpcHNdPFZFSwoHA0snI
MQN8ZXO7yT5pFX3qAG7L9qeXbkfcSQ5M6kTU9k3tynmI9O/uB77Si+RMNc72fXIB5wZni6LLMW0+
bj5mUKzmAgMgM41vxFszxzb1AQRVnK4pX/IqY+gJLZgEJldbUwp1wz+xtI4d5ySTCaoMP1mg7mBn
6rPfV4lSr2FOrBOoiR/wn38B3shVbWRqHFr9E++4h9JOxdOhRq2Jvc4Wlko9Sdc2pgHA6bFfWiMP
+roC8kCB3Qzg1yuQJwtgb+AYWLc8VGk5Ex3EOWamsxG3Nh2WNDQeMT3lAZ3E1mlV4Ha975e2OEvW
r4q+/lkBI6cDxh3JTJQeCD+cAR9Xj+3InZj/6HjCsaPEAU+apNZ2BXYqF6yE8tgkJzXewDpJmK/t
5fvt15/YloTuTUV06C2KZib8KMvYxSc9PVYjKvBVIXLGdZLkt7240H//Teltv5GFgncN7DsObdz5
3M0EHg9vvHsTG9MihnQjjGVSIKUNqJgOa35N6HOayjIRB38iu7z8+Moq4mn3afjGJ9qay1ZIvoFa
+e2dhYbOE6/iCRjVOoCTHzimQCuWu/o7uRZD3HQIHvvo+Xlx65KmM8kIvqpQwQ50fAqZAVEpF5uo
c1UMTaZR3gswz0nkyV1ibnkjFquf7CQf1JmL8FoaV9V5fTHBUm/a29fRpWMnRVxgZ2M/6cgf1FAM
JPutfGJprAob3/pdrhsaIY2bvQj9cwvZC+z0tR+FvjOFptLuYOGKIpKy9DreJ8VC86DyMlSTl2sE
9LrQn0zB3LV9m3Gy8koil5ZQoOeiLtmQpU2kwDEzso601LibpC6hZtkDN04Zx4zQQBb10Xhy6Hgk
NtI7JGW6jMarqulmPLWcncdrDltTxHRjt+kmTA1+n+XHG6avK3tgW7pHZ7oyg7Y5VU5LjO4GfiUG
uXU6iG3J0XVw1yUEVx+3vJw0VNo22jqH4HPWln5h3SpFOHCeXUdhV5O73koTY81eKxAIa4Wb0fLA
2wTmW/Xjapd21ptIo0mE5ke7bXW8Bsp7/XDQvCtvk3IzvYzemFbGHiEkwFOCZpWsHGjIqZ/ORvD2
n5nEq6Dhx/04UroUvK+FzqC63+FK1pT75cbIsv3T7M5/ksviveovR5WfQ9GXgzuss7+HoNg+p61n
zdhxqsx0AokZUSckmYmh7Yvsy4aJ3/TYLEm3/XjcvgdD1JZylv2lZ09ste7wszdT2j+nKV8YLt4d
d87ujlWolAbwkJVTH/YgZNLTAX6eN9o2tcevMhT6bAqMEpi/T1fOT8t/k+wTK/veEwpt3ZEZPhvY
DfNHPKZzLqiuZsNf2dq569Z/nuDGgfkdtv+jP310kFApZj0tsd/mRPdUIVWS466lsGV2800NDo0p
M8Din+v4ye0eNXv0yhUDd2FdVLNjO9VvnDgaMTx0A0RrBYqsTTmfM+dcW0wKmbgp6doBlrNRGR7f
T1B0FMHY+i/HM66mHAfJCYAPQveQJatuVfDj9WYxjIusjW8yTmKl2Nrsk92QneLveUHCOIHf54WO
H4rFwcfYXhEAlDhQwrzaQdztFW6lJQu0jxw5Q5uFEmoNoOJqva8v9JwU023JvvSt8CC+cF0r1igN
wl+MCocWSd5Pno1viBb4cjF6TvP2VoQi5xUPbHi5q+998VAaSUJCweJcfhK7//xebzXKD0LC30yL
skXQtvlXOfMf8/PI0hJj2mfDljvUpWrk5gmuro12A2gCGXpDWHcGziZsGAyagXBtGu43VRoMuYh0
5+/ONUCQXrGeL/mZLGS50aPKj+55A+g2RW7rRitP/w7tY2nDNqBP21jOTR0sgL3c9WqHeW9ow/dr
81quqI1+gCrNy/cgWGWRVQP8XmB3pnhbaDf1ADZmwyWaKhEsGds4ic59GEYmEzFEbKevfVctSXHb
l2dPn587jd92ZqvdBnGs/QVNfGtOOGyetT/AUgQeD3IwB4SeVXbu2gk5Y4xWMT9hARtZobXSWao1
d9WZI0OsQCc04RYTvhUIpOJr6DZX+rXp7Z9s4tKqHYvYlRYL/mIHK+2CY8k0uHvK+NYPywvKOEwm
RmB3R/I7VIetSaxbZmfm9FvZHpKYAMGQCBggCb4C4VzkE7+LvAGqH87XxBkpEo+p6WuVuaq7MzAD
csTojYrI7mhuouW8JxRbB7XEaKCzDxwGnymd27t/UFwX4Tj6yjaF4G+iq0O/Mzl0+GeLKBfNMaUq
OsE7lRyC8I55e4hCYhJ9CDG3O+13tdz9z0VL+LEIiBiodoBagH7GwBpgYoX3CTMSBaK4A59htnYv
lDUtfg3npCyyQcjanabPF6d/9y7/ZJRHHVizW6sjC9IGejns4izSETpWlslTiaaqWNhnvxyJlXKV
Vzo2gJuRRbAiJ1u6788HvvhCv6xvR/d60/leyaOf6ItHZNg6DwNc6BpQA4Wjfpnwj9DRuTLxkoEw
4Nuu/20f66E6plkkEAFTZIAjcIRqemFsUzkOA3uaVLSfrNsrIMxgBFD9xdwNiqATFYE8FKw0S7E3
MyScdJ6RxXFRaP2qfrH2gH4SjyNP/v1YVfsDpMfeh/dSV3Sn5TVD1TA9HXnOCCzUbzKhczDNsZIX
YjbBKiTj+CtzcUzx7p+GsIo/zBGkEke1K1qsm0iBhkEHytairmPeAltXHsCLTjjZSKfcCKNHvEyL
kpMzk5B0jCkpvmEGEXlm4fglUih/Hfj+CB6+1wnOiGZD5/UD4VIxJF31mBpfTPoiXJmotOOB7oER
KwylxbEcauYs+I8lxkNOldJGrKhEWHEUop74KigqSl/7ns0RWNhz/nWwrkBwTMU/YkxGcGYNmv/i
WCyrBYgdo28HESU76Lz7Lfopgm9dkib2t2TJmJ/L3i+pHF/EyikdQejuoYogjwec4uirE6ZWFqcv
BgzDtDagomavUViXYXSgjrNdLHcY74lCAH56NrHRCBhsUjcjdKTLcaGnPnU967+xq/Ao8024lfW5
Ckt8KrEXEDq1v2MpiEOOa4gS3n8Ndet4LEF/CxG+VSOvso/7lqUgssErU1U2Ff2JVhFYKKT0aDjJ
/gqlNHd7o9/KT9eWk24OX7S4PFFH1/Ij636Sn9HbudPRyPeQSRvfmNWpqNrsHaWgcatPaBzKbQzJ
a7JCQiQZSE8NfK4myZ78Dc3fxRDzehg0sJwpFz4oCe8yi0HFwcBkBY5ev4ZdNJqJqbHSaWFTEBjx
NEaRMgPmZsC23VJuUQaX0pPpIBfC+dGQ3QfXYStHJwVONPeY+MjGnrb9vNlQfYKTAdu3IbGNRxg1
/5IiXXTYyd/QbsX+VW8GhDjLp5BfYSl3M7MqHq8l4ZZjJZdZVYGJXvVtsxe68S7CJSHnGk7s4FfO
VJE7pubBUXQmFO+Ohvj1Ll+FODqejTEWvkkVBZy6XzXrr7WkulIEY94KIfc1GTKB2lADE8GyOpCS
7ofloCsHvN9am+AvdzBDW3kjzvKDvCbWQA1jv1coIheUd4nVge8pHgNgwzfBKEnlc5aj/x573Si6
MbL3XYeu90OwWT9jprRAEuWKBd450BXD65Gn/fpfm0Vxtn4wTXRSJ0UmjEuHKcRNhOzbABwyv1v8
qx9tXwX/rw6cVNjaER14q7yqw6YEoq3dQpLl/8sanX+/h10JulsQs9Bzhv7PEwnXM7t/Sg8u4LoJ
/LQ4w1e7b8fZEnIbSjhQcr8N0lo01TEacfx98PvQYgsSSgpd74skK9QN5rChQzn1d7bXcgOth22a
egliSwQzsi5stxqCJHMxH2yDbgKE32YwziCDY2WKi/dJDHHdhNp+qdMRNfIj4GRgd/9A0i5aCPvu
lDvefvrHT0W5YqCKTodgECvIGFanJAnet+0YUywkSaFXLCqIe45RJZBEH6uYfNkued6wb9q45chs
5kIu5jovtRvc5fejy71IXiQKYMK0+rmlRSxkUKlLTvcnyFDO84ewpIn5nkvC/ptS/uDOqTZjiCNi
cus4nGqVUjyAaMyhrcjchSfSF3Y8fnidr9Xb4pVDzLGbDuc7l7ar7+3l9K7aqvUZDAFlBIMacHeq
mVnf1K6wwSccRGc+GedyQPgM6xm3Yw/3KzWZhBfqWL12cAr7UgPkLXpcRMmxHqb06Dc0tZewZBkd
DiOdTDNzk8E5DQ4N9liaj4S45Yduu2h32mm+XP+2wYgdn67zP270k+cdSdgTIx4aslxpaBrCPdrF
GsqTIQYLZ4jVclZqb9wQlrC6oLY3iye+btHoM+jPUF59n6KgRrZDX5FEe6Zt6/pQBEH+QHCAyHJD
bI9S3t7aCMQJP1Q4w1EYcO4Jwt0no+nYxCDF4hftMBT/T/WGDGPieMCuGXxpwWpgSg5YllrXKHj+
1UnIawedV5pslmTgRGaUmdouNasigYCro+veerBrtXySJ9v9EWkdRg2jh1LmBJtdIbWRjMBswuyQ
548B9/6c0ua/5EY3+xHsg9Uua/gSJkp4ukrSmM9CC+IlBmPq/hkUjpdcoW4ZbODgOaA7mQ8ijyxZ
DaSnLKjfEd88QzN+oihD08LfebGisQkNIMfaAgaoQ5N6eoloZQvyF/7QUK1htYLkTozR0sqZ7aMq
HjMKsDxjwsdle3iDIQgwmi59zf+szOKNAEq1fe0lz/K4BCvBEzfYQu/qHXrR8hcoDrpsjsURLskw
nP0ZJtdpu9Hrx/HwRgpH9ZivHdcHYm+cDfCHv0wl9H9fDcylzPtzTz2hXGunW/ctZjS/vlY4m3l8
c2oV61IPB8Uecjs/AV9ybuWSFI9IYhtE8Y+ukOJRV1IdppNixFIT264iVcsV27EHLPed6XuNKJ0V
y3HnXWV9Pb8gQiYer3qLEAIhgPuujMkyX8ViZtdCfLlRJIMB4FoNrGZ+dDs+vZKA/HuapMZP9/Hm
FxLevZOnv91qolwhWcKzkRATzL3M0c54pqIPx1Cfp/UaEL7SKQh5YV1noS5Bz7TNV7EVYbqXi5Mb
clS9spmFImug0X3ZXAWptTJu8v3WaeG9bEmej34Y7H9hdnXCYqsXgBhTkDjr43YrLV57UVELNuv1
SU1FaHFQaz/93UyMiJvMJeC7mWsrJX2ZG681b93uxiJgQtzmu+BJT7Xx/jHciJ+ixh7eu9o3FwcH
JOvDbqGXAmn9p/et1SwhArZ7kvpAMaUQIK6UXX+iovJL22JodxyeiDcr3NidH1RqtrWcVALC9yKI
oOf/KclOm27Hbhc/o4WV0b5cqjla00sOweWT1SZNmsSVKmx/BtS2e2afLxsR+gEZd3RVwzP7Q9Cy
5A1l6iRkqTTPNme0agJp7f1EbR4iwgz1uVBE6stpLes3PSUNc4Vw3BElx2bprQlIPrwRKMtr6aXI
US8ES8TxRbt5jlfakdIzjkg6a90nyErmDqvb7iLckxvTSKpHdxqxU4vlrfMFFgI0FN5GPecV+vdM
DwfrPTj21AxEdZXbin9ZILGsygvvJgPAveU4+dzPC1hzQrC6+wLsEyrDWEZA78tcCCsvOJFetB5I
6y2MBDAwjM2tIQKMHezFtwwh9DTdidENoHNeOpiN1gIJJmZtaKVca0nk+yc8h1kDaQdXpvfVgvim
g8rCblPZbNH9ZP7pXaDCSXBPJ+P0b0uGJwfrRwxVvk1znmsxs/cCFH026C/eJdsHWCgJ5f6L6thQ
ly4O7j41qi3wX9JlSZYwms3F+8l8a8KlBFdo6gDKuds3RqEIWcV8BWihHECqdVIGjU9Te3jWdqAY
+p6HfaF0IuZliavsZsQi9QZ//6/WgCPI7rHMlBRGj4HlKvFzlQm+ygqOSfiLeWf+F5gtEXiNWHLO
mf4xiRjlCqWAtT4svwOB9qthdKk1Mlqz38tsTZzkdUuU9x+n86KYV4bOfP02a3fxVTd8hL+p+WKA
WHcl+wFtqaZkYIFGFQW9wa4kYtAUjksl3MK/ugG7rwqZbtx+NiumFEB8eMA+c73/h6wj6jMDlJCj
R+w63NEXHscT9cjKofqU032DH9bY5St6L5X5zgGL+uIR/Qov0kH+HV3N6ljGRekWPhtCUqEoaBq0
xpmWltJ3pFNcfOk7bAAqpnPTjh2IRtFQ7E2StmszHC/hWuuG6RzWX+Ge6aToTHYqaGaka9m7zQND
3j8PDwx/V/JDL6BKIOWTcNXKZRqC4WNFQqW7BFjzBS0+77wVFgLn1XpUtRhzVP6GopAot6BKzaZY
qCyh8MHlZMKATBHfum/OSHavVQ5tz9KzvC0i3VGAkg0151DAqSBwJfxikIAk8Vs9AyuIFU/PyW/p
OiYV0EeNSNYsGOEvnnMydkOgqYiOzULdXvroAGo/YxOBPpV7S2PyIX/DId5AtpFae8Rz3ZrAFnRZ
BzyaKVJ0y4zghiebAyQtRoNRg5/OGcxsvDKqiD6nEmajXNM/WY2hvGvUarHdH8Pt+c55hRKDeUrp
E4HDhwWhxPvwkH26twKR8CQUQ7vj/fygbGTYQ0nqYtZA05iVJ6kIexSljZ9FZXxcund2JRrV+51L
Rnz0AC/3xYspGoqflwhXMywhOWZEcUQ3GFPFR/w/eJhZuJqPYwfKBuKG9tE+fmcgFFf7gxhoJ+HL
xUNXiyk7EcScgkWEwK9hY1b6fE2ZhlGPOjrSeV3q/8rr/ITjIZpDWr04gWFm016qja2Z8+1si5y9
LNazkseXOl4kQpIAUYOvobvAnf03QOWzlT5uwRhtn/7Wvo2Vw64zrLhiAw1MVa/aUwcz3q/dWXq4
mR0E+49w6Ymzp2Y0XSUpmJo0ehNYsx1vBMWggYbmlf8YH9vbNRjBeTvkB5xRs65+U2HMUY+3U6wL
9SXEtkIFt64v8OmR8nDDJ9y57ZeOafaIuu+NKOUeiijBP6XFhz3zzZMj1nY+fnU2bV+A74KjXMpA
StWppuWwkxWMirBVQ10XrHkCNnJyL5Qp+mg/v7lXSMhO3CREh0x71cVotAYtvTAA6PuSouiGw3Pa
77QnOyoEpHWrhe13Rz5CQpmJgj0lGN0PUHyp40dOeQSzL/Be8XUAVsih+vIQ/BcYshpPMsKgEo/1
FGIqa2ZNy98gsAC2EqOOTeU29Rm3YRcS7E01ppeksDlEdsNzEbJLklZ5NqX3y3/kSS3ToikS0Btd
BXZ25F5RVWxWIfGhqtAUzimLIRPzRY/1d51TEtpXH86hE9e0NQBT+GPsFc9UDIWJGbE1DZ29p7Iw
IZnxux0N6z6knCnj3H2JZbe0nHn5JbsbeOhyV+NPZjOiStQzPGyNXc+lN0lrveMup8PmwBsWxGXq
V1q2GEHyr0k/RIsx1rGQynSJN2EeJMidZsD5fbiTZaJm9Gauhnt0tfMZe6st/qjTQiBi/ZnWxliz
6eyxCkCOWqQwdwXdw5fGnDWILXZNrJskg8f4lAvCXaQj7DHJjMN5JBk4kjx3taSp60BT4zOdrqFZ
0Y0Ys5YAHMPdum3TQvU1qTVgKMIBUQNKE0PX8i0zydnpij3eboN9rV+lYOeEKpJyYdm7ctOFHo9/
GUwYoyuwKCRxO5MCH/cBWJ1wov+BoOuk5E0+8CiyTPsjU6v+J7hcEr6nA1r0x9yUOmO/cC2cNLNi
zEGHc9EraV1FCzwgWoA6xQkOi8srTj4gYxL4niIlWhRYTkHN9N27INZmD59KAYyh0NT6o6O/2tMi
VINwZpCAE+58cBxmGobge91NYKA95Pp0fXSudVvxOdLJT87n1S0IqBlR+3n03P8JTNwPCOrsr1zC
hceApMXI8OFNOsjox5QwXtp74BimRCFnSDvNHSEPEqRPYJe3okwyq+yK5UsNiPYlz8CVZRnUWn4+
F1xqjAtngRxLkJ5oIYHJWbmXPIinlx2XlT2tsOxSfrba2GPBTJ8VabDr75GM4wbQugXYQwD9+bpe
dEoyJS0RZybgX3uioqs8CyWUEqGGtwPnxycMwMPw0E+ZnSs9/rb+g0kjWeWLvrwOOHqe+G+qTPRn
0k3rXiVhgAi4OC6NuSp/ferFoFoJjPOO+CydRDI+F/yMnuasG0zXljLZV4PSzMUEYXvAOtgYV2Mb
es/joBRoufZUq85ryCr7AXnU8JAYX70HZKG8MyNYGruFpOdu3uf0tZofvnBcYhf354ZngYfOP0D1
DVDDZBWb+Tgp+f2P+L3C/JnjnkasKjnZqJKP/+JnmSzaJzAn+inf+C5FjOlAdTZ9LFx3TDU9PBlk
4ql111EMU7UfbMq4DnXWMkrVUfip4z1/Zgx6Am1BmSEuUaOwO++2DBal+xyEEP6P9bXzQ65fTIXI
uLSgxuzlaT9WLF3kfRzQu9hThJcWBYDAaaSc8oamV0lXOhG56V9LHe+tdz7xB/CCWj9dHRfOBdGg
seRp4DIKeTFhPWmo00i7A6ql3rVacZo/JlmzhtzJk6+vdVcC2rNB+sZsgu1l8QIc195IcnWssH18
iVbO2L698Hc9931dZoOsyzuXEoPULcH3s/1Yx2l3+/vPbOfqY3GzZwaPMZUjpEU4hriBMNLwllkg
bGgm5yNErNoBtuDsTklZARXb3MVzD1NSB7tw633+4WI+f9wxDwHYqwBxywaYgvB1wp7cE69Fgdu1
TJwicRTCW5WjbHec6kJZm2tF0ACnZx7U08yNH+A2RRruSNpRXIAek17tAD4Td9rwIqrx+B08a563
PN7EOC9XX67js6vPXYRN47XSeotQkIPc/IWKvfiMoXTb/ncEa0DfBv6j7967hOf/e97VsxGFQuID
a1bYFmNuzkJvy+Op+Y2Zoo+k3s3FCi6EMUdjhjevXTUjQ9Mxa3dtRhaD2RsjlHn1bcCxe1xSdGXe
mkttHrYE16AWz3AZ59Pe/h7cMx6RAzf29H1lzw4q+CDqxn+cd/KXVGWhRn4nAknePHXE+nTaRjRe
eO6KR8CAawZHEXzb6DvpzHxEAJkXLaSfZvsFR/fMV56ynTccJtxwtyiNtCG49VryRM3vX3jufPZo
EmZsJ6Un+yrFxxYkBNRhOk5HDiI1mH86jk+erVJ/eWDPFLAY++GJt+134o7zIsWr2CCjQOZLWwlH
VaSBaXNQ2hMIOomokeHkiegfqGS/lQIzcpGuntBJEPPXQ9/4qXBoC227nSHxO0/Ke58RTuNY/b8c
+kgSvE3mEfG/D7xCiIsVW9u1IgERl9JT28hylOA5qGAvlMTVn6vbuxWslV9F80W3scaXkxtxgrLu
chKZwduYETk7IquWYk8f3ISd5eqd7ApJKjg/myIJoBNdGepSIcxslYchqCqSo0Mk87A0YgVomDkp
cIFhJwO5z+Gswk2SAVXPmyaclA9pU4TcfF1BLyyW0peW3UaoKgbFOZW0xYfOnTGWUEUHbPK/uXT4
rm5/fCq1KGuSUIk7daKBJvrOSIpnyGQCbjFvrDKFSOIQEB//1oWhXkz24ILyftE1s0rr4w/VJX2+
JyEBtMXGiMzMPI1jDneLpO5jCtUb4vKbYVT06M+dN01GTqXWOk3m0q/JtoIE/4EwLbzOKXPFESU7
+1a9ZZp/pc86gRb3j/VfX6mLzw90Jmux8nMClCBpbcJ8Rpdb46cP9jQ9/8zOkbXEYCOD1mTG3T1q
Tn6di7erK5TzKmr0xvBnTZk9Yi+pqjKhnQrT7MxOTiiYCHHKI6m9a65E5yZnJ8GC1PrTzLdLnpE0
VqnbXiMdTqm0dXzVDcFNJwOpjOWosBvy4RbT9DJJetl5mYn+voZwf1WCekp1aVvYeX0VYk0CvSoY
xRJL2e9+NRVDc5weMGcJL5pIWmc89yzXh99fDqtOVU+vIUahAGGkw/0dJzc5XVhlKC5ZiWN5eGOO
1+Rkt7vEQaodD4ExEpc//NtrOgxwf/Vun9qO8/oJCy1VQw+QSrcomr60nld40+zmDWI5yxqiob/g
fwwBHhhQeIv59vaElV7oSjUYnDJnNWlY2Bp618/WFpUnZR36b/HYE3sEU8auVawtc1dhx5yV/e1u
wVdcrqKaY2Tc1pxs2imdmruVWIAeXl1ac6upIJWJSmsYmusxxkNst1LZihhA+BlAR0jvpFF4Rpob
7aBO12wsOXYGw6pa+qmlmv8HtQhi8Y0PS/m1qvX03EK5QVLCptjqFjKvlEnttQ3oiA7RWzlBh4/R
4n0Q1nMj1uwVV50asqRc8GPCh/FvlTvqU9WWn2UA1gJHxOySBK/TGiQ5v1g2rBPAqKEt2X2ZzRyr
7n5siINCvkmcoHDnlPN2emjTAp2y5qHCBgU6URLtbAcwmd30FDYYod+6octmowmFpWO6pw0L2oyn
30DQAYcypdVdFw5nlc0LFGDvCt888ASaM8a/zpLmLYSw+FNRG11/T5pGqBksyU+/qztjwKVM8kBz
M+n9gPUoE7DBH/RtWWl3jMb+8wRheVvy71xQkuyylD3u0n7OyASHycddcs3LdBA2aGowKSK0XQdw
YvVkovXtm+FYb52qiTD9jr9OdqWHLjdkKP6TO0v04eGz9PS4gnJw7v1GjTUPQ8Ts1GxI1CxD5UfE
CpuCaNoZBU3iRMeAzRgWJ/41edSgL/qWo7ubXuLyS0/ACwXj77QABaF5o+6p16frBrEeFzP0sgF5
fJt5ZLUzA7aZ9U3kDzF0fvzoQedOrtmZegq+/lTZEhvJ73tpP9btWh2kYLjpMSHf9K8DIfrFNutY
QTO3CI69yiciK7bkSfAK48L4Or4bfRnGQLSMytgEI5smK3pbN2SjsliY7IiX/M+TVmmE6XuiAbtf
/pYzs/4MVaUJSOnGobZ9/AYg7BTcmIoXVA/PjpzX8+BZpUgVdQTeiyZr9ZxZGEJEmodFAxpdnrO4
AAxfWnTIolaMuSL8TjGov2AXNhDSVEOQjD13x9eZOlh+qnywesctzQycXx6mKAi0D6MG6n6zQcyH
t9AwFO996IrB61NycMiWD2pLdSylb1lSu5nVzXUeYYtvH+Hv4knsfzm42dyjUda3jZPeSOUgb6qT
ybt/R1wykO+s2Pm9DQSOuv4yxd1wJFg99Q9mbJmuelEeJLcHHiBvOBQSa40cqsGiDKSE7kYmNZYs
um7DbJhF5CbXeUjiPET36r9frfiXJaqP7W2fXW6qMrKuRudks96e7/P2oU8RyI2N7KxwesF+61Ys
tqezypHll1O5QZorPB6CHvhPSDR/3fTFV1M2Cd3XVVHkC92nxL+TrixS0wZDbOsPYg99pCJvZ4nR
9f3Vxl7juA5Sf/3+cFoW1YnzeVHLUO2d2VUFsJ5Psbn2qUoRNjG4I7TDQ3fPCXWvOSXdGuPyc+4V
XDIXFrTSPM8pTizc8HJSlqllOvK6rqhtZdepQZEu8hnd0jTbDW14nGzEhxBoVfVhil+JPDseO0uM
RI7BcDSR4O1HIqG24OMDmrWYPIR14//fpzu8HQprawJGZgPakhppZ158WH/8I2ijbCQyrYXSlldq
iIsvol90PDIZQaFOYOloLrP14XptF0Ps1cdAaRi12ve/t3AmbaCsI37u1TfzFN0thtziL34tG081
rZ/yTzwRnCFqnNzGWVJFBYxCWG8qoJtUubwtKSYrd96szODwdvhZkVXa2myFpZzMtH4YhMXFtKhU
7uDCYW578NM9biHZ3SITiB3nNdXfCpkC/6qdZ6LDpqsL/fkuo6K9LTWhr1Skwm2c19g+5YpKJ27g
L2rs/Jh9Wlp0xL64C/16VJqEDRcnumXZjdnjCYkR7xnDcq9YHwBRCEokbISk7ovaUmS/+pyBxLwM
XG4xtE2zRGNlXrOo6APBxl/0ebCXJgWZM7LwME+0aikjBL1ffL4rtA9D7g/jzsIEXNrWCV310HS4
5/jRhqa72nSWMXJIl2sq5Oc1GEsniZuVolHKbvbMCWw5fg1ycAGiqhlkWDGFc2QFZKpkCC7EDTDx
bOHyTa7VKtK/2G8TlvNPvaAF5+BEhe+M+2Va6uR4T+IKT7wSgmqQ1Mo7ucIFdIdARULpvsjlOsdn
oARSjYBEMiRRThEmOURk1NrSiXJx3luO1PzJyYf/tiZ66K+ZMRookkHcVOH1sWjSwSodBaN9qG/L
nFUrr2OMy8GnHvoxw+PslgoBoRKgswJ28Jvrc0cZtI0dW21vA7hlgtTkCfiXjlgebQmDwQK6Xj1Y
a8Kr/8jrDQKm1EpNkq/J3hd8NKbrfJ9dm2/UOCJUcz4yslsh2qkwuulv351dPI7Qz0LggYLyCZ/s
cdpBqjS2WfutmCE0QcBYjwnnr27q1CnjbA/zJEOtXzSuWbPfdqrrafhsuyFpzeEp1YpLVcesUAJ1
dIAIwnqaR1ZzUFkd+KS9IdT52gdJ2BUMQhBXgICeKrvzqIFN95T7QbTA5hA7bWvlVdNseCfFCz3k
Gxh+0EJn/BteV87ggry+FsiL8tMLx6CsQ+AtLyr0eTnFGCBRnMbfj0h9+ucOoytDK6BaNiMHSyWV
9QY5Fqk0zmMk2pYTX+uvlVp6PVfvIuEj07dj3ny4HxRcm6nxEDwEdnUX9KkeR9o/dFN+qDCScXIB
oU1pAGAPGP7Gc4KNmDszoTNvaV82BtcvPLYhdLtmpw/RM//Uf434k7D3LEijUIEHVw6Ub6c5VOig
VG25FdNz8czT/rSsdXdYSaeQ69AQIRmq6BIdPPteoYzeZiMUGe3EALh2u7zh98ows4awxwDehP5V
RId47lFiRs1gUFzvgba55YgAxXgyC1ESG98JuhylxJEL9mad3R/EEGiQmttRHwXARWy4uoiIVXE9
s7Cy98SpG/DA17AmS/b1sc1A4Mle55VTUCBuJo9GWUfzf7wyQhoWyBERZFr7GdAO8vOkrwJB4rIi
KxvrkTbbSLevAVuYUMkMPHfSIyTJU6pdi1mNLTzIgMQbfjMohy7j8u0zY3AKEvstJUPuc43xdOa8
kRYEtHR2kZtkQxi9QTU+vikf2s0e7uHU47DREDGJRcrfAokeRikSnsKNIAfNDIl0lA0Eh+afIrZd
n0HKM+SzGTVgXiULma+LvTs8cGestfKLfzQbcBHDVFgIDMad8z8hUwK6RreIhw7e4P9EMuaJv8LZ
Phi0mDBX9YutwtPI3X0bklsor/UjT4r7byATSagICioCJCS3id4gYgz/VlGtAxNfE6AJ62PQmMm0
cPr2dw8wqfcUgUT+08NV1V52On/52pFaUyTh0j00rP5+ObYYef2+JAIV9cnfg1C1+GtNkYOnQJRR
MU0H7XzNnf+7iyKjJgz/A7nT/7vIEBmH9FiqUxU2WbYZYgkOEj54JX0AExq2XhEJuUkYYmuKxVX7
+OE8QNK7g84P5UL7XCfSyMPSsFWpnuWadidmwyj9Epw/CJNLLR2spv0lEIpejLOOrZTEepdc1LpH
Yqy81QmHXHoPhV9TELLIBUFALYTO5LtZQJpXmDXz/l6z/e7K8q4VXr3rCu4LVdPzrfWaTzxgz5an
GOE1ZxltBSK2N1tRiHHS69adGpTIFkvLvF6XUYfPauYR+Kupc3YOKd0x/x2Ei0+4fcaSeSBv3K7H
ZwFaIbszIKrvbquMVFxfWd6yc8czE6tBzlW0l9+rmQztvKiAk5BJlSMsY4yXbZegRBTb8l0r1wCK
2KZgSZf1ZSHrB8Izz1BPr8qmxk5NsLfYcp5dpQFaoO0YGeOsx19mSgd1rd/ASSHmOjiqreMBDTqG
r3peWKs7aNEHJsmWZCw5BZSCbSs7Em1zIuRjaFLbtGfTOYoIiIAeua7ZYBCT0V7wZnM7RK7Y90U7
361KRtWojbWsRVF8KRcC08er/KMocLn5mYA0HRRTYwS1ZqPkSPEBWFRfPUBWbitggXVeYoY6c+K6
5j4kwNtHg5/d2MU+XMk6/azAPFSImPMrVp0e4dSB4xrgNIT29FXYgO7Sb5cj2EtPG8q1ASPQyOI6
nr9768UTqEzCrcxZN9IHB2nWgHY5CjMkdRS0/HZhmb6ZVpz+f4qU07QLuXdWqS7uxb6wKJTAe9x6
rFPn9+P6kI+dgQIba/t4oJa8xKJTx90SRGj/oBtlHS/mczAU3XA39674+DtVPi50WZEEjrA/FL8f
iQ7Nej73J/H6sQRau8leoTPTXiipsLP3rZIPSvZhzYuczz2dvu3r3s8hF8scr4WYDLfq6jDy+vlM
mLlhzY9sRw2iWmMlePekAxajWYHI9uONXzY1w0Ccsy6mjgAHWZwV+QRD8s7BzO7M+iKdPzTSYMfr
6lMkpG4J2sMNMmUGJW/ivIylx3PwF6ukDQod7ZUdO6wUbXKsZ/SxRY9kBGMUIemTiRwnRzPiPoby
YDIUxeF+mHXB9wYljazkRuhHTbriok9mM2nzuAoPN9LbuItbkPuv44H6QAx3clMzl/tTw6M39KBF
qhsfLuxk/lIEQZQEzeRRsOgg8DG845XUrlI/fiLpKu9cyKdkHUmbxp0aSLaogAdFsIz6RvOGMQrq
5/xjjYMDW0V15gMHHvJSYApCqoFtMovnLYRpvRDe7diPwgGL9lETW/AfazYOIvpADG170duXTxm/
kdGcJFcF14X2ltJDoz0TygJjrNQ+gpREbTMBS5BQ3bh+jBgWEi6d1MHbXw7KQWklJ2dMfEsxdVmf
pzi8B+0ofxBmf5B+bqJB5DvtN1LYYwl5LrRJQg6ySKiUCBwCOoR8XNZXpb13utyaZF65hrSE4whK
Z7K/eAoblmFXUdICCdT07G5ZurUM6/Z7ZzePB26nM5bREBru4nf2FOPxRf8BguCJgtUbvOKNHWzf
Vni606Ydk3xmT15Snnpcxi0czESKaYF7CQVfuAzSrwBciAU3rW55TWaJPQkONLbGO/uTou6Ua3c/
rDepjMLDlhmLLq6eMFSUo31yvcNfypGayeGr3/fmwIq+FIvds0c0aTVFpBfe9bDPAQtai/8Qsuxf
dzp07H6EF1jqGQjrjxN3vsLWbkJlxhYFgiv06SxB8btMpPRTseqk4mPiTe39NywZMxWcWB4DAJFH
qN5RbAIHFZ50RmGmLvIyGwq5rDRUKH6fJFeNIx6vwwy9rIyerrRyrslNI2qIifvuNCDOxRNax6Kv
3+yylhKGVboPCA1hxmBym3CQCzt9aRoAXAyUMIMGD6k6DEjcRETFubOuSUgLgRNYAUg1DU8j1/Sk
68kb5EVbuQ6S9PGpyE3YZsEYf61oDGqHzLBdMrveSVgjzauLhNpQe+iVY/fNHVOX7DfXZpN4PQ/G
QXeGN6YRiwwI2Yqdq4t0rni4n6OOPz7fv9+JibovlaOekxb4fmdBtrCHIvdsSNE4ad2SGyQqwM2r
Z9DooKsUP8SaCiA1cEDB7P1WdC0wY5hP0pb/wnN/TGiYleXFMVwLtWE2Qsd443gLU8Ez/2gpstvZ
+YlzGATcxFXsDJgxOQHAgyrIYv8aKC6+idmQKKkYo9AIz+BLwv/m7TP72gzUA97f0mdRZfWugCmS
kvjoq3BDZeg3jb8Bd8y19YmtMefL012JzZLwyz9mleSlcB5A6x0YGDA/x8Tu0M86YEu3aA5fAcD8
6T2Adyqo9//NOZyDCjyGKrKUK+SMdxezb2R4fW+icUrYMRBVMnuMdZsAykXkhoyxvOX7bRVbFGVW
H38/UmWFbFux1bT/cbHYtRcfkWegjav8LpcqpRCK1Vaw47IdfiKwBKEFwapV+1YAXzpiiG8oeXIl
Gh4mTWWSjFh/lHTuaM1bxhUu2VQ3zoqgXeIcjwyTTQ5B+iFqpU8QfsuqJohLPGo23zSjf/+PD2BY
LZRfsMr5Bt9pcY0s0W/dcpvHXUZ4drLuIF8skT+kp367MXf0LZS69SHz4UmCyOjW5QJMHb/HiJs2
secxVuVlF4i7RD1r/igMSWZC1HbxlRiyWFUnWPwhR4XkpMl0pviuPltr3rgVRnIc/WMxQQbWbpYK
jeX5G+bq7SfVH9w4hdGDQPXOUiVFxOJ5sGuY3q2gS64ZjIVbDZhSsvpznEU9dtIZ1esNBAAYZceH
qLf+MMBYtXiWJr1cvDSKh6RXvn4nfRpnIfaiLhy9QR0L8FltQYNk9f3aNOXgaWH4snyJggXqTh4Z
d1Kuda99/XYRXm+h+/aIhii90W/vYcosnjHWQop7cmJIH1ZGq0YNLWlyEV5EifkDoQA/pFRbzBG4
cjEu3+TyaLethbX8QP3DI3XBZ93raXCedCGCyaSCdKK2BNOVjQpMN+ARRaFiXKInR3+YBjpT7zMm
Jfw6adVuydkrwOPD+6dvjTZJU9kqhhk7nKmhS1Q1kqZioo0fuB7fLmUvy0JheMG78692fx0f3mhu
e6ED95qZQ87n2h6qRaWzPthx8OTif41H7Re+1BIffVFOdHnTzClHZg4STim4gDGCmiaxZXfsP2Qp
WnH1F6geHFr4lShD5vSL6AHgwh6i8u49L1RL/C3fRvBq1XKZVgRY7QUzvJldlc4rOl1lNocK2rKi
flRS1e2tQNpm1ZnR2xTN2EN+tWv0216Cd/KJ6yFmODM8tLE6LO3CK5h8X1XCQqQT1L3CYghW+jvi
vVFm731QPlPfH0/F/9fDT7FUTEAGOCtYOIc2uXWB1kknvbDKtdsyq9k2TcvQrywoirwAencJM6lc
9LL19v7Kd3MirlDJjtFO0Ky57m0Gt6NUYu5QR8dIDC2pfWRFY2/TqDl9c/Rr0aBlS4Vu5yFdIche
bwmxjv1l1Kk0827c5j4GZAw4xffd1UEXU+o0O/zuHnMqZMq4xVEOb5Bk24P4+SSO1IyIPCoKRwyD
Ab31C3ceV8FVxckGqculRARu3T2334Pg0ft6QkbvskW4nkQNjjX/cwjI4gQ4H78u9K0ZceNRR9FQ
R+2OkoBMrEGYDHza6wrcdhdkb8iaZX86T3BQQ0XetLjqGrvJU35Rq1x/03+J8gGVE8zsxxyqlTgY
VdKHhkFqRqOzTrwoEurmjFINwxuPgl1X6L7bjXhDbLFxK+8hICzokzukR69yhMSj8v4r6YWoP7Y7
7T0qVho+jeegL+HaGy4e8fvf+sggQGjWRsT30bYPHyGa23gyV9dkQTvGOUN1W6O50s+SYOaPL5qq
IfQBdUIv1w0s3J4lO1w1PEKd7IglwzonPd145ko56aGBsD01TqpwY33Cl3g6MMWb4ZU5P5Y2QGav
pfz6WnGRsJWBz7WfT4NNUfokTAsdRGrhWTX0mtkscMjjo69dwe+/juU6aiwZUn/ETz5qM4qPs1eO
IAjH71uskL0ENZDiyjpjeedB0LDX5YojrWRUzrTB/y4sczI4Y6VcBk5kDdoLVjYDiM1vHM8kBSUl
2UA+2AwoUyoLQ/fgVTb7ABY9wgPrRaH2K+R7+kXcZo6icTdMK/tUpe9xTODCdk0UhC3/jme0rdq3
Uwzu4hugZqjaomMbN/4tOrCricmEBu6sOwOyrzl6QZPGwzKKURJL7sw96tdtRtfGDgA3RjwUkdqE
HTA8sTKgw2UYX+YiFNmNlaSvujJDtOXQNNoEWAXM6JuxvSrZr5P/9BFXK9a6SvZgxZewzgM6lqxM
JfPnfrIGk8NUeo09ZUX99uKLIVQRxBE3N8lfPENf9H4/uOH765LjlB5Q/20gZjJiFSQ7Ve1bK/hv
KzVm5d7t1/4AZcmCjRhr7+j/z6/0etu9LGtIbjGx2iJmtaFRN9gDciaCNVBO9H3NU1aUO2lnqwPf
lzgCyZR4dNtBskyBw2Wq9bBERJFw0Qg4FzLnIcaSWsQwIyGSu0lrm0Dzlu+AfTENi8KrD/URag6n
q2O+FQnmULp3BLj2Rwt9PgVmJWJoPE3BxvflqEgys9DiOXMeIs7Lg8vaI/fBObQQLP2hAfGhGfat
xYIj7ypvgCPt8kQZqKYopKzk9pWQfHtgIsZFONQxQkRoFhj/SPwxQASycHquwZrUV6WYQOIvPp6J
pDTFmPGPPkCIgW/ttC2t/lu75uc7KKXTHHUfsK7ipkD6jxsVL9xu3kuJSfETun+LZN99+ERkmIUx
TBlS0lm7DCd7WXwzJXvPQ1LFxYS8Pccrp9E0JIgZUB6T68aJN1pp+vVaHLeL8EQsG55FICPR7g+4
2rxJfboXb5biIbGbtXOWF6Y9gS2iWmPjHlHRtZLvcPWEF1T00etK5Ybut1+KkGsaa+fT0IOJtGUX
RTZq07iCIYQPViwsZsXgZnHTgHMMD/fvDO+9TqTyJQHmgL7T0iDRMb2Q+xxoJ/0MeQbaK++HJ6XQ
xkdEBbdP9+J9we7Rpey5AHqoVg6W8uk1B49fjb8dLbHJDZeCWPlpxK4ECe6+6wpTjc5LPBKmB5Pd
sR0sAT+DdiQM8PhYbOiRcnzKn6LRx8M5SnbMWXKTVamxgAvbKT6+b3Qbsxvb0nv8IngRTDMIT/yX
Bi1SIajR/4Myl5QXfftRMrj3lQAiplVqNN0bhdWcnbagYPL1nJoj0EoGmp1zH0ejDycoeeyleAEn
rKuVgWdXcvoZqDYYV2MMmp81b6H5QKO7384/Cq4hqN8naXzfivgENgjELVdadirjZLTWonqKyxSv
aQgHFjdwL5EUeYJshT0y4nuTVMn3naQYyczz+Y1K0kBdQyeiy6NcQjSI4ZYQEC4fnKS1xRzeBSEk
OwcqwQKc4AB9wpQPgS9KP5NloR46RJhC0WKP5O7pim2lYGZ56m/kN3JxZaFB35dXGUxdE9SFrm7y
VmNeKjOdsX2xanFFemgAF/VIn/rsMw9+7C062WjnRdIno6jcsoK9g7SuwyakezpSVdKX9hxlDuVO
DzKKaF3503KC28UU6VFJlcEgigJUFQTfa+GiSFfIvk5TiY3Ewdx6WUh2CIgoLbEX0IWVTMLMppYE
keFDGrGFjljzMJ3jWHlm7VNhcGt8+zhKCaJsjApeOJ2x/lOMV4fWfoENLqHIjNQCA3R8bXScVrID
DuhszTeRXsdvulUe75DFVOyiKNmRp5CU4ULMvq393FHNUnVjNu2fgo3Gq+cBGqy+MEOfXXmqS+2U
+oDThWWpXKH2PgyfmZTOaj7pQ1MIs7UFCKr3O6iVVA7tUMGeth6yJMbSpqKQ8WF4akSQrbSzpciS
7OprBCozKPPjDFSO6ElNa5+s/cphn1AnKGG/gX6mZSbT+/H2UHX06u7R9zdNb01kU68Ugw9rTkMt
YoucEYzxynV42uillITtUlAZKoTVHgw9tMcCF5lLwZDluVCKSDmH8imYJZ5T8Ot7h/cGHUXLrziE
kQJymrj02s1NhjrsLGXrXivFGsE2a8RTfMSsBYuUmOyP3qc/vXf0oS8ErKXvr5/Qj2CJBG/QrsJ7
Tez4zuaD1/2kkF0yLIYqEvUrs38KT12S4yKS6tiabO9qIUgnXeXfmLuJapDWLOkQrWIWmZCFGeiz
c/QaXolcPjyQmi4WL9qSjfHT+IwtHptuJCULu0kbr7hevHIAqAWaL+nKta4Drbu+9Z6CncwFJRss
66Kx3a1KGoYkhvQmVYCdWMNF8BIPqgbvwxbqzq8b7mBbUlFuWLMfRL0fTmWf197PQbRc0uAva5l3
KXCzcdktD2iIRWjlGomJufKaTtgVL/kd+NUnKDeOjCDrdJ9miYU2MUnnXChSFwv27VW70D2a3ouD
oCkkkTs+AG1EtLTHjG0Pv1Cz+eJoY7e540IXL/PA58mmf9T3DImIvvLVix+0vV1i/x/vK4AGiIoS
u6QXkn+ga9/9QlvMMho5eS6QTjexDTOW86dbnCJcb8IJcCatZxrYjY/KGlLXqn2r3dhRgfla9686
hD95wd3lrvp8ezfDjgGlX7bBKoNHteNghgzlVMkppUqHbcS9o6XdexoqBs1B09ckPT48a5eyZTVb
4jt8ykWgRVaSoEIoOlS5t2vevSY4B/eACs9x4QlvrjA2M2GGuAtk7bQim7/fGf+kkKN/j98bk+at
hl7mXc5ABPcLyOs6E6liTgpAySYsLv8YRnUJz/gEuPLJhQ1BWc/LFt3DXeyRCMcjbDikX84wKcau
zvWWlrEc5ihch3KUkPaMSRvlCQPJBsxLaP301vHMxumYLeccg6t9YVEEIaLb23SUaWiqCj8nffBE
JPpR7Mom1h6vC2rzTPbOS7wid3iI2ix2Im9Z2cg4I6xRSLkOtg8jeOf4g/Em/mT5aA3/P98+oVga
CVlcALL6DaDBOCzCYDG2OaJ3Rkp4G65Rin3r5eQGDwX81omlvmRbDMn4DHyA603NK50HdUDuf2rv
3cF7TIqXn5dyY1ZVvPqwstFbooJcePk/ChZObNRP/MlhD/vCf1KNjpu41EQS+uadzAqWteHoKzTo
MKypm0yDz0U4aG7gpwX0dBjPUbyAxcM+gYsgCPiOyWxJe/MEKQejApuYcNI37jCwe52o5MAjxzbB
3GtCnjNOEE1VAofntfWH9zBJgMEb0TGSlWw6X7Xan1si25pgLQcocI/8sGg8rg0k57fVUFrf9QDj
oiAj9eKm/VsOi0qK0NUerrnk/ExARVi8qDCFDnplJyMtBUhQvsTb+J/gdweY+eW6tS9JIXZlpi6L
PJqghuz3l75up80D2ahOs+u8J1/memPk+uWQ9NHlsdW+P/RHBjkJrpeL8ZjiI/zheVKF6+DpJP+S
02QKUyGpSgeMWMjFqw8POl5vu4BxP6x1OxMo+v7hknG4mxtdGSGdjE105Z55+TG37m7UvUzsU60K
I0Q5+8JOImcEP7LPOA7xIfCoeeZMzzTQ5yY2/3mAQjpMdmHoXiLpSg8njaU6GomPy6eflSWGvz+w
aUL+TxQDBZXQIUpMTAbb/utuCnvJc4TGjbNUUNU+kOfQ1NlkBw9mgxAiWVs2OygkpicXSLq4aF47
A9WKximQFGPxHrDfEWnoShSL587PTJx4CgiTP5VrkmN9Eg+d6Te2UMew0MY3S9AQonhBPKBtcxml
O0kY+4OfodSb78FZF2w1tbSZS2Q65lApHpaUvnzFkgRWBiCVMizCB44k7fZzOdHKtD7VCpAPJnwR
0ov6dtzg+BdQJhwdn0fxsjZBG9RTuL6Ykg5UYRMU6amcLzoH78QEW1qLecJSJfMLE1/NWJNXuqE2
NbnlMUB2QfrkoX+bNXGqn1RYDWunEcCMRlGV0hDMOBrjspBV9X8lqcnhIN3kex/mhNKRjyBr2Yip
p831jRvCx7+eTl5Y0SXgsKDMQb/waQONEOtwRFBolr+kRK5zKkQe5JdWovFiP83YsDurY1j1bPx3
Jxqn2oaeWLdv73dTuzbZVNlumVlJVNP3k20blyXCB/ZzwPjBkbcRMec7k/ukA4Nnb4m5MSGAQW2f
bIJoO6OIfes7fkoVO4ptZa6ocduN0mf5lyrZpKJKHNA/ABVKMcN9DeyYmR8rooCC1PDyBfasQW1K
1erJVoEHp0MtgGLnqO/yxSPX/aZwW55voZylgLyaXohYH2hMd+ti2zyL+o8UtCmIUyPB6KpV5odH
8u7YJH2PNH8miNpxd79rxbEuBy3II8wIJziIOZvQhujURbJmGnAg4sl+wikpgayPD1taYMZ3V+00
uL8iTJI+YBGtOnXsnrwwb0rlW7LACSNeLQ4c9q2H6qQazkjKUFbsIzboTL9JnM8C+Quixp/tyEqU
+D1JS1sG2Jpx0l6zK8PNwwyrFXMwiIpghnWpxfwWFmGv62cnwSm6NHwQ2P6x7Ckl2EWseGRxevM9
QmRPDtw9sH21+qcpH7Lq7hAVS9hEC72j8dcw6X8eED825Dmg8dtZ9ui6VmRr32xC0r/yNI9av+BY
53+jCj+I+OA+7N8vEIYXipgBd+4yBBKR2EP8+nf6xYZREW0J7WZDdKGBT0q+mYhieaxSVmxpFGnO
uISndT5KJ+mvCSgI5aLJdiQoF8uCxJGzchG1C3X65bwZqArhpenTbOKh1eyHsr2hj9h2TaHm+zkl
Zngpq0X1wF8Yyru4hYrLTncNIoplobwzo0fmfGDeXa6oNxZFjVbdTjcMOtxCY5ycwh8XqipBXBGH
KOuJA2ekhCeRnXPuDJzL6Jl69YsSKDs/RTRsRmNMyenWYA4Anh+QPdc1JCs7P1pCIbAu+vvSBVxe
0PTPMCpO3N8CgM7yMMA7FCJ7ZweEenPFYiaFzvBzZ6BxWOnP/rDO1Nqn9fVjDohVN483Yfp2U+VG
o76OXqlBWbazYc3xupuGs5RNJE3Ao5HNer+nRMnPoJVrHfti9Re1wo6R8Z4VwfO7rBYMJoXy8RCy
ooxEcrcyI2X6iFe0eANYifPoJINGt98vheMbKnSX0ChsfkDwyW4cAqdC1a7lwC/A0IRYP1Ol6RNn
LTyQkcy5u3oomS34+Ord+GwNYr72CHQNj7tzfXTBHZ1OAzlLY3YxQ0kr4wIyugESOo4ZjjOkeQQc
sI9ha2xfj6IRVxgz01EtEx1Si41Iq9OlW8OBAG6O8yT1XgSxMPslg81GkErDokGQ1UzvQM1G+nR+
W7KUQeQsYnO6mPApGyEQwUD9ud3O3W2rvbhIy/+xRcc597dVmfI8C3wB6daToyhAgrdedJGybUbc
0/DYbiDEW5xO2gHqasqkev/5KZE7bqZdv7muXy3cADWJD3nfcBOp4NvLOMw8HZYWVxqXsNBi3jpA
E1uMtVgDIjjBGbLrHkMpPZb7Qhikhygj0zkknXzjQICOLr9Rap9tiIeZBPAamIwBmLK8Jg+7vFTo
NCUOpKEZ281DeF4gGSN+/+iIEsT46ezfVZp9nz/W7wdliI/ze3mPRgUCw9XNwOAbhgZCZIb1WDrc
RWjh70MIxBwBZqIzTeiCysAN8i3Sh5buiUhSwkHrMjaUz/LO+0fpTaedAYGY4tgfo9ZrcieLBqrL
oMxsL44wrIseca+8kgKI99qGo2nBlsMJ1BP/LcRdF7ahtr11qiKaod+bnwxid5EWLfS+n44jDtdY
2MEDLQn2dArdWMpPjXYcnmmyGwVHCDrUbjQmxs1aaBqxnkVjY0xSHnC6xBHl3qxnqS04PVk/aetd
OBPZPwVF9Iz+VJZ22Cqgy/sCphz7/gqX7LChRijcR6mtdxLSRnH2JWQvrmtHc4uO/qBbfW8du2jU
r+ukm3JTpVcZwv8gX+DFY28XTpXvMYJWS3qWZKTNrc3sptwNXIThT6QQL7QpfgSWJiog5TQEHOio
LiIU8dOXvCfNesHQzywk1J9Igr1gWHiMZWNuZSLktqJXv6LlTY+33B683z+CpIQT5qe/HFWSB1ZH
YDQZxzgOkVre4TBdtTj6JkOjh9SSp5i8J3NFjsEh24XudOC2oR6uKPFINc7HtHKZFaC1bXqfV0v5
HeNzVBcW8bQF6XmOvebovfWKId8wuBlQPb+tGBmjcle89aX0/HCqIVqQnTzvUJaKjY1otVrJJhdf
qhIcmP61+nXOHU14rmUYMHpYJsf7/a3aAFGCz9tEq4UeZF2md/R1riHenLW6c3BpuOZHMRE2nLo8
ffnW62gBtL4qx5DHRn0BSWGue7i4OlhRg9W4XuiKvBonIny6xooBTrWBPcbyXjsGX0YjaHwLJOXH
FApMx5hmds/P6OfkUu/nt0dDrFJ936Yh54EOkAW8WUMSav56BtzL0BaB0+U2CX9q4LjTWv0xXoci
Uo/jyzvfZzmNWRZTFScJIAOKkU+/7RJrHPMt2yOFN9i9gOGo9Pl1jZPwgh6FWV2+G0jGMbtnVwnq
f9p0DlT/qMwXBW81jUujzRNLBcrAtmoQawy6GekFkBCqPzTIIikYl6zPWdxvPHa2ZZ6RKf+RBdDi
O6RBE4LBegraB463MecEW4k3LK39nDJyL9rMadBp5wmUiiSzeYMS9K7rTa5+nelrvgaFZS5tvvTX
6Zqv8Ij0+dgIh9AVRxvKitIGrTl52/HEY1dXI+9QTD15FgPYyV/YIPGG0C7XOy+LX3Xr1pGdLmUW
IW56pRML1yk94HXeV2q3mvBoBxB5O0RVLJwd3d+bn17aWZv0bWgzKTFREfau8ymJ5kPT8fx4Fjnk
7rjxI/E7Ch2l6vX+O5DZ8JekKlx34nASnDR5eSR1HEcvmQZgT7QkhRcYQCgTH6iNRReX1b1DKJhI
e9r75RSMsKge1ierE2aD/y1yIMXqO4S99AweK5yVnKeBbuteAVDJKyjj0VoapluAhbgQ0NayfTOs
Aztp1Q0M+f9+Ne4f9js8JFsR5m8uQoa2XXDwIxHcFwJYGDSa9lkc4ORlckEbbkx+ekpaiiLW7tvd
ZpYoUp0YtwQYk9Xl6bTRg+KMPEy2EwcdWv6YSOJny93LV6mP46SAWYisGj+o/laxEJwLQgNthCgR
P3ugmAzVUb0RVQBpysQ1N+GAoFKfE4+1N4H4Kb/6FFX19XP3kZ8bOjCC/ut99w+s/wFeVQk314L7
ZbKhq4u8mt0qGOy4IcvOHKYKzqzX+/d9dXkJjecYckykWVQSMrfYa9JYvrdVMkyI34TsOwUlwswd
6/dza8RwRHtPdLVDY6uRaxXJN0GHiVwIwqqaU1vtjP76uGBpJFCYr7P1DdcAqvu1GZD4sJOA0bU7
yUxblKVHZIH44hoUUw2FFtx0kd+P0pAjblRnvsEBV7NNmdhZJhCDrOeeDsmpMzGoGv3XbA43d2P6
bw+jQ/QP+LHbyzW85XmsEBg2ie5gGaR73wUjClSNts5NHOWmvscyMJCTu0LMHU+pakHlzYAF9uhh
sWDegakV5plVMrmeHnEHKe/ju83Hs0ICiT4f/rkYHvR3ryjzZaoPUGnC6IPBmMXYRTdk4YupJXMb
DUPsyEkLW660IMNe9G86BQx1oB3/pNHjq5KcQWs2ZnpU6hkJyLi8qAIV+3I8l2pX1uXclvLf8NIX
xJ6ScA6KmlR8F6mhmbGILUKeypfFJld4yL6lepL7HU1l9FgHMoftOO3GKMJy0rB88+JbiZ1N+w6K
qBZjfq10EPtwGZy3fywC5aw8tbC0RVtDYXwjy4bExNYmGPy9qJg7Nd3aaF+Ac+h2hAs5zW4oo1fz
lB2vVKyP2vNFKFyw6EfVmDGrnlnMlKz1d4nIJrfjM7KuAWEJnozsavBxw/ptDVz4a55J7a9FuChS
ztBouFLm49Zn++KddLSKa2qLA6M8NlRNP4kSNIwbioDZDGCyBXotnF3tQKqS/z6xZrRAxCfzVwz6
W5kC+sosyspgZShslrgs/FIpc6HxJA5Y+J6d9kpxDqoo8EjcS7Np5UjEWZv08nSAPVqvlIi20ooy
ej7BFwneKj0f9/AazY0QaTxnnGxgs7ETqoU7HjH1JCdkq8npTb13P2K7X1fIuE+QvtGe79RW4aic
L1v4e063K8b9XQvr7KR4OxYgg47gJMj3TTpwcUyUC3b/XfWXoHS7UnZ9+p5ajEgrNh/fDvWu9fDo
X4rwipMVGJT1/X7dAisatC0hDD//JzJdoDQRbjdPX72EkGgkpK7jtUzc24j/iRUy+Qnr7Vcfdyu8
MYfKOchLsEgF4rYtEfBGK6idCByaH5qYlh2kVDOuXiyhY5WKOnGEuxl6fjdZfk3XcEdAuTwR+owq
9wpfsR9+qN2LUNFZpMbbTml5JGlF89RWw8uEd28lMfpiCA7scqv7ZJ4vSSf00BS63LYTax+NoAjZ
W46bfoUmK+sQ8YKFMAp946iy0N77wbH4v5p8GET828nH4SbAUpYbws2v5W5mh4TjVJGoePuG5MAz
N61wMSCTOGTnvwlZmb+ha7i7lwKCIzQJEW//BAhrFvj7cEQzpeEkaTrk064kW/7SrggM8d9jtpg/
VKV2Nz01tofYH83roljL0CGOgbabszMN/yZ2B/UTyMqUrgiD3I03o2MECYo/DRzEA0HTwTnRleBc
nSbdjx6QjS3KJu5jZIG8mPu5ofhYTtKPOQGt2SoqWPIqY+heSy/O8Q20FzCV39GOjxEAOJUj/e5r
QR9lBATFIZPOnjG8nJ1weOsOQFvjA1BaFl2YfJlHp0xOPK51TGmqb0hy2OzcqqmWAlQAzJmTOCnu
vs6YSk6YwHwpTo7Hri7TFk/G7cS86Kz5aNRTBh5vaYZkgOGKYkShNMIN2j/O6jOZtBJRUx2E6+Cv
g+Uxujhrh1/cpmVqShRyHgregcbTFUwaY/YMHHio8gIDTT6CUfsdjyWNi9wl04fK2L9oiPCQGVSO
xzHEmRXaYHXyPOPcIcEBe60OqNHN/CNiuSpMYO8IrCb5oEsvVc6NXbegcF3kHJbd+rBmzS5+AU7M
Goj/BbwaXonjS4Q1kKlhTfCIIc0vFLiN4TlzrLVuc/70Y7RFU1ZYI/bw5ZYYqXYn3gQTbOSRBLE7
iqS+sFpt0rLaVpS23hCWAhZJC67R9ZkwNq1IGakW9bU2UFQKsEtWCA8uL0uY3G3ZET//Wb0EySQE
AR8v2TNva9MG0hGL4mDw/BKgkHeWpSqjB8P1cNssEbAu+fVQtyoUIEtIXKiB5nsUr8fI7mymg7NH
ve81Zvmn2drlaFt1ybUAFuiAstc4923oGo+aHVNuodOKgmCqDbw3hyaIJmF4Sg/nK2QHlk6ucgaj
mZWB61f3KL9Cps1JwSty4DqegtGQHjx9dE9FcDfEkWyqCpRPCZ0KjQo3kvc5Qv/QPD/GOhvhDKZp
tnPzEtSmvs1a5cJVxkJQr84mYkPqElHdLo59nexu88wKTMXFPq07VB69h1xcnagpv+h4zhG5d0cM
/LzpQD/7+ZqppcpTp55nFD/aen10aA5JlPtLweZ3YRxDAMmvH51xZF69SzPlmXeM0ogRX5jEIYwk
kIFND/CwETJEfvPEvmEe5hnceJ4KjxI2Frse6OSOEb0gyU0qTHwZs1edKhGTT2BNuCYz8LZCbm6+
lRa72q82tvEzOApI7BtT0ILpVWzkk7SnS6KFRIXNkp31IlmF7zNZAQlzCzuqhiMOoANET8pPiBPh
CBfjs58IwQyLR4OOgPJumiF0OkoaBHMrRuZawQXHk73bspdqGdzsZHNdUGXNtWfbRcZybi8Uajz7
6dWpCmOT7KWkGOSQtrlYpn9Kt6bKOyDStpl8szvCZVVk+oElCpRW0u84lzk8k2sIx9jIyJc0ssRQ
79WuzCHXJe/dYUl9QpkdSqQZLIorlMRphzlcLTTTcIeoeT3BZJaaM8WG8Q2auK5n6ptll0vHuwIk
8jlXRQi1AVcQpcvZ0h5lsbO2NKYlS/5nZvoSN/YKeM+QmdBb1LRQ7o/G3eDtu8eVcMG2ZO/tvmoB
ONINCb+/k/KNwUc+ErRqDq2knJMDD4rKumaMd/QbCmT+vECYtzyF9r+inNKLsC7rgSX/JIOt53DX
vM2tnUw2sI/MOz/hf5bqkBJ1cr6dvhqLRuYw7s2+3if/izW8JFXD2yxyQsADFGMOzzOaag/gN1xA
7smzC8lJt0k2KFUj9q5XXYIWljgRSBy2JT+/ck25JBFznRvc5BrLM6Bba8se56moYN0Gw2vopbNg
+k1Q9j/nB9xXjNcSNg7JsX3s5Ob/X3mrsnLLvYd4bt+nfKN7t/eIJbKbirpD6GzA8OtWMxc6aH+3
uhH6fhM6iTccyD1p0iuym28/ICq7wolYS+gZM4Ipw02BOztDxQUlewjvfo/TjG50xhbOe/+rnzQt
qM35QTxoDqPXXtCZwoTQ4Vj1FZbSGCMtQDGMHhlIT/OLgSCFWPOXWvumv+/ea0MR09z75iqvjN8r
nxPcaDMmVMj2Xj11t6loTwtgzpjwi1CGP9rDD0dL4F96QL05WDmj6wpA55fphTemYc1gyeMdLk0g
WNNPv0HQiolY4O4oxvgWWu+BmVY7NxY8zTELaJJ6Msi8vgJJV+e/YwhWaStYlscm+qMKvodQ2Hcv
b1Ms6YkDy1JKa+bON8QU7s4h3/cZNqseWLNP7CvkdINTLpvkk/jk7F1k+WO5nrA8F3Apt+z9lH/R
QZeCCve5KPpSd03CNdmShW73V/Ug6PTIdYl9BSnRF8XSsPKSn8TeYslIWQd1EVgrjzQCEnkqzvRe
WvlhH3aj/QwLL0hqozYHYXWIcG3UErHE4H8SDxQV9B4dyKhoc61lEbRaylYsOejOODwh12YPfL1Q
06GNkOPChPsmNTgJPIvV+b2aDUwaPU8HqzSTTFi+Gnr0Q1LB874bMO6VmSOe9RWouCzJLBK9ZTfC
OwEZREbJz8nBd4WzKjUgFO3LsmQ9IZt8czNgmPY5jiHEIODO33PNL/FwGmgNDlIUHRC+HVLgN2Tv
YXJUhT1rC339U+IfKHbTIxqM6go+mS4b2+SiJ37jA6kt6yEl3hVmeCuL5iAkU0t4hTzKWG8O7ZIU
Z8v/Wv5BuEnkZUeE8964GbSb+IZQGnesI6hZ9b+NoCwiVCGY8vXSlXoTUpY+wHzvQLcfbVzsjXMZ
rZ4kSRZwivkKw4RyBBcgY3glKUZ1Snmfy1Pe0HFFeYY9AC7c78JmFtcWgTmsG+Se7RIV6JpERWoo
sCkVjK/gHLNuM7b7vmm+D6YlNaVNlX9N4lk1DtAbFxYdolsWzBcCgOaEb8YoaMgZdldYpHdSfgvn
n5phLtlfKR/kYXcPXSHIvu/2pEd8+y4j8LasP4sbjeE3ANC+MoXZYgYadMo2jcp7y8hrmTQuQ9BP
31F1s+rwsDPMWdsZ7XuywBRO0G7fjWjbbqOasP8wOS3Qzftrm90uIvUSlUr7pHHArHx9y800iwxX
J9rW6jsryXR5Zf+VSXVUvxamf0iwHlBrmDfMgWdFd/24ncYhiTIxEm+fX3bNWIQPNcK+wrWIcRRc
m3tAvZz8qnxPVxebo5cb1GgVy+Y/Jy0r/4H3DrHJpBqkmbcrH6aDsqCvjNypUBEjE62tOf5SD0jO
IxyQL+xrryMo6M1NZH1U1YEtOAsfW4wix6OrDuGrJrAFfONKLdY6ylCGSA6p8U7qTy62ckSmmgz5
o9VXJtY45j0GQFT1q6C1BftZp7gWDdoqlYCSfnpT75/1Q7P3Uyc1wrsAvVJCQW8e4qRZLSfH9atN
JUiFoyF1X2MM849LyGVrQAoTvBh3VKIjrFvMSH6/ik4/OAatiINHe9u2p9bTUJCM0PJgevuoxN8k
g4AafD88awA6SIBS+ThIN4VXIgrLt67znI7JU58niv0URHZA7oW7A13GjwH6n+cZ/xd06cMuhYSH
JS/HuLoQRnoJJwxGMDVyd9UEk2lywmAB1bYPYSBWaY/1VNxlx+WlOD1jMCx1diPUXvUgxmWuYi8R
sMzOkOo/pzq9DaVaokK2olP2IRUidg3RWQi/PJg+knabRSQ4waDBz4nHAlaFxLOGtGuwgEZMIll1
2RMUEd4Oismui6QJ0DGUK5Qz+Y6Fw3uW/vS8Rm73oEyybrzMJ/s5qHUZaGBZ9xQGLgxN1igqMCI7
b8d1nUZsFgLYESN7BDrk1f+oBiU512MCvUY82EtFKt6pBt9anLOqH2Oh9nVCmq58CI/TnQgRZR7O
h2hRfjIcFpL/dSsisQ9z9L69zHIpRb8qpEichRVC1nqXsSe8CZS0LOuLXKUBFI2WPNhrwNwhorz8
YHJr+b4Ib7g+6mYf7NkLgulW49mBj5MI7y9aAMni9C7mPn2rB9WICoYneE2aawFxCVQkAvBrrWqF
t4F4LKBIx9mQ9kZBCWq+WK3V+oK1sayHlnCt/aFtaqBt+klFZE9gKD/KXpzyN758UaZFhbUOfp99
Ev4DBAsp/GKvlrtPYmi5c1S7WLDG8rqR753Rqx4Pf8mYI2nebo0U4LW69FFsG6zie7BPNA2U44kx
B+7esyAIxYB6pqVwZARF1ToCc2MutRLVcWWwcnV3+43lMaKTGMFej8XQqnYyDB1/oUyrmqo8UldT
YbgD5jPsa5W4rbKGfl+lPK9VAz8mvyi2LmbwHkUuWgR4SA3+Fk9G7piBtR3ydK7VZ59+1pJlNPVP
Hh02AcH0ybTzS7oP9RetfoqxurhFx/AtTgiSlYBqPvrgAdNreVYRJydb594TSVsP00zK2jjonce7
q8DJVVTgaUoHMuEj7qkcbCWfX4wFJvgJ+I/C072RovD37RQ4XFeKzDR4pStFhujhfc/r7Ay6rI0X
dRUGfbqer0jH38GgnvLImULVHM0hwJwHhPvpZW4IyAqxTN5Gi3hebv6xDVbCaCF9B02a8yas/bpv
Rl2JYnggWdWf9NMUFOM6htxGSsmjqBeCGRmGUm380bWua2bewczHNXdikTzHHpKXzrliGp8AKag0
LVWk73WqXx6eSwf2ugh3POnXmqN+zdnL3fkB9tJFfAVT4MBLQrxnmR2grzvmsUjnMupukSwniG4x
QgJVpYcEUBw2iTacaH9KOpCM33k6kP7l4JMQyr+SVtlB6VUTfV8Zi+qb4V+reVeDnbTuDBahpjwC
JpVdWvxzX/bHtnUmYjVCe1ZqKfqhH4JPLqe0/mGWTyjBTvHXymz8a7hvKqLfD6FNrwzJiIBFl2EK
mpBrzNK68zoQB9uDlOL2p724LrhmEHrWPAZqwRm68+CP34pvRCJWsqGs2J1QXtytUUwfe3533k2K
rLw3qwXhdSAoYr1mk+eRFghcZD9YsI5buC/YZjyc8NQXBaK6jfjTXwJx+15If3beP8vzoZX35iAv
qnkzpjY8UZGJTvotbUXRn/G421iSfc5GkNkfROnFSnx67A9uBFLfGA/GHyPBwes3LA9DIP4GcKXE
2spYC3s3VZprB69Ln/44MkI1UCRbfAAkKjzFEbbJboexu5Fp2+UfMqchUT+tvBGaLhdon+7u6bSE
9+LNha4F1EoFNsTDb+o4Qd5h2Ot3V7PDrlMgSdnQG8GedT5vlfzniqJVADBMYXJ3wjswGw0HTyKx
FS6AITmJT72pvioRweANWyggyKigMGGgAvXcVogEaXUC5wBVuZ4hxklNSJdPrEt005w494bqu7ky
2hkTy5/nQLXaniXquI+orW5hCpF5LXx4m5yb9QLByZngZ57um+ccZ0AFXslUYdT5M3gqmZUaSaB/
fQmwD+PZtuRKE4V+Stvzo40HqRIclwXdly1ul7Gw89EwHD+QfoJt9jRy0McPoDH2/aUY7lRNLMQh
4Xrd00jV80Lj6nkwb6pD+6An9JpYwRkGr6BtN0AQfOf5IMDAwxn/Hzv6c1hiVspiP7+ZlBWSjLO1
ypU1+Xs+VxLk3a7UiaXvdtjlVSvt9+Tr4CCir8/OwgB9ga1y3jtNXZ/5bsOaqrlYUGVInDndseMS
VKIahDPcy10Xf4hgAHwB8r8hVh9830zmFyzUzi8xGzr8IPFvx+V4rhqmKVslhDd0i+duCraOVqo7
r8TO88q3CUsN/9OZ7uL2pBhvFLDs3g37pj7J0KQCzd+Ap3p0OQ3kQFwq8wGzlKNTf55izsnC2qas
zdWxupG1wDlJOFunQ9N65JTcF82XD6lB0wrgSLV64hbdwQynkUPqUNQrCyKvJFXZGyQ7wmjErkPH
rbqqCWEGM1HAyPV7pgLJrgMX7yYVu67ZtpM7W08Nv7qY6I5JqPNTrdGc21Sh2ioVukB3rMNlER+q
aC92sOite8gWyt0nxKCZ85tVcHW5hl5iEcCgHRjV1p3nEE1hWhlsIlOdv/xtmdvhOz94a+pLSFe0
MGcwBQuAA4tTr+xK0LOTSWOAPjCQTC7AVlskMwKJKef96jZvfNqARSiYu8W0W09K4Y3TZ1FTz4P0
uGKXbBF7J9xZQ3wjHrmxmqR2yQHXvZYeMTNClt4A3D82j3OCEpfsGL664jw/hz/CVh/x0L8mz7Vp
8UvhpCE0jK2Xn0mNaUQDLE1OKHKA1YZnQd5+zod9b5x+Y79mkhw2wG837ibIjJ92/+8GoU3IOJBF
MYqxHTpJjEtXBEoZmfjQr5ve84TNmx4+RoftU90zyNT/BwGJyYC2Kewpr4+eBTtJ8LEvf6PG1Atv
02G9SrNqGKRSBAa8NLk35W99up9F6FLqSrHidaaECMovl434+HrtbfcImHJE/VGIwKCCd5kyeNzn
9LlGRVH+drpVAQ0ktAkDaYWa7Hh3dxFM3AIxFul3lohpkiQUeDv2Gb+Vu6yDAnk6C29iv0T3zWzy
cQWpuJ+Q/CO09WhcQIfjX/v5Y3HPp1E679op4YB8y5L5DTun5MnCSkf0eqeABzM/IO2eIf4NJpBf
hEcO20m97w8lD+19oP031NiZ+AiawySecMqpRyUKAr8idD5+zuLRsxtKpIb89iiQ6pYbqQAR+cCX
sIIUuA7jknAb5VRQIzs+OLRijKAW3GYvHSjZg0FWj3SfrJJL09IbTpNkt2+Wg5o1BnGKBdzo7xXn
wa+t1oxDASSygxzEEEoBhnEMB1b6Q7GqUXCFvDvlnmabk4xiM/eCRSzsGpb/DcEXnNNGv7T8UY+9
yuir0jw9juw7TQnPLrhG6ygJ/EXCvq6DVlvozepcCn+NNOhd7eVq0EiSkb6sp3GGPi/t8bSlnaP6
bNQ1kpblRA/sfrXRuACMPtSB/3lpRu5bbzZKdUPvlV4tWvek5LL7KVPQVCOTmyyKHSht0+Ym600C
UgRqQtu7ri+Od+iUR2a/cpy5V7is8E5ZwQ5glQOPCMpDuRa3gqG7L8JTqQPs+nS5DeJG/SOGbIPN
HIi8XPaOFf12D1gkwA+UvhE8IdS7IGbt74BCv6e2wKW4kegz1lhX/s5CCn+u0E3tv1DuCWLh+A94
+sERgYbv7+Vx8dlJz+Yorx2Uxsl/whKLTA9NzzBv3H+v5JlkAhuHWXGr9yTaOmPF/8UWPbHFbdmZ
qvMHc1MitQu1PHzPq27BRSboVJ54GwNztqiIPw1pvcWHNhU/UDXq5QyDVqOWCN9qc7BTp3ruRRim
iKg6tnyQrx+zeKgW9AOG+9p0LVinH4aEwr1PFOTRmjB/ljDaJPfmwFmlVXzNBnodc1+enz+isF+w
il/rbU+AiOhXPdO5htbWX8HtLK9lmzFb+yp3J8UtjjeVuUk+ympvADmaX6Wjsf2BUDvPhZya+PPM
wItcIOs4tlV825b+Z9h2LJXqoYj1UtsC8PHKp7GWf/lPZoj+sAWE2vBT07+vsGIaXQlHIW5uI8OO
eORL/n/fXjfFP+mRGYOvq1AySOCmfYro8wyvRtqEdwqwnCFGZ3U648jCF/4eWHsR+HK2UhOV+6D8
xSwuFbqlHT9O53tMVhA+1/Lee6XmlK1fyU+5lgb7hvwkhv2Kafg2Z81nt1nhmoV1uFHVcrB8XJ1q
eAhdySqexJdPc8lI2VWkkzdO69ZmJc+QqHBAOeLWSTSCalZso6Dt5VEQVBhwx4MDn5zD5R5UIfay
OhMkSouE8VCfX5xMwW9pNqRwVZWm0nDakA1ZDyMVoZhYFnlvaZ6lRktmozDjlP8Kc2RZDMwrDNHz
hybuYc4tYZ9DicurTnqtmq4WEbQQ9eNE7LSvHQs/F5YsuEVrmpBPdgV50SjLzz4f9kZd3TubgSYL
mIxF0D2hv9ZHPAPLaw/1JUjSuevga511k+sBWrlUIMyC+S7P03xFBaXSzu6l7hr4KmIkDRT2o1+6
KU7yuJ66JsPMWb0vd6/KIoTCFpPq7ZCHO6v3x9+JdtTG3FxcG21U7DoBKdVgwKJ+yP4PUkWCcR5M
1MbK4CSjy1aBdYP9P9mlbGBeGdP1+jS5ZMfaQuAOFpu6nB/sZKTAbrMPdo+Ef4bZBirbcUOvexKj
eP0E2CRa4XABDk49SqrZHOm1bq53IXZN9nlwzYWqWIl+dyJHo2gyqISfnJ1vfGy00gwfbPMLUz1Q
5kIwRH0EKadPcwOD0vCdrKVpPe57uM2J6VooxjgBhAeTyVdy/xP9idlfiQVtSxgD8+UZHMWm1eMt
+DhSHD1eWooO6UFdC+zTwXGyyUgcxv92ZQ5izhg1bOVlrLLSmaDsOi6xij0qjOOK6lDLXV8EN1O8
wdM3Iw4llae/9Ua+WWGvgSPDhSEw5UgDeuCvIRIumMLMtHEZrmp6gDYzl0qQdsz9XpeFa/moARGb
pkaKeKWto2ZeXVd7ie5oyCIfsiraYaStT7C208D2iOBhPc4bgvvuGPNoA3Y7H09/GHszdAe43+P/
5aznWdmctPDgMbljn/+Bno0Qfd0cox4xNlhdTSn/zD3xeM352RLbWiRKFMpyTMrLXFWZ2M04UVLT
yhmOpU+BZ9gLaiWxYfc6p0ExZxvFG7nY6t1hLh59sRt0JpIeN7mWz4RIuJHQ/vuYeHn2rwRKUeMo
LAUB1MH04GCPXk7NIIr+kmOi6O1hb+AGNU6Y6BBzWOjOu69IZO5RSRpdC28/YZb7PlX2k43vRH2W
XgCS+xrB59I82UOy+VgPsCcdRRq6PSz6g2mMyMzrsD+dV1MySbf9A3A9dLZQd+8rtn/ojjazHTUb
A3ycK9dZG8xivewLqF2GYR8aVgrqhqifr/+mbUhyQTjvGDOx10ZQ/R6zpDs8+6rW36EO3Bpt4fH8
8WBrrd4HSK5smh4khjAN3ENqj0mHFIe4wTf00BiAM8Wmeqbqs1sS6ySuDNRT6xDTC0LVx0/0Nwb7
/RSJSNaklmgAiuPxA/SA/oTOsLJ3OlCCyTzFSS7+ahXFhuNSuBdejhNrzeVXztcWMtUA8FeWj4rr
bC3jtIP4tcqnLbM2+7St/u+UHIBfzMan23bfnXlBwFEmuI4/3d79Uxlw0H63du0gYRhNtcgT65fM
1n9Yzop6LeDXUCEFdigyJEu7Tu/GymwlmEgCqtJ/xqxEdCwauYVQx8Q/1FcbVkb11srSamu7Ogsx
iJFflsiSA8Zaa/gX0UY8Is1qcSv9Vrfuj9SKxoioH2E9AZutrXwzawdSl17XPwxJw0SXIk8dIBFC
dt7YrN/WVJHdDxM5KbwRIDDcU2Md5b63olXKsrESRE5WGpAL4KpZ9oSxMTXVYqOdxcn6OezmeRAj
ry32ck+cCSryouYY6Vb3DujyEg8LbhHSOvywIA1qdVJE6BtYO4RjscELv8zFoW7ctVwxM5bvmRtR
hAJCJBN77bNwHeq6fUqqh60XnHTp8dcDV/9v7yC5rh2Mq1thiO5i2nxuLf6VOCDFxAo2MAW9mjSE
EqT+GijlT/Pqk0ertm59GKeZ6gsf6gKJXWHc5rTGa7yv0Tt+gaMFdAWNse7vo9qcx9sBqBMGUMZN
x7D/Oy7U0gqcddozcuQ5JvR08jK13ksD0OY3PO1HOTL5upn4UAw82869nGG+TYZuYP6zh/UAhZZ3
8W6KE3WbPTHisHBShZwMJ99xAWZ3VWOfPeZY7l7OcQTge7xGVPv//VSVM+f1EbY8aB/SZC10ofVC
AxvQn7sVzVzGbMvOcSkA1Vb+U0jjt4kw+iI0+I/wiyFL9PlTQUGqJWSUyA9PdtM9L11JldwRFL/u
D+NfkQ+ftRWi2L3++HED18yeQYYp9NT7cpLbitRh3S1uMI+pjPkG6seTJZfrgB1TCtsrWgv/dMRy
7QXAPJ4Sqa0o3yXRU+YGeWyKfFL9KZ3/58nU4LSrnv4KYGgczMikhveRUugMD630rR/xPAyCDy9L
3mbXgw+slJDA2IQ9sTRUyAwEhx8NM36lJW1C70XPvodhaPu7ODo5NbGtwjHCr8+pH079HNRPbuqE
UCUhGO1EXSBxzWPnuKVTsWC7LLCIbDqSaUHMS1N/nQuhmBGxGko4mzs/gey2BIFZYdy/BAozSzPu
xmqPYGySsap05evoj4bTFBENTZ/ZBVi6X3/1/Tel4t7e5UmdBt6AxSg+cm8cRtIxpacNoNL4Ug29
5r6TpTNcM4TnIYnD7MSJjFWVUPj1g9xEnoGJVdMfIPeQf1ehOIzVZBTfAOLaCFxLWaeDC5WFg2wU
o9fDGF1JyTT69CExVXflWOnlj4wRXmODenhLCeTfwqi5kAI2V1FcgZRC6n7xjiGLCQxZxP+Voob/
+sde9RwIAlvCY2SKFZb58rvH6dVbHiYqqyLU5u1q2pJijPsreToeIu6S+qdWTNDSvJQHQHdu3x50
LEVYiaklUQoAz0YWRhXxQxxz7kjtQXwtSG/KBoe7n+EMWxqnfV+OMErB+gYMLkvgFb39goHgy/55
HrYwNDJSyfKm1iX4MqDRHgA6clXbzFwTDHOHjfDa/2QV46J8J+ftmtocHsIO1QxW/VqEhdSaIfd9
clCpvbupZ+osmCGutL258S6q6BLPHLRG3Wb69F/O8nMqeR49fqmiPReeuU5AKROCt8zVv08kvQqc
ot1PIG/WZZLSkXB/ey6CAg24BtNsHAG8qkpLDmUOLAdCNMhtYnvrxNO41CkXVgq5NyWAgbUBLK7N
H1h08g7uR3ON/Qb5IHZk8t7aSb5FdDZi2n5Jj1vffTbafssSv9qqdPm7frxoSNz8wX3isRSULjr4
/MEzJopaB1gKCHAJMHSRYF0ful5JfDDLs3AyZtuGmTvXJrof8NDrm4+FfCrgDYYtGXbI1M/50DZb
NgE5MR/HDBqDS+cVEUontFJeweWJ0yPgNxePD8spVqE3RKE2WN5SY7c8Sx+Jkv70Cjm7koCql2uc
Tn4s553idR05ayHt3IJLMhRO2LEJWJ6XvFdKyPjaa4bQxuYeCMh55JqNRI9R38lnY9rE5/I5D2em
u4hX2QYvuODOY9bBILwx34U58Hci7jnwWpuX7JRu+aPnZ1Y+J73m7KIMX5JanxwB86TUqlkRRXkG
Z/IpHOHlQCX4PebDeAoc7IijAVEZhUVa3u/d4mYWtskwqQRJVpHgg4SFTcNlyrWE80qPv1kPSsr+
055jz2AcFUnBxZqmymiY1CwqEKTI22LA4kQkagz+8JpJalUnbpRR6Ktp62AtTM8X4BGbMWhceJcs
bsmwZPPxNsHaKXd9+oBHLa6N0tSDzUknJq+W9q3Y1EydOjvGiNbv9wtnxHr8s47jF+90FiWedXmU
ZeFkM/TWsMS5xf87nrtb6Kk4Ifs6li1xQlGJ4NH+GoLEWpdpTD2XA7SYraAnYa/iAvJJxRiReKfw
v3MfcNwdrQE4LWULDN5lrYQ4QcAJAFM9t9m1rpfCwEeYl3n/Vh1dw38NFUSgLs2IYUJMcSHJs2jw
SZxCXqi0eRcJr1GduGehhf2El18e/RiNk6MWe/EXQBlxiRhCG0T2HMNp9rdUAN+7TZLbtrwjQX1I
4QN5sb2efMSeqJoBe+ZcxVZxT0TWM3EA32i2MVQkY1nwhwa1P5KTgj0RLGCupm6T5MzlnL0bNZP0
a9LmXBv6K6T6VwhOt01THxZozOYnX7QhgFApN1q0PsA8YMMmUAMHzrs1t5iqFOcQPoCefKeJKYhG
OwYG0Sgp7dlSs0GY2A64tXya6Vz/wdvugK3RZRxeMBgpFViqegkK6F1pGHyf/BxsO7ToLNYEwc33
VGkh5fLdEXgfdKZgSKkJS04VM6GO/RXA5Ze/g4BPBMBXTFjjUytNIFYreYf6vLz+ecpfzsz+p2d6
VEhZU5lojJoIrf8v6Zaot2NldPl47HW69sLUObOOArVflsPn1PZyndvPdVXR+hTNOL02F4lFdMPz
43Q3egpY9cYvvmOqumvAeaqo5mwFsj1AcsFbjiyLZ4JJWx0g0dIe8I5EepsYJF65WKSWm+TwZT+R
sPcBfXpxITjVCavY3cgH9GDbGFJUDw4559IooB89ByGJNSt9GG2ZbzkP209CrQv3LNvxMtvxv/Kc
tjQL+pxAW4dfQVq45icPdIewErAStXau3SDEIkdnABkhpMal0tkIGFltLqPCQbO4QkmBTWm/VSw8
BXlmQAV9mtjmQTl/mgwWIJLj5IYbg+TJJ8ARad1f19+TfiND/ErQwU7y8DAJsMisrU3gGKfSxK5M
7Z5Q7FCuOuhVUGQKV7GPduY8/T7a8DCQPUV5xGL+wYTyKV1Osd3XvD4MmQsYF4Z71HWfWNC0cFMX
bX1ESlRZRsOQmFJbvbgz3GZhK2M95IjZH+4F2NvGm4gwUHNDqMmQH2VjmxIZZuRRv0S1f67hhGdI
WifC5sbWOAFQEGKTnzovPIA+3aquJoqssdTnnkj8zBkaYjHGZvfPFgEBz0pD6EnJHGWrFx6BD+x0
xOsDsVSPJkZsHtbEzxDJFDZ34pPBtH4s435LRyg38GpBAjrnVIz58AugYEj7o8DJEEHCGK55VPJC
aYu+BN8dVwdaqY1XGiULNil7jom42JKkb1pAf6pv9mD2eXzSHMnOnLzwf/2YYlrYzSvczQr3MOZi
ABzO6d0bzTd/2jjJZw01Hbzn/x1Ydc+WrPlkx2acz5xr7plB78+V3uPWiWPhVuzazbiSrx8Weq8F
BvotdyMoltQS05OCfEayhSet0ts6OK7+HyxhtOuOPLH0RJoMolQsAHlxGsGUAhLQY1vHc9mwPEte
lKySuMhTYyq4gL0qcoH1/kj9TH8TjuFXhlSHv8a4M4eQ4VaacT76UK/jiUjBKxIIoyyVYNPQtj+5
z66NvfGDTSRWbGKMq4zTXvjlf4XRAvHaKcPI3ip1E0Dv9LaGWO7M9NMbtgFkbgyJfTuCRapYdrfl
/NxhK/CTkUJjtQUDYcUmSy4ddTyDUPrcB5zdrBHjb99UzYMgkPHS/3ZFNSButaHOA8oR8xXqYBXe
fikevkb2gFCdtOM/inaaOAShdJjllxmSvqcgznbAIYLKdcgL0SxmDHd80liaL1VuAK7LmVDMwz4H
gO9MXvv9z7Puynhw5PCG5PdgxPHNNUgZqsIZ4+g2WqddKAWcp0HXcHYHN/6wDJSO3RDJPixqA6jQ
BC7qiCvUMRkisuqbbe+Yjvx/2I8zpJ8O7Co8Z4bB2HJ5Tfauw6VJTHJHVhIxj9I+idDc+seA/4v3
3/vML9EOsASlleLec391eJeWYuUm40D/eCkuiiYgv/gkrq7MXl6DT8esHW5uX6CORzz2GSz48njk
0SUAPjT9xjbt2KnCmlVzRpSzQ4V8tXqwJMyoAsNgBsoKBJNgLcn4+89BIYfFTq6n2eyROXlytilc
UPEh3pZBmd4Z2zubamYQldUSQFzl1IS9oUSdvlFZAv4ERbIub1KmWRU4whaDZmCPRZ9W/ApkNuup
VJb7KlKhSglaga3xIvp5ZWu16c9RHNtnWNFI9HSon8EK11tJdGYXWzxZ1epyfe194a+j9vAO6Klv
9wwKJA6LJhYC5adA+17bipeY2louBQSFEE5yi7wD4Afp4+Yxz0928LezKh2gr4mKE+Id0SNU9AlE
Rvt6tP5t/vhRX2J0HzOaORTmvN7q8kZ/shI6/sXXw7jCP8aakstMfMgsgQEah8QO1cn+y9zaPh8G
BFsXfD7zG+0K5p8UFRZcO+5M2t72H11xZ7YPnuq1QPUfguDJJyr2as37K1F+H65pwXrqd2C4LOfm
+RJwc4ffKCyWSWhoJtSVeT3nRNMOVezL8oP+ym/ZpOsPT8dXYIY6ygJyZxKr1jSLYVdySGLpizhY
vdevXQlBcue4eGta7KvWWNZvhPgF113VO2Fx55vYOMbEqEGwIgFqWDIXc3cZ4LQPoSBSt3m34+Tt
9AjAuAZIZSuPtfofPi/kCRg5nOLDO1rk9PZ7kBZ/5nKTqb2J26CQ/OtjA1KkpfuDy3gar8Jzy47b
Tivl5BtPV0texby3Z5b4cLYMUXNqxgSW+y2Ic0D1Rxh9VMTDdrAEKLfP41F1p9mYSnyG/iSVT55h
4tygrJTvP33dRxKw5XbyOvp+IwooEJ3nfA75eAp/HTlkYkNxpLiy/VcbiTyFqXTB/xHtz0dWaDOE
g14PHXBRndCQMfcfur89ZDC+2mcoFqaMzhUQboNM8Do9RVO0zQMYigMbBe/5fJMYXwOKJqSz4a23
76GoUrL0hQf+eP7p/qnPYCvx3HbPkV8iuTFe5HYBiAscftDuGmaj9lNE0E9/1NI26DJf0e2B24Jn
N3daUbXmj4Ju5ved997tb2BAuh5pulxcL7nRaJqcLy0mHUBvgjldJvgv+b03enAVTMUcfTVjzfmk
qsribYNeUjDk4cyR1YH8mazj7oRyubJZK2CTXmcvytWsT5U8v79NKIaj+Oe5pAuFfYxpjUphx/t0
7+byYg8600Ayx5Rw+tCSEhZ8BWQJMqEompISkXXMCykRPfRmqJlmZpSbLpr3hiS2vzypaDN+gF5A
36CzDfUBggpG+fBLgL7SYe+5I8VJmIhKLFNwTlsYmSrkWc+YjdMnzK95PLkAFE1/g6cz3H1vmGVj
1AmDwHuzazDWxFdkE2hLSpD+2dXRCa6vqT4LgCbNZV9/63wuSkMIRrpOSq/PV0eKQNKikHZTyyoo
bxoZwh1t9om410iugvrL1GQKhJzbwQurnHng9tvbvO7tJif9N6ewPEBgfWoSCoshqs46wDHoGFA5
/nCri+dWGinUqeYMgi4EHuLK7CyKQ/kCgeC8JzABmyA0o4XVptjNf3w6pBX6Q94OnsffsqSCCDA/
CjH9g04DDh26AtBpB/ES6cXYbsDWxhX160eX1cMet5etyyW5oBNVK3Bv+2gOinug8lj7ORq1msTv
Ixn7RVehIpCHJ9L9hLSfvM+FiZtdkOz/TRXg7khTk75rXPwDgtV1RUlnXarEHLReJM0qoLdOl6/l
e6wPugkimyYw532AFIdIAEiGsGZ669vM0178wY51CxidFbyb9xdlnE7xdoCPI5I+j6xEv1qCNDxG
tGUUAlDcXx6EYi9L65nG19NFKMJ7KK6MYFCzL2CI0PavInovUAG9/nx6vwYD+Mye4Hv01pQiCSi/
lCHLPDE17xjxynAB3UvC3pmxFK/FPy+xAu4xyZc6SBCbE1hbxBlV9/cO5aZBPsZfwmsII/8YyMCT
+PvsfkCeePMEGvps/GiAOnARRq2ZUGe0QJxe02XKNe0YqinYwoAVAKfzt76QoPToY5GJD9C3Gsmy
jPtMV4UEn7be+dhrojf2HV9ldm/OPVoFH/QAkEbKGBtJTLUauzaJFRJCXQx2+nM4IvVSrY5blmY4
Wn5uHt4Iluuter81RE8pC9ak3jY4Y5nZOuH46nKKt/p13MGEZK237Yck49HbbTtq7b+njdRtbm/a
ZA0GEqIBGdyn+3cs8zm9iUJPHSoecu7zlbMB7HVhX9xl4mmlAbXXuXq6amAdgqZ4PsUY1ox70st7
5tD72UNZy2OmPFHsFcHfKmRSjtX15PIIm8LpH7ra7Saz8KV95+IW5P/EtqAmZs4fYpGyDnoZEwF9
0d4Txk0QLIVZBS7PeeSch19CaJJGTlZ0fY6tLi5JTnYM2QjtQJjVriSAdn5b4qhH1CB7CTjc0S+Y
ebYRqObXb94v8ZPpuxTtQ+Jadw6MSR9EqvZqRHYKEDL6jqW8SXkrbvb7F1gBa/kRaSaAXdmc6iX+
5pUCMhxdOvmdknqI+sJJfTjiRI7mArqCC8CGNz2vT2Nl7Hfcvk2qOfA5ePm7T5MdMRkDNuOGyH/O
B1oyYalN+YDhmjQKOk/yTfHvDTGuiHEDWivexsnSK5nOoYizi4jEsWtOQgXUh9jkPmlJWAxYbmjR
NP8IOcFKg+OoPozeuRqXFSicm6t9cOsaYybWN0w3BKqzmwrUv++SsLOLlBJAXH2/KnezOKzpOYNP
ZDtCEpJYc0E1AcDqT5s12ZBfa7el8dGzg36GeMNw1Rcbx1yr0+ZIrMHYLAgZeEO6UUYwKeFCXJDN
cvRv9zyLg9+F/By57Wy9rEJcLVOC7cddG2hRVBrBTByHk0Yrj2kEP4eMjJ6yFv4fyqtzvpNqTGHo
Wuf/DUZEwiid34Ed8sMjlx47crC8PW2n5Mc0FEQprHbSuGLBBSGhlBvg4kdqlS9LctSap7C42TfO
sG6Om0iTXSW4AvOKhWWIwi7orrX85BrUmGSx7dhCzzXHEaVTe9qrnzTDeoCnkGlA2nHEkxaLlCZ1
NmSO4RCu/+94+9LKg0aprpFK4objWujTIKP1y3QnFj2iChF3rdHHB7IPzRZhE3AAHP5Ve0gHVdH1
lMu8ULUmNUCr6YU34Uq/Fw3fqWl48RnZ69/CyWrVs6OXiTGo3qx7rm5G1iLt2Fj45tgUCisJyO1n
l/nF8eJWgEt9x0O2p4Vx8YOThgm/oxNpFzglS8TpHVJpuJOhIDUUku+ybvbFR9GczifqwTY7L77u
PTHwS3vxeUUn+8kQhy4t5S1GgtnhZ84Cu23jcnUbj+7lneDTZSRF5BGDuzVMQ+8QXNdjgWKM1NpS
EKMaKqZI9ToVZ2IBs+sGvomkcgUKjWfaigjUn+aXGRhYsVaClQTbclD6c0ACCpCR4zqVbHTggxjk
ITchCmIfWfA85/om4B5Yd0/rePl1M7oN5aon7J/na16RlA4OyAs1f1Fxyu1RBPXs3icbCtHA44rT
5GBQ6uY4VomTa7vXybmG9xBPBWNwLDgyAswzcbUnLqW1ScotznzbDMbcuBytPCFulXtt3zrbxZvh
5C3xBMeadyo7u5mRS0ARI/ABfYAO7uMz/9bsdnNA+gMhMvsoZ8wy6+vIrgSKW8/MGE45Cs0lHsPt
ZdiGs5/gWivmfsagipVy1LRdDZs37ufEGAtcPQIJxDI5OIvJ+N7u29V48QEm6tg2zz/kLYds0Cot
wPQ7NaxpSzK730WvYmhZJh5/AnhxlqEyEN6t/PgY7hshfEOni6IsXI7jFLvAPncwgYuCuE4Ht2dn
8sy1qsER+bfh3Qhe+Cg3s5Y8C5c8ChiBf6Ucrtn/r0hVUpL6YoJoxyfNU4ESnRlsKPtRS9pI16+M
zFsEZZVDgCtpyxn15ikYf05uA+6td6E58s2/MIK5cm2SWPdad2GC+5nAU6J9VdQLtHXIYcJFzAnr
T5+ebMukeLNl8x163aSMAhmIuLPbkcgHQA4Yxrew1blc70GUocPKvGW03Uznn6VayNwnv6tQVdbG
NCtzavejpD5ofScC/dQZY85cuDbQM8CrltHFKLBa84K0Gdfxo6CeOIBfQUcVH7/d2/CkinqWtk0i
SG8M4VklUP/9GYAVdySkU385n1v5WTP/7O9EDTBPGQEP3unVjPJBDB6eufzxp4qTbZOlXNbAcx6R
dScpt5C3vgcroGGG7RCpbu0MLdsW0swDrAguHpXcuwcwB1Sza05Cf24xu1GLd9unoK1+b1n0ebP+
74uVT+E0Ucce2BkwP9yduBlGQetTjWH/Iyb425fymKLhNfHC+/VDD93SNcNh3Re/0NA1xlt/MimE
qHnaEfOuwcViwZNNXoJAPuD9aQnjN0I1awOuf3LFmt0lqXW7dPL8651U9i5WtTajpn2GB8WRY0J4
vT2knMvWDsAzHcYYZMrZH+cj4ahQ0+HGgRhV6dHmQFpwVzw0qSvTjHg/ja7gEfK08FeiTZaAFqMY
Ekf7FirAyM3EGSaWFLZHyl5t3vwQ9fa9Zl4ZCXPuzwgkcjJbDvR79d9QMFanxW/vpejISXrSIVSH
zfG5AuA/TgstzkV6etVao/wPVr5hO7YBIyM+t9Q1BEWMv+jCjktImpVG/3ULsrTWBr215Gbki0+/
D6ijsQz0/0LB182oDGHYfWhdycEM8lJpW4rFI0bRx9tOJ1KvRUcP/kOXos5ok3cFsgvqBg0HwmuN
cmAk9ysKpdkKn+Qu/RXJgCpSSFX7kXtI35n3bXKo8M/mSjSx66rcx7XrdJKhk2bJnDqEI9nhZeZx
GehHl4zvaIPkV/XJLQr3G6eyA1gJ14wcul0QrN5vQh+XSBy9n5Zgot8A/tkZeL49M8roLlw0Rec7
sBAgi4LlOhBGZ4B+EqkEfahjvXFlB0lHg3bFXRvKIISpm9KoIiGwH6WTUkdn/5T1ZhxmrZr0Ry46
m9BXZdu9ZkzIDAdL+I7btBIsFeOQHZwIDPKVsGV/yBaBQRoYpRV+LhjokjW/lwmE3+3D7S7mIT65
4ffi+kQpDEKmJtctMHG+mwk+pS+I4WnLJu2pZSrnnKzDtgOIhDYblvOoAE/wt7+QuFQpW441u5n4
D/6S9JLSEGMLDjSnO61cF70nE9ko9pkyigTdaebL1CYhf8Dr0E4Pn9oqQoCJGkGjJUXy2UkMjw9o
s0oLgNALgn0TEXj7rtkCvtgSBVZrZCI70CXhx8A42xgCZypg1LHR8TKw0GJzZaRSegVvV+yWO4R/
BCK0/P5yy9bVcjLYx4y40t0bperBQHbuuYQrXm71XV/7CnC7LxwbHUZdRFlxFCdY+Af1I6afwuhH
mKWpYH5zrd99FKB+mvTCLCJ50fvCQOxYmrmOiypq9oNGjD3+eQdKcXdCS5jz4fRJUcyQvit4z8yk
wc9kjoyklzwMzg8QCFBYhhOYKbednS935n/gsaG5jZgW6SD973hleYkLIHp8eYKyS7cka/PGpLqb
7K63Ah6WZDCNYsyyijiMdTR+OFBFCljo8dg1+dN3cGH36Ho1F1bUVmVI1wQb0AsEFMv6GfZtY7Jy
l0G3VOYk30/ykhGW/sLcHg540JA1Ds2zy8SWEXMDetABWzwesHY32bc0u452Lp+B8da5RNp8Vhi8
Ufjo3wZny1K35G4cqFwKwvlLTo5KfIT+RomCMaTfQeMmE4e1PcL3UZkiRkz659xfo0TQKs2Y00M6
ZmOgCglHqLMKIGcDx87Dm1xnR312WrRaF4Je9F7K3pGbo9kMvq/kG+E4eoMH5jSBLyGzkWapWtMt
DdtZrUSH4LqQdtE0VjOE/muaJkWvJH45W0RBmqVxQ3NAWOauCibJJihCcR9of5oMic0oaM5+vCM9
hFURsF3/v7anLNnxWMrc9r6724ykGiq0uBT8Uh/mcOds6kYEdx+cxpqhoLwoRyjjbjTYdLHA1cfr
f6vMroWFO4aken3CN4SuOX0LcYhbwdwc993HvL9gtb5HQSJDJr0WrZ0RuxnGblCzaCwCt1fQC/5d
YOpIgRYsuS8GTaAkzdpE44T0WU2OzhAPuvJWefhF179ccfvDZ5hR32o0Zvt7zsaW/jIzh2GsPXQM
GVDs6YClsLIWfbLmRni4uxz9x52zZiS0znApL96eAM3LrUZRXp+yf3TCuEL4h/QzCQSbab1Ug/+U
qU5emKInLV3FGg0EEyqyDhdLMackr960A9YooODW52Yf5xGzQpehae+ln99LAYP7YgWiSvzaZ8Qk
efs56ErqISGjxxoBk0I701en2KvmWC32Pj8QJ5cBq88pHBnCZp6S4LzF12H5Ms6py82gkGszHO6H
MnIyel/toSr90M2dARNc6I4PFRjVBe68+43pBmOJiGD9SmmX2A2MjlA1/PAOoSz4pVNWkn7oNw4X
Mu5UYIPMKWh9x60QKbIiWjz2EhtD6SqDUwVXehNuVNu6uEwTliF9rsBeRenw92+LMkvSdeYif3FB
QpCM05FC3dJvOdMbp3GGpxwsTRUNdrW7F2JqrgS33gWwZxM/5yp1qQxnO+lGQnfDcO/a40OVrWVe
uX6x8B73SdtBUqOyMK7eqxJToX/fGgGccFMiv9fs7opo03oKRUeQ9VleDcIhV1wLVEh50cM227rD
3SILRhNJpcVwyrltme+osG3+ZVz6Hx8ZBvruvv5i2BLtzINazSr0tTa8Om+00bmsL1vi+pITv3r2
ExXpD/XuT6ertX/qSs6lMBUm6aHyIL7e7vV8R9vDVubdCc/iO1d2sOSsRKQQZV6eKHyOkKBJLGk6
BPy5IHppsV3ZpV9Kj3H6Zgo0F3V4qz4ISy583oMLAMXXkFOxjFG6witGviFXt3zPNL2767V2ndQZ
9HGMtjcPlEA5vch7PjweQ2VDQdyVxVPShVW0uvienZSV6/KQbnEQlvPTH8C5ziKn+t21rWuzSpqH
nU30XEcpnHJIDXfr2J3048dXTfXvBGaI7I7soxdOA2/hR/btlMeJurFZ2qDvoXFR0h1CWctb20SC
ArU+GIrkWbVv4Yb1P7rM+TiFC80/m4qGqtgBI0RoUNhBfkhSnsdBVzL9RfDa7gwehF8tO6IaPolY
rat7iJ596eWxaZCaccKmXB+Lvt3AJGB5XHgv5crDVaFmsLbApdkWPbiFYlKfrl9UFGU9U7GG/Hdg
ZbMLNErr1rZXBG0Ld8TqyxDxaAsTpcADwmtGMvEDiIokiltXT2C5O19xeGKXB3jO3DXUNfIPv6ZS
ap5PspafbFQo6vTwKWQIRIou+kiF3Hnpi6v/Z22NPtBPBdjHZo/dhUFg3XDYpn02QWy0ft56Lsh7
8qxpHny0B2s+XrKOn4Gbhsv+Ns2H2bINRSzFG27jgXPtkpNGZytMTt7RU90jOstJnmYfNSue42cH
KdTo+OyE6d16SeCE9yWKvR0/Urtq0Dnbw+KKZbGvL+EnyFICcpdE7v/gPaIpoQdQ0kHTjN2BOlC+
11oN3FFSB+ppbIUidwTMRJtCFSIfPYklKx5aBe6L0hqVw0F+3sTILYzn3VKCTEWzI2Bi2defWwPl
OxUsJByJnIUeY/LQa7oiAlJjimD9G+lrcCnn+BN/FiJyl/T3+wFml4TDhKTzkhTPzXiDPYiZK2/t
/bYIwwapYklieVizuztwej2cTa1BLN6vf0+F74eOxIURRiD7/zr7YbxfUwaygp54CCgLRG7PZnnX
u7J9TRbJrcMuqm0VmhivjbxnxnrDNtmGO1QuCVXmqX5NzrvaML7hPqcWvhYCAyhSs1npvptAAybP
DmyudN4zH+wK3flUUFEUUEjlbXKVyxRro+Z7Zvct/ejd7ko94jex4IfYhwDOyIu73UyQz7tTeO3N
vlhFJe7K0nK2HdZYe8hYWQ52DKfZGYQaam2aUqdgpGEKMKuJjClagBfbBssOjoXum4sapfp93j5o
A7ydvS8hdqC3NSmG7Jo477ANhmI6ZeR9x2QI8yPePnt2ekwTg2DvVQFtzi+pUOKWUaaBydro0RO7
c0h5K0kRyUCB7JD5syw8iIKwk8QlocA4gFj3ayxgzaYttzKT6M4z1gbeWftC/24NrojeZjsdavyb
PhuFYL8IwCavoJqb7Is8bY+Arl4IyyLnD+ty/eEQQlajVttnpXX3yRCyjvK9E90AMt53VNE3WWxZ
y/kF2/36L+gF2TUoNKleV5r5iwO2cWrrg86VxwXBdw7i8SYKyGo0OoIfq7pA6vMd9VfYXCXKzd8C
pANXj1LWLegyZfb1V0N5eVGqbD2rLUK4OyHxiZ0ebTM3qwVW9rqH12tvzUhJrjRr7YQMGGioDrBW
W8bCsxILLNfFnohD1QpLyrE52Hg78BWsb8RK/OfuDik88gMh0vLfs1Nrh5ZFJViX5GhLLyNesRcQ
MHXLDl9f5ZmsuarWKkmneRK5QJozO45qjVmhszLuJjsTaBs3cHYkUCRbUgdWAHZeirJY1tS9VxeS
PlxgI3VBv4+GYzBRAgHcphPNOeoigi+GpWOi6rwZfigF4d5UN7iqLScg2JUGkynoG/5nHP/9r09E
PUP0804raiz5niA82tRD4BSa5LDygGf8+OjB69WDrcF7+Qf62bNd5jEygKBBv6ibxj8C2FfdyGC7
tfvL1gmzD1rVEfr2WkytvViTIq5hrAnURuKvNu/ZumweCitnqD5pM8NBZGxNmPAVCMn7V7YcbGLb
GxUDEwFxfqb59Uh+H22UY+0IWZ5eQUUb4XBqClMrClANUelqKcXr7LVa2lf6LGQ6j9pUlbUApFhj
YrvB49eEs+FQKYPQ/TuqlA0P0gwwSKjPioQPC5B4xQeF5zY0MGMjhHqZ2UdylAqtrV+aFiHXSm+M
wAWde2AOyxQ2SsHWT7A3obUfiuxhBZ51QNjNw5mTt5RK4kTssUtKodNJ1YO9L+WozhnEeP5+urju
JMMx5UkQX+zasqNBcQIF+36y01W6jWRDXxOMGFKC53OPxJj6l4m+UZreukmZnjIeI1H1aFW/ls3m
D4DPzn7nkX4X4IXhbqcZFn+bkzSQQfZhq3mw8EoQvugQ3e4Y828kdAigy3LQHjxkwaYEB+Y0ImRo
vRdhcOh4MIYeSaALgLf1S1R8FRTqrT+Mu9pGGwgOr3wRlXNQe1r4lfCTZWbh9++eeisqj3DZYMze
ZtvS3eNqYYHFzAVYppe/GXygk6TL0s99AinipNedwK/Msc3kDr/F3lH6FjXd67FCrFMMd+onQgKG
qfl48ft3hn7EkKhgY2gEtIG6FkdvLtTrwy/mhFk+9NFG6mTefoC+lQR/Nz23Aut0Igp6S8BdQoHK
NHsHBNgkcd6zcmjEXPs8FlbZnQA1wJkbYt30OCfOHHmpKgJHLsGQbaKZNcz6Tn/0C1roih1jf6+h
CNyhrJultg7pRGqu8i17TdqNW+DAmazTgvuXttEDs9GQ2w+E2BfDXvmzstFOCNZ1YmuGxaYA0pYj
e7VIkIdqq4RTDZ5OYVC+hvJgMZZzLjVzchNFwyD371G8ZI1pae1lBeHQCc7mxcJ3B+JINdRp9ngo
yM+qNf7gRMw/D6+sXXSK5CpTQ56MUNGbQrA2OPAh2bmpfvSf+Gqdmq18HsaZYXidkik9pICbwiop
sW0b9174sr6D73K+NT4BypiviCoXQl3hFHDeGDNdwcs+pMsvvl/2NtvFldl7mD7tgGQDHhe8/zLA
Hl6kKb3r+xvcBDyNZCSgYVc/vBIHhqs9vNTWLYPbT7Zr/gbcyphYl5iNMCeA4+jhG5SW8UIwsgTL
FnvceIc+piZUHBape1OhBUOLwmRlyhKE3+T8SKefc/i8tMEisK9ldbPxwDjqeMQq91tnj4YHTBNI
2heELhVf/q0EJxd49jwk/Z0dqePxRNGtv6TT+kk/CNy3khaYLo7B4mLJY3e3L8XhYSTJPboMYZpz
3XE+DI4GLguUjh9uQStcLq4f2RCFYEeatQQaAjkKGosMNE1+NqZIQ9t/pe+iOcQoUMje109dlTJ0
Elei5QU374qsdgXAtwn+LmwS1InNAtDnXpP4MNwU6q8VhwealK12Sqjs1ICVQknakjqJswmaUiX1
6wJq0U821jhZq3A2dZGoReClLsJbjnn85x8Y3gQbBuHhRt1EsTqsA+8zNtVw5VdQ8s3Y626JrSIL
CaeFMac0cHYDbz/GbwdeIkE5hJ31ClBV3vb/SD6KTNUGPGzz1soxE/de7CCXMDp2ySgB/+GKxFbv
mRaiUVYbvxaSdoTUTFSqy4gagffxc7z+Nk+clMRE0lXBcy1f8Yg+KoygOCBfyBeWKbjwOzBkUetR
omIZRQl4rH7fd8SI1xhFFYYoltUzrt/dpejZRP4S0FsBBKXlEZlfbkfmAoxtoB7wAjoBffiDavVR
/IiFYV858X2bMc7/jPDPFtnLGknvT9ll9atIhWdgbzQcZEHa6olfQtYkLVQcUDegLkjglNbMH4Ur
BRGTsVBJhpvZUmowmxMALVDgmkhxaOE+/gPSsr0rY1NKs/guDB59ILLukzQejEnsGbxwZL9x/B62
jh4y6Eyyhu/yXUFsFG4yftdyO8M5sZsH9fvhI+pKYUNWCVuDI8yyR2m3+ebskQpZUW8NKWjoYDmX
SmW6gVgvf08sb2wr0ptPygYzhQXZgIjFLaJvSBPEzrw60O5Ij1rLXvymPALzWrgpy+IrjmpI0RcF
3INnYLJLesatKpVnXj+t6pkGe/IRl9gaqoO0JJa2L4QE5H1hs+64s5tIUVFM0IZ/CM5xOaapk+PV
M5aPuq9jd5ZyyyXG3mAjv6NazRgQvrmgpkuCJRL61SF6vGgB/LZcoJzIXDl9E8dtzeR7hxQ+F+gC
Hn7sj9bs6k55WiQl1DxHSQ+O0RsZ6ncvp9qTlCBUv3pZr5HduX488kDlqBhiZHhCtnb2NEBVG95l
2Gst6s0HjiM54ZNY2LyZQfydFO4/qjqHADUm8HFJC9bWT9lXI2igA7LCYU2LuHCQFZk6Sptwyrhj
kto3KrTrpfhC835CKL8WbbVxNM+mU/GxNXnuVqn/eX/t5BeaL25zH55ljQbuSEupkT5RogLANCK1
2r73d/2hnIWtZpYNYRQ04YaC07zBPNzCNwgJ6wT2bPtdpjhxgrwh+LK4FHX0MVCWFSGvACcMCJUG
QF4Dj9V5mtGqkricJoq/a5DMvRJApxBQw+D1rEKtmRXA6ZmTRQzyUa/GVLxut4xVcFXDKHCsUzo5
QKCxmd+4lj6ZmsV8w8mjzoE9J2ib6Pwf6g7ouII3oI1UEOKPqTK5uuvd4tZQo9ygl1ARY9iBKP2W
ZS4qql7ByJiExbsIKe3ejKkmiZ8UTLeOV7BcC6hUgXeKq4BdmhNRptfbVdlvIg+uCtdf5YCHBa6c
4zDF+ByRxDvUk7/d1zbAU/lwDGLiaT4duglGQFiwN+xh1Dmdn0LOkwm2jfu6aqtZYy27KewvILhQ
YMEix5xG62ClzYNmu7A4qWQoaSp+IrZENFgPJ66xKpylMiKeNVfAYYDJO9DR/vUuQsxGkJZb0/ym
lRQjvg1mTTzDZT7Mm45amu6JLdYr4MgiSx6xqjcIzQLzT+Q1dj4Tcgom4bFhw+gtlNIhragrpVK4
VdB1ov2GIHI+P1EzrNIPs6eeXIU+mk3C/PUbhjnTTIRCwdbEeRP5CRSfl2FnM0pfq2oEeV/EYVeq
zycx2nHqKRqa26Cc9VDIX8kPmyj0MqEnhc+LUQjd9jPdskND1SMz+rhGsN/igOmJPI/+QNMEwtcL
KY3ZX3JAK5SsxMT7zBT4NfdB3qgH9LSRQ9Kl4jOYCokiQHHJU1ZnjDTiZgIXp92gTrqG/bjJS8jy
YMentbfnob3kSS0cvhAjqcIRqxDeIB62PV5y2sk+Wrpfa9oZlLwVIL0GfDA702SRuPNrjHGffKxV
lqNVHxPBhee72uO+zZ2NMfoxEIza6w6cHgA5Gy6D3QvKrQYEt/mv+Srdj8QSErxkAQM498bJS8ja
PRMnFpXen2plXp5mQV1PYbmBD5zU8mURyLF8/MvwzecqlQT7BlWcJU0iV1wBj9lej4uTrjs/OrI6
28EcGYNZh016iSyDeEUH3oTAVPNvIX/o11GlkJdwJ0cJ3Dv06bAnQCf62MA99NjW+O/kjKi5hzHW
m9Ko+BIk4J7o7TM0PVvkmjek2xTFetx4a7ehLiu9lUMLcG+hs9lK6Vz/MBrHYMcj9jSIsQkwxT4Z
fLtbTrorfdlO+cVYaLeSwD0+2iiaQb6HgDF9FyfPjH7uLYZZr/316LnDNVTcjrNUwHPxQAlxTlB8
/Jf9y/ZuKyj3ssuSv11//z6o3LMueLmrTO1f/JWLkSWtZfbMMMUOmLK/aVLDe33nOQorv+j9xOx+
PGDx9pV21llT+9J7q9up6nMuKMkqulXQsZhOnT0Jfj+NDqIg9feTNPBObtEMRUHbzm4k6CuJxboT
d9c8uGn4Eu3zs6+oOfGPUWlQrsoDEvARjoZPSTuvBzM7fB8MMACprfqyej3LkYxBDIVOHYeuEDfl
Xkrr+7jOvkD3UH3ExwonlqrxGOXThFsSY0DloC5qLtGvCdSjwfjDxfiRrFr2kYJtznofBVJlSeO/
KlFEP7SmuFpL4y/24bjix2PvrHn3HhnVil7qDxEZv+i7fau1NX5L49IYkBQNGpve+ui2jqlA6xbx
vLaALB4qm5oElI3QWk1hq7p4p1yfZnuP3C8TcyoT9Iq301vbhC5+rxDDWfLeviCSbaiTf54wowJd
iNqUicQ7/1N+lb7qcOnnBEM0Fwc+whSfwVywxJBXXg3rqVm9Ek6c+YkffSPzo+yS+ngQrNz/5lPr
OTOJjoOxOGoKxyiqhZpp03+hKPXkcvdY1gPX6VG191Pqw572Z1fpkJHzAdcW6U848I1enhRvzTn4
WptbGBpLIAkcmUxAyWkW3WXQmgWNeo8bmFMPaV+AChc+KuvQgbcu3XDbhDv1M0CQXRRtsSHdX06n
7RoGHcdvRX8/N48jMwHmZvVOpqs7Qg2E9mnRR4T04Ib46n2DDmMgLAEi/5vSWNpUg4X/kO4x7+td
M5rl810CMBsnUmS8uiIMnE73vYzaEyhC7CILtxTHFtd+HHm0iUdj9Eo2435q7ZZ6YC4SskSedMyc
rJosF1HY3FSmxr1OI8D0tJJy9GkD7gL1ub8DAw/G40EmQA0Si6rTeEnEu+GmHceuDWF8OECX0dWX
ebZXsRXPqpq/VwOQr8g5d9tXs23e/JmPI1kW3UNomJ8hrmJ+qcNk4CEWjUYcK36OYL07BHO3yWmC
lOatKKushPSh+rxnQxWSKoHvHUtBp41pj8ekdVXCKD1ixtY964mU1PidXXY/MULBB3ub1uthnWNR
phxLabQUuLWL0iXZDDX7MPcTb2r7ysAXogIzEBX/YuOLPBdzenW1uu9WlwB8KfT5BuVLLp2cUspR
R7H045VqUc/3uquCLmTdDByw+udURd2oWkAeWnI+LDmL/0BW15OfBY38fYwHHHdwNje3geanbGbA
SS+V71fszuc4Xen28l9nmNqRiftwojCgoQ6ANtFMEssd9TjyBvha+pSmaUSVHcP25H2UAXus01ZQ
q66KaGYN2mECpXUzCWWwW3m0/riCZ2uZbeUPgI+naML7qr6a0bycmm1ZciUngS46t8pFU9KDS156
8RCo0/542fsqFCO+J9/jIWoNpFEmEr/OLf4MLFlOi5JucVdu/XWqjidvOHo6/9VnPFhnOL8eGt+s
1dF8/1dnqfeRyCjmoHCelQ7VKi3QuMACEEwYaxRHapozoCUyN9t2WVXyBq0NyHsy6nTl5lzTrRLV
JpW5XtyxCILAOsfn8nfPQpTOHSSnSlH2tGFwLf4FwXadfoOKlHeaCEEcn9irWWrNZGO1prJF5pVF
STKGq4hllXqUSCqXlFHsM4ahW4ojmcZ0E204xUi+9BVs5AzgPgDfk7mI0V+WoVEoiHBfBidv/fR+
+Jjf4jbrPWcG23x0oLtv06CVzCT8MjZbzr39jDP/20E5UWf55dk9onom+LbQLdJx8PrVhHbrSCi/
PfMsALuQ09STuDiwamxfRonjwSOjt9U47Ifk+pMJnKXjyGjZqgTCGtObbHHPmhHgCeJZfE0mIxL5
yoBNmr+V2hTf2prAjngj3+9xzOyJ8iTgxQw8LejYoxnJEDMLEhn1CL5N/hoQ9nN7RCvDzYCeDqgE
ocCAl8oX06oh53yGqEeJhY/qKtTOsC42IuAN9gP80R13sZJ2BHcSqsBFwWtQltpK97GwKJ4MtvBt
Y+IR4VpHdkebBMlCTPntJC5nHWKxqfr8tk4NRhJoOuGehemUAAYAFLxMorakGNDxRsSf4nO1NUl5
ThVVZZhgRfPq3JmMNKRwmCQ7ANfWROqDOSWLN7obcuhxrf8dVuIFNB1Pp48FYB9H18qDEzyEozk1
xWXWIgAhlJ3cgXN8xot//lV8Dfob3Tt2ISRyu/CkidgUBk9cBiGifDU/DkhQvjmIFz+XP2gLJqux
2nq+ITpVDuiL/LC5fUt8VMZG3AZ+IJljfqSlkQuiaTmIEx6ZXR4xXxTGIMQRUjBlP+0Vtta4+WNU
B1QaAkM75anDLNGXMduQKxkSfqqprKfbBmHntnpeO4uo+05KM2YsvYR1GMS+xRZcGdVolsyoWyr/
Pp5YCkvrQM4fNAQxKP680g4gWae4M5CVG3NVuUpqV+S5IBIiDqaV250oISydSj7teWJ6lArf3QmD
iyQDZBu8athCDxKrfjssOrE0cqyAuYOew1VPegeKBtfpFuPZrQKcLZNKZdG/cFjLups2cvfQRZ4j
uUuFjGie6m0S/doOyEup5esE2LevWX+oQVXWeEdNme0BqKmWs0WMeOaVnpim5Ia7bx9y8EFofRY1
OH2nvwtrgA0l1hntzxtz2lo+JqyzgpC8eeyXx+U32ZTtUExZJit8Z1h1XyHzk5FKp3QaXRXe/LUw
eqI+oJgaU5a/pdY6LNx70hMmCYyM1TnNkLynyVC2DzqJiTzDYu99GDWkGPF49bd02u3FaC80notP
rq+py0edIwRstTfpraja+G0NsNWY1JZ/2Sxno/MErzmpEGVjnUcNXAxCSNCL3SdJzujX0P6kDT4W
Klu+xOLHfb8VPBYcQzoS0JUEwDZZPkm8i2aC5Z/q4rgc8cUDevoudgC36w2sj3uhZqcMogvkgzNT
DFbt8rwgcP2hX1ef7yb6E4RCntyMt4evzL50SzPQpBZyaEnjS5YXR8UdQYnKMTEq4O0urHusRyNk
ezPKXQ/gHvoSOPjGvk2qzHtv37X9VdLIEFY/UBLSIrEazn1F+vLFARvMjwguneNXkcCo41L4V2jC
6nhOIvmeApfVPBLLnID7TF+fM2M5MTla15YbXxmJiGz2VR/BBtuHEBwK70CJOzcV/sc4d/2zd9Ut
X1GJliNlS8CDEmo5nh0ME2fj+burnWweLzH5CQZlfQuENWHJWnh8VT+0k4jioO7+Eviw66JBcnNC
BRvdXrnEYg2Oj6Ct31F6PGeZ5dnRba1sN7e1c3XUuIiIO245XMyGkNePocRQ5/P+NEDRj8Ue9p3A
ZZRt5/qOASD23KscQ8Q0utz3uwbGObNsv3MLnztc2BsLqyzynHgpiKjwj/D9w7FpEn/lvSCvfzQf
bmvTQE+GTsAtyWf3C3e3vLSEHOqazqc3F5l3iDB7sGHimcmXMtXOA28qPwHGMZ3YVZGQX6WVxjt4
ldx43cO76/iSeuSuEGfRGNzRAsjajD2gkhCCzN8z/TqWXm3B/4otBGg+1or1xCI8xeuewgCfCR59
5P+pX9FeFYAdMAxr/rv0W9pSDCbboVaNLOAsxX9/LaaBPjL1kkE4E+46ve8EN//czMcheME7JiwT
iBeW0VjnEusXcXCIodzQGS3NA2wf1+IR4nHBoWH7GpocDPZz1uo/5ig5SwqydLUhSUSn8myOVli6
8vwEl9yOkn1ZMoxZ8x/zjaOWrWNuTtq8Ev3yhi6uW9dJjWkNK/p6vGax+KSyNJ+IIWWZ06cCc4iW
JNmIr7TnfiMIWDd7JFr9sXjO8fQy0tB5pEUOexXENkG60gCHKlPMbqXLhp84tPP9OdVVVSqJJidn
b43DJszLITPB3d9/1dqm2ZXyqTNIcQZHjEA9SQ7OSZ8vKkVUdaT1EgZ9dRcJCU6MzJoFpcHG6t+y
EvxmGwBSUEnKT+O7W9u1nFgiUqwfJ4eCUfdLNR2LrOPZtXBvmAH+XuK3qxaN5+w99xucual9gL5F
g1UIZA4rFinsVvfIdzsXYPRiQDkuvIcHDBOwq/HF8aFXLVNaWj/NJ73RkoNSmHTzh5VStqUd6mxR
UG9TRxjjt2zou0NZ2XKE4EenUMJXTMy3XgFBJesBSaQKSo8PWv1DYG73bCyQJ/0QSGYlCKG6rcZP
9/r44XYSBxjGZdn8iCMURxEFG4z60y3aNuVnCS6T3mIFTdeYeUuQqA+u9lWx2dGxClEzGES0hOpz
RLK9O52WwzosFqtruUp64Az+erfk4WlMHP/KMGh/0LpjJCjnE2i/iUDMyJ5pCqe/gblZtSHC/dVM
EaA6OvLIed1QWyQ3RZ0KhimJUBzcjIYsPVRQb+RrAiBEev28l/jd8rCqebrGOhZV0Io0UETJ58K5
xdDnpl/rXTY93MPWp2d7egsAVujfzdjrymBE5TqzVzaGpIt3GX8HhR/nih8hbySFMCXE2Ru0zx3e
BIzK4uGobQfN4FP3x4ZK7/CJ+sSh9ZlpgtCi0edL5Y30eKsXrskUWetFC6asqJYiebnTBLm+kkou
rzgvxFVPneEwC5T/YYYS87hCRlgVy6tsLj7xY81tGk2O0ilm/k4SdrRXP2PQTRpxzAPxWaz5smvr
NR5pcpPxxjqOAkIPNkdevlfMZYk1p3DfgfOVe0XaeCRAKt+QOgykByhTe/475lwepLf9gjG8hanQ
ZkTbu06sQVJWPy7VFC9NsoU5zg6DROL36k5+QCqZ93dz4fplspQG8LVLkuffpUgL2TYrqDYLFLKE
5sqEWbjk/0SuxWH4/1m8pyZIMUUSGHMpcg/D0gofiJEKsov3RNHgiKr+51KiAjCmNg8rIQORecH+
L67uppXbTeQUUGPoYGft+hjTJUUh6IQFlDK27VEF01AQHpx44P+ztnqJvloDHBTl9pVbf/H2p6pg
WPzqs01N3AVVK3L5icj7HiRtN8DNn1bIrWlmE7DY22OvrJ7QtDbMrj2ujJTG26uqMl2TMcAWoKe1
kDIeUhZltnrshhk83r8mT2qvqUclAAkIagYNGD+UzJGxqcjb+eBlC5GpM0D+MUWaWMDGljo5YEw8
vON39XFNciCkJItgQDF6TamOzRvEal3o7GMkexfKLuS44IrHd0SDC6xK5c766L/Mc9wL2UZ4xViA
hSyCrE5574Bgva2ZWMG99fw0w7aQi6ENIEVW9ZEmXym4w6iuXzWynV5qJ1djg3MQiTwtBTtTdMit
NVGLAeGq4tApILuwNgPyWKb70D2Tnq2LXP2RVS9Ozp+/WP9RUpoYLxqxl8vOx4Df9OcHs1hI+NYW
Q2akEMFzSUdGHuvCLXp9hhv6BgtFr7D6KiRehZCB+YfUewokQk9gEULvVZqVajP2uanXdz6QgFje
hpC4+w+Y0OaM/nRjfSYWuna+V67fl3T00zh3C4gDp7cZwNghS4WwI5WrSjxSx3LzGTsIj2eOIAUf
9+VLOaZ04ijxc0+CABwhowi5XbxL/5PxXXEGBZAfrraMPfrtFHIyIw4ZhvbP1eL1SEUNEF67Ff8B
iR+JaXSJ9M2tJ6rfhtxHVoo/a801LQxAYalpWOJYEiIhyg+yjw4raTSpqMbNsrqklLCjciWQPOSv
gN1dFPqryofFFXgh933mXHNgeBSDdK6s4JiC0UdysOnuSDiuPONvh++pozi7KsaWxR5WfBNkHMci
p/276uHxX4lngqYSMhNFU5NZrNZLMjcHc2NYAWNrgu4Ie5JWGe+k0/qMUm2YNgritffYd+9yuDib
iELr+7vVSCxNdhSoWGOsOp4h8JTTaOq02JQrvPe8g7pbN5SpvL95y56p8zDA1RJMcfsnNw3sgHIH
PCCnrqgiCTS8oa2UBqLzs0H0M/F5TqjWbKN9SufFJuzlVzLphefgP7OM1bIg+Gp7x9HZc9kKFmZE
otbOeSijFHW7VKAe+zJ5m8buRSo0USmEoKt3eOXoKX45raOSOqZZyTkDlmsMC3BEKiltuRevtPXL
BVTm4Ao2bOMgUVYpC/oSXq8TVr4BZav/+Cux6fRKRNW6Qn6Bd5icRcNZG9hGL2CeNXI8eHS6kx0F
L6GaeBqZuCl0kNPhiAEB/weh5A+1hUWdsMyllbZwK0kRY2zbq4mRKzjpWRwzAI3hUn8FIiWRQWGy
0oHOGXAYR2Y1OSTP0QtqzK/b08Vjhxlur3DrLdrnmXiTUMiF+4Qt9kK5eGnTaIWjfWLzQ4M7SLlK
zHAj+F1En9bX3WJzeNmsoa8bnmluXrnvNpeoFUE+yXGEqh+TmkMSoa9rLEmjgMJ3l8V1hfwtb8BP
ICyrWRjKG1hzFlONlWQ8RrkZzccS1o5IP36zSXFzHbNfO5OonktTAHFBsEVobtlX4xWtsHCaMrNz
ae79S2gsGPvFmehJXurDz9ok5U/kVKoIdZT15RM+Bni+43QsICEVig9k/kFnxMWwzcDEF93GM4iR
8mR7fLkuYy8aF+JZoT85w77j43yQABR2er02ar/diWO2oL37WstL7mUqxG6bbUQhmaPSaIHOQ59j
Z352Vcysd/ZkeM2W6AaUlAbw82aD4BJZ4LYFiMNknv+KsW1owi0v/vrXXI64rWizWOyOql3eXt8f
3AjAKMhDXxoI/6WL7OgsbGl+bUmELPYahsJVclPGInZqGGU+3c4q/k88of7B+hQUt7VUYY0f0rrT
uAKbqeopyvUolefcbK4S2vQs8y/qXM2I4Zpu4QFsiFUP+I3YVpp7YyL3KSuFdxFTVlBzelLS1wpz
FHchlTEV5XeMUiQw59W+34QY1YJz4wZw2I/Ciil8gRAC/5zAJ+fYsxDLf5H5XvKZP0Uhx8NtjjxG
H2eqyI8cAbZEA3fobEhN70wrCFF790qnvAgDu9ss5+AOCBCSqOG8aHYYsaY9zY4m9vH87R3jM3qR
v+DNa+IAESh1mAChHv/HOWRRzCiiobSlDQu2YtG1BhhvSx3cyo6kNdHS9JwedqK3PUtLXHhta2T1
UXKeFobb5+9NanTzi4d/QqyFs00SsYp5JPlrMB9NkgysKnCTR+teGfx120NHzZv/RSZM5s6VLihv
NaxqjihpO0+AUdyv+ibAW8J8Rw4E0/iQNFd5tGvoC6AMEizgsyLXBkLt5/fL4ipJAYQdBL83/+QX
0+k9zARAoTbyaE/E3bHstBjdAHMtnKYxF8te9gYB2x/7xP+LQtQv24z3kh4cAjv42IR1Ep5Vn4a/
Ox6a1oS0otrB8f1I3lViyWxRlngEINa/iLWkxasdd4l1Rhe/mlnfan0p8SrFyW2HAVzhc4eOVegj
B6/MsuJde7A27gEiVXkeeqlNsJK+ZP0ppZ9KLXU5+H8JIjx6OVUM9NB0LsB2cZaZC0q1eBuYXOZi
bFc1fzS/uBLpH/IBxFojps5ssKJfZGw5DNT5gwyZ9jyjBW8f1JOhmcr4pNE8Xe44QGFsB6olhJhV
rCeM1KqEq9ug1CdaahUrskECrzrBf5jGI8EciEe4ZdnCJwlW02hSyIuusUdopi6nqK6UIZ1bzZCz
+hewq/AvV30NcJSMXVBn+Oc1TCDMv/xerj7/X3cVaTjboREqlOPOqgX05p6pJ00cEvAunt4+N8Oz
QebfFmnSCleTgE937+6E74Ofp0Ji2gdx5WN9lPhCzV4iHwVg85HlcYKFeC37JmQDuRbVDypkPjEc
uG7Za9GaqlKfujCsTepI1iOHLX9+2eukWAmDgR9zk81hVckcy0A4poXqZL3F03EpozIwLFUXDtmA
mE3o0ZtkRbMKWzLWWXhc88fWy5/bIifXY+Im9mPDpR6K7YAUoiIOiqu5hURJ2PXcclj0ixDLoUp2
IfPHv7J6kF/0NfEHOO1AO+R6ZAvshLJNoM1RSVkk9ifdrAOyuRWavdw+BD+BErR2HhyXXLYvLhfc
eD4xPBDNRoJH3QLD7W1wnb97oeuJMYwn3UeOZ78o/KH2ag4uwnGK2xvkWk0AcJNuNUg49oldUxjC
g4/Iyntb5SVYWn+EQ3puwVkADtkzi/1T2HhQeaA1MuGGcIynx3jkxROgBtU8CMq59oBLiMQLBG0O
ec597b31kqRcj6TkusfaudxJB8MPpzGtrd8c7Btzjh8TPtxDVHl0DQlHyHLF/ANHsPig/dGjwzB4
630wJLMcln9oRDtQppgBFa06R0EFXpH81Xc9PqEooqwwjMHH7ui6WcJ8SxbspRJlwn9TUahMk+Ma
zSNF6G8No0yIx5OVKLKEjJ78RqMO0Nc83Pza67vQutPjxT62xyAoTI8Ag3cg9UfTJP5pqet6K7Oc
21IC+b/5b7gOBnIg4gIXQo+krlLXeVbQlp/7x59TkIMcGoLfBwXDknwQrG/MuovspSiHJZA5rHoM
kRS+5m28gwOUosVviNQ+45l7tlZi1kwvhnDt/dpSHe+UgGXJN8mcBA5sOwMQly4t2rkOZnV6cJ9G
GMcCCDkYYZ5qrvAq8ZmEM3PI4+tncXP6sWEWfy4WD9F0HS2AeteK0XZdbqPlAtsd7xHQOtXgBHmS
FDvmzs4LtqAjYio0zysM4djVMHl2wwdnGLUMs2jpjCd/DuWtpPjgXDJoQ/yWIlE+Wj87P/ZjLD6g
M+xVQ/TJAOVHmS9z/O3AvKj9MMfPpRHje4d2CyBOaD1+xXF4Pt50P7UsBu+/BMrpbS5tHvYRV7SY
Auef8z8QgLmTdQlEmzdaFO1ZtFNVbesWFzSEYSYjd0QUDjIKuBqXGA2QO80ktu/TU3zUPCMWPfzV
nE+U4VPfMxXggkqmazknGM3kjwXwjNkhePf5JyTILyP9SIbzjl7YFTwcpR1MNaaRoKfURlpOLEk7
PH5+HxDTMZwR9mmgwZJLiQNeQHnxpAnS0I5Sj92s1XAEH/ETVo356XsMfdgmyKCFOPTW3Qj8qFYL
5Sxl+7QdozceBx/p8Ox/Xl9O9KulJjYr8L1FbKShQGUjKl1sTs5/LGbAVUTSMK5wLu9Op4DofGZx
GWUEsbkWBRQEGHEukItTJnwJgTKSuOY5kuDhahCZs3sYjEFZOHRAp7n9rNk6Q9ZRQ0MEk2/nyNzp
3xgamIJwvymeTX3FJ+TX4c7xWoq0ACQKn1UJt+FDVp4qIkMYj/x2Ht95nDBXSRf/QHR3gHac+YkL
MudKmeyXVslvdN6SYcPvNAulCtcBnk1MbBSdKu8wjiC3Bso7AV3EwMjWoAVQBHbwI7Hu1KTrE/u2
CcaamxqOCjf3xiLN9cmEIlIhxI96OIhEO4HNV5KaDLotwTLth/MFXbWXDH4ejzHhz5gXinOTK+CK
qPf6YD/X9JwMchaiR0jGWrOUv8yD+8Ld1w+7AJ36tEMvdnkOB5IfEzd4GFIgbmzChwp5iuvat/es
qD0RjZt19qLTQ17CkmHYgZfz26yPNV7P2ao8jnW0XqpcEBp45/FK52M638WNxRsqiR1oN1RX9L2m
QnkWhhso3Tj4gy2a8M/YKx0NtCYGVEUDuiQoeUZR71RGUPPgVPj1B+j+pxjA49fYslMIqJPTud2Q
ftEWAfnQjICjeYcRXg6g+udhQ5PzP7C3CUvpczYhGKr7cHF/+2BIzu7ftlftpXktPMDxbu/rhfNc
kiC1w2b8Hg0ii5BdLIEZ/tgyS2Hri/Iw2MqtDv/M/S4PjomEhX8riFIKMco4NqZUPiP837QNwmRI
Lq7d3YK4P9bmrOKAvATXUfFMyFD8WYBjSz2HSEJhi8J6tq5cS7K7h22FKO69O32IhqyWckCki6Z7
Wq2dqVLZ2R6nF62L1A3+OBT/E+OhIdoxjzPOYH/fhJDZvfUXA0dWmk8opmMF1OPqVmgoIuFfiwhn
Or4ILs9l0DthgB7r7WYXssh3ejKTZVlWxT1La/NJcaB4gGtJcBxK998O4Q5dOOuvoHcWSpuBosKJ
+XscYlock5MvOvmys6BTk/bj2Ost0nakUBG7a8/nobrd5njkSb8TtuKF6fgjcwqyuJzSFROoRYb3
3q4qtl+2wMeLzRfVkzvmov38Th/ncmUSUII9kK9tY6B/Fhj0X848BEWVvazjIajFvveq4KDdSHco
CnUxf2G6dUP4JIFvTQqfIip1MgykwKbsCNNATsoLTdONvHxr4CnX4xL/HNgJD3nzpDE+m/Wu9IKc
TdRF/ny9Evjt//CQMNFSyN+XEPlI9OPxLvSRAauNJaAg/c6T3sJEIUFZoWRRgW1E9QmZvBEc7ifH
oiu3qppWBdhQzXCtgN1kY3WMC/Z8ibYmnzsyvC7F3VM+pcIm6+NcjCiv6dEpv8UBoOEaT86NeLmj
VQdp+sOnU4WIqTrH2s0MNY1gG4fYj/kFTUPRp9OvqzcABiPHAD8ZVh3nOFUxxLNFHp8+U3PoVwRw
Qy3FBGDs+jQfFIHPBhNp4WfEq4T/IVGBjuKD1kyG95UGRI+kBEkmttPTevt7WbVDCnSWF7wD5J5W
9Gqc3O+zv/lAmNZpjwHixnC6hI+gwf0k1kvNgnQFfOsLKZQHOxGOhgxJLBQ+qxkLmLuPOUIpR2AV
9VykrSM1SwEkZhd0olxQ7KmtbCyFi3+J/81MzjHeD0++JhD7WSpYxsSPRGZVFhjRpr4pL8C1nv/t
U8vBMca50em0atCMXyr3hHR2boIoM3JK4oTND+NshYREJAnwbsEsS9enMWlxxJZQbO8xmn/Fhwug
15HVlg1s3chrdnqdccGzCbUitY2gUOpnw6nHrllRP0U6yL+UM3py/IrmIie32IsnjDiinbm9gspE
smOXfmio5F1ai331as5nrBG0YPnp8sM2JyyYWLI3bwdNPHoR2dQj+rOGCCk7TBXIC/80LXA/YYO6
X4Wvf1jmVWbn9tWiS2Qe2FOh/vBTHMvDqCkIOwgqSPE2NO4sLV8I9M4ByVO4SHRzhocQ4GxMj2kI
75zwnh2068HvgYWaR4aqPqj6PGHukisRuxEMGxlisqR9R1IBHy2LW+b44IZXOrSh7ujmF8FgFVui
mW88LznzaS0zYQvNpe1ZhUBTotezPzHqUnWkAbmgXN0OBa+bQOR4Z8+AB+rrHnmdcXESg7553ClP
7j79VtIj6zamlnuUCQsH1sOhtH6u9lIsv9jsf8FjIR1nSVTqf2MzciXCuxn9wYFbE2cADB6zLcOF
ekknRqX+ncVKY0gqgn/C2PaymEq6ZsyEBDksHWQ6UZKCF2hvPVPn+SN3IiJ/+h42ZOdF3uXgJv/o
7D0TQb8T4p4j73E/VG9zEy1wx6v5goec3Gqxq55leWD/bOPMZ/6WmcPsPMzlNsyWZIsVebNMKDla
eIZFga8WQ2+xcH+CdG6ah3LLEe/WIMGAh4la/NNOm9SxKLI0aqETSMn9cilxJHm4rVh9AStV/npi
9SR6IpOZZfyIP7R1Uiot82q+1y8xwyZtC13Hwu84SZDX6itj1cWhpmHvKUsvxii4gq8FY5Df6McG
WbZeil/KiFZTxId+LwmDd58+B6yc4jCxGRYhIrc4EUehEf6HegBt7j6Ag2h5R4IiIRkoNvLI40OO
KR/95aBKpnJBVsr/fwSshcK/Qa58TGII45IaJegBukc6OHmBRzrXKMYYeU8mL878Dtx/ID4IR6VA
PmDPxGZpjAvs1tkZGpwLwjz48r04ciyxbVHchdG/5V1Ifbf0ELbqRpODfpw3j3389MdS4EKeNKHb
4LKmLFZ/1+jSIGD24TMMvjZlfUaCNPJO8hKJe5FoWWpfPI5vM7HIiuHy0WXEqNBW9jy9s1UON0Ds
6olNuKbN/uvZAz1X3r/HlU7/XI/b8toHunceTHbWXO3d4dMPdGB88jE9TAsBtGO2C4BTFAdst1p3
VQ2gDcndOe7YaD0YPV5IdjW7ru9yFMU/WUbVA0HxGiRfEcPwJd6E+Y0aHtCW8IaFS59wSKY5ibCg
JrtDDdWvMYsQSmY8smAOstm6oskjH/lMNpfLnccgn3N2NC61GvouKpcO05fTfMtO1FSVIwizUtzL
6nBQOFBOHKgKY+q3cJb4aKnCoS0KxxvQoHdD6cZMFLp5IGLmbHPRbvRiY+GirRkaVa4ydXajLBKQ
bG4ccysqBd8Sd7Uzm5iv4ENABow+VHRx8J2isuVc2lcSxSBfiPDgcWrdqmNHu5uvIvzTfXkuk0ET
2hFRBfA16JhBwZXeW7fI7I7wi9zslwW8hEJ4AtU2iXQ9mqI0+bIO5OAu9JFSEC7os5Y5tiQbvONH
1Qjbvrm7d12WNPSR72UqnXusFAx2Wb4kNZlC6XrOvp+zrWXIKRtKH8nmA1lyaLlLf1249XCGuzg9
qxr2hbiL2weFUqWSvbRJ8NeptzM9TV8xMjH1iG0BwXLlRfynZ2X8bTP+H+ZDm3+XkVmrK4q1XJOs
dP3ajIsCkEJ5Awv5GbP7VMWSJNWzfR0qXm/uCi5peuHDrHS73OQdcnaIYjhndwPvSrBDAzDgyq8J
KvGBOShVeXzAuYOvheK4w/wKtjwEZTpWhIAM+7LxRR3tTqcy7IM/HIq1aWwf3YD8z7PFSXq6CoxW
vvoUUSZnyG3DOVXTPkszYWz0DH2U5G6WnqghEP5u1V4ACqZ0JVu+tLTrfvF8b3Uh98gX5VDU+ja4
AOU1+YU8oktfzN058I5pRA8rTQwxrS7JDtBuAXgTHs5VVKr/XQbgO81YaQ4CJSVxltYw0O+bfrB2
LuRYMX2iSzLAwbAyt9yN1f6Uci9fhumslhyC+figopvByRXAkWl0jc3ktI9QKI5Rfz47CB78tBOW
YHm8l/TaknrMrU4Yqn2MVZvEcERWIXpNyggIHELItj3hzFxdzh9ZHZe+4HgXhaMhNeAxnX702/eM
8ZAZeDU5eBX9u9QLKe4w2/iLIVZ72T7jYsSRFf56ZKTnxl0oXY1NHx8nYKxUV4IEH0lIRKlBJy3U
s2oZ5T+IaisM5+zfmbSZiSrfcySvO2LqS88lSHtIbEnUZ0wkp73b181W4myDtc10JlmGzOJ3mZfQ
JjVZr7pESTErQTYzHcmFTd1B/g7ti4eGLecItS0H6f+D7OtCy+1kpg92LBIpZ6Y0xWAeqgn6PBz/
I153IlaNf6xRCwGaF7DT0UsvyvPjTafIP8tXVjJ8H6eYXVSaVJpkrMYRR0k4/uZXGKZ+bpAPhXoF
1fZaF0eAEHaNEVAgS9uTtuGnbZtF+7sZBFM4ROeT95X4+BjCvicXK9CU/dSQFfNFyWGm8iuBce1T
Su99pNTiaEtsP74/7YIOAElrCXu/nZI3mjRWx8s785acYUjT+dkFuNPaQA+75KaYyffJzW78C82g
1gwqaKr1fogL5twj70ScrXz5JVejQQO9+9LNOjtjvhK4jvtz48TwEtqsBME9JkRLqPCBb8svWUGY
aeZKnpl8pfFFhkzIexKmAqbmBoGhPd8yAoGJcgGVy1wq+i5JVaWz9HeMT7UyO30hH6E+hvErGxmr
dsUGlDyWysDW1u6HcDJew2CllVRfLkrLwk89S9Q4jx9StFplY39cfuceQNaBeGL74MRpnOVmS0i/
BSNOvBNn87rTl9uxchO8kMQh+MW5R1D4RM+dvU9jEjH6RTPGqmh4txJNbgYaM006eWOdYZW9Bb78
yrvSmevIIhjxshZktSkVozwedO/p4esTdIpYUNBtpPugOYtFQi2r9P981sOT8L8WefLweU5La+rn
R5gMZZXCXTlWvjRQdciWLNBi/Wf/lwSW7uHnDjktOOdJEGTLnL4kt1qfKY2Rr2hLM70goBzOp9qz
XgtttxnYXdEPz1lEZD853RQcnWj8kLylPI3ugdeV3HrjoGObqVFZb/ToRS2bnnJ21ycHJCTAPCZb
H3mPqP6S/b0ThxC+Km+UBQGzucUjSw4U/6hSfotU7JyqejxPVFwz2oL7oNnJaWW2wAcELYzW26HJ
vqkTvwbxNscjSdQIVvVQ7K4JugjanFWQxhE6KxF/xLdSQOQEqfKM8tFG+VzGmwnFz7RkgHxy/XVX
HvjG7OqLDycK8qM1c4kyAZbd1OGaI55wIYpcvrlApUitzf48Dsht6IWK7R3Mgp+/ChCWOT6gvWnF
1N+wgVnheaKmp6qUW4SQ9GY891smdPToHllOYA76RCOS3HYEbdtOsWf5FyLxL7NOfOfeHk46HAZI
eUBVIl3vWevq8XMYWq6RKQjL7UXqB3DMJxfM116S78WtMi5DTTGsPy0XgRBR4GP8O5iIZZ80L9BH
ppNsUui/CImU+b5uf+cUXQ4z3jxKLbUaTJb2OU6GPke41vCsxSD/qM99oeWonkYYDmZpPvVmeEvR
qswff5ChgTl4fcFxlTzmUcn5P27QDAx3pTdt/ei9Ei2abjEGuLVZtO5VLvQvNNr2NM7eCzL02QCG
yFDV/QXNT+M1ClRq3meuAC10vEqI6HRRqKZX5IKac+OpRLBdI7WSjlKhHaesx7iRrl+TiBjcPYhw
gaEw9dUtKfFDGqD6NIj28sVDv06ldaVXg7OsLq8p1J/4j8fS+80YjJXlI8iTWXzjMGkZThBtTnvK
z3MO5UooGl8XuDwOmzTUgZLFhU8H/XpG+J4fwxe3UE7CwZiPV7rpHeKNXFR6OL3GsQun1FEehgvE
o3Rl8IMPVwEjKAUwViGFRjkiUv1+b2oTO8ByntvQDrsFyKrEhcmnzzct5H+LmC99hVyYJbTqVlIv
fEkthLGMtVbYFQia2NpkmX5XvgxV9yTobXnrQPpdLQvbsb1MwrdqX6rNiUPuX9oRBMRhOeogYEbE
liVk3I7gPvuTJFn7oTez58WTk5IbJWNZFxwbLF/i0LAZdX5Nsp+IlA19IkO3P8HAdcBTjUtFtfOZ
dveQ5pZ9mcnHZF+VaX6BKQsS6PblqcodMsLCt1vGbtZfWgtgOkXdlYBHkahKfDi7avbTZScM9xB5
6CIUWDdc9eKtddBt1dxEbYLsuR/0ZRN33/hojJYMUnCGvFovXMkbeu1xOtnxp4Qd6VYjvg3Ypfzu
vKifD3/aq+8l6Sdqfd9Yoy2yBSsD1u9lDPmwOmgfzZC3aq3Fo/n/bSiZOIZ2CquJbp59yUh8V38G
0XK1H176/S88AJ4FvfwRIgIxhSAKAPTVIriJMKgNglGOhKYO2Yq8gxQpJaKDQoG21vtqBGRzVjoS
x+vEuctdNdid7vedSuI0knsfS/tO4JfzsblsbG30N5pnOn02RLS7Ak8ElB3Z1Rvh9AURG5XWuC7o
xJqwoPnGoQ7Dd+bgXCwYDZEt2O/2JQmoEY8Rkl/vj64iBkLvwVAQh/ZN3m89Xw275kNREV6KHI3s
p6w8jw3fPkSmqJuVc7uERDrMV6PeCr+wcE4QfyUiqizw6VYKxXHS4HLqii0UFhyML2L1gJSjKKr2
vXI0mC0fTNjCOWcCCX05dIcmwkcafZ6lZcCn6XMVvmxNUKxjSJnCJ0pVAMifkdeVQLbwV6MMckgY
LTqq7qrlFtSrImz3uIYqtebKTKbYGduuMaaaN38RYyGnqtGjQ2Byv/SHgt0xDi5JU3sM6m4l7IKS
gI2XFj4Od9cm+smA4gyOP/1izeJH1o4UD6BSwQkOnoDmBUQYx/km+3L2fI+6zh2m3vYXMmx7SFii
mYASFHa+tBN6aQAO0bwmZ1vavWynFDZHxv5ZHs5pQcs1KVuHXQ6XsvwE1pl3JALvrugSPoyIpoEw
NZfBum6rBN+8f7/Wi2E6CjrRAlUd1dyGe7XqR9xg7mavRs+yk88VTIRewuPVid9MFFTga1ivzJnn
r3doSozcRKuMfLReorhX6QkO5apzf3ucx9U8PSDHpRQx5wmT42GL252ugMY6JOX+AQXN0GcGoqX3
iEeknSCKnnc6FqLYzsQ7jqvsm5hxX0pk4sJNUwTo1/qxkqgqwXJB75Y8ee1iB0jtYp8VV/dNx8sc
Mp9LLHMx1/rWc1opMIfRlhsCryIB5lsr5fKulunTd4AsmXCTzwksBxG/lQrjqB7GEN/L4YXhpC1B
fecXbeYGW+cPGqs+9mjCtdIJG4lxPxT8eGYpfWDv2//twKgMn5/e52qdys2k9TIVX2syojTeoI1J
xnigHiZnI60vj4cWWRrAqJtpOcBXkuWObxaLzUkO85iLRiAJbgHqIs1Fd1quLotI/5XESuY0QvZ5
A7ilqOXlBxpY99JBzs//BzVGd/xc00CD16Tz/AP1VIDBKCNKxZy+mnVGbuSf4NSnk2eAwVsBRv1s
a2N8xk3NY1l7qb4IBCfcKspZhsRJ1U1Sdm1yVoVB39Xdz1Vka7tNJTbbpvX8cnJ6uD5sDIrRR02f
Sxu4JCT78Rzz0Cy83RIEnb0BwTh9JrmL9+tZPqxhsorYsKWXdPZoEypnmEnwsVZKq78nXjJRTHic
OTKWPl2N23rXdlKZu2gP39n0xnhq2dIJkaE49BUkX0BIlYigd1w0fshKx4cNv7+sUIxiuVMIeQZM
AWcAovmyNmI2rPccXacgDVjugXQc+/3ERl4aqeSAgPAFORyqlKIEBat+5jrPRIT6ao1H8W6FNXjL
gz7lkEmJhIzMtZXeLV0/bosP8FOtOdw0m6VHz+NXlWzq4Dy8kBPRuYmzcNmkvrRR7j+GOIi40GWk
/sz+yj4Jcfn8X/UxvkIvk5ZUZdkn15YTSJckViojaL7V4y3+2VoXmM8vkVunxoi+YMbBzRghewqh
HgrgNKSGRLycpFvR3r+feQJ0XwWiUm4TPj+H068m/nmdIHPvJ/EFvYyBDxpBFC6Cl3FG6b8fQK+K
YrIa1fx0nM+x+58OxZI5TBxWBdFE2u677B2neN9KRlRj07b5zhbVLtcW2+aYYQDUkSVV7WaqYc0P
OWuBb64lrQPDtggTGXPQ7cWRxGUNSfN/n2Y9KdkoiuxG6hI3lbRMshXwjGkaUvQ0919AsoJacfQu
GZmXBQ6zli02ilVlj9gwyQd4g8qrH5DBbnqOhBMg0S8w2GpiZOgNfb+oc0JL4wpw4T8y8yjGvCcr
VlH8UC0Kha54RV3IaLMyScr9N6MFT8LxcvjJRCWuoUxHJQ5XzyoaWh/6d1nKllsf7ZCAurc8fKmE
yGNcnJrhf7A/m7rkYqa83lY1jjKsvnfWvV2L8pOx2MigKG9g153/nMgBhwZUM/V2BJPpzZ6fR7wi
Bt/OKCaydsid2iAldL4g4/MKR9zRpFqvKkhTSvuxhMzLCdZekLENCcN3x2pMUpyBZBK+14ur/F6e
xfC8KKDvYdfBtW10fH/7dX3jefI4PfdMc3EKuziKbFKHn0cOOzOLCADBjwCrA6gppar9qhQNzgvg
FJd0V9WjrtHNuyxX4xEOL8BJSIGkyf8ckbNXL7ufjqfZbS/H/AqogLxkwqGSqh0Wc4M/c7G8WOZ7
pzWBjnwQkoB0fBDavlJcV1p7uGMfqR2OozyHwR4KUu4oqfQ58sF05Ug+OSZmjFpz+TGQ+cTzNarC
B1Tol3MnZBpd5cQx6kvta24n+smrANNeTknsZN8VmGBKOLGvQDvFpAOCGP+D7unRy42/GHy3tFZ6
OztQBi8ENZ7ZAYXFscONu085gTyO2yN2vqD9Zwj18O9lTg60a+RfIghgWlqzYrFNM64rrrk7EUKa
9LakZMaoF0jrrwsLhy8HiInZSpbbrXT5GGSa7qCM0tbugi1zd87lz0UY8DB7vdf94WdDCUYJAGMs
R/rDkNO3/BIfKDmiMI9zTyh7kGnruNcYOZ1U0kRqamYT4w0/hhmj52b8rt7Hs5avoBrcq0Vtcbup
YdiQ1faGdDn6xIggS9bjmrKj1t7mIkRa6UZAIyaVI7xmOm/3AZ2XYZjL5uF1VoG9fyXRotAJY3OJ
yoWFhka78W4ybT5c15q0HpVt4SlxsYQuNCKnKIVNKfcLfFpR+XIfXflahr3JgVv6JfMoDfUqdZgT
l11nlB+xGGFszYJMW9geJDgnXku3DtHFc6EThvfX5jUN4Pgzk4lTbM1+EXS1GFhsBY5oa+mQrJQw
ASGvNO4pwlxv5fX0sjxu9Fa/hzzEhIOvhaeD26aCz25r5RabmqAvo33lyn9R62yX9QslAMhjDxtE
EE7yUkSMeGfln+lUjhAhT7zfFlr+u3S46Cn13uEi8tGG7bTPpGn8hN2G3oAGpCWToEGYSeyJBj5n
8bWwTIoefTA1pQVLC2Ke3fa2JUi0ye6DqcKRvzssOUCRHloEpw5u1uj1xjVkYce57UFXgMkW+9z3
rGEBCgFCPPqTSsqPhbxjCAXyISaGHWviDLMTDBshDQ40ZXuFuzUVJXrksxq5hS/6xbi5mNS41xkh
HPDCTevcldv78A3RWyf+OXfrjQim9sbZ+LWUdRqa6cfXXh2Ih5XFJmMwnQnNxlNfqrsTZzFSJ4KO
WEsE+Mn+t0cULP9geix4k7MfF3QRA+8IFXbNlpixJ+N5o+g9/RVX0IqvvLy6h5sVYvxtUIwxaZYp
NS3I0aH3b9r7SIwTk3RQRCGRL3+whyv1C3PlKNh/sXzOHr7osStk20RIrP3peU3LKVRGh+HCt4XZ
3Y546IMe8xkk2qsuqe6arenJIfL85dTZik/V/NCOL38UQT8XDkIbG83ix/1mlLKPeA2GD3srH4rL
jCzBNnEoSYOvwGr5OEtNt9PT5gqvWPh3YrKklPt0pxpMrQ7Pj14KVajOxm86/zFBty2/hHe5fA7p
XVBBEm0RJ1sIf1l4fbD6glY5njwBfCgn8FObxHKtSNUDKHow6nIPMPn3IV0ZENad1x7guOYFu/uQ
SlRU5kESShvbybuhWe+AN0x1maIHN0pagufA/W2iLb0ay2zz79Xclu6F2GtDLKN6NkFt97HZGSao
vHdsE7Mr33bXEqiE6qJz+kyhWL004EwYMPfQ/9MGxz66KrcuWFCvn/WzfE/HpfPXtVMZoGssUyXu
0kWdOuGLLmV8jr2QK8gGPOggSYWWJLOWQ8+eLLW4ile8UeC2TsAvEIVgPiRunsJCtkj8vSZcWe2A
/7I+qiAU5g72fxEpa875/1BGOKxi9Q2yqA62BP7WsVa9+CwJYK7xNmQ9SqKgMoSoHCt2B2bgBF0x
NvxH8yPxGq47WY+GM4EG3Q3rPGUSHCp8RfEjuHefdV/gxweBp+4aTFckehH9fHkcF8w2eH12e5hr
cgVAN7hQ2Ccoz5xVLqRvRZwJts/N9r+z+ukdq8WJP9ajjYmCQQlviPq/J2Nq4jJho7gWs5KVMJ5U
bNUA58z9v3e60hhvyFmamm+eAA/d3G5urWzNakgaTAbWBCEQE1F1XeZfg92d+cLzkS4z4ryf4sPd
YrShJ91NOAp0s8wSpFeRZSfhPIoVsobnZ2PpaYGmxMZ9A4jnlJR7/X4HlRWu5HHkzTxX04VpLc1h
Bplmn1Vxic+d2iiGRj5xp9l+HX/JKPjoCDE/ANLDqwPsHYp7IYKXv9317ce1b2CF0aJvhf0/NTp/
hjgbkG4wzC3+wa8xFDVFD82nRw8pEskn7cs8e/0FRh3aaodh/uJrw8CA5JnrN5c86cn3pNq+7O7m
RhKlQvyN+DXh/OROdS7eZlr9/rfFRVA80XxqdpbtB0qGerCcEKp/AY/6YudYk4dnujgq1zofF7p8
R8VxlG0F5/VNE0XNNjE/tuh5duylAY1/uqdXF/fGInxCbmg+cpA1M6O8HeoyEsqDSIatmct86Z3y
ADtF8CxWfuSgTgn/QHnEurbndzh45nDzE6UmWCshnw+uwUFH5K9KzbfWHzgUTy3Zk7AdZlWaikvB
1ENr4jdps12WQeKnAbKEq9LLqSREYqtCi4BpYntrseq9FhnyhXj56r8066H4L2NNhW/eFMzC9soZ
Mpy1S5pXxLj0MOQe/3YFzCJpq0vSkRo+uN15bye1YOAHh+VwsPAE14y4QbLzYHM2IgQfppYbc8Rm
eMNUlCW1TgJM4m6VqFVtbujOjXHDpf3r7hMgoghPIE90N5L0mWrQNX9TT0aBEalT6RsMz+DO01dq
bIY+p5Zae7tUszCthyAVPbXikg9ZZlZunEmOkcOWoi+0hx8/uvcgtXdabMXYppEAq1Yn++PvIZu4
RX/CqqUscYjJvkG4Yz9Jq/GLFn+uxSgGqJl7ITIBMxnocmgJgyGSjwA+F3koTKMUlovLjcA7NPO9
1xNTAKR0rqbkv1nfeAZIvEiehh9IASPt6ninsqviSUpW6kcNR8CZ0/DboT0ef94skHzNRPAQxvYe
8eRDivpwW+3ny0w7q/Jy1yfDv3J42dL6yDxGarY+Y1RGjQn0HrEXlQPsvaiMra7x094WKGa72Fr6
OXgs4c9fN3eUaCRUkkswGVsUzl3CMtcY8cNKvmbG9eohRB4n6T+LZYKSGrLWYr7al88uztnCRdDc
4RfQMODBiMr4Y/Ce4j0whqoQfwtLeuRUIGe1j4+Dz9QU49Lkn2AUplh3wtQ7s1QSHHs+OCTEc0lv
n8aXVfelOrCnHS/neYKdvMSUimVhdjqfDoG6FV/yFFo9SKWmNAVTaI8h41C7uHC1Ou+yVit/hnkM
Qqj3iJ7bN7I3ZhuTbeT4httwpOrDl5I/aD7VZzrtmAxVIdF1y5Poj+1VGh2gCs8JgafFO82wfaj9
sMMOTpcMUW5smtxtwZVDHDEi70feoMH8/RQOejNGbiXBXkpmrHhiEFrx51orh3wQz90+qAnZNhnO
dxdkfycncb86uAqkWoxjPod0L73PFlaDhMrzBwbPBgTdEABF0C1eusaTPo1mE1CORSlM8i0mlq2x
yqw/9piPl+jH3WeTilB0tnldTBoloUnmLihVaAMYG7u96WrW5ExxBWM2b6/RYKd7Taihd++4Dxvh
IbAn5dP4ppq+pqDMVACBPEwZ6/I9RuAJ03emqGY++Au/4m0Hh+qHvsfbYvtAI+HGCQmk6zrPGPw0
RzFQYXe8+DQ64HeOkgNRjQFGvisNM5IVM8+Am51YAQC4iUpb0SM5jQbzZ2kMwmM0aKmZDGB9dQv/
Uz8Cyp7msMmw19Pk/b1AI43RjsZgG7ZU6eI2dz5XNrfUV1wyMZeW6sqICScQePJ0VZdqlkYPUffy
55RbyQtP6o238gR6N1IcBFG8TcKoUf/PNtTZkjL4r9tbXWsQZoeVUHHCwek1+S9wpSsZzYcobGTb
N6IodTV9NyZ1DsASq06JVCvWf8sWPeZz+caaXQHathbpmfkS3k+4NefqHH8M1zCsMD+EB19wBoJ8
e++JuN94ifFePV75kSchJAyHF9U/T6jFuVCgsFkTyNtLwJC8ksoNToALRYz75q/eqU0FbbWQ8y5t
rrHYjAOs3eymu4r91eFi4krev3tuP0l1Du8cQmMtEAmBjgwrdopWt3CPasEIy3u5gTi7DTr7Bpi+
eCUpTxPFB9YorNXJvtQ5ha/IC/gJrjSVAPaiNj4YtLXGLDwQto7Uaqh+BGZmnVmY5Pv6mIn754s8
Cm1gmtz0Sdjkz1Mpe2cBrtqidTi14uZgJwovEEjyc5qGF+2QCPidilk+0UrRlbCALuEVCcvC2dgA
1pEZs5QC59r2KdLA0sTyPrBrsVQonKNIH+WmOknFUAnmk1fDnxZOOWNLLL17bEenM2Zkpk0+1wsz
PGEw5n431mG3KjERojip+JvXVWpfpBFF3U71YxNvYX2Z9CVB3NFNvC/QCzheZ8B905Vio+v+dmP0
HuRVefOE7N6ORkaC7mNL7xqXAoFA8eOUBGYrR7K1DEKnLdXzlmei2uCAYjNPYt9zmddTxqAm/gDX
RtSFXqZMeozGurB7PsyhQeMtAuopRcEr02/0QlxRIAfh9n0WEXwsuNIljPkLVufbqF7EXy/Wqfw3
70PnYLUpmMbmoDEMdjHKDsqbDFtdTHx0HfrLiofpMmyIw4zsNSQz/ENPIKOFgFeDk9wXJUPfVycr
+6vVgARrx/VGZqENiWB2bEcyi7G9luHVl055/aW71qUoz4SGn1JvR7JmELGt9+fOM/qfbfwMZ+o9
hlQCZYoY0FRC1WsmpM8tpz3cWk8HjNqB1qipWBxR7RA9OtGhJ/0+bkpHEfk2tPCBwlIWKwl+ae9e
It2b4YQXWJiu1Kd6WoVfilRZnrenX54lxuHrfYX87uFoY7EssEhYNm/Nn6vx10xCGT51jiI48prw
7IUHP4R2jVIiKhE0zjQ8GYcXTLmgm6ul0Vq+CFrVXXMRUrz+kT736IHMyYg27FoBjEA+uVc3qGOH
zNPagkRos4JCukCVRDqcmCbD43NuA2lsx1dww+CnkzdwJmvU/wIm5iIxXIFoQ0KoRAt9+f0aef+N
sRBd+Ijy7XPRFPbfmL/wAGqmUW1o1rVi+U6P9nDboUGJuROKbRYynFZ1DGeCmO6sQT39ULlQ9fSw
9YzeUr1RC5/+uFV63CJ0nS4jkT2dyeNJ9hgvP9Vrtg7jwXLY7oiz8O9Kv4d7esfI7JEOqCQoF82U
3eYDAa8rd3gSW+Zt7TPGA8urFgzqiQRv2PSPQ/mjs4LpSsCjuxv8nfqn7vl++GWWbnhkuxhVlyiS
5RsGwNLO4FmLBCs+m84O2ussbK9dBXpNWwk1qpAhE6Qp6ETuhw0IKzuytxjisPo0jxBmNGD+PwE3
gyTD6KMMZiJZ2NLgsB9hvBuUPBvFMARTg9/b11WZdUAdWhWryRxP4r1EWUcnyCwPAlQdehiz9odF
7V1rqBIUoYGCk3u5VnirVixkNAT+Dho76PDlis0xqTqD8jVemaLVl2bi4mBbNex18sQhLQ3YXOT4
PStrqM9KjySlfxaDOd7qlZR7zZ2VjY3QA/s8fkSQvBRQZVDtELUetzkFSRA2npfKW9LarsbN0Vd1
gt+FFmKoKrwu6xlvpLC/sbd+Sg4mfliK94ByjGg+isiHPF7dz1+ikd2Xg70QCibsUm+z6HbYzOA+
rM0k6dnd+cpVIN3umXe1fce15r4GW+nL387VyNsk7C2SQ79HApgGIf1gQyrccZ18yIMcpYzmMidi
lgKmrciwoIkElwDrRr18aNz+gPxbAOZLeXnv+g5yK8NRA142q3DiuVHQFSycmvMTTRYhk8gKe7mq
fIzY87AyajpHSifjR6Boog4iebgKZf+DqLupXNM8OMqdpTesQkAhqau7lymKTT53rX7MVC2eAwfD
7xd86fJqNU3qv/dOg+osu8TX2Bbalepp4Rhz3rsNLQ7zT9PN8PVieclneA91Jiw1B9Ejt1KOc1Am
IrT1/MemxNjnt63aK2tgFZNW/0MOPWg7Wo+aktD+6jtht8zi1Y7QceqGebNzUbDHWND+4EHd7lK1
uWsDj/QpxYUiqXEJSi3XA8TsaWGrmrG5CBs8TIsN9BmlReJcvRPWURrqiVnGuf7AO7K2leSNVVN/
Hf8t0174qucKg3V49f+SM4aqSgTPBKF2iMT2n5RjoZMIfnTWMZx3cJ94PMIYL7W8YcUKeVciwbtx
WUFjUj8a5FXqx0AOyQYyTx9dvga0LKnNx84VohTUHqjuFsQDDbealGxO+MXDBZF/twq8P3ukBPht
6oI7dWFeDa9G7ZFJ215nLiwAa7F3I5dbCEJeDUell6d+iQDYLX70NCm4GJnBSVsS9Li0VkR8637O
22xCV1YZ3dK/hDXuL73yFRsF4WFfYU2PUVJj4kzaDdeg+s7L+rqCHvSWcEvVTMyX/uZiUGonB0E+
cgouDW6468GKRhrs6VD+aaAKDZQgzcUDGpX5oT2a6H2yWbaSKm8myi49fBq4u4UVXoR4njRzL4Fv
hWbyyoF9kcI3a3FQ3Jtaj0kUgvBbTCPAZhgkpdCVqnZq4UPyz0XGc7cUf2eQv9PGaZFBZgELYsRr
/mMGutREE6Yx2oWCAdrm4zu096GQgbWS78CcTWwzaw1rNX9LAJcCXh5/0pbTR1KxWDioGlnuzyIP
M/gzMQf8sr2rTv39RaejX+8RrQkwp88tjK9i3i9VHtV6zngFM0SuVjPyL1UFHFT34hAXQQGGDSmb
ixMjHppkKfDuBzlkGFCwqXvzf3sBtzyciOrIs4ERvuFZfEUpbFjEnqLEQBHBU6u++RlJrEMbRaXD
mBf6zXcF+42hJ8D8p059ltvzlVuwuLjZkMIGZ6bQdZrtxw5IN1V6RqJCCILN8EehqTgaA79M1qep
0yhgNuL3EqdrIWXI2rvOlMHdoPhbfVKrF/l92lc31LWZLERLCZfrm4JqM9TrJ8+UWpR8jJXCDEkF
FSo4xErKFP0YGN7z3ixCnbmEnzlfzl3bEEob8SaSgwSf+VjSjpRy1tQ9bnV2e1dVs3RfRhmW60b7
vGA9JXFC97BHYH0Vz2G5HbaQpuk0WRVgdLC0lyVftopg0ussxJbQLax4E8BpuLEJ3tBLj+4OnuM7
9KqQpDrxYnxSgaRu/mALZ02KudV+0aYcVMj9AUS6/NYq5+71si1Y38GRymOkFCKEF/fXUTkwO2+e
cGV9VGZnfXwE/34gThRH2GtUerIW2Cx16StGxZeqiSHmlIZIaXJ6xAQU1SEwBQ7ugW7XwWPltONr
wbzKn94fTUZFQ7Bho6eM7s1uapt+Owywu+faExVphPyiNJ1I7KdMuctm75Do6vECQXosZN7DqPL9
Bt18kda+rT4iqgy9UXQdjgE08QAWPzavYAT9aS+4RzqiuKR2AUqIEFEUH6GkJiYKRwAYIPEiXMLz
1ub5IhYb41CbfNoym1ezoZBHcMruFbFozaSROVJVTS4WpjBIuwfGD4yTWw7gDDNsExe8C6LWgxU7
ZvNNtVaaBsD2eL/MoavDEYlHZkYC0EJkV8CtLDgp3baaq98amqoVu1JbGl/5F/GwHuU3xX+tvcZr
ACmmvZltkJTjTVE0lopBlWz17cND2hL9JQDX0HPCp8Ena6NQwyFmbXHCiFkYEy0z5Y1fnqASjauq
nFVBYTUJxN/W2o8QMa20cmCPGH8lQd1RDhFY8BGQE2AnmHDzIGI/AVyKCLPAGf+wJCO52B639BSZ
bH+ekPrUb+jgRbeDQEQU4d/cvUBcViOhR7k2k0LUulqFQlUgUDOZUE/jlgxlbf7xKW1bPeXT/f4O
kKanP95Sn0+vvgpcuAiIjh8E4aCtPPo9wXvZFhC5fqYn8hyXTntjBAgIt5tnRhNBYNsdNBqEsrEa
f9GeqaG28VvLX6Sra28JuYpKGP/4NrpWI9YFNS28QrixrBGih+JuVdnyqP4Flo0YsDEFSaObcSnh
ap/G/uY+OtITHu3FyHpiJiS8Xz0MNxq9Jzd4+c3ntOppwOOylAEcgzyVeTKwuuUGyV/p1mXJWPmZ
Xl+4E4lwfTPN5SuK1Irw9YWYxVPzMSKniZwkvEo0LMtwI00526wyljoBP1ctmlbUspcnyeAbLv3c
nUpmq7F90GmyF8yYaS+qbJ9DlsYKFgae6C4intqefEaE9N3Igliba5Qma+Qi3rYBvh1SLIa85mct
1EOBxxGrGjUThnoBbXOtpbCSh8/67SEBN9gsByimRTBlxfZ97ILETlN55NwuRVBFuwYeSYkmb93t
rNNUWzwyWJs179o8uClgHgSGv83RKjeXsCn+9ee/rfwyDWxQu4nqo20z7CTgLoGq8vGmBzXO9ro9
ZD25l5VNT+YYMGqK3EiWJ/Um616QyQrmx8lNnjYXbO50KoooeCQwVmDe2jarhdVE3oj+bkQb+ORf
6rFuoVwTedeK+4O4w6Fuv1alXIT8k9t70bk+60tE3DUB/LscJJhszXz8Nj7ruYqX0j24iIdGN154
vhKTjFFolLXPc37DWnNAjfVrDT+/TgUqq6LHeEBA4K7v/dDgD/5gsec27u0tvmzK6kkffwa7O1m8
X8YSmq9a+0ElzRQ3Oblp6Q40DIiiOOMjmcVz9riTdnAaBeffTrq9sZJwzdIktapsSMvb9wS4NHK9
aNgqq9e0wrGlca1TVAlTj+EPBmW+OItgzWfB8bFkd5WrJ+G5YQNQG8Zna6TaPWN9CWsIp+6apFLJ
lH7pH/GDjUxiDhd525ZJ6t8OC/JvPzFgCbJsqJy/0+N5t/gszWDHKvumIiQLgXZxlm1Hu4k7d7KW
l95B86/giEPe4icAYtQW0lYOBU8U/1EVrdh8LiMepi2kCDSpkJvubGMjzrDz2cOtoKcetd9fE/sJ
jVB2kgMyrvXn2me6CW77stpu1T+hUpkyJBmYSZhCBf6Xgo3wo+YKymJ8A+MUHeV172aFLLC8TbLQ
mJGX05hPe71bV8po5HXtDZK6L9+r2j+ZafuyBBLh3BRHLuCHJVM86PxvcTt1zN+TNQIzhZzizgJy
9z2tUS4kRIajCN6LxLzO2YKUku2phaBztoWb3+E9YyQr9SaIQad2Q0dwZqc+0IM6shDEhSD8er5V
yfoJuVpSvMq6rqoHkFi4Fh1rr3cYiPSg/68bA5x1jaQuAbigXCJIOvRQJ43VqpDuDqtkyY5hF0Ig
u/rRhEq6ZlSrVzSuxUyVE2HyVjPJsZASlSP2t2SINo9FcMxI3RYE7x+QVo0Dbmcd4CRIG9bxo62d
XRhKeiG5L0KxZG9R392xIslhMuK4xvyTCA0ZOwlA3BQOAuDeSgYyE4Cal+PX9Belu1HCMUWoXnpa
kiIMhKNbbruAVMIGoUZEsE0qROhlhnUGRy+2s857E1pM/QGdu1Yh3jU0dhveFjYeiX1Pey2SSCju
eeZ7hoVS4mibTyTZotNfwfbDj6Vhq8a5vtn+83NER7UsQYX9oRmS8ptoB7IoIyL35PZLeWghjKTE
4Oo+PpZ58h5jbSgqErplJsYLiN8Zvy02RbKyudczKzFttRipzDQ09A9/3HFueforO3zIQKLZlbJp
fraFkPjAvsWqqolyF6u7Gq4gGzMgriF+pUcD6u16lSPBzaed4POaBEmWYPQ/A3LZSpkCguKv+hs0
1tx/froDoTWGQWCn/RQfCYT3uSr7DFmzb8z2oQtSpyvzWZbUX71/ibU3/AQJx4MYbiUyFcet8ZMH
mlzRrdOQ5AecdUpstGQOJybZa4g0GxVRzpS8kjHiTSTf6MR1igu+5EuvgMbttFBvWdXgCvF8b9DX
cJZMR4+MsYn6v0OUIJUP7B7Vap6M3OLj/vSL1lF9vP+DDMNsLviNurj2NhVbdxL9H6Waxef3SaJC
AXL3A3Qs1UvuQyn8Lvnqxj8edLKFkKWtiOLty2FOSBWRTEBOGxGcvZQbLDMaHBuK4P42d7/uDs7q
GKLAWKjaDqAk9i+LrOHFdpiGC4HxYedA5anPygOEwuXdT6WT3NukSJKDOwrpxhsaXcUmX5fc4g2T
VoFrT/w0EQVuWGhgv6kbThzGZTKc8afpDxoaR3ivUkwAPQwFB1ZjZ4qZDoFgRMlQ8f1l9OeK8X0e
9wj7gPvX4pZ8R3XNSVGKtxMvQUC/53svtkbXDX9CEV94da0mHTbhlUDWqg/2+sVvTm9Yl5BkFPyk
EVm6rOUNpLg8X4o+RsrH4pWLCwulD7YxCPRQWpMG+stPK/evlxwEsTYpy0dT+qTtlATM6aXb/OXJ
J6xS98hyIHaIdf2rPj0eLzGE5edqNjJHCqbx+ukRZcxDy6s9LMkGLW+OcY3vzNtAQQe4uX3Kx3vD
R5IyespjrTl2+XTpnVXZ8H9vxSrZpYC6cfTlVubSb5MtTLvJNW6oOE2E8EaBIPWc5l1F0QZKXxmd
EESIab/CF28yMmGDQY9bn2ftt7h2UdBB5eKA/KKZuFB2W8hK4x5eX4wbV6JvrC07c/qaa6v1j69C
wHtN/ft9NHnrOOuAafcXgD0Zb2fRhYtfM7T7XES+bGMj7JEYiAD9kaAsIdRapWTsuonLI8KSQoXV
F9pOwZWVRE6IKPjXOQkn0o72vEgHsYOTI5ethz7GJ5RW8yhUhfO1ZT0ObxLJBvVzuw+Z+Ud92Fwe
RBV/JSZVzV78ifl4BpsBHt79tysaNHfDDFdaL9slA6o92RqU1lXO55CtizwySzeE7RLASvuf8tTv
Vbv6TELWctppHsHUpC9fuT+66LVG/xwvhdPeghuGVlCc3JektYH95/BQQCXexTmIE92L6lgUBbFw
+2of17lX9wpfJF6qxR3YXAShf0IvAdgVb7EFfWSzAD1bTkcAkESVIcfBMo9/6+8K1LWaLPe132RA
Ots3sTfEaUIbokkJpEDTsW1oao7EmWrat6fQ46M285BTxJBXYB8vVP8B/sFKk8ByBsCSatY5Wdw+
bTvO7WRnkZxf/6+rN8xYOlGynbaOA5bmqcXczObvRpEZ0hyDN0Otr2Bt44jBHh5iafi8z06El6fG
SNwwmrfTNERuW3rlv4tb2EWX/48wSvBRhQyIWQ8ufW9E9xfynsgoAkyYOVrzdS7QGZa/MN3kC6In
2yS2GVcEmW9n9S+2ZH29N2mr6X9TLjDDAQJSjkLR8t+9u6uFtHLjZQwcORgrt0VCnks2Pn2uUMwy
vLGC6YabbFmvfM34nF3ZD7y6W7Jl7XjyYGm7DNYExYlIzQvNFYnZ387RSxxQGJblNJ55ru97woK3
fM7t17XWrs+7hgh9TM608dGQzJqdmotw//l6Q14jC8y6od9T4V4+wAI5WJOBqARKkGkcy/k2MJdR
YunjuPPK/auayKKez7WcR70/0llJolSlx4WztukB62DUhPX9niwaFwdhkNUZNVUn4oF7ojCGIZys
fAZ9QCW6OB6x7pYofMwy7njNtdD0pRgu8Vf4poOhE2OoqqgtZv6Brc8L7VL1v0E46VhgZoO3T7K9
vsrtciA2hN+2sN4hNT8CSrz68/IJW/VzVC1G1O202dOTtrr4McCZZzGzG+6DdqLYrgX8nuDj1uGp
U9hC1XB/wH5CSPLDfcBaNnRZfYYbptQ14psGdP/wm3igNRkcgzNnsjcQ5iEKWAKqDcaMEU7MlScK
PhntpnfIbbQsnDchyriJAGs8wNv0sh2AzEwsFXVS76euRErqc3gMIU8/mA3WOtJJcYYn0KhEFiv5
0EAac3Sf4ghn4zZjo3QKDGJM1OFYpo2n6bJxr63uZP2gq0hMdEUOMTKN3Sq7ERQq5vKyE2ic9VXD
wffCC9hCvZRfCO5lsxwpduBLBUoeV1KvctuQZh6D6uSpjBaL7e+98UIK2gDbZkmnYOGe3CPnPr2B
CCSJruSTFwRdofaqo9UvDU+TyUaQmsmHPjI9AqSaxO8mLL/moFor5g/eN4g9yZMYS3svHNdqnaf8
NXVSb0Ukryr3TL0xp4pNrknevoVO95Rmjd5HgonKP1yGxceJup/w+J92802mxxbFUSUpmoK/q61X
fMEtOWTZgwv4XngqomqDLVpVAXOqXrFRIfXIOo0yJx7Vg5IRn+3JLX+kgmtndntFO+7whmTpjYIH
JIY791GhxPX8KW0+T+Mu0pLsRDbNHHnztQCZMrdeEy5Piu7q5svtVh5QUqsBdwb+jac20gx6IjT6
8jkO5MNNKViJasGUtWsmFB6LPMLJeejOgf6Sk5myLsVq8tQTQVZroVpp8NIfT7c2jBlykGjEAqqa
jwqIlJpbAiYP0Z+eCCJv0l8E3gS6eLnnRl/o5UZ4AFKh23OqUbD4pQVFvrZDNvVv/G0Kp1k0XcVk
skQ7Ho57ZY97GyPiNFPjmeUHXP8WddviUbC7tZo8dQJLi5nliwqD5vuw3ZmmiGJywMUrtOKOHToK
4JPMlld6xzrhMhIzLHsPHYUmuF9ZXjho1XwiHGDVbHxud8kapa8oz61cpvAGChcFOrkABx8DUDdR
LKSX1HqbGdSHK1G57FnkEwDElvU0hTEycrywifxezM48sE5iLnO+pg3eQsaKi4wYojlhOQr6OcVD
iLFyz4JSqojqM0iyZrC4xTMtyFSDy8qWE2IyM2ydoV/gc58piIEKhMjpH3/6KjUWOLhti4EMeKkz
/mpViZiZu15USlbFNalnojPmRDqW7B7IG7UxKGxDptMS1GNsJdFZA7J9iN5GOJFyzkDMdi4QKltw
HvFELAs6Ro3NdXoOsL81FE6RCJVC7D6IFcNA3fjUxy/fjhFuVeKcbY49bTb7ca2q+/Rv4Nh30z17
AkNQ5f5PYJbIVLtSnftChRw8qSY9IWxWa1MeV6mROrq+C5mtmQbhT9iNXhRQNHDihgJYvy8V11OW
o1Fa3lkm8zGxNQSLiKfETC+bYFlmzbdwokC3SBSdTzrCEp0NwqsFQQyu5EEMAD+M7Z8agmVgKuyo
zy6C3ybPcI6Ne3E/YLT5eQaiuDzf2DLeo91du+MxMA9fsl5yR5VVhS+DnEQjHlxB9XVsQKAZRQtE
UmWfvc8FiasT4Ks3iTAOIu9tX3wkftWeFZYOIfhv2eIqAT0sJvBzfMsaFogkns+/x7UM22/130L3
KoCuU5adV69mvOVWHlTuNgPJUexO3Wh7nzFL1c7DnKd+FwM3TeX6k72P4hGRxXU4o1bmAco2MH16
J7km2I5qEhhMr52WAGPVuRzvpCfHhLzxQawCVluH4N89LbMCWRiTqaLiguqwZbH9ge9Ia8XBIcEy
aAD2v2BjNZW8NPgLrqjMfGp+ygmRWXe6vdQ7XGXatWhBdbDLZN1fgHmwUSJfIPGtc9l9zoz3x8EX
0Jt9xDNf5LmZUSljOiln5LxGkcffen24ulKUzSrskBuK6GMPICMpQqYHHzYTwFYqX9LaWvUef/bX
+yl7GRYelI1FdUKSGZ8O79WDZufYLTP27ji1odeq1up4TANbDC1KLVYbkE95UQrCOiv2UZ+r/vZ1
P+UFIAybLT0GiPc2tiKi3XzB2BWdVhbhFL23vZGAax0woOVh45K9Yqu9dY8TKoiXvkUt3zkZpBB/
GnCfAI+Vys8QO4/pCgBZ5nLZitoCQSVBXRvBc5mK3nDQS1aSygLfMVQCPlyULn+SBOalvLHCsxPK
gmo64MxVJwODqukIabtQ0+U4smlPyyy19/nQ9RAZCTbqDv6TmYsJ2AWBch30Fd1jo24mrVbGQPqh
VomHSBbk49ACLIRan6dcHm5xsSQG56mQ8rM4QbSrU9RzWWG4TBbJm6gTo0DFA7b5t7dhekqSWSn3
7EIaXIChqEuoOv7yqbtSaM9ZomJUmG8lM6q3WefE/+sxuWrXL1vWFlo+h2VbGJUHaK7Iy+A/bTtM
WGnotTdku7jaqER1iCwiUwuz9WpPpjKUKLqscxD/bJB3PMR72UAug5gWJgXOhQnDnAMA8KRDGGkw
i7AmmGJxlO85MJ9DCifYv5yuuQKfML3th24eNjREaXZlOCmah1CWIvakqNpSun/IOmcX2mF+eKfr
8Q8VgJI1MG6uE7b+zZ7a/TsMo7/60q/OeHqAQ/ux9QlE8eoUxKrn+R3p0Vs0MdXxJ/rp1PmQ3mtx
22ExZVRMTB2fJum/rVJ65KvklTSTP4grgVYTVAHM1rvE4pBN2kfC7EfO5LmgovTLzYnnVcuDtK8P
sDQGfAIqO4ksa+ePQ4z1mBIqmtUY9lR3RjbpsUkq30sdrRNuKJF6APtmcfx7WQYL3PMbj2kNpmrj
gBBVh/w1E2gNmZICkd6Gex03ztIHunXNewhnwCRlwU17OaBsQH/FmmL6K+EG56Q3XXn5ClTl7EwJ
nPy0u7x8dZ8K5RBOhFqYf6tfP1TEDK+rB79lg4SLoVH3Erhrz18JQgWGdX1sLHpY/xSP9g9kRnGa
q7zn05SQm7gBlGZPz5rhZEcwc6XakqxLcWf2tDHSw//U06wOIKfHcSPkkObhu4O6fMD9ZoDNf9vW
DlVbs8UbVYe5OAOvZLOBJxPqCEeXEQY9SFgc6eme6yR6hylBoDPlx66Hn1Kw5MjHj/Tn4uwJ0/IV
i0r8ZPwtNqpi/DvmSPKeVrV3qzLZHNYYttpCqHYylkUxLzG2IFRsKKdGej7D13KtrneHTjQ1lgp2
WFxU0ixm2ZTZxnkaCjV3jZAm2vO7/UwwqIPyRPok9BiqFmP2HKuXoWZdxrq9b+kIhnng/aiqac2U
oXiunfMiw7M8lj0pp6dTEzDnbBDnwR7TjQisxlfsBJ4AcEES/MeybZrxo9J5YRVKUGe+GpeB7zOh
QzVBHL/yWLzqxYKI2HVACqmD9D05MfZr69672mch5FIO0jMzdtcEgpI4BFaATJA3KTeMVLL3Fp3V
uWZ2amtZnqkw/0Mv8lydbt7pDb5C6Vldv/6xxAyCG/353Du+S+MIdsh+pmKb/8CZmpbRHGrcC9Gc
mwbsgDRbyUqKFOvRm2Fq5/bI2HO76CKg81ORLF7IurFe1CwkAAHb0WKvBb/S3t3oEnx7pr0gRrEL
OYw93lRQC9agh/nl8QIQ5jxPDexvBm4bUsp+gPpBsZbMrThNNKZ7+Px4oEm/nvl33Fwk8kM2a5xd
7VXXh48C1CgpNrjq5QSFjGj/WX2RNBnI4zJy1SzlCyiCqm6oL13muMSk6OWJWu29T4bcR/nAAFpM
B4m7ZJZXrTNtuyPItqiRYudVeGwlHaKypunirdZYp6SrsITyKrKF+5eJB8+fvA9YLMRgWvbZYSc0
Snn0GptLcFq0f4Sw4FZCIBdlK4GkEwMTvX+f4af+BanrD+X0sk1wUVuepUcB77hegDJHnDURAB5X
4hbjn2IuMwN1DWfdCX16qGtCmp87+Ns/1KHG/wOiokMgqrOtD7vBazTnGuoP/YQNLdLQQAlJ06xu
6mHr4aWmLmhu3K5wliL9SPx/bmhl1aA2Ze0Vf/3eEluYH7uo+nLR0IOq81gOXach1lPucEMRTiIz
6YuYR+QmjpO8sqqHa2oH/QHyX6aBh83hVTdsnKjcdXo0geq/F2py8AXzz/qRaywbs8pv8Xf1DPkN
HgSqmKkpKWmi9URSjCdX4Tsl+XhIv88hG+wYLPsEpFZ+wPQ2rY5vaV2NYCOyQ7IePZLNE3l6KnKK
DuST5COcNLMCA78loads0k0tPsIWMAHAvHsG8MA7p8Qjlp9UDGRGCCIdWH3gAya556L9FUvR6WIn
jMQd5MIrTCo6NN0LwSIBWY1qqe+eqgNFtKqz0b0XEIOoga0+MbtA+yI+VJvehfwL+FTCruE4u8i+
NjlnGNLHX9Il5q/6/tyjR30ZynSY3ZNe4pz/4FOcaTSIwIo74z/DqVxt/Sflq3qWCxdnRTz5Tp4g
ysnUk9JiKjxvV415scGbH8D+qJODwuafpo7RfkomApdZomKqmhxqlJr+PMRX+gtNeG5eIqwGzZ0f
jYX7gROQk2I22mNG/5DkCFy3mb2o8WI7ig96d8OKTUOjv/qVN3PUn/EShToRy7vcgPtVqFk6LWrD
jSblHraEIurKFeB2k407P/uChBvpvPbULwxZZiggPuJ+/CpL1m/N3SwKP0K3krBIQqiuQb4UtlSz
Z/OqZ8xzNxAKt/if5WjXTw5wDZD9UvrK4K6y5cEW1mtGMA0OWHifCuK2CNdxNWDyuYHy/eXn6V5u
8/RNFYx62GD5mnHtIMCXr4sR3oECLVP5Z4EukFqJzJHd3v46PFchQWJp7n8PSVil4AeFrjbEXI02
AHJ0sG7Pli64i08oneBwrUZbLbmS4wmtHeqhh2oFTUzz/Av0NbLOQkf+3d8Fu7d5Pgdb3+92fYML
9yQcinukAAhphilHoC1mUD0RGzhSMGfsrAiNkz6Hifg4xLrllI5gZ+xvwz76mg43Zw9YxOL8Fm6k
Y1QsqZiIdPfBXCGMa3B572SPGRr59eZszgrltiz3lJEASgy3DLUZNIF4gfFpJdhjdNfsi9FUnFhX
RnqDIvj36UaR4Wg49fbNoaP9ACkQSzG/eAaFBW+D7dgCEWrAzPXgL2cymnyT+RWC16Sy/4kXdIWA
a3d7qt80MMyiztJudBy+pumW+Fq+PEHuWU0pgp3keWUqEo66pY3MCnfn0YDvQPbin7sqRyAXNci9
EK1M/3vYgqJUPBGMZ1HxA0Re1/3YahvU/CiyZtjxanQ4cIQebrJCA6/4yYe6Vct0rkE+oeexgDt4
62dYOkf7ktOf8MWBd3lygD52CJ7rApiR7htyle6iFAfbQOg26cDq1Vyg58I9mJ3cmc5S1jeq4vfW
RnsGpOjwVX3e1wxQKQPFdUfLVcb/xvFWjURh1eyyi5Eb7jeImqyWSsB49zVIZ09LLN24+JbAUGfG
M2LSvGIpkZvTwRoLccRoEPi2fsy/Rujjp6Fi8G+SjRf7SrEN9yLPmTHoREJIuFP8xwBvGEa8PKP/
N8+EhROEHEfi4NnaonTDJKbE6SbUBBUjXd/2eyptn4kpnRBacWdpA0T1r6xiuGA5l5jH75GH91Id
p5YgGfG1HBtfyz04VifbU8b4uHcpSV1BioI2VHrLI2fgC24Gzm0olKAVTbR6jCJvNvgRltZMRtu/
vWJ1CypGy/vcmgHiR82kULEMgSNs1gTU7hoTLhOBYJlFoI5W/zULLw9G2kJ1Sfjx3yoefoDnVldo
T80vdDd9+tcYpFsHJqYlVt82ZqVH2z2atoD9WHi/89P7wHApugtvvIsdbH3qoW4MYJUu0En/5F8J
7QOkokPaBKz+lOAnsOZ3IrOyjI/+Bj0XEiLKFubtqTRyynAaKYnSrFM7x9tbHTUxeV7S+BnWX8m+
5jN3iWjejsjrQFccDjwXFe0fSLdNpLnVreCThSzxyjMN9libYNUENsseiIkdzxK9ZlcrXxPMmNDO
JhFtjyz35I9jl6DHi2xl8B1+xgzL1KrLWWpf5JFWX0uAKUeovx4IlBPaOxr162LuNEWJxQGWhdhi
aw6FCyhv4Jedqa6+hV7ZAdIlZ+UmKBNgeJtcj3L2OF6uYOzVyRIwTHYjOy+Wudff5F/FL2kw2gMK
ZaVZNBsfpx08i3AQ/W3kRfXm5Lyqk+8Ma7mop5JyjsTkGkLKRh9q1mLCKtX7eoKW4lgiiA2Dk9ET
rEexCzC7EcbhEwqIcI0UooVETKz2yAa2LGjdOHnorewwD7pWRSMeiDHTcTqAjJxMARksOcHRxw8N
8XVzN6hLu3J4YxxrkEK39yBjsjMw1KyZSJNqTKUr5h449mQSNl5t3ib6KSLFp5AFFz2fSG4SbYG6
zjs2wu56QBd75hc99se0SYrs+WdzJmf6LCwJy+lpYTKAD8F43tnDuXpMCmn0UTL0hr4aNe7NaTnx
YISyns4hJ7J9I7pkb6/n72X6EFjPAQI2AtCWbmk1drq1XeCqHeYWE0p8S+XXPf+xefeagitaldds
UcBIhAIV9FSYXbiluemBVh/Z3I6w346rKra5Y42we51Vw8JOxEaztArHWIEzjDnglhnte/Iu2vlz
ZIXsH/8DC0KmrKple9W2q3MMOZBKZ22jehzFd8sEyaqAypvGoBlABlaYlBJ30gF3i6Z8rtmrc30k
oIQlyA1cCLAaqRoPMomwZqUiDMLEJ6t8GNwEyD2kPGC0PuRmmeRbcxb98mq80CfQaXiLFObjFTBe
lr5/ETS1m0vC1H35cPmI7DFKeMvbZxSpttyl3yKWigtXS99/s/TAQIQZZ7nBBOMm7gM7Y0lldAyd
ZZA/q9rJ9jsZCrkGvSuhk3rbRZcWeDBP3kMcTVbrjfvjHPZrcVWnvuuq/C3C2wZcLxP90TKtWolS
ub/jme5lm1Ux5EChMU0KfEtp4ZtDDn0cQbPrXRoxs+ePX1wT6nuzFTea2acwJ+k2VMTKpYIbiQep
DlmYSyuRleaEAOMxmVZP4mglwaRNq4r5sZjH96K9qneJcJxTuqqPNUmzy7WfQLQvj/b+DA9/wIdy
iUdN/FNfqYxU59tR3JnIbadyD4IgCN/p2aKXIS1r/YL2p5g6PgrQcpFM+1Qd3JWthgask+oyUC4b
L9C7vqaMcVkt16VDmbfYvK5KYHXx6JTxAZP4SQHlB123/Wgx7pgadKv7iBNW0UuvJNDO5r1FAkGK
uX+RtA6nqBm5wAbTUvbTzTQOIORZzC41dS3pEDDJhKopm8121AyuWdot9EIRl+71jxuFIRPKY1NY
LwDufmzHTnXdkC6s+fyPzeJZP4c8T2qkPv7nXhxB7C2iOhIz5mU0UXlXMJpeoFnN0I5wBphsIIAt
xSZhdOY4LAG59XSSUafsM286eSz7QlVGauWOiAilc0ynEbRMi1FQMxUHT8g4HnETlsx08MOU4rn+
E4KmO82W4o1sFfhaL8prRLR3plptw2PPOvpWeXvhn5bWpbQ6moloFiVf01CRuox88iGHBUGIYsNS
RNrmMKzRZSZ52QVHD4Vxc99vLGOIXWB4fmYF2fDeiBNZ7Q27FCWKpheIxsu7Wi5/ltHPnw8FmmMv
Om7re3GB5M8Nv65QEAEyA1nhd7/+T31CwdOwo3p+YPMuoJvHnlnSN2HxhlzG/pcuOWdv//KtKrnd
dnqo/VEuiecJHVL+vS8wkwVYB5cGs2wBzrvQgYr82cyvLM76mrpCVZjwvkQuO3PAGFs1UMlPnXKB
EiDy584EAX8M2dyka15J3ehGG+trgG5crDJjd5TbDT8Pumj4MDGW6spLNAHKeBmCT38Ebt3B06sw
67NwUwBupXuDXPvDgMNGeyjUzs2TNTawnZd4ezVfYoUjUN/EdxkYRavSvdhEAcOTYjxyvsRQ6gOD
LLcC5+aYRPemrfFRz+oEhXW8AHG7PJeActt8a40IoOTDdXW3blbCBCQFyGZLxhEBYlOqvTPoUiZq
zMk+utdRCiM+sB+4VbRng4T+X4LynvzCn/kNdLkT/H5N45XGu3Eg9/T6+zRvkhOYmTik5nVg2vrj
zptc58okYiDhDqaAIvRb5ruqCgsa1S6i4gQcdGhTUBoynIecsoISUohX+kwVE/S9WPkNuQqydwNC
WrU74zm4zHS4Wq0yEoapWgObyTwb8D/ORDCqzsh2SzxWOobr6dACOrHHOAIU0h9PDc2RQC0uPHgy
8UM61rB4PfTtMTGWsphge7xjkWmtcqwQ4DPSd7qvtC/OUFdQY1ilzkGuIBKb/QqzpU+sqFMNeGIN
h4Q8W/PWhtWMeTC1mPEWhgDQPEvLhuMZTUxUf+1WnVTlxZ95DzDPI9tU9ijDH/4XTMlZU7H8az2H
+m9Ydgc2haKdz0S4ngoUp8Y0eiw75H3CvK5UARSnY42mWiQUbkkprEhNp4RT4QoRlS3sNDDGv/mY
dT9Nf69DmVBFgzcz5ShYUltR+bhdqYXaxud48i8T0m3aG56PWsEbtBfYnOc8yVc1d4s0GV5Vwke8
F5tWxJTy4eHbkghSG4+K7cbJAqlfj0Rx6yA9iQ5JNfuzzoy/ENJ4+y4g/oaln13yh1CjmUJYZscC
Sg++ViKOotZM/r2ogRMytnq0dm2z98FAHi1DT4SSd/7VO2eW/scdy+HniEZNu5mVaUFk9c0dotCi
qkgFP+ZLxTe87SO5H4hmX20vaUpmm808T8bDcwrEuxPkoh5fOq8gTDL+ww6Fu3rP/5iPdSc1uptB
sEzTXieQs05N+uDBwd4sfQoYVfrzp9emsbfeCQaWQGhyYdFrzBuhaFenJ8qQzOP5AoWKzAd6D5Oy
auxn3ul8rzx6Oo4/KNIEr/o32qrKrO9FgwYRai+EuOnWCGq42NADiCMAfIDDprf+k9OeUm9G2sn7
xbwVDQKHHprvC++VEVkrCHg4COcioBkguQ3gW8IXJ6kUhpoN8dNh8mHEnIC5x3FNyI2UnXKk3QEt
TsTcl7aZrpyBVrZ6I/U2m9IOvhusNtne8J1LXAI3bXQU6AMMtuy0YU2SiBC6099v8tWsEHw1pFkJ
ZqjSHqXAOus7Yf8uInBE6M8tqZNM0DtRWkSwAaxJUIlVrcIa5cLvGTXdmKuzrPegGkEsk7AMZddW
jhxcpZJND9sg3qVyYieTgnxFcn8xyCTmfFVZM8QQVMKkWqLMl3tgqDnYa/nwzgdKQ6h1UnMRSiyD
xtNUNur0+8EJyFfWbaQBOCldeCTWbLyvqvSmRRB8NpRytsJaI5XOgXCxGG/efzMlbJlY/k0pOqgz
ljy5gkJzfgIsjtYCua4bUKxr+eV5bY0rAO6kFoKGVPFBDXwaEpQvxLJBL9s5bwagppf75KM3OJeV
2j6MzGpIm3Ukm0wQlfqq8QgiCA2d26tRrNpTyy+hpfmyWMtWZflRjTKM6Hk4R22A92jlLAFgJYCu
0k9dKQ9dlEuzKC1bASp/OdyY7kFEgYA2rlDCgVA9kY4THB/0bguk3RvTO3BI9oiTxXh0jsnA36lA
MC9YjCmS9Z48MFZ9FDNIRJ8aDokQQJYT59HhZhzL4kQAHcAIbTs02RgRUmTb3uLSpVUTVijwZoVW
IvWoDvMTWqSbTwm07ohcfOhNbWG2IiB5WpiETHmoeBNwaDwleboaoE/gw6wPj2WJNt4Vit0Zpwt9
yB/VwwAcg/6JdFx4+4rnkbUCnhnw78mpO6eXScnrOz3hU2XcBMPKcAsnpNfekag4wjupcmwBBuPn
rbjUsfpVia2u0jz8L7bUR+GeYNcwJw/ft9uyJ8jKHEejorcTuWAsBZKIzj7vzNjM+b6/ZMm7CRao
J46E1VzXIMGXfFpI6xVyFzEtXt65Yzmfc1TzMkX6KvAAifMscJB3g6ukZ2xgYNLAL1dPL6RBpW6l
8COLnMsaEgXYFd5JDWP/2Lr60W3vD81O5k5DUJdime5VN190wLvigENuqFVor772uxMH9A0kv+/B
/FElYpf5VnyXHJwtlUcZZh/B6oR+VPMo91/CpJcvjLv9yC7f9nRYC0uk6SzBE88Reo5q/6UKUNpB
bG2hhHwHy8joy/Yte9LRwnh3dU80qlsy7g+xXHTlIkaK1FtUgW8dj3g3g2VSWZ2opmr7f2r/bDcm
Lkj93Ej5jSN9YgZCtkUYkEOSCG8QlliQxDML5V6RDIkZOq6NHCNEHOClYahPgipTymQRZQ9TULAl
bh6lDwhuLBkAzRKfLgFDfeNqGENA1z8r+tknCZXXrqK9IVRFRYyZBMCIHGJIyY+eM7MpzmR+RB7h
S6rwYcLJcanPHDBUhY9HsVS0iKi2ovtHMvFuaNX3MdLcq/5GtRLGvSJBP3yfeIDIu0M0hRvrFMt/
q8+Z9Y4aiGX8yMcfoPF+OYLqfWnkK51/DhUlUP7kgf0eIp9iRwztCcEXcsPuZaQaWpX42B4CFn5k
Xc5K11ot6Ii6pbZHiwSnWByn3ZfebzhHLbwFjvmwsCmk3aYjqEYuokMoThlszICOSKMDEnaNFzhJ
Yj2HaUktFq4RNrYvHk5S+76op9ftcdmycz/kD9q6TgBi0EYK9YhdZZNcEnSoj0J8WCDPczYcd8c+
Zn4HJYiwVDJvgYI2V5yt9PqO7efX8u6W8hI9BaZKsgNi+zrBCZ6wh6tr2ZJaJOvIUdnj/UDPCzmA
n7cAF3Yy2t2HvV3tS0eBUJDfcPAgvD3HPwzjmdeURSe3TbTw3xDyX7STV4hmWza3iNcEoMCQfgsM
eJlmABjLrhZiaNk3e+rmf5XBJ8Cggy51eYF232Pj6vJd/Ow5Wc6QMIBAP1g2+/06W4cs2i28R86T
1Ri1kQZvLkzN/0xEzhWPUE6pep4PNDOPDNnA/9XdD7f+/VWMkVZdEZE/+3wQ18ZvaEaANZEZcmbw
XMWR4Lk4oNrlAkQ3sRSjuCuWhe4nd+auHADI1m2YsvwCAgz+Yogq8J74NcjCeqL0uUZXe34DKB6L
HK5UbeeWocvKq4eaGRIsT6myGy3hC+jjP+MVzFI+khrkrM1TEqBpaJC/esIQ/KywK36nO1keP0/2
rdNgwUB160dO78K/h00TRRGjhkt/e/XWDosLVMCkPlMECvTFZ0X8xzG9aZ2Y6AnhGQhwYvU2hDKK
LGU0sb0ogCArtVTGUkyX3niym4DFJ6NzJyvoRfWlrjB8hqAPGZIQKWGt8dfRxNJcg04RCIGSGHFS
Pq5+Cfo7ksv0RvvLi+ZwOI2UNUzbRAznUK7xhlt02TYsIt6K5se5XQv3PVEIZ/QZMC2oLtTuHDDS
Q114gKV0pIQYnIG5P1YiqKI7yUyBM/aKAM3/iBDOwbmpL0uxZBfB7gTUMRqZo08pyUs0QHJugjZM
vodOY63b5gWZg7HsVbHP9uJy0bOtNGacirztL2VFq8KFN+3gtGc27jFlFJ9vi1hGBWwCeJ8/w0w7
L/XeMPdRJWfzZwpooxDPF62wrsZ4dQPCBBlMICfIXYPexCeCXoAUZpRtl4Kl0JBpTp7NWo/wJIu7
Mbw2N2Sd6iAxW3ffwAVGSCuijeIXA9Q3n+Ek7G/cDVNRueKcthxML4ePS2NB/FWdEAscROgj4PF8
ZT2EQ/AL7RmiFBtlIXKhXOO6kK+MSMl452L/CdiGH1WNO9r2EDT0Siycz5bP4wSMHY8Wh87N8Zoj
yCtl4P7gS+k4DhAu5zliWZ9avKsz3KPb3B/T5Ospm7dK1CiKV4qXVFNwejOYTA30mk0CWqQYdP9f
BkeIt+cbn6Au78SASjzYJwuSDUQ3fRc7mc6Jw0zBULodXurkaHWc/wvv6EeK2OJmk3SgaUVli3Xp
PHJmGT8t5POUej77X3qT21ZKLW6uAIItttdcwXfHbBpqZIJ1cV6IRykwdeJaET/1lazACRRaXxsP
eg0qf0hKRydvVQ2fSwAM5MKrHo1a2+EKeI/eZnAnOGnrgtBdNd/TrUH4b6FoOzrk3Fp6ZkgovSOT
a2X1B/L32OJ3XIRLl6PXF92MqV6Y7CZvej6/oYG7mOApQgm743Eo0mHbXmBZSV2EZUyP3yTEWIJ/
/kfdoDaW2LWeuHAcmiuWJ87ZJfKNytVhVbX6FiRZcO15pImHCFOlERzwOAe/Lz96HSvnXm/cjeXd
+P/nqItQEfN4PAYh4wGhnSMxAcdsem0UsPdwfMKc6ZdH0VRA0Wouno6vA64nFkn/Dtcmn6zhD4E3
86IDLKGbldi5tXDnmokueNBzLCb8IlEHQMt/9yQoyqA4nN1wOWpuk+oRBAcjMimk3RM2tp75LXQQ
tpVA+mkGovCoqQ/Fvpmp4p845tEc6kJrLlCJ9GUIk3pZDjs/m4oKrUNMKIKkta4rJ3U/arGSwMFX
ss7GW34ALqjEeBCXkjAjTfS6cqyiIr2qAfY+H66GXz4eKDx9UpBPp+MhPqvnM6Bw+Y9CU/Le4yHo
PxXk6Gn21vhJoxDBVYNQ7FRkJngctNIhADMjaMAMFF4eU5nYUQI+ztY+tgucvR/h0kP+2OpP/fbk
BWapyEegqDLezWEYZ0azGDxC4JQsblOg8RjtJF3qANiOznJpQLLVOwp68uZLvrK7GTrV7ip4Q9ye
0DcKJpyrm4U/dtQFzGJjf4hCUGgoqy0zZ6e4DJ34LOinzcCes0SHeZPmd0IjxEFUDlt+pAxyY+C+
g4gUcJBws/zVP207yhEBgDsxq3TE3hZ3VXGaptCld5vFgS/Ec/qNFNaF0zbpcVGRS9ussYEgc3cl
XQQX4B6+JSy1kV4xySmIx4nqme+Ocp0XlNbLmVAaURvIPtdZ8pHdDyEJvUxCibOx3A1j4odqfL9n
UukC3Rz15JtdAIib1CklXeD6NnyqS3t8X5kEuyPYyEqT5+PssGsN2Tg1uMPDVa3lVnBYhEiiCaOy
16bcMfK8VG8MSZD39/iUK/z1PS9FC8x6pGeofUNo3gycaCVdMTyRo9L2sICllLrBd5VGAiAIYH+T
9OJhVAjURsdHPhMGCI5UMNtPWhHHG5UP95YikCxcFL1MsM6Tn4NGoQIiPhM3g2odAnpzBzghnJwD
gZSOFCLokVBWZ+QykKSK6WgCZbvVTqPXqRp64fYjymOWIO86FuYZnX+Lfcm2w8kGuIrLCF1akuTB
2x5tPj1NQQRss2ZRBs0t2MvkYCYr97LBeuewzB5P8aaBfRukrl7q/h23b/lVYd/ggK6RBzp9Ob9G
Gy7JUri4nqbmCx9gH1AwUY+KWAlOz/AQVFC8+GNhzwh0WLPaIehZ1gPjGz2fxsNAHy03fRL4fmxw
F7GTS5eQ/lD1UEyh2+B9E7ltlCHKMkLR6DqUFWnAJcXmO+lngbJzzeoypLLcWEd5yWPgy9iUijif
5s8wTJJ8B1Hu9KSv2Qnz19PnOSl6tVoPeKIxKadTkJGSVkHKhGB+5AoRk1//IAxzaGIeeGgJLXhZ
vLJ3CGZPE6jj7PS6Hne3hpMs+MUdWsVvvf2FPbPdHakGKNNQY50Vjpy6qqE6LkkQxpLK3brBHPIJ
/iaudgbkS2FlLJJ+zisR1tLmPOPWn9unzZjI/UitnbT3NSaAsYGXde5ZFse/5SatQ4QomS57iAzO
3+d7tD0+KHmCHYlWepwXHjcYqSP7ttGk/d5JHulxcQsJpD/gX/TxXUPfo3JbLj5QEtoJGvgxCYsX
bS6jlDbLPmG3oFt3QKUFaZBRNtXymQvJ5QH6SyWW/n124FO/JEGpR1um/mFcSwxaC/F7QQXTSd/Q
7rVNlKk9UEzbdaog37XBHyQ/vJbCsIzplecv7YB+6m2t8EXloRliIvgErQZWUzXsQo0gNDze95Ih
lJqbcGrVxjYNh79gmnfkTq8E6+/RgjNwW9ivcsSzAf5X4TjqD9FSNwS8QTLlXtsy8LsnL6pZBwDI
keYu0D68+zjBqGPr482XtFA/e+NYE21YKGnXGDYOVlfyUZzEnyPfDO/yQTeXDMAv/tTj+3XtBy/O
ottyba6V0j60YRSNiV9Rk4kUxAHCBm8t6JJFMwGjA7rSO675478T8En9kcSeXuteBqp2V1LrPlpQ
wMMeMTgdKAhHJzGrkkpa6U5StmFlJHeHw+S4oAyp1kbwmkVUJjod3EIhQlIdrhi9/edabiDUoDeN
lCgy5Od4NcapY967qFIShjeRPQLpim3t4LhDGztBUQyLjqyvhQjwVJ+x7PtUOKWVtXO9rLO7KpOh
53xZlrBgnXUFZxf2WJs+0ggQkuXR+kc0hXah2yvxE82TDcKMwqZ3H2YoYGjXwS27cM9Th2hKMTxK
Jq+h2YLQAtDG1VAZ0THT2ioxSTB+YRopmtBLAMKccxCoECMR1yj0DaGUogB/CWPLvw8Vk+9hw1nh
B4CMoyqbzo6bg0+9ET8Rjxr1XApK2sImt2T8OoOtNlQ2mZaSxviGX+Ut61+ST7Qadw0k9bWCgPgn
+8xbDTsnR9/e8pMqcNgN94hcX4ktDtNbOgb4zl9HtYGosQ8lDI3A74LPDelXTciK+0rNTdw676hj
HXpOrYZirX2U56I3G6POyfliCC+YUqQVaBg2cerXqk/pxe3OQCjGVcWz3tLHbSo+CvEc+girBdqn
0uB0sIbyhClSYRBZWQuXYtwpnS0oi7li+yKk7FJdalXnnKwbupSerI7FyPC0cXkWeoheb8cT/23r
DuSIj1tQajbsTpDT4uzxjS+ff3NfsEAPLkBsOo0dJaUK43z9J/ilDltVemyQPa+dtoBDT16RhESw
ii6uBgiIh/w6/T6hTar72RpyPm4WcBPNrA6M+jrMg1KgTKusjfcEuwQPLNWaC9Rh1SQSTi3B7Snm
gkrFqvsl0YLpy3ODiyDxMKLNgzJn+dOwzE29iRIgcrB8T6xBP92qr9pdp8a3Vv8gRay6ajD2MdhO
PmFVN2CyIHWAiMq/ZxyBgdqudEOfVC4GFCMjpGBZsWc2LAlnEmtFTiIH+BAwJ5i1JHtZ2gobR6Zi
wqtHH0IFcCShIUDfZBZLu/Wi56hAmzhFC41+cpgWR6knOYIceT/h142YlifteTV4A5A9xQ9qrcA2
6xMS5p271j18Aap9UsT+u+nTMSk1vDr1gHN1RSitWsQxwq212hZc0PQSX9NBNh3nGVzr87uxIqv0
NgYyrFmUICE+ootw9nY+BJ1U+teAZeD74LqTN9WvqLfZI3gn6zpRcnrclmhajiflqGRgtE5E6TJb
NwS6Qt3hfpU3PyjLaG1TPlTH7sOGcLZmAk44wplbaIzJcOQXUz0aGiWWaP5azyWkWDd24kzfujYT
yo38xfW/27Q+uSlLDS3djrfAq4yaZZuD9TZrlvifKVFRlbgbUyoEGfQTA9HaWx6iJKrbGHRNDhOv
7SEGDHw13+j1nF38PJZPOLlc2MGbmloykxwUMIH8BW2dQ7coEpUZphzEEWz+ZUfK/ZxAQeMBo7h5
mATS00ggeM7SE5+RDABIs4CLx4XZPVFNk03DpDApgNN0O4yfuxWSCsNLbt1ZjaB9AJvO/l17SLkx
73ES1UcNZTlXq6wi+/Az5qoglvtllCvJtQ2ho3sZvhqCdCJpUjGS0u+AV5izqkD0111bmJ6kwgtm
07Nq8sCh+zx+qozRuospvBe1j38b5nAmN8V6k5biQ65Y+88P3YrfJn56FwLyDDlBZge6s5bzQ/g6
QG41pmK6zEawwnjFaTAe0H/D4XYDTUuctE6ZvzThHx6wdyR6nNZWjdYcqjj9YZqqslyhuY7ZRiff
Lr1wmetooFrdOcOGSW8NoR3VtB+s5dIcrLlef5Q08jb3YY7CCgb5sgCSmEZTF6SVm4PqN44WBza0
7PC5oEdOjJAgD48VnH3aZYXHHrp73F6NovZrSvBtqbvaUCYpXwbltb1GcEFaBALqz3kGRngNqhdS
I7DzvRzYr1EuhUZn34haWm5F+hLomu1fxWuLO5DHoV4o/Ea0Ec1xO2zo4Cq6iBu/4J8wYazbjNsA
4TwhSqF+ZzeLLmHDJgW1QObZP+Pm1RP4X1bLECS3v1M9Oc/ry2MvxlV0ExDrGAJQ3sp4cV0+r5EC
qxD6Hjh8uoDfrCavPRnStop2rmwvq3twdAoSpEueW1EtdfgQcNbIM97gLnl+2AsUUFilZW2dRM+2
nT2j4WhoIVv8NQXyllOtkpUotlBUw9vBl0mcQ7vI601uxyYCYPfpbi6bJCtjWNxG6P94zGk/uWaP
wwLPOdtgtJVAfyaWSgd65bjVpvnUYK3OPrMshPxe3jaBBfR5Z3hJNXpbyt0hD1+wm1wGu8u4Kn3K
2LhZfaiwFNWjUYSi/SeaVMXyQunl5/gaKe1KaEk7xI/r07reBDdjo++29qdUIFyU18/uNJajM22Q
/Ws6/5Z37GoQF4eBzI8wMSK6QJLX9QBplH4JVKVOsyxR0tGiYtNoOl1z4qslacLbOdohXTeHMI+1
emSQYf1SzEezvUp3zweTZkqPpdBXboygN8CHpCAo1EFyjK2VGIEVW/i2wrC5VKhsFIUNlb1x6ggP
buyE84iv/ADlEDdEgNPplQ+TnSmnM7RwcK/BVyDbQm2H/kfScJXxrQ2z5aFcuYqK/Qqvz+AkimHs
zVKOkdjwMQOW3G5H2JCQknqeAAIDhU90WL2FlvKZX33sD9Laqln1+tlr5D3URtPGV+YqsVYjeFIt
M2zhuBCFtDIqWoprXViV7JYCWROCDUGblwd4Tll4CTaGkY3x0amWYL6LFgzCcmnlqazQjFbaI4aT
Z5EzMonXCkvMVfEURDn8dxggVCCruIpxGzB4OCPibGvr0noPxU9wDqHq/H6XIcWrwdZBx9EOzBGI
ATvyWCvyE5KcI4Mu20eFWgcb67iPHplecdSvK8Y2Vz+NLRnwSIqhHphfs2yKQJ9nCbpJLNZyXkVy
wYbaBzMyfOUKUPTnXLXjrCRFwfOWQGhHbAVxM7gcA2CPcO7yeMqCG8TKrIysO4bLIfta6mHsW69e
7Qx+VxArZAvWHa6Glu5XfqE+eW8SC/GAEVqatRD7bvbZTJD5xTE44LSHZTgvjKR5sLN7tAz/7OVi
vt6ino7gOeCFnLqinR8/d5rTDRecLYuTIh4XwaKPzJQXpuPCnEM1xllt0XdMOUiwYa9RvdfmRQej
HVySA+8RGv3ZMEw6hD5fC2NIALunXvqN6iNBxH6GXY9lxezT9VjTidYrPEo8uoppMJFTJbtFFgCH
jeWeH6YHMxCIlS+GK3wn1x/r91w8Oozfq5zMHiLhWiJ5I9zoBzOJWL74wCueXlIfEsSKOzxWoHGp
qBLYRpCXZhuRka+Hqi09OPTgcjijNI1cqgpO1PcRfBXHe501dy0FDVrJWKD18AG5gu5o2u8mpcJw
VVLmw9o1bG6TFldXfkDt6AviVCb2aMp+htHjStyQw4TatBFo9dv+JIbV9S70TrqTK26KBLRP5tPX
OVObml2yaSQKLIkRbPRbB1AnKiwQUM0OPbyBqxqqw3UJlU6kd4HAUo8fBgxhdYxm0uj5JtI2uKWo
qVC5PKdRKuGO6I0phQ+hljLOUQXhH+dXHpj4nqORCTPyMEgz+lVxxFUyms/HjUcecRK4Va71mWq1
jiP8XFhZq9wqBbKzVlWfLctjMnXGgJQCyENSCpjUoBCUo/RlBqLhVGZxSUiYWlPvRMSotcv8EKbb
gRfwY1J7gQP6s1JEQEaAg5bpMw3KwfcKCLbu/5SWjKSMkuYM7zPd8r4IURHZQgDQkXHUEVJ1Yhc+
33kMWc4Vm3NShLsxXmuoz3tlGC2JHfboApsJb8xbciQU37gy95tj7EchSP4TH3g7bQi0I7XZXTl5
twPGA00DxEQJmlycJINDmD6jn43UFA9mzNY941+0Y60ArsfksqdgpcaDX9ZI0VoQnXqlmN0xASES
nJvI+sroXe33Vg7xtqCnXywcBqBQVm8BrkmwdPde/a96Ox04JVBYcie8+5EXWn3FDM5fW5Eba2kW
EpHU1oEWEMM8pzCyumwRpBFeF7efIl1m09nc2aBWSFAj5dpLJnU69GCr6iAPzOw41F4/iPHLw0+x
m/Dqod1IiGDWHTkjaFOSeqKbJZZQSOdhXbfzCfKu1O1ZvnEPymVsz2sngiJDAWg/WpPVr2iQJgJC
iEB6o2xQDIGsfX9S6U1usUjEd2Ki6KE9/a8c8rMg2vbWdbGlArmKT5KApPh3XW6/czwO5nteuHAD
1rbCeJLw/yrLWvdcnSG5O6eArJpNIRClYdmdzXOsfdqXwg5eL2SiARN7C3dkY1uWfyz5s7qg0S68
A7FFjjxPhpiJaoDl27U4TF5WzzOiq5VwjIotV7DtGDVSuSEDQd5J1IxnKTg/MPPgu1NYRQXscdQD
P6gwvYbf9Qe2unLm50Pm3d4Q9yXnOc7uO0Vma8xunKnVmaKNIrd4n9QzgJ59Vz7LLUE9qKD0j6nY
EPwyTBxZDY8W54fledZulLb+z7O93+FfjT6l0cq1gEEZVqlFos9xxvDHtIJrANKBao6QTYSwIqDp
lSEzEe5XliHKEZDk9DBOt0wvjAfnQmF8bjfERHwJeCMxNRBndwSukA7xxCrD/QoHzZNQvi9D5kGB
LkPe/V1s3DKo6RqRo6eZaxYfZ+ldmT6fvktG5hA971Dmfoaih0D9s4jd1AjKgIzr2QWRr8ptJaAv
oCzPOidn6CdSd/vOZzYfUjqcElurFGeqNJKb5WmL8X/NbRK0M7yWF4Cs3/89Prffb9Nt08DShwAF
IpN1M98j4Vs9O0ityqF3m+CCv0jLG+k2FQJ/hMila55MfkMIOPq/u1armGHFxDPiTpWBnPHVY2G3
+VzxWIKvq57CKT9zzSPmImFneCn/gQjHr+JWPxpW+8IgFlkoGLxlYE7bv3I9E407w7+IDFxQ120I
jEGejhLmmTx3tvXisygq31jdSbNQjvaTJ6cPKLKT6yRho9VzkG54BRfMl07Xoo2oiFfAgLdaFp/T
odHWo1HLmaYfV5VG1DqVux1Er7fgOUCwjKrxbGgfoF5U0xGXjsWGCqD4Dibik4gJ05G96RD3rUnq
FSuyC9S0AWeGG8Rb3XtGUNievbMidzbWk1c696VJWR+ZYtyK1GqeJxAIUidh1A3d5XZdXTXAXbs9
jH8XaFAwJhSllEocW9gI5wPEAPqaf848Hc581i/RryalAdyhZPoUYxg2DXeM3wxFd0a4G2KR5b8k
49YIr77qtWGCffPvcnmK+6GHUGL/y2uLkzymHdZMagOvIQQE1k7pCnY9L260nREx+rBowKTVnPDo
MPNefntr1ap+4mIahBaj0estDTFCHVESWswNm4nyDLcmtB/cZiMsvvPaanSHb4wMxz3TWJB6krGq
PmyUFRRUN0PPpLo57a6c+LY7VCgZrQZNhEvElQJJvbn/AhYBAhh6YKI6GPu/rK7issPBK/ArtF0K
GCIKTq2cpAtAenII/IbhlrhnbFGPmXmd5a7zZbi6FF4i7SzNMT3EUp/tlv/hyCjVL8ZxNZSRvZm0
MPR+UAnywvqfTyL/ylyQgmS9BZ4So9cdwobrKOSwYJWiBTMikUf3GhHTaKcl11JpH9i7owOQzgcp
BztiSgyt+uifslRQhU1lR9QVxuaE2t0ICkj6hT146Onfe9++WKdxNaz3iq+GMg2HkfZVr4HPwWHV
sYzRnuCXilvrWfnkVJ2xqavA1E6nTWnbZ1EmPYVsezqK89aTJxn39+rEuhQ+zlo/YPiGRr4Xo+l/
XSEznPvzLsgh715qRNEke1tYYmD6cm8G7GEiY7pCYP1NDMF0a64Rjcb8py0zCeycO/M9KxtB+nDG
QS1BExy+EBaay2r8+NIi5/LaY6jiEkJv69SXh8a7lERmwCPgXbYzO4OIjJ0nTyvGks1PqFNhFovC
86xRxyupmZXIKTrTDb/KHsoaKiypYkXAPn6zYhFeasbBThnilcDYlf0wLWCa7eT8HqovOJsRckxB
VjTTrsJiGBueSUt3i+nyhUYsAtKTuUku7wohYcInn/7tUXf/n23iViUtmW1J3MNuI3GXA3pxbcZ9
vRxUX2gQfdYOeCUGR76wQG2tweFtOfOBFA6/deWDOg31IGJO/GGAAN6cDSw96VZ3ZzuCSIRgxV2U
H9bGIbEawYvVmi0XXuEaQAEEdwc8qdjbxdGbVZhMA85RDouei5l16Jc9wJLHJSkWvAes05tfDxlX
Z7sRmS8P3pvlnWXVo1zM1eIB8g3ou/XXXmB6ifT4PU3kROfZJVrAMl3qFkHMDZ2/Tozu3PsaypBV
iYE2VvWxLDLgPqLv5AcQshP44wgg0wd3aokqPFIafapwBMNhTXFEoO95UuvfpVPwmKw4BztCBcOC
idqNV181IPjZn/6mGHFghvIEb2rm+rPJEN9pV9h7Ad1AstBiEooCncoOMU8OXps3lRQbWf4/QlJj
U3j9kJcLlhFIUBTfRAmaVGnAGMeTY6anxTxuf+hALBuTCzSTqBcNteA1hnJlEx5d3anNBicBqY0Z
15k6JXkNofQDnmxe74E03uQ00u4sZ3ORoytMdG0HdaW92TFXRoPYlhkSbAXfkrbnXfgxu+DtOKRy
CCUBEC8z3Lx5neohYxZJr+GqP77YEmapAt1l5eAie9b4UW0cok4FKTPjaVIEfi2/dBD14OyaxuHV
0McPaj8G90qudYi4KFKOcTl0670ogu6RMDD5oFJx4gMeG5YmEBItSsv6Uqu1pL4ofL7erOYM6MnI
HjiyC3c4YppqR/z0UUNmrj9W82T4NuwLuab1ENYwEvB67GXkyMjoDEW3TT67VO12/gzt8yDEznQD
9gR0XMcWXPxQf6xeZrXmz3FMFKVnWEkoOvoqqXdRc/HppICJW+LElJRJ4qktjAZ8fFiSSY/O0Da5
FWwMO3dA8/Vec7Q4e/p3pgv/Xf8X0bYEZXAgIC3J9PK7R4XNQzI2YYpyw4sEHi3wo8I4qG3ywak6
Cgs+gGVnnuujqXImiSTIyYsC//0c4S+WspatV4Uh0LtAIf4V6F0LcTSvMa1IwB4eE648iZ6LZGEs
phdduDTUe4T/3/HpVqBoZsMI1N+Udr8iNRcb+HFYtmIgN9ZV7N6ww/3VgjFttrAV84yLoGMy1pbh
Elfp2YGQ+LpEu9lPlwfpZzEuMQ5Eio3ZDe4rHUgfhPemuSzhWWeL/HW5+skyZv1IpHO6dhK+a5Wy
vstUg8YgHkC+Bqgj+q2S20FQm/CjnSuIuuhoGptqaJ3ncESpnpqmoX7E5TabmbCw1DcyD8JQHZGz
dWbgEpjLqHB8Sd6CtiR2sKmgxGNgDRxxDm6Q8RCxTThXquNWLsnNRnto4h/X+jti/uXWAfvJpJf9
pq1Xk5/SmybqQH+XPlvYcGQT8KxRm57DuqGgnNi3iXyZmHpbZYPtYLD5WjQJlvoncx/m5VvsxfWa
NZVaPjfVHev6zqOK+pHCJvv4XDKJ/z/+QYnhOBnmLC43mbDn5IPlQZFd5/UIL8PP/mLAQypaBLuS
29HelNh+rAXBxBvPMkFOR8nk++vOeCq2lYSR486p2gznBT+A8eH0c9qkGkSMQgiPXLgLv4Dj08Ee
LsSwT4Z2wElolxP9IMATuTnfNeMIxIFdGewxGE8td02Q05TGHOp8nxAayaR+Man+kySknsTVnpcC
nTmF3z81weHPssleuYT9xFJUWDZrgLuwBUoQgMKFFpWwvJnq62EecgE2l2ZQQhvKwatifDzBE4cF
P39JBdhFsjHS1ajPGbePZbQ4KaPOb6lufd1IlPn+QX3i2Xn1fpO5fVdXLYw9gKITmPvDrbDwLIrT
MTtBpqxEhQl2SxqVsYPUKNEhMfb/BPEB1+yAgUf8opcs0i91TmxlcEyLmeNZDpuOemQvpkk49UTp
tbRjf7jVON+pLTO3GFh3ntKc33hfbYyL/h6eMznEuUBaE7+agl1VUTa8NgFOzlg6ofNluFun4O9T
54BxbVfNV67IBykG2k4MT5xU/tTFALb1H5g3J+LrK0oU7Of1+HQNw/Q6t7vD4hGa2AjGr6zoQiU0
J9OZBIiEHIKBdHb8iU5DH8Uzc26RagfR0Hdd6HAgfX3eoXzUSkPxpfnJ/MS8s+y+h5Tswndn9LHD
eKf5prL0VvwirTPkpv8j0VMRBSE6DuRW2fw0gvEWZa/8NS7BmyxnF6866YzEq9BBwOJx/XKZqSxp
CT+UlFrCcR6+wfWisUXb+gOZDTw8FEZn7k2QuhYgDaLS4Jfa2FGA7D2GaLNmQ/L6aibbgdvXIHOQ
nOpaYrZO9ZEs1CPDUxBGHsrjC8nmEBOY0o0akoylQY3WdZEqULBtUAZNyh0/BtHhJb5kZZoeailk
8KV97SRo/PzlYLqAf6qGApDGy/OzCmNWKCHuVKizyCLNq65kN2ZwWf01snE7110J2r/qJHRxJt9m
KjeZWOvlFkJmtusdne0x6RAxyHdbcRBA4obJTP1Jg5CcQYB/QfeWecYiHYf9fCj03mwtwqOwJqjI
yiggtkw/HKOXo5xLgX1PaqhkFBG98j9EO2ya1oqn1lBc7Pzpi8omKnqok8pWYOKbs9vzMjh7ZRpm
2PQa9uZo6lDgZBlvzFx5yaqtRqrmWAZcG/9Qp77st1NtcMvg99Lhapz2cH/C1LQ1hpI0CY0b9GaI
4SOpuz2lgdkwcWy2zbsNP5RfMjU5Edbrv3zhyEbKm4HZaY/I8669kKkomaNvRuw1oW5M1thdoSrm
t8MIEF7gjGNFjoiEJygqXFiTCCm0yDkauSqvyxpJYv9Enb4sPQG6BQyuEW0fnIMeb0stkle0pQFq
/KYwAbvDazAFnjnpDNF3kc3zm3vI+3sC/sJxddd4BuQ1ClDbG7rS1ckpy77s65rUbJXJPvfavtim
LRdl7kUHlH2cG7fhdmHuz6lMfUIS1X0CxHSMctCE7f4fuB5Qwe1S16lSuMxCb3a8vM89brNCZqH5
5ilT7cuMtmbZW8BmtvozgzmmKp1/r42X5QHHYPDTwGHvlBq7ltAVx7WG6BQC+GPey8yoDD9Bf3WK
gyWAY9+jv9IvxmW3nqD4fbng2bpdjRB5/tW8vuC/h+z2qMN0CSnPYuHam7UAsezueE5/Y5+1BaAd
t9BrisQ/QlJfrN6mvLhYA+IuvETTU6mEZ8WE7OJvR/QzbDqpyGqFuC4vz3CdKJM9TQhEsD86tKMQ
ET1Ce3VheN7TwC7mKNVJv99wW/MfwYCyYYfFwLe2vIYGANpgVaoV2kS03dr4g5OzQ7dS/ecQYKew
FGTiYqk628ZQURfJmwL9meRNdDzNZ8PvkCh4BPuviXtrwBkwMgk/izP+RIgUdnseJzAKmNekcFZH
LV/IBmvZhvPbD81JrlXTknRvGECZBPXU54ZHBKe4znUrHez899u/JDUBcgB+pZ3tcmfJ5BPFQvvv
g44ti9fIQ+Tl+9E/hqeXpREKSogB+xhtLX+w2puUJOZwC+ZJhkL1u79Ze8b0NeZckgM72ggZvNM7
lyiXiQwWhOeXnaYHRH5JrZi+Xkpy0uZ4DPmEHORJzHLNjsvGdaV60PGTzRfqKPeukU0x30skXbmu
bCzGDY7lH7PXey1XwOZCzjfqI9SHGfeMhzrLKPltsK6kzhjqTco+Z/p1xjdbtFAr81MW1OHz8TIR
5eqQVbAcRFup5YHfcwwxiKQElcs1rNCA0pq1GojXWo8YQQ1deVjBreixhoZQoLjW2D05dcDvG/j5
emATBKmKCEBdu192WDZce4KN+aNi+YKg47mNudawUKb851dRXOogkCWf9wcQJSRloUFcRdmDSy5E
Sc5KFgdQnaQAx5Cq5y8cTcF7JB27jC8wSDGjXlMXpEtO6BNim4LZypdFZYVCtVkEEA3ZrvwOmKm+
0nnjM5xm9QR4vIR6vlkkDFADskiWcmVU7R5cqtW5sYLs9wFu/m2cbqU2FPMwhhqyCIi8ePkvx0w7
C+eYrlMjpNJDoWJe3vUIktn+s9OogAdcdJB0rbjxpTZ/p7y7kBL70TdzoQyVp9iJ9PZesWBkiY9R
eBf6pK3zRG/I64/IrNr1n4i2YwJOqUCXFRpZoc5gZ6cnlgewRTmXWPgmfkDIavVq1Bz4MD4Mtnwk
WBx9wpyzSreHU+u40B7RYfHe5keGS1zGyf559q/IVSJJhLLgJ/6nJDBqEaPP61HXliZ9Lc3t39bs
NHzPnu6S99JKDHl3XiDHtEPxAYADyfsJYgpFE7eBNyUz4BQ9EuV51FIJiOlGIM9heMN3a+axF5Ru
gK149wgfuyQZwJv6Bedgef6iq3MRARiFEo0S4cA2/4ic9kYg+KfTqa8lN1CQSkQ4gSVmjrgUwYbK
ih5YccZW5gjWlBOVWKJfEqC9FeNDNrIfkJPqVsGa3Gdch818XLrn9JDTsJAG5qYAflvKq/dXzJqD
ogPrd34fXZB7r34rULKYGrFEgEXPesPBzttqTuoIY2yQy3OzOtkuWFR4UQ/8mZ2F8Dq1DyrrkEld
Wgh+qYGK64P+1u3kDci5bijeiDLDdxGR49HgvpxRUU8NMdTrFhCG6i4T3STP6RnT2CRawWdupa8F
StAZYUXk0OK3yiPOU1kSf/g9yytTHGe10N6V9M/f4d5dWUjit4g8kd8QvNdl5YmccEtv0V+W5iWw
Hn3yJWgF96V1SEeJ9BR3l/+BAIULqxe6nmRUc0mRgSyBo0WSZxx3PbGPuyCUdCEBRCqqcO0k59th
RF5ROSgGnnwFt9b3eaXwWEMjM5WtMcfPnOn3gcLNhzWXIj1u57RJ4bmzoCMz/TEESg2FObJ5n9oJ
jTvguXFgUvit9ABYGSArKOYBdjyztErlyyafscq41vdqlf0tl3gpYeXhgg+ida3LcniYn+HR5+5W
Jaj0nIKBtOJ7rgpwudJpzBScjzq4fr2CxTJqj+RCmkw5PU2y5ZOQD82MIWDO3baExvqdAg0U4ifn
bmi1YX2xouMfOKyKf7up3fclXYFuJjSORzAmo3dXmsWDe3bG+gLOvAEuKtAmxZHSHH1hJqRSwarN
lyQaq7LgfqzVP4XMYC0HMUzgF8uySI8EZsanqQg7soEGjEcn6PwKKllOuMESDvZrAGREl2OHAtIB
ICKHxjUJVMXSFHabBgzhccQjMhXfUd33WTouCw5XyfarAkKCEOuF2xJm4oibdtfpxIYyi2Brnjjn
cNDx7wTP8JMGg0gYjRlc+8KDF+UpUx+JWgYaGn2xTsWptvFyHLm7xLhY0HWiVZLLPygNxKqQOREn
7F2G4+QqkmZnXoCp2iQTW5QPXzlKYWC7OurBDpuQSuq5ugd0qDg0I8fRSqth82pvdUzDs8QJJlZP
Ir6Zw4mC6JxF9P5zpBsaY4KRnSjy+ty5CU485WFW/io61HlCEfwyvrhGA4DNRTCG5IXl/ASGudC+
Qyrq8QovGmUNiDf915zN6L+PviEV6NnKes2TeetNwHZdEdY/tCP5qMJklSvk9ziv+jQnfLg+OURR
h9s1PeGApSdZ7H4eS4GHSBY6jEPXDO3szjkqVmfOwkXSmRvvhgh+9hVAGlcjC/gvwP40CIdyAgzH
QF50gHqEbF6yxREu2K330IRT8Asc58GX3KKPGCgi8xudC73wnNGhX1c3FUM8mdgvqa+q00QRw+kH
QC1WCIyICgxReXper8GpL/eg9ibhPO5WQkzz5ewwBawIE5sOMKRONnovwGmaAauNcooxTWsycdd8
YNXDkhYph1m9S9KHxNQ2iZvCu7Y6s0ceTmG807m3nXlASUdgypQMZqcQe7iX4f+qtwFwl7nOMcIe
SLfxv7CieKjmnxPw8SLQbBRcypOWNxMtdDsqxDw3XmhTtTtG6hpHlG617aGdgCf9M0AocwLO+E0k
A2Hz+IdbrWY5c6YSLZwTwN25OmzlMZ3gT9hesWoREaTIP1ErCb3WePv/owJLtGDD+78G0up2LiSv
ahtoQDIcU+7FkRawQP9mRyeIFieR63yXVSXAES2/TjKPPOv3WLUpOKkSqZfi73qQviFB2k/Z1U1q
ChHNB8H7K1cYXM3GpdkWs7RYr7G2ZGRmSuA5CNCfy7JDha1q5gXOjqIwT4hm9fnA8mytHF2UzSsj
XcQM1YMWW4vJxTOeH8Z53eIQuq6/HRcSGoj19ngfykgdPOyP8v8O+6MQ+KE/gc1QCebhq0QT5+el
9D83QwrhDAWZQ7Z/A6Y2H9MpZMSR0Lw4LvYKPLg7VDeVgr24+1SM+QVszj3MHIJ7YiCrg6171qJh
RP63HoekT6ltb3TgZOHPIIzV+t5awdJzfdivljJOYZYVlauXt07Qg4UbCvReNfGsnqk61yknPTOg
y+pz8vC8R1oY1wqn8N40V6tGbNvQ9On+ztI5WFWuw4Z7F6OJpwkabt2xpK9P9DPcg4/yshyzKgQ2
EoOpTjO4/Od+4Q7QwFYSsiyWNcaEImNuvw1CL5NzY447Bux8Uell/0rghGJUigKOu88+/7wOei1W
Xh6Q3udUxHWhC52uFzcjbSuuCoREl/UAiXjNCJ+HK91SEQDRfdQ5+pkBiAsG1pT15cX2/laxg8kc
FyEgaRR3XWBoiF8m68J0OztNPiOWncW+/YESCfqulEy1uiT+hXpQ6uXndwaOzYC0i5tCTCJcwHGP
iezXzVm0SAtbD7+H3i3btAMeD7QBoGxBcR7pnnVFYQPOu2TrUCyd59GqV/+WdH6Y7CiR/CL2YvQO
oVXlNuExb1uhCekGWRUAxSOfgM5WBEpuYDISwI/vgRTUyZA6JqjtJ/KZ+xqDV/sT1tPf7E1SnKwH
GqJ1RJKI59mwEixN8RgNzplx/EbRS3tLr9o6hBtOlHil1fk2kgtc8opdORjxFEhjZmnGnnBgMrlL
eR2zUnio3XuWHv9Bm74gqGdv6bgzHl4tZ8W7Jf3z1Vsqr6HmKAFqyLpa4hjZ+eU8W9wW8PngCvGo
xuJWvHwOopUO6BbZpmPBARYU3AxbqfI0e7EsciZI9M25MYsCTB4Bxn+CPmWPJB4/sUsuBF03rviJ
ZPr0YJF7IT6LO66ezj3vJ46vNu40D1f99o/Jc0/39uuooh5GymrhrvjBWwC0rsZO+ljZ84dQF+Kf
Fh1Hw7fReVGvoejYwi0iEnNq99dRtjL639mSsm8U1Mtba5EXKFLLMwldvtoI/9t3/grLBLuBboEb
V+Wi/Lsg32cR5+8gq+WBfR2/sZioLthlKXAkl5m1TMq61m56R3BMyErhhct6HFm3TRS7SLuoLL/w
T2ouSBni8asyfFboG21qn+CtrX9YhEKthmiwb+9Bq1MZtqxBDGKSQ8dLwENqJnL+M+TeNMffvskq
CCBZdGfESBBG5MFpusLC9utLGS5eXMi2PaP2UFum7KZbFiOdn7QbRp4xjp/ppGZ81wA2uXfanSO+
XxvWEgpOHhjJbRH7Myw0uf1KkessDeCVoWx1RctGsAyU2xt+0c9Hlb6ryh1TOWmgTuUfoyOdybFf
279ecwP2OI9sgzpfmKl52Clq7rD3QeWT/dm47q6JFbbL7ejsZiGE3aAkViOT9anbE3iM7v8LPPJD
41pIO0Q0QfatpKvOka2kt8H5/+R3FlyVxaD40syPe9lOYLn40xVe6IloxolpcFWX5IfrbSUUIAMM
F8eNg2W7CqSQy9HhoJBAMpeyL1ZYotQrzan0UXL9xDh495ctb9/4ol72PMjCYOEKEhgC26phdWqM
u0gBmWeOBKknMfoqmvy8z+2T74XLWVJx0cpFTvWL7utvmfvoCNrDdEL9NZWItkk2ZdUnsXgCxsEN
Nk7Bngq1HJw4YwyCQO2cHsS4KaEf+MQ788j1CcJyo5GXgpgLYoYwrAq+MUV6/tPJr02gqfuHL9Bh
1Zz/K1UpEyWNzmig/mYS1fKdYTnfas1XRbkgrQmNHfdgJZbrbmDGy5q9Q+aTAzRBxxMOtuMo9lv3
Jiz6akctVBD4mgrRIbn1cxWrwQYD6MKeD0LvNhdssrSEVojoUtdOBTFFSkTuRPMQMKSCo6lAjHMV
garrXWLPlxUUNDge7+eeAZ4pbdFGVQ5zBW77nmRRT2HBxaY70PUiAbacsCWvW9Q7nxRnt9vZrQvJ
zam0oCXSXV/1D+D01QG9VMr8AK9tZBoqSB+yxLl70o/gRS8uQ1Gdl+Lox4IXcvppxC+OIFIWLHES
WGiiqhRuwSPFr4uf+CwRHMgWKgiN2C1W1JcR3qgx2b3opUyFC2tkF8p57xumFkIm0zgLPHBQ5MEk
H/wDc90oe+NH4GHwUpUT7FvrOymgMEWxSVivUATTKkNKEFTFVDs+XsLhKAOUeCOnhRjXzBUgksKV
eDD6wBresF4aD4kDjlF/mIym+Ni1yKnIRgdgl4UWCbgABW9C4aSoPLkYi8Sk47BS43iIsV/UUmYI
RSsLGQaeFo/nFGF0hC4IGMNt9NSgwrTHis+BXBE92pX2lph62bWzmYj17Jc8Zg88AXWjiZ3fml/B
uJwWR83JCdt/+rWoSijlQjk8kR2qV0+W49HBuhKfcryHb3vzQ6csTEbqg0Vlhlw9nH7QBeM92CfQ
U5UX9Om2GW3OzDURTXNgRGtskripOVyitrRNg7OTOsxaTz6BZsb8syrS5Fhm270MYc7Ps9QtCTff
ZZUOFnZ61Ra2Mrl1gUap2mi2X0RfNW05ZdEepsHtN0d+S334Il7KbKaq/suIlbIOYZ7wRN394Dug
WN2i4WRMT1Ey2H5yiRgmq8tDAYNeKnGuhvpX/J5XtFz1bIgXj3BNkFUi37rZvv5dKpEQuE8HlXrP
rsUDEnn/a2/jrKUFRhZZRBsT6vQy7hWST/taVC8k43lQW3FlNsMq+QdUrJZQbxLDjs0GV7nlWli+
S+xf1KIrOfoKtKU82RBaTyyTyGb6QyyzNy54NiCBl/j7xPZr6bbNilOKEv/E2S0yKQNSAsKbUl2l
Zx/znhVFM7tGFle3E+Xu6ApaZXMSn4cyAFUFNRXCMVZzNrgJk3jTDy7DTCzQo2/h+l1iFjaTrtlK
728CffhWhegC45icasgRCpnV3DR2EQC7Skh1Gt1VjcyaqCQYzgnhORcja0Cmy2ineK86DSdbR6x2
jN8H3vOOdbfRH2Lv2KpWvQOEePTvRjqGubRiDFaNuC9BQfTvUm25nBlE7aIe3K6+XCW7Eiu2Uphj
JlqOdIJ2Pko3cMA/XXLzuOmr0hf5oG+dMSZIu0z5fKIYyz5nfmxNmwGkEJJCubzgr3gbXPOA9o/a
5aw3OU6BBJWpCn8tAsvdFWAestfAK/FFLUQv2ilqzDI9pHyNfs0+GOawhzbicihenqDOtd/LY2qZ
V9Iy89cuDsArSjqpf/sAXkbW0x3AFT5fdqj2KWcXlrZFxV7wJCC3g5rz7w5r+c4LN6hjOmNYEoc0
9CBwlFMKClHKaY1UVVcLFgsQOLtKLA+fLXzmyt9/r/euGOB6h+1v5Ai/5HFBSH6WuqO5jnffU8+t
EKm1mFN1dh1Bg3uVe8q3NFWMpv0RlLNvvmfGL/3wq3aeGxb6cAiGHdFbPK3SH9zB/3paV+SANOvg
NA7JQdZyhHsvIqtX/DPEC6f9L/9xOBSxzFPhWPHpkabVBgrFeLSryPERJjR9T+NsvDyO1hDC1TkE
jft7PnWbkDd76hs7aRbDjTnwhU4fyPiFfTs/2EcxUBYO6wp/ILo2uDgWmUDvdOfTw1Uj2dBWmr3e
wHwcf8FTJut3m56S3b+DZ2k/yUz9noxKAfG8Urhw0iGRvPbhX2ML27oG5BBckcm8/yP5JoGBPZLD
8R5Idi44579Ni84SHlCbz93aZ5r8ZoI3jTpYvfqc1+aZGPkFRk6/GCUqkoeJWEmtZbo6voWU+o+m
oQOAFSe1ZHIIalAroZTPzCqRAzqDWqNzu5Xz9e1jNwyGi3TMhIAz/VL/UIISXRZ841CkGzua4kuo
WQ2cqEFq+HjABoTM868OJECU3xj+TgfBXPZVb2eeoixBTUakeVaqQLi967J9nTysopm8YnX/VdlW
cxZW+3MAUFWQoVAhi434niI+CkGOf0+byiigvJbntnqFb3g3jWgc74yOIpaBVLhe8ZLRl9fy5/wc
YafMvyEEQLdhPYEIVufY7z8BL/cFsgp4QYHEHA8gqPGMa/98LK8w2jf662w3ibuuAC0Ko0HfzCG1
dl5qg1ztbAVMjqPNC5zmyflUzj3YnlhPrger545zU1HPpk62a0hFjWwZ3sLzNjXe3aRaYQiMVDJa
ZSRAunQiMHahLqNZ2/480h6w6F7odLxXhSxQr55jMXCuuBMtKa/95CuOvsglCbrlOk4j/mYLatB5
tYyGsjuEzgxj1bunWWiU8rBRIB79vnJ6YCVCMDSE1pxTPJU8FO+39sUqrcFOxZNRAPJ1znYpih0Y
ApSejmjP4oLmgttZhd2mM8qukO3eUfh6u2JgP0DrUToGZ5eUsxy4D8A9a/+99CVdDzGbBB9UowrD
A7CmZ5CpbMuasy1duwTPq8kShkJdUHquAWyXbOH+6mCZNfROqTmqxNI//iLDn9T++g4hMsos0rYM
SvYa+QejcpPNzWSKtShSWqEuV3kXOgRkFeUsuwc8Jasa3FFZEKA6rtjdQrXMoDlW3tTSsOuY+75I
Ny4LDy1W+g367g3wl8I6eQEZVQKkqQYshtkeOXiQxbZpfkIwxI/qc0GKwuKjZ16GBmc2EeKKgPE/
esYefyedfeVbDHV9wyQAhQDebHCzXYEIlybh/nNOi2gq+tnHdb4uow5aQXuv+aBj+sGp9eeEi+Ci
q7PCrLdCiAQEGa/Sde38ious7stPOhwf+xtjva3Y369bpj3zvKtEOrwpdS4pZWt/nsS2Ag3ufbRr
W5IceWGTM9NgB469K9nPneDl6W7D8m36343BSiq8szDtIdINIufVdZf6vLDWgBxdOLAeSf26m3vv
tYBFWgPgYnL7DsD+Xd7DnaGM+fT6IdnWHG+KsFGDGvjTC7Hby5VVPQpaciKLm6p1Zb18Olln5F4F
B7PRW4OXQQM1EuoDyEhnbopOe1HcEeZkPLoL+ddi74odmqV4n6aQJbnNuvBgYn6lqBvs+OzoSQR4
K9V7oPmcCEvJSQacYQuwY7TO9bRvJIcZ5eGJyPUuBGTU8KPOIDalbrgwBjqsRYbvoDcExA6Enw87
wCbGPprvg+FHwv/hiynRI3hwWoGaT3bvH3VfJqMceSwhtiOJVXcGhGTBcForfFxqhK6SgPVPHC7r
OEbd1hSUX4Xr3gv4+rKZaxmtDOxVrXwvBMQV4ZMHwplgf92g2ndaFjp+MMfoE2pfnXwlM/VT3PvG
xkhC/c0U9ZnbYClgwCW2PqREKDnOjao6uaUNOHihw9eCnbBL7328ntLlQwf1aJ5saN6Gr6bvNLrG
OfTWTOAjKUFpkuR0IUicT1Nxt4PoKaQskuYC+b/jrmHYYF/kijMv6lvSI2PdwMonboPQbIkKJwiU
3F+hEBTlnqjF9G/G2gvvFI+sTmsXCAPcloyiQ83ENePzfgFbPP1+wYNkTVLZWzc4YdeRxpNFKEEh
BckE4Sn9Wa38Q6sNgSKLGOGdJASlbIUnXojYPbfBaTbmajAXZ3TnRgk7reSacAcrvAz34pMum4XG
qGpb/FnGMnNCCUs5vQD+06+YxFyJDUq6iJLsqsZUd/RDtB9psD/4UkSk9b1ESuH3kq9XrEZLNnor
0hkaggg5MeA1XXCDfFXFju1g0+NiNaTlbkjMcUWGv0pxDt1HZwfZ5wjBC55Fhh7TJozP6xhoKnqR
OBkLDncAlvGvq6kJV6VAmhHqnyrVhJhCIXuqJv9ZNujWZqNVUMG6YbmI2fqWtZwLb6byV1MZolRC
FTYsAF/Y2JMR8fNUoenOYHPFfrAv7xG1Z2KAgH/K4Q9pz1iEVtdc3JqlC094yhdT9n/j9WG0KXDh
cbxnbtHBjzNM7nxbilxIUlkElEWCrWefhEa6tXsxMASwppst/50dbz6/Z9PW7FWg0HfK7x6fr5Ny
HY3KFCnzyi6P1QxYmRyhyU7JIz8m0PauwPiMx943FTdZNC+pExxuh6JW9aDxWbBEnM+My0YdtM3d
CWpL5Oloei9evBqZ2sHuWJncEt0IB3eUHyyYwPARcctfJ2FMASLEpoZrCddaA7SR2xtyVvoJ7xev
kHXSzExhDgOjxNIrzEC1V84rSx7XROfz1Tkg5g+eWs2lxPn51Xg7NVi6u63ynOVFpgeY7pilguPb
JXviVfW0nynXBjkwfCiR8kirpcqcJV4TMKVvvxYqL+vfku2C9rlEQhzcc1HurqaY/WH79jT8tX1o
pXjEd2tNrqsFoG/EG2UdUkr9PKaWI9T9Q+qp8373dH4vX8SKoygcnC2X+ZPue6WvrBkS05mPpJcy
KJtnKRFxD1AbzBjrA9ee3H4xJ3hGQ+gpEQZSTY5iK0djh6Fagi1jE6kjlzfNTEq5UIvefPuyooQk
7zxgguh6FED6hmmG8kWH/h9e3UURQnYqwvVS22+2Bnyd+Qc6IBawyvP/By8oIH7/vdMlgLWIFnAg
Hf4cWMRDT5R/HlxvS6FoxAi+0n81Z1usNooyQ9qbhMy0FVVgeH49BoK7NWJwZMxBTL+4a4uFvD5c
g9LikWWVyqhirmF7DkwD1H2HJqvYm2Zrz7UlfNMzCd8hFZxMzPGpdoeyKMZa5PWm1VuhuVAWFwNK
cSNFXtSDBDx3Qzp5Q2s+IUjG/9HmUBLIYIFz+3hXShfs9w1nCtOzBbcquPI3G9URc+srvFF5guFm
C4aO2tdFVxvCqWvbYoLGmo23dZcI1pQBOkKztrOT3HiBXy5SzJZJrgPQ5CAqebwGbYlR3kqbZcAv
ozO3zRE+7wmvsW0ZQOSPaat9Dknwc5cKcIdRMq7VHquJZyjYre+5uIrU8nIQxzaX7/aI3OwqyZbl
b4q0mLxa4XzhEQRg1R6+LKZWK6edN1PGimecn0QI8wtPWlURw3ngTqle+2YqsUjGCz7Hg00CWnjt
adPwkn1TNBwXRuUww3CT0+4SWx4XlxH0D4mqn7sW3N7wQT/HrMEbD94VOfMTba0gWE9QV4REIgqG
JZ8dtHsC2FjUUfPjadQtmCBkqpLIZmz1Vhm6X8H6i4sB+8p7zmbUqayV82K6qUkZzMKApZc6AJUK
PK5DlNCeFa6qGggEBxMIdrkFQjMSoIlrPrjJrcND6TDGQCvgDmd6PLLtCZNLDdNE5egZWyTZ/AWD
21PmFzzGjVpIBp6zb3sArcF8DRdqRwioYzK86Zg2PR1Xv8VBfGwjjiASe1GYyi6s7eORV6955mGU
f/2H01PRAvYriq1fIzn08WzzGYzjQlc0tMvxJMytRbBIW7ujxB6biEXEtD/viXiLKIfibidszHWm
aELGwZbHidObBbgGT68Vnj5wBxrBilGeAegLM9foEDF6MRPaCNgRSxzoBaIF7wpp5WlpjQbx2RHH
G/07BvBjwqt0hmLk/1IYHJnmS2MKRdTOeObT+fpnFdXMjnVFyYBvEeNTH6qIYjnyC800pcmr73if
WZROtkXvs4dZixIObhE3OtKEizeVQIOeeTkiB3KVzLrdBM1Mc9+f7RvqjRtpERak/evDcCMwVF2+
yb/TssOptqP/s8uGiACxyFrE72TnWj34v0KLmfwhCZMMqoGeXZeAagHSMKOs2mGQC+2Mf8+O1sp2
BK6iUo9b8thqSbi4cl1lxVtEtMBKtBYlsU9xZdf3o5mt4Ct+9v32dWtXuZ4p+o5vfcTKWiFSbttu
c4d/lLxx5a//3fHCx5HInBZxnBGxHI+xxs5KDzRot2/3UzjktkrGxdt+GfAqL4UKQkmpH8n5J/2A
qByOepZfydYRgjJx4K3O39YllAws6sRYgX5nf/f8Ix3mP/5Dm1evcKykrH+G48ZAiR9zuSjF3w1c
T1k37NYC/5kuXrl+3y9YeE7vCKXMe5/XUStA2ZUni0PhYCeWCiLUkgNX4yOqxA/Dk3t50bt6jdG9
S8JzOkvYL+EIrH8r6Yvr9qfyPTteDA28ZmlILIJLcCO++o+5PP4QOPCPN234eiWbx0l9/D7sBTwj
/DMvrBI7sVH13Mam882t69vt3d7RVahdMvCG/tf3MwyKwL7kB6JLz0q5aafyMgMAtGfTUYzgjxbK
s6gxvURuUG/+0uldEBdWgSbGnUmt6MQ5HGKkZZ83uG/uVpCoWJf4VaX5lxrfV0WTn3BnnY2mmGf8
sTIiZixY9LPlSuV0mKQQM3NeBLEvvxJ5D8FTvFkORShJaZw/6+x2zkBaC5ecEk6Z1PxKyL8hsT+l
fY55uqvbm3a9ywsXi8Rrtt5AzoYxzp2x6w8LJKrvboEuwO37ezW86JjM0d3h2qO7y9NH+8/V0ysM
A4jWWMt7KcyXMxuWoe+WXfYmhdk5ejhAyAGKhjySYw5RQ5x5W++MjqBQPRuKBpvPhNeGvG7jz+AL
b2NrdDrz4ISs8HcZgMFbpk+bfDynd5Br8bLLmwhqlWGYZCBYJaukvnzEStu+hh3IDEhxGOsMxgWE
tGAw26H2aozekhvqwFcUxPxdTngsMDpqLs2ik5VZDc6qgSwwwx4fLs2/KBUVoCrGi8P8KKsTzY32
P3UwPJmsfHIVeINJF6B1fh5GOXR9+/6k8r5dlS/UHRJ9B9CIPue3U1To5Q1wRH1JX7ESSYfMF1gz
Hb7duHWCTCWzIxZKQQQF0Z4X2pUZ6auflCJH2ETlb8NQ1TLQ6Ty1mH9EpLbzRVlDBd8HYIuF2Qaq
C1SUYtB94tg7mL3gh06QB81dxe839GMa8ryJAq/ro2tmS3cjur5ooFJ7r9gvA6tXRxeghyWo4jGs
5EWPhD8b9Ijxpcmr5zaezf7jZ5zNkE27BYC5QR3oVfczKamQtGdHVQVeCs5lF0cMdZLD5u/2Hs01
OZAbhDQv9hdskrBW+f3NGAcxpe/1wc08a7Pq8rYR8/sKj/EQT9UI3EOIoLceqtkrGTVZH8wfdsT8
anlc10NzTVBgID4aChfiLO6TGPB1c2qYlAsAABXOq6ltkm+PbjMvq9TjZqJzDnTVkaKVG90CGj8U
5SM41JfGFkM7kSHWlmVRg0BQ4996nY6jblZv3Q3lcDxhreG+y10iVlNtHuVX8lJEojSSZwwlfuoH
JNXbWUGKG37jbZov6kbjahiRpRN+CKpXxzupgEvXODyqKsm77RWI53MOpb42oBwAAtFskRPjDF/l
Pkmz7pc839daJq/yWE03L1kiU2JI5fIzvLAk0kqHdn/jGxn3dZ/ukneHaDKhqMaAYQ1Tkv+quixE
SU1aQiPf0oy0xcefa8NdeH//BxSGDSE3AoHAz6qIARBH+OCldbDd+31KmSMtHU4/ctFooSIVNkI4
NnzEZP6RM8UMItNCbTakqKmJqlfFUGMQhvop+GDbHJb0nuqPUUUg4X1v3SHX7iu1Y+GkOWuh51sf
cX28TiA3u3Khi83zUe4OpumFIvVz06OthmCrK+JQNYEhX+5gd6o6xpPtSVnZyo1Pq5DXJhbvQRNF
LDNJLDt8ECH/dt92fegkIDqOe31gZf8LxuXoQvx1yJcGhF73b+9XZaZaVaq1NFJjGL/5u5A8h2KZ
7IFE386Wwk5Nnou35zihtETQwO54XsmprFumN5qfebIvXUyGwRzO8ByaEjOrmveMRZZsNmc7c7IM
1merNm8M+eCqDVyVS8IqQDFC4QhuDHpSdc/ohAQ2n78AbUj285puIVM/V/7xUAjDrEw8+yMLQlr5
63U7y0UmVAO0VXe33/Advla+Uy/JytFlmT6VRfXR7qBRNeBLPyuqg/04fFl7plseKiXlP0wdlRxo
QpX3hio+hdDFeATKuGu2le9DyMIuc6EdPZ8dgMoBkytgettITlVXx/jHh1zvevxSoWO7NlxbUdEJ
01r75TkST7ovWIfz/j3Ko7D/xg90l75UZGC7waHXdwvrsHEU9W8RVvAta3R1nzih4z2pnfUx6Zja
svYFGKRERgQm5JJj+ntUbMbcyiUloeob9xSLnbargJ+Tk8D6ZRU7RKGx8clRjgXKoPzOmwziH4vD
zKVJqyZE25iPybUdSleT8zVKfVG70ll2QG3l3lLfOkNMQ9qaYZFFJzp6QrUtwHoNDDRLSi6x6PEf
w8xLF2SxHVhUAB2nsqImLheBJv6kZX6UYkW6AvrFcBxNf7AGuXxr1mS3Z4aFsad1j9kUzvuJc601
zyKWuXJUeN8UULAYqN/X4EE9WUP84mriECb3XEx9/A467uFempB6qYqUPwsaVLpB+8hm0MQl62Mu
/K7vvHznQOM8HFe1da0VwllwWAR5lXT9bFiXVL4GL59rAspj5PS7+mMLthWqGZYXdRLckEbjb7YY
DKJzVp+P6liUXxvfsDKfFX2wkZvQ+wMKs4eeGvQot/UpsuZaC2jOMk0j0uB5BopcdIpaCdmrwu8W
jS1e2LM10FgtBdgKBZTely6G1ki0Iua1LY5S+WEo4/zif7r3/UoImtZRHEy5aKdufDFODMF96EIa
jnSqsDdKZF2CAkrkFsVzWPKoihtzEOwbF1ciCPh8lHzNtRBQr38AXX+DF05sMsK7A1WJV/qNq0Gf
FANf+kMiIgZAauD1VyTaWr1JQqzi0ghK3uITyRqWWK5EWNWETYWgrhg5rh8uI2I+H5Seh7sOG4dr
aOJim8CV/FBeAQnfuaGqS3flJWM4vv1F/cK/kraX+i8g4+OPbQKbDkN2D8vQNHaHKoE3ZnSOXgTC
YLjbRTNzt2dSlfxXYNsh/ONCLxBZOfy1I83B834y+Wd7TOy5HRjD4rRP3nXkOOS/x/MyksQf5E0Y
2H8jV2eKXgV4DVnDX+DesCenyEh6oE9sd8Xf8Y8KQk5vJOg734ypzj7NEBBl2qnRuKv6m3z9W6Ao
8kTMl8PxAaiGZL8F84eDiOES6gPqtZTFAaWZYg6Onhd3xD2Vn/AwdZ7/KQcUZ5Qo7wJ7/W8GIJSa
M1f5BVXvrpYsoQlYqmmvJfh5N44ux6l7zXZAPg0c4j6Q583vpZnrwkF2A8Je0LOKMEwgbKUjcSWx
IX9eKtBeoU47WXC9zTOw4PNuRZ+Q87DyYTe6VC7hagFxcZ3/ctknZgMAXak5MBKgFpBVdHmhYtEu
ZOIWcI4yUcJlWXqc+p0KKM/daYKs8qP3Ylen/QoouxG7lJkilGqM4+9wHAqWxvbMUR6eUGHeBGUr
pIrVX3UEyrHC7Z3eOpcTlTtelUbUwxcQgHCoLRS9Pxb2qDCZnxcbW8xV7H4g99U9jBi+92MRk3Oq
LeHcMuo/tA7w2PV2L5HWKaIv44QU5T+C0xrDrS9xCofMoM/Q9HPaEpFekC445R+l5Y0BDzZubh5t
zRZ0qq2ylnrlowSBbO0y8AVDs+cgDolmyRaP4JklPr6DZhCG1ZachDkhvFofpWjO1TRZwYm3AlME
sqZCp1vK1HnPJ8W5jR3QvH4FjKbh42ujQ4fEHhqUY1z7m1cf1Jv+vzkQwgJTDuykUHX0Zigxn+I/
f3AtSA5pjF8z/TV2dov+E8RAWl8I9YCbR1xmJQ0uuJxTLhzuKycc1dMxgSP0PYXvUyzyjI694dj4
vu/9wl7Kcg3dbD8MEP3XKWRmYYKfwvRJPgbI8xD4u454BD9kGQRXp+6o+k0xm+HdLRnT6EiJiqpr
Q26HGZtuEdLaw6ZeVIB0xqzZp/cd25Q3/5XIdhgvidkRVR8peB7K1QFBnhG1FW2Wtzl0H5Jr8PaF
UC9GmGl7u04/InmABJ42lBSO11RRrNHvomZJsZlr7UpvgshVqUFzzdKyoj4uoYE3ilCm1Bftz7Xa
rsIGydrgnxDBALZW0UdF8o1xJ+x8KY2lEP+jC6YYnafNX73xdos28efKVbpqV4ovjPH4dCVqsOZT
indE5bFS1RIMXR9mHb6FED/fN2kvyek7yu7chLCzHdLHYJgRqvDSvQx9g2dRyJWrxM/MohO69/kX
5yfCd+SmReIJ/sEtJSvYrX+g5w64cVho0iCnWKJzFX8JJm8cfh3f1wI8Dl0GXEJwOB1eCPIovgiJ
vLSBeZckVjzOdMvXrpjqjvcBDYRGV5U+s3xwClzkSIltu0JslnDdFubqxi+Mx4n4Ah0UvwHDoNxT
C1hARlbrzRCczhj2FsOK018yz/b5SLnYyaC5gYijsgt5fpE8QcZGddf6yxH1s58SHEsbncEJJqNH
SA9SH0onnNjuvK6ICE4e8JgMkOHFW0RUG4KoYwwNcclJw7ZTDI5fmBTj4B4vH0xvYJUj5ChFqxIE
ZkFlpPAMRffF5/HKSuNjlDJeHKXdf16PNO6OWlev6ok5+O7DVsIJ+ZpeaIvWlwVAtrIhJGLqXaRe
8EI3GSYlbF5ZPUHWTw2qOyPoiQzxuoseqWeTqiXsZcxGJBTDQp+X6UOvlF+TfJMrTZ4A1smK9FxR
HnlWKzQ2S+y/Eza48Bm7MyYcp62Rslgjcw6JbsbVIRSRR4aPqlILnUYnGhgLeGvI+DBFVk1Ufc5+
PjuIh1tsyAQG8YgkZ2hXAliV4H7D0EQ/v/AqqXBero29Hy6zQ/vhZLWLkkD3hPX34+aGRUwGhK6J
t2nTQzzc565AeP/wL4hHUESjYcGX4hVNBNU9Imx/Bs+LOwYoCnXr3trzmuf5IYCptFcFX3naHX5E
aZTzQdQwjZ1L6SNEmz6796X5ypyH28JcCMNDrFZ9nXFx/sQmrpqwuEvhUCGtX2TMfIiT/VeVAeAV
+amgvt/+poiw/vbur5jhmzHz3tRlzBEnZNKIVGYC1f7iKEWgUQ+zWUrXnDylNChm2Vf4J2NAZbCE
3EH0uVndnlXtN2dv4+jUQKtwKddE91Eez2bdHQwjPHP7e8xS6l+C0ox01WDcVOZkFHaxrA7lTUxH
miiV0K+FefEzybZHy7llduD8Ej/H8lHpFtxPAeu8n2vg03TL1AGaLjmooWZHeOeH/3AcYsDH6A3x
WvCXoimFvthp7anYMkrGtwhb9ImMEOK7Vr2xhNc9GCGxG+WTAFtsN06LQvq1Ifh8lzLz6lrIo0Ub
ewrrERsQrgxobi2Nxaycyisxijfd6gYPFS078yKq68RounnRiW1BKr1eddLgt9SEXrBEnanAH3YC
avU3QPjejkC+zCGxXJWfJDciRL0OLMq5/fR5wuUg2ija+4TU4+RQl63ROZqPaha9TAwS/1nCVDqS
lXAr4yRbUSUHl3YnBmoh62/uUV/QUobA3KZvxH5muYRmP8DOQTCpWRYjV3N077qq1boykUlGRjvm
0MprYla+K3JmPsOnJeOZgwSI3Y5WQgYy6zQLl45bDII2SChs109bJUvxUUQAYgPs4PB+1FwvyrMt
ielQRsC5yWUtIz/5lBpO2BrDvfG7Nai4RSx6cusWqgFhDv0iWvSoTfNEkp9zi9mO3moGHr5LBtYN
RJJjX89MGe73Xn7bsU41YiGnRVlAISt9Fp6u7eXogEhOSAnlaGNfkNMd2wAIyqukrKHjgiJTSxHB
4Qob81e9IS6ZGIzm6C8B2/eRywayS4CePcAtSEIwuI4ompeFq7wC3ewa0soya1jiSOXGCrEyH8BY
y83gq3uvikNvycMWTk9fzU0TAs8WAm2cgzblQvqMxt6ob73lG2dwzO/m7t7NyrZnSGHxbiD/qUHd
T8l82bIwH7jXNTAbEiMjBxMl7JTHctVQdu753Z88qt7SgjCLNMnEdHYRRD8GOjDAuP2dBdPpQRDJ
5XRO4/gvgSD+Ym4e2kloZ7y4iNZ8CRZ+iTGaHwhf5Bmdk5NFdr1Y0ti3d6cVBy5CUc5y+cCJauqF
JCeiMgji3QgbE95CXGWJpc3POk8T8F49s+MGR9FaHhEp7E+FP6zlAIX8xinu7Sowceut4QImMsiy
JbfxULFr4mHwscJ49bKfV/NQwSamvs9bU2ENxmQaJQ8DE9TN/GB3pPCUYefjScFg6MTCmlkjkxSf
3zw4Xyz0RzQTsDk4GiLyTiAWbT1rBWujDlNofmI/spAcStpAVzRztpuVHhjShAS13CwM4Si8esNm
64X+9STPOqDtCQLwFJHL6hTS7B1i3wRCMnzBZC7O4685lbSnCSkq1chpvPyh5qe4urvtrir1KFAL
4z7pA0GfV3TlLJIJG0xgwRHlUfY2v44ZiAOTX7/HKaHpxSJoxD+RaQQ75w47mCxGeLq18owUMx3s
Z9ORgjCo9RfZnlVm57H672khr/lllkg+Opj0WPU+epp4PtsTzRN99hC9nqKWtL3oX2ToHnQWzMir
7ryS3hU7XqpRyAVoJrOXey0mnp9uA1c4M2FJyrX59xeqaR20rZPSMrcHfaTD+izcubnEjPxECl98
2CrC4/+yNzbyJvvtSSZS0EbsNu7rQA0wor3uRhAe2Q54hD2rDmmGnkHExTijQo8u4FJP/t7A8a0h
2BPSl7hhwS4qHf0Z2aBc9TNB4RzsN+IVBWfOTxWYlvZLK3q8yj0V0AVw7GmcjMx0Oj8oOifkCPCq
vdrh4mXDg84/UHs/QRIf6t138nuGXpaIg4LsV7S7W7MM/vEEz2GgMX3dSFYxmwQdmcrJIBKQglhq
ZtH3fo3VynfclkvERFb02YFQx0sVu1qlSM1maitw7gI/g96jKmGmAKJZd9BWME7C2v1yE2x8phSc
t81Ry8wxaX4Znsxcq5uB3iC0oQlnEiGkaXJBRYf96ke/FaMwpfGWFJk0XumCZlJey9rDECj/TbBR
OgYl1pw20ax39L6AS7N0HgRFJVsUxxUklncnVk/jVxSvtUPQ4r5+X5RmjaP+plFIDRNGv6wYi28T
yiutwJKYJySGSEFN9p91y/fS/rAEO8Y8gwggV3bQLMQsA6Bwyj7Iwk0Xt3mMJ6iGWrzoMgEH3dHZ
4Ou/dItjgdzRSGtRdNEIF9SChVF3eR9YaRBZUKnpEjOIB2/S1lDudb3rKeDjIPCILcK3CIUeUkx+
kowWea+adctOq/1unXDqn8AZRkLYyQa2REy1rxW8cqUWHGT6HEdxu8DfOXTISenWUbv0qe6Frqbu
9yBBMJyaJj01dU/WdMuO+Vx6cJvNz+XmnJu5nmzBuZ3ajpPhhqDpZzda3WhRiDZGKAQ5vLDk+fNY
b/1gtAJEg9UAEQIw9A5/wpnIrv4SPtqmObNtmyRc7GZDiYsRFTH48M0lQb81jocpWEyESlGqPUxB
WddZMndnWnVGobNeYYOlvx7/hh2GKRtgvpPjhqp9dIMxL+pZz5Te4TBdj2SUPb7dx4vlJoZq6ToW
iRnDrUIq3d+xiGDHC45DBR80yLItK1u9k9Q4otQn5XO3Lo5sy04uVkUrqFjbuXEE3H40YWGfiQ0q
+tmO+RNwcy0QbNC/34cyocCRPSo2ZrmL6l0M+owMjHDoCR+Lk7A9lByha7Yd5XYzXnQa7ZS7mmBc
ipb0cMcJFD5/aw4bQI+pqKWQ0vhFDsRA8glb136coXKiYyhQYDDoxPVZgtVY+/TiMmo244bw35XY
eDbnydV4UUfzYnRBvWB61ZFXJPFsfQ487Q9nimmlwZya7xU3vB/8jfCu0xI1IIlL/g9TRNejFxmp
1Ie7b5alPMB/JOurE7eOKmQy2OrV4oZn04EuKrImMgyW9uR2Yv0N1ob5TVqVjznxmYbF9o1OjGj+
PNfknP72V5UpoZb581f2vbr+KzgRg4s8o59B20zVJSkEeP4OK8HV0qDL9NL+9jXT83JafHZrXxMK
v04uBBKXr9DRqDLet+ipyEE/98uXIPCkwS8+b/VWVFBESmyzGc9gDhXeOXLIOKCxQ0Syu9rNw78X
NONZ0BBaqzIqtfhzmixw4aMQi4gMOM1hIE/vRZsWkPQ10w6Bk5Y1+k+6a1GaU2AP4IywrQvNQvq4
w60Pel38zmUES7pn4oGkaMsByVkhAaXpFlct6SVBklGoRX75KOg1VKizcG8soaeMOzH/w53R4l4a
pqs9P13JcX3BzwCol+INoA0CeHi0z4NqBHRYChcbH2KPDB/LwcCLMJ/DRxsdwL7YSZZVfXZBITOF
1/877vHMOcShd5SXpmCFD8kLDsdOXkBi4okygaopUnuC/OYDJQWCLMhwxmErYQFvne1YslI0vqt7
ijSg+XbUckU+xh9xfkJd/AcXrcFiz6ctF4S8wrt6zm44ZRmwTbQWjTzEXIWX225HsNUaox3MUt4Q
zRzsZs/WoEwJ3YHWmY9gvzXW/Fhj2YdGiCWn3U3nSItOT/b6RynDHezoQxou31rdwkTaiRyurppX
vg9DLAOqMKwQVCrk7RofUdLQ+3xrE2cgXpBD9DG/d+YC7ND4uT+8JWejnCDYgmGojbDuFcVf54eQ
YatnaB4ZBs0nAYqRzFWkQkpdQzoUydcB3vE+2xD0phFSx4xYLceksRbfSQd7BJsKjVhIU7t6X4Zq
n3DuEyT63uK/iAaivyn5MkOtvPlr+L9WX3pdYC8pM+yuGUoAVc38eNTDykr0gz60k9Dki+Ff/DEY
dUVIcS13L9rCqs9u6GsfhXbknk+AwjECFsFQIYx+Uc4YyUnYNBiPkGwjKLtgSz9o2+bBXZ6oKjdu
Zo9H9c17KTJSgSTOJVY3yKblUUKuXpumm1dAIk1PJtfwm7X7g3LgITeBJI/J+we6fZMYJrUicJkZ
MLH5lDzGUOzlLsNbjNvO+aIMW25TOC/TXs+2ItJwi1mHNbqbNBwsFw0cNQdx8QTDeXcGEzKQL6Yh
UteZTs78tO7zCzZPh8BpYJmEFn4aB0Oo1Pzl/gSxp3tAmsaPco0xXLt3kw8KjNgiXF6O8A/2Px5h
NIXRW/EDHfRQpFtpPuX1kZz6Oatape5rFGOlhoSWlBlDcKby+3V9oW2E0j35o7RpayMTQT5fA0Pi
I26s9HkUZSvy3dIFInT9xe6qHvFnsF45y2ETHd6lHgITOqg8XA/Mcg2GGzFt+Igm3qes94TgScBQ
pZ7RYkQQLh9zCVo/k+rKbRPxhmZI8LCU0v1njQZD6GQm05HR9gmUsBgWwiiK/IfPmwse9SB3b/2A
vuHSie0Ibm74lYGNRWqgBIt1MKgLtYY/X9aDwtiBP81Hx+qzMjVzNhxxHN4Y/eYpKM32+okxxGqJ
9Q74E3WPZZK4OlpttOWx1AZHoOk9bzHIKimCQvrWh8ahx9kwFupq0dQprAUTCJAGfaTJI+wKtsTj
o+W+aiF9dbJCDihJzc1zWW0SSlIxLw6S7CI/toIo95GHdFyeOhhsuNeJnbzZxyESYeQSO5ClyqND
ZnC8TWxjXw5+XKCU2yrvgLhe+ZFIvqlKGFasGPzPEbN3UDG55zY3CxHb2TxUzOr0sI11OFFUZT9D
Mv2lDA5jDtNZmhpQbhlhaYpkpXo2MuqOBKuTZ0ic++Y4r2eiadaWAF4NEz+db128mKW7Xlqlzygn
NCRGilFepJ9SpSHtF3Qn/Jph4oOTl3y+1CTrPTeKcSyfnOsenoG+us0A8wzBriIhFKHujKTLNpaR
kBV8oyKwpIAaAQ0821TDfQcoSkwfJ/yhho7P2M6ySmBayjv1hiGB6pW09HW5N68AJKNIRT+YaQVf
5fxodg63sOhuOKy03JaqTYhYZUf9O26nahs/IizHApYdGooC+v073IK+7HU+4BOb6lCBzRF/bxeK
R12YaTRPYtxUCJg0L4bwohAk/hUVWW8ifVU8fjD43hTScycOQxwOiNVpO7RWLJ9H9Wf2JVxH0qd5
omRAbN66l3yF+QpONfzIWBzW7pt6uf/3dg/lBklpfgjib2xQCzhXidlx7ktYmyMb2mk97aHGZkHy
tAmtAy7VnK/JgY31m3WCzKn+CAaSAkDFe2EPxn1LFtR6oSmM38jL+9wTygToZs/xD0SCtLxHNASX
iZ373bxW1rcpvlMdpHAHT88HpsBqY8CChEQJhQOy2U385cIl6ck6vuOINyl/ebgCbhuuhhVfWPe+
rhzt9Tu3Zg1ZxfRHpjxTHdaJyzTrcCM+rF0ztiT3jCCwjRvZoDKBYGUZpOwK2nwJiP1qG0STco96
+wqNi1jb0C2Db6NXP4+bltVsf9pjknLcJWrgLneY/quxAVlCqnDXuDdm7aAPwrONeTiq2q28u5Hf
+Y+qtU1tkah22x6zepa6wTKrN9IpftqpIO/n4+pfJYmIHNTYvZYgWcH4ql6ClkSTwqRBLM3bFfIs
DLY/t21J8aAVZR867An6OtYGbYmbh28VZBgyF/bRsBSbp2Z6kklrAGc//arQDxUXAuE7tWUjMTt+
ar43VthyVN5DUfDxivSTaK7A7aOC8+Zykwo6RmaPPYUYHmOzNqy5n3tSx2GXBPw6CmbiaAxOnz2N
IOdJ/o3gZBxjuyptrp+mfGwCObrpisELu1rHg/ZS7ijUMZuamevgbOiIHlf20tMQK84EcqrJCmqv
9smRVryvGj/8RcdK4Ql5BPNlqUE7XMvC58dI4o3r9lDWqydQGTNoOp+7EI5TgNEgY8iUnSPrkgLi
pDZOeJ0AmFS9qaJHb9sVUD8XvXUm0uTB7FGhduSdCivDwyW52ykNzzDt58TaRAnHnHkpb7gGuEGm
7uUxjxLRVSnzVcTS9MF7j1Egfbly2T31h9+I8ea8sWxXbv2oOvRDpTyE318wsQiOD7P457oC8Eqx
5CaIn0825njk5zalzUX9ZjSBP1k7jcGES+2erDxw/Yt1cyRnVbyg17S5RwXbKUUQXohZ9Kezv+/z
KZFtPziQ+TZTndsCSprUBpqgKJp9rjuouHJYPhwnrtL08juYItbaMSjImM7prwBD1C6FpQc/CZjO
/AmfLE41pXCnp8JineX9wxafwseF0Hec9b+G6i+mERhA29YHLVSoLaQZwEZXZ5oDmR4XbgHbiSnm
EeRHiTLhf/GQMyCxQM2c6Pp6xp7h/4Ixv/sa0o3TM/8P4icHVl/WvcPLp0VwwCTCAwipuNpDVQnV
OMxBS3YnXFQ68iHJmPkZ3mMT5olXCJu85ny/uzZGIWdAgUO2mkny5SLoWxhpc5mWUckkhIgmWy/D
rI9hXmTf1CfGtgGWJRNkltBV6moJk06RIa/XLdDeV4TdwO9LBnvuuuqoo9b4PLjqT1b0q2KWWtgT
IwXv7veRG+ex+P1KecsGFjELcO/4bWx5nDPPZlF2vCu+tUvn4hmmUILvGWZAkR+aGYD9EeYK5zz6
SrLSxJpi52C/F4YrRhg+Bu2P/cSNfJCtEDrW0I+VvgY4sIWJUurvH2i317PPP7J+2J6E9qeIMmgk
+86bvJJuYhqcAzsLxT7CKtSu3trNwYQSBcwqeusY5Gw6ZFCrb/eh3s8HCFDTDGZv3g/37Ldd8+CO
fzQfRpRE3nbiE8SHU/o+BshgrplPBAqnApV4H4GwSTK7gekQ1p/c8wrBAObEL60FNpHW0TiZ3LD7
C53OMVPkh2fEKwe/W+OqFmkLwxq9D1LU3PiZBfPyq3YF1MsT9c+F/QYDnqv2XaSFTQ2RPktiBNVK
+WsT+V24KwBG+z8jVs38aPivjuUgU+zskkKMNFVHujNmtDyUtRc9puzbY7kVPSnPmU42LNuLrb+p
7iNPP30LX6fsrFVgD5AzKqi6JP1X2uV1j1pa1lFanPqW/hdLyCH5S5MzJC6JjXxRdp+Wrq17xgh+
Rf5wSNFg4ptYLmvh8KsSPeFmp9lDznN3WL6OifLB7ep+4vyLTNgGW4sXDEJZD5aLLr+qpV3RvtEW
ZJIjtNQ0u9qI7MYMmYeRCAxXLX9ocuGydkk7PTyFPEAi+z42Z9/ppL2N6uEQ9gYHlwyHvVkMmbfs
8qx4HipimHX8yvarzvQoJiVfTMjp0scGrRSet3dD7QNrHlmSsB51CuFzsjA/xPuAMsj0KYjA9ZP8
6caT9Miw74yhZp+y6sHdFHSuNxnMTiUVyu3z9hdYRsv7yPwasNQLpeiMUmjpRZNzYCCR05fnMCFR
NyRTXHX1Tibf/C3PpOIZxXeOq8zWJcRo/BjRyZ3E6cz4ZYzcpj+5pK/v6PU9IN9Cgm00TE8Na9eT
rko4pVrI+yjd4DeQ+fHPayD4mws0xaWyOutIUXKf4wllu67+Fv8kGLgTR0h60oiruYToKTA4ypdX
fHiGB0ipyq9wXzjtcJbP1XYh7nfovRVSGCJpOybVkihUE6Yd1WfNQiS04e/PVRN2fuymy0CLV422
FlxZB5ngIgjmlA4Vnydw+vIKPs7Hz2/xRbiqx47p9RB728HyFkMahvkaw/h5UYXNQkp9sPN2tHIT
x+gRcmpbppKfatTXr5s68GmDPHNjKNUQBiFTZPSOorx66qnxTi6PF9CAP4xsgAq6uUDpvC6jwduJ
TGHByZ3aYfj+3mVvkzQ3LSjsyH0/iCQAyHW4DtT1eQ6947TVkHaC+89Z/JepAR40fucMwiNEadmJ
iH93aWwmwFG/ZiEtAU2OOOG8pS89Av4uCg5JTKlGmMPx3+vJptLBkPR7aPzBzev/g5gZVHfLUsfR
0yUjaIZ61EwEA9KVVW2PWqcoMG+5qFtsMOwGQQvPpTxZThsMvjd81vQY4b0oT5LY9JgpcjWETI1g
muSSclaCNUf2BJNxZMHp9m/zIjlZ5qPw2jptbyQFzis9Mzr176BjtKTrBJySjbnQ5QXfm07uMH/S
AqbzvLmHW1FW5gW8vAPpT/KdXyV17yxPxOhW2VyXJaStoXMZXUi/aoBCz7Xp+tZaSgIFA0DbzpbQ
kfyB54sr8Ff6Tmbg0/U/+Zjk4eRg8JHELTxKdcYjNHO6F/g7CIc91T+tyFeFTCWTmbX7pxqPFQK5
4sJoh7Zp/caHEG6wskfUJfnoDtLxkYHP1dNjJ5qVmueqQ98mhxzEvu5SMYA7LVM6n3Ha99xs4jX9
CIlpqsmGubCT2Lx7MB6prupaeJoZhrlvil6KA7Whk0JdNDylfRXP37liOV7s+8pT4c/ABnnkDOdi
CV3MaRC90DkyPlEytITFQCCguoVi8W0LMv7/sOiNdl1drY60qO0OVSxruOgWRo49s2ythSz4kWbq
pb2Ajx1V+liNQrACICLYETHUXd9HEMP5M4hIdkLRBdZhE7GoqahjdAVVR1lf1/DRvrOpX7aLcjUi
6W/Ii8DLfJ4WkA9ySHhmMcvhoNvuBrrHqkVIFEPa+w/1zZvbxm/MxymGDWzIBGf6TwVuG+Yon163
LqMYPmNp2AmqaMfpPGDO5uHV0TakXvUTn7z1OB46BXGKg/w4HyZPD2YJ7vffRj7BRxqoHqaX2e6x
dLDYc4WyQOZYGI4lnm7M3rS8poIPVU8Cpw+DoGsyhqNeFV4k7eDKSThrU4KtBgUyBeZE+2AmJbb/
CmftJAIai24SFzRRjO/ToGXCMIZ+0wWfadf8ag0YKclyedZAaPZj4f8Y2QbxJxWOcJzYwL/DP7xX
bwAHM5UPT73nBsSOYR1YVes5Z3U5r49mVNTtccg6PDqSi/dgxJ3HqRy067mrTv09YxhQaimxyXKI
x13nH/X3HIE93mR3GiPY6ANnep7g11jXEcjWFXBswuiNpnqOMq0B/knaPtbFiAoHzM/5Ap7sqzFS
iUVvNqCgzRU8dLe0UzYszxK65ShiytcziGrdx+paACiaOdFJKo0JtQ2bvNY3A8XMDDxEfBivM0na
0m+D9ShDENwbw47gPHVqPxuL1JnJccloi5AheOk7NtQpmp6UHFNltxrX6ESUZSw22lVVE6WviiEW
HO0KLFtMLCgMu1d80v9L3OwAgRq8J4RGYQuCx7QukqCrQ5FJSE32ZcfmOjPCpA9MB40AALqtFYOo
I3vHLwu370Uc0v3kn6RDPUcc1hC/AS0R8BiDW9iKwr6q6fawdHRhcEdpbzH6/3qVH+u2+o64bdU4
8YO0/ke+dsY8YWzFOpZlBcsSPiMXbxP2RTWa4lvfoKNH/mT0Zk+WG9urN1jUx88VxrcsdvNzeYwq
rA7Y5XT9CA8Qh3kpoiUbdlIwTNunGiisRltChPP06Cwhf+gJ87p2ti560bJfoCv3J3xu9DZyJ5BL
X+7cYb2tzo9cQP5DDEmWIrbFrhTfTBpSzXZNtExUxuiuIoTFRvevm3nRPOUwwQwPkSuojuEfXS5L
VyIfY0zu00v9JcHtbXXvCnMFvjO3fD9uM1bYxRfeMZUJMe94otj61jbNcLEAJ6Yy1SkQz6H8aEVb
UVc4xYiYKLLYo4mMrQcrsKnzAvKyEv+bk8S1IE0RFL2Rm8hBdigK9+U+YeMPrUz99tlG4rrJ1dnv
IxotpU8o0CWMTb7MfJnwbOHZ4CyeqxYUFo3dHurLLhxFbNbQkW6Xb4m8g3qRe5FQWdfaa6xJrWqx
VwYfFFqrmi2BRItXxqY3nBaVwTcf+qPVgEt0b0bjkbHvdeN9TvSl/TJQ7eZocdn2fXuMiVic5s06
TeghgB5umerndj45ql+sJFb+BU2xIKh0V9IA3hRZbOL0SzQmCSdQ75F1lG3UOaJ47AtsT1mg6QU6
ufq+bHAblGy3+A2R7N9ceduubQG+ecEMhjNVL8j8iD2DdbAxoHolpB/bBPYk7CQ/paKhWPLtr/bZ
ufsufWqvwaM1ISOwhLoAxnZJGhUGwRUb2VOJkQPBmLknLfU7/IXsHlw5O9mXnDzRQ1ZNfCsfcdom
ZuFBT07KPT9Dsi0y0EcTKwkIY8HwaNN+UIz9Z5eMiJgMPG/BTeQ+3jSpl0sNg3eq93IXECD/sc7o
+JyHlY/7s+N0b//QaLPhbJyuHe5e+sWlLccaLHHYYWy4t3L9u1HL9lusIeIvq50k4UQwMOhBjE9h
0RirY/7qmFWvEmHsGKUG+JipRrAgmifMK/DwVmoLSWyao9g9mptqgLH5LMYU5vDke8ykNXAnI8W1
pLAnY47Rsq4Wo/rx7FyrqUXVFhLxM3ARIteIJngWt/SRW56m5vOuSKZEzFdRZnluG+RoO3bW+YtW
RMDs/OiwZmL9m6SFlaPmN4cHGNL6ygifns9ZOGPE1K3rBUz//uypmM9TqT4tEBkSIviE9mcnFQhj
J2hzzRaUVokxuq09JQBzHe/L2U5Y4HanYD3pYYCBEnctIxkDOE3K4Y6/5tZh3uZb8LeIMOImQc5q
RvWflZPnnkyhPP+ZxoQGgmFBUZMPU0LdXNXAI6vlCK0IVaWzjuKo5P0V1hHFwikmuqqKCH/aVigx
jDFHAhmChVpBnH02AeoSMq8MIozbTX0mY/IFYgeYMgqAO2Ip5OmIpdI2z+HPf+Edp+arwTrqyXQF
sScgbyd+gBM/CgvFZ10Qu6Lk/PuAMXZUgWeZqLSbWn+AQmJISUYf9El4Qg6zBLrKFjiJ9MVZmP8r
CDuCeOKEjHSmGkb/w+4p2EZFJqa0a/ZrOtxqUCaMFUafjnG70/SDFKnU9UEJc+ay0A+sdyuwXowg
cGcP0X9QzqtzjScgSf9brD+esabmVo+V4N8lebbGOwat6tTfg4IxfSGiz7ZJ4JVgwda44aNazPy6
aPtm/bRzXs4RenFjCKlaOjQ+VvG4u57RhfqS4CjcefUTyjiao7zg+LDD2kNuckOeFpQ339Lxhp0n
lpFM+b4jshNBXgwOYlhqd0Mi81qDWlmZBINb7ApxFnpv3Lf45js9G29iZdQkfXhSLHvQZki/gnHJ
ndkmi1vJmPKIt3cT8F/lt6oBZY1Mj/g+v2s0akxIld6RXXP3c5sdmh5KiQBX9E/BmWBKrOf3I8p2
H2SQZ5p+E0aB+LikoV7h78EJQGyUKZ4UDHydn6Oc38P7UV2PMXX8gZsnLZ0k1gt8fyT+N/7nfD4u
AhOdem1UhMI1B6ZTyy9FZxZ+SSKg3NIQECIlDYJd8q5Ih4fCsx0xmyqnz7Rck6NxgBIRtlQnjPXI
DRbheSpvAsGbXBuk44c2KYeSpCLWf52U1w6b0E/SUcEbSz2SuUvv7lknvZbxddXGKR/7rILHEBB3
Mh1t2slhvvvDxgHOqlwoU5Ri/dv6pJQWzm0LoBog5mkGkFZpAskhBSWMuWMGTbcovKBvW6CmNugT
t2Qah+1XhoxoTMal5z0zDlOgk6Fk7plAfZmKGpq0ysChH8iphMfCbVsnsF50kKzHmcjrZKpv4/GJ
fJUM+dPLPlxDP7ms4e5fLNguDRMjQ/kaLh+AawWHWZj6+cJsi/rpkNZYO0LeKBxH3PI753P6HNDr
cF29fuTRyByvnnfgW5YV9hC1XEZQgoY0EptI7j8vSawb1s0GSWWzun/rVNpEEfNoY9pMk48eLr5g
gWlo2FrcFNGa2SB1tNZZBkcYJIoCIzxUewOB0JlcvUAMajVU4v23IF3refDIQRFKw2xvTy1ukrAy
wU8AoM/L5lKvgJz27t0MyPJbYYFgCQaBifRPpQhecqTYBw/S8ONwtOtZAC0IJfYQyXjvR+rriftc
0Xae9Ro6uuAhy/my+kaZQaSqKi+cbV3ATlXEJFa/natre/IUa7E/IKr7haLn81c4MZVO+Tz1jMff
m22HLXK5YBaZnlZny5TOzDtZZ70slB7pGvivuvemd7UMjJZLm8/OSVYB8xq15VZ9ngQgQNlpvhtp
aiktFCJf9/55jzvTwJ4dnogYIC2o58rv+QUeqPeP/23cHc3UY9/QNSKplTOI4rSu2Y6ycCFZDDBt
bK+wUlEW5By0JyELS7YkxIHh3t3aH3i77IQrW9XYSfhI1Fa3GRo6qSuOOQ2EjKnp1ZGnTGhqVVd2
G5xcVJDXn5poHTZM5OHFd3flJz29bQF1D7WemrQu4GthavsVzSVaP2v0tiF4ZnDGGdVxIY5sTI0i
k1ohBbaVHzhmWoFBIQbrnHFLmWuyghs0Le9Nur2y9yVDI5ZAYP8+dV3MNTldu8i/CvjFaiSuwD5A
5HR7eQFDznWEVRvVHtJd+JBtLp1Lk/oYrkirmQ6Li/PwL5wIZgUN9qrEmnRAcbVZyYdIh3VErAkB
PeQiqndSxUdifyL61t3EQRRq1I2BpLUQLIRMezJhaTRRNCI0N0JGgai8q9URTFzD/g/yiSfA2Imh
yLMgjwVa63lGpkUGcU3qWQoqKpIvF4Y0N2Yh6RDGh+e7AJi4aArk319KrkLHfRewGsTvZhYYPvMS
9rcWDueWy1QUKIiAwIWQ6LTZLEIl43tdPpG6sgRjS2cciAubAB98HL9up1JMttQ89fCdcaQJwGXk
XV72EYDVdZOu6L7E098Tp8d8LhTzAuRaL/tQy4uEpTBmfRlrshXVaoi6c3s39nP8pruJJtciV6xp
V8bnqsorA/O6v5F8tUvOeZ0k4lQoRy1ceMddX4STvHmAeUYpBtoKw9YKiw6AUF3boCAdUvgn2u3M
OsXnb/Mu+M4OHxzQxQy7RG0Vdu8DIq5PP9KZ815EIVqil97yxaF4CrH0LUXq6VJsCwd+C6lejo9E
uGcnf4gvodrhferQbXyEq3mpaVJiJiPECWsrgtjU3l7HAMjYng8GiNOR0Nggz34wXjyCnziP0+Ia
NujjXV5AVv7oNYdOCpVctPhNTGyOtsT/tAoB5AeAA6RHqD06MnocECtOZoAw7FQF69PJjbGFUo85
aLrWpM+MDbl328N5Ie71gebIISdEvaW8XGeEtF8T7p8biCLCiKKdE83oCDz2xD7cflhEsGTqnBVA
2P9qFsUC8U7Ofa3O4GFTsPfUAk8itQ0DpLnEevsYcr9LCIXszav/5o44TvVyPNcvij6tb4E2u6Xz
iB1Bv4wz+JnmRni4MgB3H0yYF6Z8C55LKlKwVeMUvHV3NsrQVRMPO/A4QVEFNCbkmIBgHjJiimlP
aRO7s/PMhmkamT7hA6k3vy73JD5BB09Z7a3CBQSVuryDkXo46bNvgCz7Q1iV0q+GgIlfRAJlhOba
UksPd79fsFvx0lKXeOFBZJYfYSyyuXTsSMjsUXiyBHibrDAxZGuvezrA++C1omakyQjuJL4qO2J9
VlLEdyHP/jZ1L/CMON4lpv/wnyfSc4262tg9AxfhQWEoxsGiD9MhXS8COw6ZnRL0a8fJqRgrRX4T
ypjye/7S3RRg9J14ntaaQ90XndSWKklZMiJ5TGsJ29yjxSyACFj73aE0r7vsWr1uQ0KIAxskp8Tj
AwefolkPK3nFFfvfJ+zjr6ziTkvhlThGZNyfZLUviowl6Eu+y98jywzs3Z2PNgSwZ9DEl+cJ7yPD
ghk7KDm1yEPMZLro2AaMUEiSuuKAGY4BEXREF9ZG1OOvNH8zNX/DGZ+99lDQm+bGFCRa2bjT0hE/
VSUGEMRr2Q3XSDJA1JmqOSeQEXQAt8wkIwb9E+HQLFgObjNi2974fI/DvyFDKePT/+yMo8Xtef5G
YfzLpcS+vYO+1lWr7H2trFCHdVU8Hj+JsXxwNu88PExaYLJxwJlHEx5M1NnVqT5CaJT245h8JHh5
f+9N9M1gPiJb7vf2/NtBvjewWEsduEPbUI9SLdbMUkrlVz4B6f/QZJqLWGk7Oal4c2le0ju5gYtp
Yp00rRZLQJ6u3XP0xKDFf7/qkVx/ViDOX6VoqXMjYPA0aOc+v7GnvDo5ZE3dDKkSFylQPrjzA588
J2JLQIibjQw6LbYJXFDCu4adw0WSVpKV3oaUV8DJCP8ON2KX1hBfym0wWw4y4IGGqIUInjVMlEU3
t++OG7vmwknYZ0a7GiN58iaB6MrbKDyyDYAJzuVpjDYZoBvEPSNHhDs5E1CZv3IIOCZFqXZwL9fQ
tPPsyvdWthuTWSikfLp8Fc1uQe2lSFOsXyh3QAp+AUGRfoIsIGrWPBGGec5+qniZf6gLO+MrELiw
r149zqZGc1O85XXWpTU9qZVYHEku1DTqGeh98+QMCeWYp7ryYEfjuvnVX+r0DzwFOqrpNyc9Mx95
/mVFZeH95KxUkRZuASXk9Dl9scQyN0ZgZ1IWqXaOk2eNXnLOIlDDSfpwYT5H7iRNUGRrmAWd8+sS
IBgjAU4tIreQEVATq141vo6m9Pym7bOSUYmrx2I3uA5E1Rv2DzSkUKtH2PH6kyjHb8N6hWNxNzmj
gAuF6gX3NqlTK8OX3zCVATiMjdSKMV3Nm09hBNLW0CGDRSREX+XpGie6FToQr7qTx9R11iN9nG+3
jmlQ7jdAevIznlwntsCjJYBKIniGiggrZF9j9ji6lh7EMq2UyfsNT8AuhBIl2z/jPNKnnIovf9wb
/JqoLnOmTvM+jq8oGdqsAgqChhCv+MJ8rg0y/l06n1RK4/m/JVxmSQd0fF3OGaaWRleXDb4s/jE3
kbpl7IKlsXheA5qdGaAX/0Km6Eh0gFzUAAXXqkhLn5EMVDwJQD0DD8ZYxpA8RuG54d8IlXlGtBm4
rHpiEIrQ+VMHGT28HV1tdPO1gYWyoV2l9sW0uB5Zn4fZpzHx+7cSav88KgtqKFWXOTCI4QCDXapo
1eLVNhx5boY0OUuERylyhaxAvkCz2WkXLvBk0IlHC3jbtijLLkkoBz13CTNsGtqxPiihdA3sJhd3
TboWkchA660v+/btu7ZV10E0hUu/TNZQ7AkHIdx/lGcHOXNJiU6XtUU41Gmx0ePIl4zuPf8MML+v
/rNLswcTh04hwzIsaQYCFKnGt7BA5HbaUX51lk4i2WV0QWN9B3/t7Nos7+vEKJi8afjiEfpcR+tK
yCCEbU91umTNICIc4BWDQ9w5Y5QWFEQi8pZBmYk0qyOGBAHW7mMTh82x0cGgfMVNpoRoeE/nznNP
UzBwSd+ICB5e/gnSLU+eWn4lx+GT4mp+0h8KtgUGtA5sNjWYcgFuWUhR5lDIbPH1fODDoWSuR29b
/yKuzHsatcHev+vxcW4FvNl2D3EYc3QbUnjlpMCnEPiW6GvWBirVoEw64LjkP7rYGO/HrjGb9Eac
FRwe6shoXPIwXHSNGzL09U95EKPslABhmwd+YxujZNOSzubNFAt8WSYvfX0n8Cj0LsMcyIz2vmry
qCJbd3mz5k7W/t7/RbeY5gYDGWRF7/AFL/+HjlGPPXCNUzEKUk0JB7sKneU2SZYSVwk9XFcYIH3T
wYhwBWrf2OCi5tb6mevi2uNZnorFnmsba0socuOsJEuwHWPsYBY/ms2W7YTkNmLKkeqB8XAJZKhC
iuKnX9cUXY0srqbRSihmv29XYI+Lfvh7/5Ts738X14TbmcT8PnbXEY3MSg+xVzSLwJCqcQ1ODG64
ePEIOAQa8glflYmjwoLMpWGRDU7pyBfr9JsMZax8Uu+BPoOL7hzcUBSgTc7xA06+3ndFqjYMDQdb
0PkSgeaDaWaO0yCtYneIcNvdYjIAqbX81l+HPMSyVoR4g3Q+etiqzPbIX8zMX49aSfal7xgYcHpJ
PdmWNYbduw9I8UD9tPVBs7lV+nT0mElaVYXeP3hTkb6HKNNB/mX2jsKk2K3+p5v7JUH8U3yitbGe
uFzMA7YolBA9wGSuHdyKKmxwYG2paDgEmrTWtTuqahN6Tevule1OuuyaRJ8QG4aZwkubQkqX8fOw
Z6vbLOfYklS1/RKnPAa4CC7NSBodgcC3k/UzSAtMjhlIdug3ehS3jyPj1EvNbDLu+vti4dMsujvt
Bn8C93MeriR8bC5TJJppwyzOz0+YnP0Zy2frimKNzy2et6Qxq4aJM6cZA/tWnMbjMRAwvbBfFnoo
dC8Tt4hRREtm0MAWXbXfhH3ayvPPN1+UMTnvXdFSLHRCpu8dp1IHmcUCVW0N7NuTCt32pmX9Eosi
gkToJJfGGqXzVO+97ph35rKf8LzcUUOMtxYxTM2WzQVzUtvVWeAhy1kBb0Y5QKVSkoBBGRXkHGzO
eGj7tO+OHNFWbuOB+NeF+RwSmfttcDJlQmXCOOkiglK0xpDSxWmsbY9nEqGn5L1lGM7VFaB3bV0h
5b2kfrPCR5rNQSADR1qL/sGU/tK50/l1CaRUrpagkMl5UpjC1QpqBNzfRQUVSnCf4PRYSgg/lhhj
d0G9pbz4yw30dpo2oFrs9kO3IbQscHmz1hio+O/NCZcUa6FgIetk1VNXbq4LdtP5WkrncGvXAlGJ
ba53kfvc74jlT23uPsU0EwD+WWIzG9T3obrpbAYy3IIZztvZEatUIDgY8LQDc8CcIiGbq20EBNlH
Hr5RMnCMEjxktOLsmIiqJQiXKqfRA2OGKNnyeV4ygonKM4KGauRWK/xnH/VBx2WS/Utw1XK+66WM
m77GfOQqsJF8eF3lUpNhXV8SA95kIIEs9uCx8kWz/csmFZLW29sHJmKivgh1s5TGqmbtw3jE210X
HxNkcTRnu68UUET6qTUltV/lnyxf2Z/gWTlLk5sZxP1uSQ6jBKcmTREXNaP/nPdSwsIkMTml3g1h
qbPhCIx2h2GdCEKoC7Uqo1qL4IHQu+gXnigwhaeEf5C0cXNF+CeFkqGKu27DjWbxxW5xxtqTXFZO
0R/PmIN9TQeK6jfUT6gKAcLS2gPISIGgUADmIUUoROgqHeOM8yDytMbk42dPtlCK8YnJq2zltW79
S5ehk9gI0n9QsZ3HazFZUa7y+ecpNHcGbvhEPXS+n7HeOHcdmiVOIAjOPGO5GXn3sBjjjFT2hVwA
Gn1/+Fr7i7wSR28eGe3+yH7IahONHXrBeIswKm4JbVo6ZHfcHgZT2W+uK2tynM301gbK+fAZgOe1
23AaaW8S9RwnfatTO1LTxi5xKd0YSiUSurHlfibljSl4Ps4feg+6KU/VUcUKyhOdad0TfbkZaEyK
U6w7pSLtO/D3byNzHSIPogHF5RBBncaEgNW2l9If/ZT+wG+ha+8sCHJxFfrzpVtfrtXROUh6ZmEt
JfJOOvgyw1snV0bBWMn58LpU/bH0ItSqylWIYBkCrjRAcTgq0m5gqlMTbFnEqovBxe+E5kwjS+ke
u8QNMuoGLHT/Bt8TJ4sfVSY/5ch9a5Kcx3AqY1Hywtkfs9xcg38buj3jb/5aP4YLpjEsEw3Wl7+Y
ZiPv0dY4oO/rB2+BcWJBse8Voiyi/uVu5xzyEfOpvJsPwfX/JG1IL7nnu3z8uO59EXoIwfZg5nN8
Ugcte8TmSbwGQe28C/NG+1rp12jI6l8ent9x5UNYuFyyPh/3S89nrWQaxWUyjWoZjAdotHNcz2ru
jYhYsS6bbUxcJS/MqtTHmLvAJh4o6tJuvBBthUnaL96ADxsFAupXAetsW1CO8ABCsM3AD14HERyW
z6NPYiXXOYFPS8shDATgYrmQHDvRokdQEB5I/sVa8MPc7mTSuOafNUfJL0SAmfg20wff0fi4ZN7G
KSlQtEaCR9PZNMMy0UhvKppL9h8+27nN3CJtbC3WnuycY6G0bjQt5k/K3LvsW7SBalMWLI6X4XC7
7O9amNWiSIJewaTNMs1r0yv4B5PkB01RxXuexDllDzOzCUSBQAy2lxA2ZjJeCekll2jeALTpoC98
w/oZiFCqmKqhEAgbpofAKVAaIYEhgk+SP87C0C2fBkmPElFDpvNLI5rbIIcinFt5YJjoIH/5nT9p
HBKa5rDMl5oj56rLatfUYKjcX9NITbRxkZjYP2SxrsZM1OFqEMB7q73XXHI7tG9thBOtgt0QgGOQ
UpnkLneN4TT6TLZHaGak/4XRHlbrXgFrBKfAR1NaxSnegAz1399+tf00FIHfuHGIOlEXXa8Mcojc
fIAaJExXY67Qlz7BZmfMmBllxYn10q1zFAegrFjYOA0Kt1gZTntEIMzHNPqlP6aHAVJtbpZuQz/a
upZY0N097reSVqIDginALi3HQ5ej6fGx/kOIaKFYZP0AeOfCvvjeSD3ldn4eUjcRfxkC9gmB5L5g
Z/ycSoDo51BnuGRuqxK2nTdEEC3JckHElLXGf5u4YaePIc79rHeIAcijeXATOJinVm3sq9Uw42Vn
JmyXja9oG1NUt4uZsLW7V3CyNkLlAmGtyMQbcOdyOjYd5zodEijlyqa37tGnQxt7vU+8p9s0tdbN
VWb3wSzcYgor+zjdEmQZznv2iE04TGGFLXEu/RsZCZvgJEoR3XSAoMnGOY08The9oYxJLxlLgHxu
w16VXk4mA2i2pYITTUCnnT1lPLfu1QyJUvCaBNt+yS5BnAfL+HtIKE3oSg6WlU75O/05bWYw5bHY
H/N6OhynmpKiETXXmv7SJyYRVogKTNa4cY5q9B/Cm6nqsrD7wvYrzHb/P9bI/LmRAYozzwJBlj32
jalqTLAilKN9PBywiIp1fBAn86yQKV88+P4op63+CNRgWB6FwerZx8o1WwbPMmtrn4P7JkXge7hp
+CNhbfWKYlSgdy/g2jNjEIB11QX8AIsuxed6SYAfyq/gFIKbaKy/LuHYffPLKq27Iy7t3cXuEpV1
y0qUCmg4jfHuRjfCLjbOAWqQbTHJe+sJI6S/O+HWuYc+zmkWakt1FaDetNB1MDQPR3Qh5TCtTz27
39hhfz764LHm34PWuryKV2wheyKCRe+OtP0fAkKPko5kNYmhZljNCBHhoWPyHUV6vcl0RITzj2H2
OS1Hprea+z0wtGBBVgC50K3VrcKwoIxpeNzXC50j6U8F6keudx2+jrDypGvcM4TaPcdh0n4toZjN
oqYGdRhMHCH6MGMg0TrMr6eYrz/hjrnQq/P0sIHzAKCGZ/fHD6tmy9vcN5JhxKx1yDzgsFN0Hma3
H+DoOPUrx9Z0oxGKrbT0j81K7Ia9Zb1lcjECIQKV5bSitSOEVI23PeMWh9G2aIf5CnNvmnM8pe0w
tJLZ45e++PGZZRri3RON3NYXWFxf/u9QDh3KxUhomsOwkKBtw7SWib/ba1qWG8KiOOtYWZ/ogHme
YdapjYcqmV9+de+nsJ4f24iBB0UVDRx+vGRHkK+IDXvqpbTFy9piOY3h7RD98deSHXzSDWognTZ/
In9CsclIoro8vtohlsAfGoBM44NPbivKz43UatOuU8OzqmF/e8k/Xul1CL3K23ZENh5WwljAhAyB
meHDrPVX9pd7ZK/4KstCajwrMgCshBu2N9rN1CHPRK5sJafpFQdOxLSe6ZCs0juFabgPp8V3+0vj
mXwKRmF/dVwfG3wE+gZoYKtIuovhtQc8MSJEOvTJJERfIquWUiwwt5YP59xVN7t+vLed3+RvV6RN
+WeTVXLAXCdTqTiKf6pkgdqydW4tEl/dkekPhSWJZHRajCpqHDDPkJmRhLlZqbwJZ8LT5oiIE2xz
KNVfrEi4j5EVzJ2uljlN6dKFSOWV6zcBnn1QVyHEbL4mmzi8hYBbiKKNu7LY32xdhbnMdOQxhT3+
nHhcpc3StS9xx3gXYLboCIiiLlgpPFvTasR8c1RZAfKdwHr7CptCAbGzjZbIpmx/1c8IJ+ppMJ4j
xVNI+H/jd6mTLZ0zMRc5ChSBsMvFZbklrgShUKC72dow5JAJgT76ffdoxT3y24gByYXOCa1it7mS
JUkYr+Ur5XPlDIF6EZV4uuHOXje1bGBZzAgYKLEk+HJUV8nufFUWqk/LchwwTgi0DXnVxls9biBa
QS49lb55/9COULa587O/9FUi6V41rvmT1pEZdb9vFgZF9z2XMIiRKkEFjexsFpj7lSILqZaxG89p
LYXXdkI5Dr4eQJLpgoMmTQfLjf4FwGVPLgEXFTE8o3iolQv/piZYvlvi/haQ1wpym3yWZAW25k8G
Ld85ZYsAEJajwYZ4qCGjAS9FDd83ZmuaXcn4QePDFSmnDA/UvVW5z2Fs4qhXLg8l0nAClW5Y0MPt
f2On+ife5dkD2YWsSkjRkDnJ2nfGnN1iH/6d1eE0KLOogbEAmC48ttlty+tmvn4AD+3xOpZ44gBT
5NF524AaEDhfaxK5j6atvDOR0u/ZvL44Y8i10zTIgolk6iGJYvku4otFAuaF/0UTPQRXF2wV2J7P
K3QnAimC5QO5mwvRnYX9zKW2nEEI88xUU3uiidkB7df9NKAWfx7NpiU477al1x8AYjsHsfAa3CqK
zNSPn+t1Rw27fRoY2hcT1l+MMOJ4W4jgoXkIjUzEhJM8h0NyRAI7chgCZQu+zAZA3y39mmSQ4ifz
UPIneXYUq67mRMc6XhQRUkJ0cgLH91++WjWWgfhXUO4YTIWf+1wX0f959ljSlClHUbaJh78ND1du
FVSUmtQ3fDbJVj4/Wj6RNp9Hya4jToq8lcBMZ3GsWHYP1OJkuGGeKBwrsK5kpmPtuYq3bJAOd8wK
SN20HQwqUCkNFADi6G4c9gRJPK3hMO/f8//gfYGp5JCwf4yeCFSrhrXsa+vzLlL82R3tvQLT6uAm
QO2UYxaU4SY10TiBUuKfT9cWJJqnkrCynx4xjUL8POB9FlcXS7td7keAH4PuO30dkOORNcVUaiX7
Q2RkH1FFcHd1jamo+KyBxjW4GquU8AQQL+lzwOhcqG00SK0Snr1vDHASLCfsLkSrT7d1IC6nb4Tw
tDMb/BAjcLTqn4uFmloGiGK1FTdCIPqqz+pwjwVaZn0G1PIs7x4nWvsE0JWoaKidOBFVDDvvjEhx
/HQC5Xwgr5AHsITHAUP3RWfFNaKz1YjA1TAUqNc8AYcOu/owtoY28Dju33GtFbz66SeQaSRArjCA
tmwZse6SxXlGgwdZXdPHTZK/S1InOBYIKaNuJfOalpSdikiS1ZzyY3imU6ODTl2FDkUXMh3JJ4Cl
0vB/SxC5S3BVmnhE9I3NOBUjlRmp+zVNc4cnIskiMyGPBiW90TzuAmMEzjJQ5nKFmXut9gpONITg
RefThBxQ16802TpK477cNwjr8ztK6+pXUO7YTMJG+Wwq4GPWUfhYAgb70adDyRuAYv5Hvn/AFfxK
ZvVhRTBMO6YORtgalKBZnQnzon70yfROU9nDAmn4vyIf/wzc7GMUiazAeUjso6mWO52n8vBCNCm9
DcgISn2kUjUwYVcLIbyyyY07IX26H8bBq7FCwsdP2eAfzAPjR+qJorPjOFsUxUB4rNJGXCyHhJR3
HjpCtLHLiUbV1gRfFtdNp6maCHmWUnzixJd4oQLTFQsWVgejkvCP5vHEr3HjZVvsVXTqm8YCVd5P
Qgn3J15AErKeE7xZrTSPl5WV0LILaELpNaQ9bpi2BrcO+DrxbblnfiPYQfZSh3fM2fPLXpno4Ho7
p5LczIX2pRG4ycnxBCfisReAgX6hPlx4VEqiHYZlvEdYKKW10EwD8/OD9ev4k14fehImKlAzQCGQ
l7x4VXEXtYgS2O2VJHi563AOpGzxE9cShcxXCsAIp7BrE2KxkAD3iEuNOQ1qLOTEbNGLOociKq0W
hO7jTnHgiMZN/YJrewg6KTFy7+pTWSJX0BQ6vwDSQQ+eWXApTIg8yi0IYIP7qJ+ywIji4xm/pS+q
ePB7weFT32elKdANQssJNL00lf1q6IB73ljoVSQ9W1z28Sn7bwIWfreGRd8yWdakY5Uin2QBqSBA
GdRqP44kVio905gLy5eA9yCs9+bM5cnihlxlGjbjls0iMQmyykgQccrTwj7JTLRk1ib+7YlNBtSQ
cKVvY3QkDdyxucUWLeKLnFNKiL/11ZCm1UuH23DyEmTS9NNdTYFpQnQ2M1L/Ce32J362l5ofsWXV
pEV9ygQcNpxAOz7+fQQH569jUsRqvYLEWCXBgFoap5P1meBbS7wZpys6TPKQUaaHqJpRmysPByh6
AhgV8Su5xDC00PaUqRuKP2UBDUXOC6S9Ig1l7jpzwWewsy9W7EKNhG8MSHXmvh3/kd4AJcCVd3rV
gTVqh3jw8h/reGxRuMiLRh8nOzUXiykHUXTNzUGdATu6qq+mkay2ZVvJgTu/9NSUFpCzH6RamjoS
npg8vZqNf9WDZPUb1/c2buCFy6EABHmwHWfJTG+JkHbiiD8VVKw1ExaLOlLOqmwMdVNCRr+UF0hw
zB7DlgScC+mgtPm+g6rrokqmyhAIyPc/bZ7/CzRwcTlRQH48UuIfhgCXoS2Vvce7TD3eBJ+KXXC/
3Fs8vkxDnNwsAf6+dxUw9+4jgcuP6DrlO0EC3rPHL1V5blEKdldbiFJiqUgd2uPY13L1MJkvdG2C
ki73p5K3qyVKekiJQtTVkqTop/Bq5SBH8KcIGyWrZH+qWLUy+NSGtVMn33DwRtSbOjbJ+OZqD5XY
gGD8M5D4xr3pY4jfFHm7xb4OVufhnaValQNAXb7SpyDe7gIIGmYgiJYOCR5ETeuXR6vuQYQMbuGS
GTiJLFOm4+LUD0o/2Um2LLswyWH+S18HTkvBHItRazobEqA13jcXWvg9e8ZNLkZ5xJxyYPnAmb0c
FsgQL3YS/Lg2GfksAm4jwvMMhoKX3kcrwWADUxRCzFwuOq2EFxFJyd8HSUDBryeV16aoWSYJjhoo
RmDzyMRgtW9YReK/u3XmcnpZmGL7F0ugwIM+RF2NYSHFudyMmsBBJGZPBFt8Uu72G0cL+I4h6Pu9
Owg4g0eaeH7LgeJdYr1dlQGpFrI89zBjXQLjKnnRy07hbvTVsh0ciTKntdZvmX0Vgx9mDRXAz4ob
TSdlxbU17wcVvZsk29MGSVvPL0Lxu+J89YPsci3Avtx/GR6FoKEKF7YcSB5hFgS0r+XSxlof3Tl/
MKjHT2jV7EL1z6OeYJUepeVr47sVQoDR8dlzl+rmicEasHTgOZV/YAWJppyjigy5Bprjct/cCFKF
XDx0jX6hR+cujTYWjR94ZaLdUCJt+XO7lAWn/MhInR8D1keqhBYYH408Kl2R19OMzJGP1Q4tuwHQ
sSHDIHLOULdVkkETezQWn1I1L5+ZAtymRFOxxijOOXixNZwrBKUHxsCOiydoLhWl+9uz//Olrpdy
rt4m1dACT6782RSbkFRTE+FkY5y5z5MrX+9oanpHa0Gq1MDJx7oCjF5EAdpozE5CZXe7m07Xh9dm
l4vah++38Hub9k3z/iTuCAr3gvO4CmTTVjSsscCSgCnaVWfO4JrCyeByJWFJEsYtZPsg1trULjMw
xviqsHc1cAm/4PBEH1Q3FXLUbO7CgcJ2XkVMlAFs1XX9Uj85H5h91kioCX4zB8xSOPeinvCDeCVw
L2xEuFznPhQDa/4c74d9CEjnZTDbZpJ6W4Y00QKqAzGf3Bni5gVLLXlHcWiVkTCTv8tTF5AFjGDG
o1DxftJ1vceOy0fKxoLzAPQpdzaOFB4XEZmf+NYsQCmK1Egd0PQI/d5IqSogz/7WkGho9urCFafY
XK8BWMjV3ct5KWAQ7gDQ1FKc4vF/kSnICUGZGMXlnxDDSkXcfgxxxk1KO0+Bq3IVx9XMkbm3Y20m
7/uoL5ftEpZcA1caAvRoIID7hJ9tKNm75h5I4cZHoyx9vSW1V1G+nUqkMqMtsOzBZ5PvyP0vGQGf
AMOQGn5ontBFtAWPhuXI+bjHXmuhbXHei+RvnBDU5bZTetzY8LtkQqq1hrDdT+H+EPSH9gJ9vigz
fCZouGl12Eoq8hsC9JeUIGV/1U3ztai4y8hJyb96WiLOyC4UDd1obWaWwOb6W/SF9ATsyz9nYrtA
VP8bzxh+lr9PxVGPwAjRNK1NuC06NaPZ7JG+dGi0lejqXQQFa3AFabNJj+4s+dsIwDu0j1pwUe+E
ciaEbLSdaXCCxPNeaHqDMdwGjMkg+Q7mgox777qhZkq6UdbNhzplCVumSRov/RmTjYSWd4QbEoSQ
eMOFLBriysX6r7S9p0FiavZtq0ogmgLy1romrJSfC42RSdphOgRsI77yynWHBNOZFmVuvqMo97X6
Jbn1wnAswUbiBdfPA9bpqCeWPXNqQEcDko5+azpMwVVi+Y4rZ5R05ToZdur1S5GWmzxMCmyXxrmM
r6Qpde2SrAZr46TKwtmGD79y9wriKIG9ESg+1Y5OCQg3hfe+p2iHvMUIZIozApbWdN+g2BqWQokU
jVKJpHzTU0M6SrQHWBARTrvINj1K6WI7YM5RPTS2NtsLHnzPS9Uf+L7uu8g0+YulDMAKUjB3Dq7V
9sDL+LFJQogrLZTjheVkCH2c6ZjjxGFXnXtLAmYY1MxLWUnZwfDQ03YmJIMXSciaTMHFyEwB1p3R
QuB1VHJMiMddU5C0EiaAGpIZM9xjZWiNu6Y0Ah7VQisCrq1OVosaHvfspAXG8b/fslrMeMpLYNt9
fs5tTeY51ht+zX7ByyGQ/gJ5CK/ePZsgl+Jxf4mWjkQncyEW0X1sD9SivFHciMuxFMPhLdj+x4FP
tbqGfhIeGyQiHjkSJiqySPqeYZeho/VtZbsSQNg/H5ZIh2/E7O2jA64tR5dxm2Qcdl2UPO0p2i0U
EBecXwgMLEFd243lNrTTsd5LOZF/8WHs1yIhInOz9EPNU59bwVfgQR7zeH11BdFXIhMYvifj4daE
qAHNSJk6RjxW2ZriwJ6EiJ/Aw+NgA8B2Nd//YzxKop06sMWp50XQ5LjhVchhVq0hV36W8rajv4XT
JIhjGIiGPPEWrX0Aw7eB+Lr6j8tzF4kF8XtuzDsOaS5oHGXTijcgcSnJT37m3MuHwThiBU8f8baC
MvLpvCClPhV+YHqqlMHqiI0hG6tZOFWc3I9KVQehwnMxB3q+f2t9U0OvBkJUdgZtTQ4NcIkdOP68
USWI0/Kd3lpx2cT3+0PQy4K4qDvB2XQFOgmgmVEIA7ddAa96t6bvhIkf9PZjpeIatzJztKrDw0wU
+wbGeqRssSsadHdEzwI49Wze0MHQSeBbr2CiYbrboingn6Lu3WvvT1FYD3YYjbaBN0fiwGnd01uV
QKLTPQ2K+vfmID0uX8tQ3XW990TXBgczO3RPRfmgePYpAOtk1gdF4m0NZa+GDcDyMcRRbzLBSaKe
3ppbVB8cCKT2p58IKX7dxXMuJyAAuZjW+bpAj+xlrqzkh/KILf5irW6HZbiW5y0L5RdkOtff/09g
SWUSI44XWB1kzPsLCG5l4wPzE9ZYUw/13McQUnkYBE8m1VXd4bRCn6KVnwnialwOulC1ZUQGOAvq
msXuX3/2XPjpFrVEJTli1+kJcgk/jwHZqsYtiIsL10OV4Im4chSAAKe9p3CFFlXu5lruiU7oDrYF
fd8gsyckh9OamKIn04XXYpsetfy2KaHNXC9LwAMx9HrM+TKpzWD6r8jKfDdFXORYCMgOf1xLl4hm
XqNjqtZLV7yne5z2YJNi65amHLxaBwVls/etI9Ag+2cA4EX6NvULDOhfrP0dGyPolRSrWff3Cy/t
Jk6vWX7TMLfYsAXh6GnJjp/KbDpcvP9ATuLwrPKV+oATQTBPABFBdPicdlZs/wrQ8hZ52+iW2nde
0yS88tDa+4HnkTgRLA5MGBDujtwcxMkv4yBzyYWyE+6QAaQsZ/TNYmNtiBUH8WP0PCsiJN7Mhmr0
XUHaiCGH5UrUzfzJ+TfSTglxeLNOwJ7Xac2UlIM+ifnE3MqklkFTBmf1adNLUYy2C7Bp9AclnWlG
LSobEvbtDqnm+BVQm6SnJaKacSe1jvQ3NaCzntULUjNNjnOrDrark4fgTUaNr5P2Ba1Vl7nzw/84
DFg/f2teVrVOEV9cUraZsLYndaGe/hVcZMOPqJgK7VpszGHHKNHHL0gGMs2NQc0r94F9jfxJXLY4
XqXN7uA7RmMhCyKTqDvPvTY4CnJ/7I8qsDOanRpoGVt9i/yBlfU6mOEacLZ07S6Kx2R6+QWe8/gX
jxKVa5H+5SXOqoZ4Iq8McONAzDEjD/V4ETeL3tFxwnOD6PzH70gFQB/CPJwxu3+AAhi8fPQHh09Q
amzaTb1+ee0Rg+YSTv0Y4R/UFzv6+xusAbn1jt5j3doaY8ZnWmFVbRAgZ31z29vJbg+WC/hhYdyE
3XOh3O0ZIKWsPNxx6fkiselJ4fAO20VrHA9dUXQwfIAr0gwKXaHGPpQ5QC0xjRKjkith8SVGmqmt
B5xin+oR4OX0P6blEx+70fdqxlwC6Yq1DBjBztYuHTvyRfyLhIHnBNod+7VDtBoPjyy3CbdLZGA1
qvz3K3Cq79Ql+FsiALroa5Yot1bzr6OtpJ4KZjt0UGlz2HvAYw3S9EAiVtGn/tWayuHYTgV3bCUu
0+iT9nieV3lfzAPIxCPrR51JQsHraUi+Seoe3GLQpsKX3pfTVb0Y/qDInx97hMTi0ThHXB9xLnZt
HrQlLiYAND4E4/5v2TejoxbXgUe5TrqGh047FTjv515KVZ6JYGOnQto/wFFh/jbtlFSpFhz8F9EY
dC4hrY5AVlDeGOjY/hg5ak5TW+TBOJpfa4KubeFFr42tk4gelj8o9x73UR8IE2sxvVkVZ1aoIwNR
I2cel+1vHpU8yrzdoHdc0dRlxyCAR6h0cExBIpKM0muvkuFKFcSrjFjQC4dbMhLGJd2g/J37r5pM
HlALft+wBoSCydjD53ogj+BhlkaSjkY1s0I1RfSbnagOLQLEjdkx2FnEF1975hk76v9U6d4B6/le
P9i7qw1hWITERhfzTb8jBPp7igE9W0qDOUtmT9mNFIdstkVpsu25X6ZK/6E6G+mZG/EtF92LqcBQ
zP6fADZU8hxWwWwBUnvwAuDVeI1JAs8aZLEjbUaLnncgLYzti5amPfPrpBVsM0W4Ug6CRxio5/6C
jslB+xKuT8nUS0LtonDOqvUzOjCUrgg9Jc9gan50td9vucZhZWXAw8KP7DzDlkk1uRi+JMvOzxLd
ly7gMIHc6KZQ+IhN9EKRmmcVlYWSd/wIMPym45mJOZzNi26O1lyspWSOeRrtprRtN0cAFLwv0cR+
6aaQL8aFCY8P7/PwwJfdcir9lK9XJvY1LwU20kf9OFJtOy8Ks3dtZKyUg9+Xxk+4BIN5QsEXgRvv
7/yv2mpb0OxgLDyUmnnTftp6UQ39GZTqj48uTc5m5+RUr+4je8YQKGHC/ZtYm6aC8UIGplxiEP0A
qK3llnfh3uCMxDcB8IZ3BiNz7oMhIAVZbCUIzq7KwQnIBm5cHh/dosg14Gf7umvl7FNDHLcy4ILx
J8Jo6d+fQ8cWC5eXwsyEfiNMi6bzKKErugxvnz9k6kK+728Y0qnQKABDir3i4ijVwJEeXnsIWNHh
X4s0ndnNj4VkWGp1nJkQNDrduKAKIkMfvTg+/MIkEf/s6BrI8EXVSkslkWlf+0gat3kKqmvKYv5l
GwXh5nfSO8YPViA+eQYnFEvqxiJeZS4u52WMp4obZBQn5DqB6j8lLLv09V71oSTNPb1hXzxv3NiK
86LT11oakzZZy9zs6ZPq4xb5mzMzpmB1c8dtz251IG3tQ3rqCvDen8BikFbxgg+3sGbfCD9as6ra
X9bHm0cU1tT3VlaWUHabIdf1m7KV4VRqSLZXFeaMu122bn3IAI1Xk2dNJZ0sSg/idAJnbLq7jh04
quz79Lzu++Bc2q3RW5vVQM1HIstywD7/iV7jRVCxJrKXWHwIJda65bBPXxmQMniF2z4NKEYyklFO
YUjXBb6ag5xAY5gBMirn644XZiHK+VtAzSiuOy+SfwcxqeFKElR91lVYZDbGnLUvV0afjowQBm+B
Pw/YQ2Y2n5Egmzl0Tbr1clnvWbuPo+bozgR/U1nTPnbzzxsQyB+NPq6cz7zvvAHB2+UiNg3R7teP
aD892kZXL5mL2eq9mE2vPG4awv7ZK9bO6CZmARrWko1toVfWG6JOqwx6OLcxIcwXEoBZ5ZHLxHhG
Q1yEhxbvmnD69Euz1nX8dR1V6er9bLE4/agKNBjFZ8/S3ZM2I0tYDIlfu79y8TVUNdKB9mWYi9EE
dj9ZAjFPMK6cMCz1vtOKtJJ7JJ05YzGZ6CDblhTJzitODtUY15d+1fJ8jeu/x7ufa1VG2og3/wpv
mYDmnZeL6J08wcBXj9UdufMHGhjJASUDU59TukEOhGm+QcSWgBfvIIuzsV7LA71tQ+5XIx7j3i2Z
0q+aLXnT14vsh0vMUKt+QGsLt7JnnhKvFTnb8uJW9HeCc1+ol3MI0DAyZi0o3apOUJ7rCfqlrZGy
VZ6UAyG6U1Wmn6Elb31K/iAORdhdobGH7XHDRPvbMFPBi8oirCCVPPlVT2jAVQ97FdUCS4sSREAP
S+k0T69fg8B4aTzVd3VBuIHO1gBUUl57yZb7CzruGD1TT+8lZbYvCobJAliflcAZLKrRYoQbMnBC
7H3bZMVQHo+4zjNc47MNe2VdmPgAMVF2XpsdQNAdgW4sODWNbNs0HvVQwuAciGTZNAMGFhyt8qjU
2dzYPPRO3jhqUpVxsTc6BJjlkQE//iqvtktBihIX7bx3O04APfgPRmnHvMrIKLt++Xj7Ax0ZV+vi
B7F8pzGWDs2KPw55BE71e00L47MRo5+fpR2KYIkZjofKCtyWcXFYF7J4jVUNl19GFWlJTIpDQ4QU
1bxmiLU07nstskVaY/MvVvGDa8UqPAZHa+YwE2VMwMJGag/BgNigdpFmRUud92tGiBn8xoaDyaap
XZQfTgM+8tyRsblUk0+jnon9DqNq2eExiixWTz2rVkE1sNo9X6c/ERl17snRZnQRRSS8RDkJlMZd
PWG7H9CNl87TReB4r9s/B5UMa43vr6mHz6XC6JBmYBWVZ/68tzV+ljPkR+V+vLiJf4Ztg/+6IVZr
e+Kh/ROQ72XhBvAaVCbhIPhXPIspBc3OK+WpYF7t52AzGECfXxNQaQqV9RqJqRn+qNpd0E2Tiejz
nTlhJ5phk4TrMlb7Dt37MxaalVnhuSM20piIXzU+XULWOY8k/ppFgxqW+/htiVEB47g44J6ZCBdk
ANR5955IotFaaF6po4nNVGVnsjP7XRBYVrn2PwIcY9fC3ZqymZUXseFyWLlA6Rq1r51juNZQso+8
opiIF25GEpFjh7n3GeRUgX94cgotOfmfkUUjlRmzqw2+nwl4hDec1Fh74uN/W8m+m4PSG2VqpUXG
UXILYEZwBVm0eJxZSnVDsm7ifjVHW5CnPwaVXcVPoP2Di9GQJwLn6t6WGoNRkI/+Q+tSC0n/27sw
WWZXIqi6L+VVMTZNzydNQRx4cAFXY6rc8F3oYA4HMS9Udc9vjxJw0qXzRdm0v2QOdMLQIeR0iufW
eKx5AjX5NIAw4lnAEpnt5bPhEudNtXx20nvLgSEbdPM1B7MjXiDRm49zEKDjg9RuYsDCCYPHPUnd
WI3xVSv/TecIVwNEzpOYFMCDYFQxrchJ6lpj2uF4Gfn/LIwbd8Cb0tF6+AjyZKW6nUVOo9ISfeyI
GG1cCNDPjAIR/WhL4GHroyxzFblF/ZGhXj1fehNIMqL9UKMKFPjFQrwM8DgOFdz4B6VAl1BFJfW3
O2+lG9ALmxh+5632X80GPK9agDPxXgTmmkVjhjyOKOZdztDxRjrOTYK1Y+w6r/VpljZBxDVbdxFO
mmsPrBqJgA2yGqd4+RnBEqU4jtBSlFe30cx9jJ5nVopjancSvfv8p1jG6Kvapg5+OKfSCDbKBHxw
FqtnU4ejxCsbm5QpQa9HdBLfEpyH0cBt6+s2PhIipG47knc+sSJeGadNPhgQYIlL2UCoqm7TboMQ
M6y4+2f9PwBELmXhOOCsZdgSaUMwE4TOTOA5fGjctJ6QdTV/UNJJO9t+FvrtxcWNE9dYCtxQ2d5s
KfsrVmNoVbh6qte6Kp+7PGUfvRB0BriWx6Lziyn/1FXSWugUFadylzD8d/L+lsVlcNXS7RH8TKAt
s7GNzts5mjdrg1cUFodM0isN/rmpx0EMxKHHBUN5FuXavqbqj/k3EWhcySosADQqHPSxzloUKzJ3
ql4CjEO7+vCextCcYlqmkkWzzcj4LumdS2cAXPSSuIAbFU8oDMvfNywr0QVOkTTMbbbmsRIuUmeU
DXegweNOawTpG8NgsJE6o00yviGAaLmFyX0JCT4o1HwEPmPpaNX22HVbXv4Syl1ZmWR+yyECMB1r
hazTCGXkBfHtZPnRCW7mjLd32/2qC9woeDOiqRFIHp89EaF5qn1fRoYopDLQo7EtGgbmZ8TE516u
7DK3rYapJw/eVEC5SCKklkxEOlz8Jpm2oz3Z/lHuoZef1BfscEz/+HVhJE7bub9euHafecCox+ct
Bc2dNiz7YtKj1YhDjue3af10J8Zw97lUrL2q1k4/GwEKyOkzhL6fn/twFRXHzUcgrhPfQANgv7Uy
SwMVJWR0bNMbIXPgZfkjWTyoiOonxVYEr8VRjmpcEwbZJH20C92ZBjJQE4TjqQMlfCHeLHdFac79
9c0gQmDBIWTJCb5P23RWAkJLDJaq6eYwTBcF4xPEA/xzAtWZgj891Fdhn1ID37ue32QYTc7UXRFX
XoP5P2HA3N2962byWqJzc/gfFLYXahP6WGZOPNgwSDuLVy6zHmP2Xy+tKE/R9KCxikjq/Md3MjNC
/SdPMwIb9BmnP/icCZ5RhcX8Sc6Y+p7fgBFQ/XEBTTHbEeTYrzv9IBydngXuMmzrQrCm2+f6WYlM
S1Wx8ovkfoupiayR058kZLk/kS6E29LwBIJ0WizVca9MLQGWYmKA8LXn/zUi0Lb9Jw7EpwMa3ZPi
P5Kcg/ZwBapBNRRfK0OZHabz9KYKAJuyWfXdBXR3avdIc4nw2uJTkHcnqGWmcelbZxK1uASPlqyE
+HNBRncRnGvRgzEeVktI383fiCRvoV2C2w/OUnrjP4Y8whE1m5ReQn8SHbEDwykE1PvcVsAaeVhr
IYim70HqzFuLlWPY7nUKFnK3pPfHabAL0Zq3f3fMFJ52aySYSOHP6rR4IXWWcX651YfOhbrcrTml
1zKyZtLloc5mb3mmymIRy+1PLnBIr3tWgJdOyaQcOLjkzkTa8fhRYxSU0GIKsY15ENYpmvdfJFxP
WnmyA7W2rqmDWYRSUo0WYbldNB5+jk9wP9RSdSdAnX/U/N7AFUk0BJJoTvDuoXRPbfFnvuYr1YWL
R7DUnUdCmuHHrDZx6L2QO4B6fGKusEKzE1jzZllwYT09Xd66vk5uh3Vv3zeppY85EJe0ETgAE+I/
Z4PRhCKdE7RggaMFrXwCY2fisYwmoFBgJRpEPLNEr0sXX9VvMVWXbcKfOFin293j4DF449RIlswi
TtzX4+Ip53Mr9HdVRtjTEih+Cz1IiaK8gR7vWy+JiZrrDF0yj8E2wuf0AfRz4MybeUdKIULDAAOX
GZRXeS0W0pFuFd5RVoqby+K23gIjU+6PLtvGyo2YmSptjX3IIELK5fPPggSjHMXLw7OO/ggPCx2o
0rEmHvjbr3UlOsxgSgXXjsyFqIQ8RWFUJI2paj+lLgY37audNctJJXQZ87kkJuMLLwK2WMylP89Z
pRer38Rlyk0qN30mLUYsHUul3d8w7digW6kH0vTG4xU+Giz9U5ZFBn06bfm6DufTc/FxUmP6I1w7
0RGec2CDNwVa+tJMG5h+je++syTwXrV5jCoLDQ1Oae5PX6sUV5vSFwb1t/jGxYQS/IEH+dtC35EZ
riNE8JINdN6TjgrzIaNqM6B/nkkcmt2WL1FbOfijlHf+t/MfN6yK8ybol6HD7p0d0fHDiLnJexvI
NdB9frkM/Rp53U9/4xyqHcKs8SiWNajvb9r4hZ6cKMpDwfUSY+Knyy5Q6FH6i5zclp1Y9xlImesl
eICqU27x/lZFsMPeX0lEaKpZI/3RTnh31k/8mRAZfcjpaU1qYcrO0hwcfDkaBgVSxXvi1a1pA83u
ljGxSpOrHMdCY4CWrl5MZqUycvA8nxcCvW6h052NWxFO4N195AqI8uefVCok+3n/SAJHAZIOBJSt
0d4dm9cSm31KfWqtbOzo1gh/41Jj2Jpq95MR9WW/sVzq1sbMPxa8qGRljTLO7NcI1XYcejUxMIJI
63qshGm5X92UooT9w2CixjY66sxcuvsSA3hd9s76bdNlhXfQ2rtiIRqArzpzKdfTIZOGn/AJdv29
RyH4GX/ZRrW+zUQZA1eoze77hAgCwFtxa7xexov74BcE1wd+YkWWMi3PnFJaPLpIQqW/YDGU1sh8
pH17gzXHrvJXYMFdHZ59A7fqwL/lJtRIYYH9/VU85Th/Wrr5Cyu0oKsgxKU2t+iUNU64gFMtEIqx
0WV904mJlTCudVlvCi2E82U9xFlB+LK093hxzW+xsZb0igy8+YnGlH7qD7IrdsRk2ARRjYN9xlY+
VJHMREnqmzalUX37teJ8tQS3qJhPwOFC9rO2sftQRvsTDSJEotuWOldmgZXm+APW9yUYNm+D+/qX
NCuARKlqMP3dCqrQYfRla5gIz+gFwTSdo7iSmwENr82hyei6NRxkDHbiS2itUdcE77pym5wamyby
pfjGvDW+qWT3Xf/gkQvuGh0X7dsHQTLsV++/xYUef+EkFolcQMJqtZGGHqi772CWozHsK1zVc2IJ
88abLcf9pvTrfMmiV/IjON2YLKePCr3nx4Zw0AQ98OefloflM+i3KNjvFDrIK+IbyGEI0fcvtGIB
iLgzvpl6bHopLiT+13ngatIZ5cJUk+LgqFXS9gXgwxTXxNA53H6AViVG8We3DGZYyUWljPn9goj3
Sd5Mc5MocjLUhu2SDnv9rKWpIQWUe0iAGv6kz2MDkxH4IAIY0KZ+jXDOEiOahKTDEOL+jj1RE+lV
4hoa0COc3NhD6bc9Tko3S/sNgD6JgzgsUJJBU5/AA5LcC5nPBDo0Tu0oYTPRlI++Rfn+wQUZB3R2
ncXYyVVuVXEWIpBoZp3zcMV/UhbMvkSlt20H62RQvq88pGRktKz0FV34hlHI934PAUzjoR8AZPpU
rNryj8WH2R3Ub6+1c9JTyWuLnO0WoKk9iYA86qeQBRAjs89NkqGeT5cgFiGJdeW87GykQUMFuGk9
MqhXmajTgf1MJQ7XA6KxIhZZ+1dEdLzCIbjRbql8lmGybtis5EKGDh2l5yKW5BmRbXp7YFnFVAVb
y8CRz4m3pIeoQgIiyncsiK6H0lL+pcCYonLnsSl8m6wyrZjB/LK9GiRBrw/jJLopn0eEi7tOwiPy
hFHP+bygrGu1Hp4ucEcS5NG9phzS0Hwt21irCVx4uST5AvU7D2XXMvbVx57s9U+1ZQ46IzljLBZu
O0aivlnmgZM7hMiCTTo7ejGBdQlxgpQB2hamhWuKZQreOk8qFlnWdwwW7Geqh9M2MYQgVhCBPiWR
UAnsWsMIFxw/5CzQG0YVa7y0VoTbk4sDIQcldujXnJkIDh3TWJRoPfbBf4feZX96drwJGROd6R7n
N/Yv9XE4iWWC/P1mPcadonCmLvc2whJBjrpEvgaxXBCmz/kz3Ao5+ZwQmlXM91Y1Filxxq2lTCx2
9GarR987BZn/hcaUpFc7xNFAIo+OPO36mqoDYtrWvrzvH3tZHgSwa8qn/rag4xee+DvZkV357KT9
jAq3UR/JBQzRv8JDsaYrM3yWZ91UA88Huz/NRzik/T+qE1nKgxv1BNqvanq76W/4nwMN9LcfmYLS
nPc7YKLkyyvrXMYkpzpK6W4e1Ytu5p41DbQtQgqtQ6s9SN9eH2EtsXdVFEqUM4y3JUrfrqgpF5zG
DE/cSzFR7MLTrgukJv7HyCh+3So2l0Zas0pNzlcYY3UExLAnk90w9VfYYIqL4gCuk10ZnRhpgTbJ
3Y3hozF8xZIvLboD0vUeoUnlsWMAvYXcUISIbKasDG9MbPIuQcD3CEVq3m1+xWoGYs0bOzwbzwzp
h/4wC+nijHJ1veuWuiiCI7baKafqmr9r0HL+yivpFdc8vEN+odY03D7qV6HHw2tZOHu+hgE3ronP
p6E582sag1ntuvDyY9S9FdizZ7JK/iPGiaXzAEhmPXgXLw/p3KSB71OMvDITvb+QRQleYlCDG8Wg
PDLiMJ9McEl+cbLqwQBX4J5oOolTmY7z4327w1KhJnTOU/akuinKTFlzmEUY2sthJdFuJfeMdnUM
jUN2JL4m8Mxk5Q8GGKrADmbBY4rqeLVqxbqbArj2Y6ThbCbGkkjzOZaVPUhI/NRf3YgH9ol7EC0u
Y6/RN2zP3oHHO8Cr6roRmI0etkvEXd4Bpm6zii0dDvYrcyDVRgwgAmS5DEeZJmH5CLLsodWKvHH5
D2xCRscCaCaTN11VQfe/JeFvudZH12Vg7FXhM2+BE/sq7aiOKzXRxdqjaRJuA+XbewWj2leljtPx
u4WgLx4t1JsvziXeexB+qcMHSnijgPay3D1QFXBoEoFJoT7mosb/lXqLBzKYDkGQhXCJhnncitOl
Ci/RsJ1rF6sJJYNjO+f89Jy/IuZ2WhgVRV1CCuATehaVwZX0aIOCsSUQwDYa7RSgz7xeirEH+alC
zbXydsITb9sj2K6fBqadfR47ItC+WwpeLOCAoxFjJhyINa1Y351OH5Mcqq/rCeHLVpDwT6CwYtdP
spQww7JnthS0UR/fK1W+gwEXZK/aLB05Tjh0JYkk5rPg4HeqhopOisZzJQ0AQM20APmsVNHQFKCF
dDmy6jtnQTZ3cVhnnDQULBszwKdMcTYJM6sdOam1MVoTBYd4FlzxferWbEWuFRsT3ZYoLSglmb6X
zsv/hCK87zYEOUo+LBItAlMgTyV6JgSCfEmkR90m21jikaGYOcNwk3t7gpN6KzAO7OYUFJcFq2AN
C6nCdUxI6hY7nFnWQrrW97lPPVWwIW4n5aDxb+b+jc+l2f1eJKkohT//Iskbccuv5TJPOBQJGntb
kk1H7MXd513A9t5UWmDKdM/e7xsYtc7TxBxCuMVQHhPnpOEdKneO2XM0DMVNt3nhYvj4FKE88F9d
N6M58CwfHtkYOmzod37zaOr2pOKXqDKeabjnM4o5dABXy8lyGgmdyBfaXtua+OJkhRVu/TOS5A6a
rpDy20+kwZHJoQQ0Pqh9kZ/d1zGLm1FiD95+oIeZ5QfKuCdFLedQnYuVuTh7qieLW4v0fTd8WAlw
KICkfwOrn2o8cpqgsBC0Y6h82VI6AYpjqvAd3FxDKQdzXyf7h8c+gCxUYaSMddctclEOZWO7B7au
2Qf43nm5KTzaZvqe8yzvCetYKKGT/Hi2U62QUhiM1YSVGrDl/VJhimoAKFmoWkfwDz9wTuvUAZ4r
qBoSsvizBxVmO5dc7shAky6/XGGSFac7YUvmAA7M4NhN7OO/MkbKSqYj0UTpcbQ3pgtLgnr/30DW
7CQPfCJxmNcHiV9V523sPV/j5QOSCjDbBViRlIZqdiN7RyrLRMXZ5R2ADeEHrACsvyKA8+jyk+wk
PsgeNUkfUtBqCytiB7m8o0cpLJBF00aVk/HPFm/z8KG7zVZOjca9dPygOzqAVGA963NjZ22oy1At
xuxt1vGp7WlIORnh9P7DeEqHaFfF1WRX9hrjRY2BVlbquAvvs+O/byBW/zErFNqEUFdeNjl8yD0/
+uw2rUAR8ARNxgOGepXO4BZm+A9DES1q/7QLr5L3TliW76joPuND5DfIZbxrZstREwAuYsCNX8sD
XPW9Eb566u8U1P3zWHP/5CqIAsIqrNVzEAO9eNskaBXFsEvJGnelsRyGVPSjVAJ4CDiUU15Rag5V
vi/a2FWqMTpyhHwgdCfxEbujiJoBiNIy+HkjJkCuwJPo9S7UtUawLLaEsEsX+F4c+PcyKQhanlsj
kraz1HhTtctL+o+2fy+8VLKDdLt+f0RLAO7g+N2IJF4BWHvPaXYYEMu7EsP2eley6gTEOW1hBv9G
ZdiBhFPk97JmH8QDtHWk49zUbiUxY1MmyXa/YPzYWhBRie7HobpsGe0GD5/Sis9RPoLbmOo36z9e
1d1rXaTowy0XPIwBldX2HplEcdp/wEX9IZuaAovfvKmR1AUAV1s9Z1tRRXW+RivpzcQYpag2rcuc
OPRewDxHxarnUXM5HavKbynJXtVQoJzIeFyebVFinHzTjxNCyFB7BY224Tr1wgDKvCdGZLmIPz+w
p/A64xUxxp3xecazs9DSnq9NMEX6y42Uw4ETEHZdv71apsOt0ss5bFng9UvnQNTDOaOE3/Mt/vcq
4ekiSB+IeTw4ABAwXX0ZR5KOONePvUdMCFKsbIJVeqVz+pjIPI8sAkdEP5VRTZzIPgS2jbNJBsPy
KT4bTgQyw+yQ//RBZEioV5lY3xI1b1YBuI+73JJ/kYnNKvZMsGBjKVH0H6rlmtkbxOD3rQvOuo7+
7hhn3CUe8GLV+YosGFMMoYqTmbKHjxpE2UxZ32r3/sDjDCVZcYpugb5O1eSBK64cmwKNWNTUz78p
979tlRvkrNEVBVA5/5nc71Gv5LQgJ+J1tyDA1iThxxZFDv6lVleB0K+cXuAG5EY8OdBCmz+ydBpc
DEZi4SpIpSTt7ZJl74Ckez2UBtGh/Rk7Gg9cSH99CJYkIPqC02Q7kP+Tnvxo2y21fB8tF6SKjqeJ
BZuAFnAFzotlPj0xdcKgyDr1B6ug5T2TP0vBC2vmtCGaqr8+QEAAQpLr0fWt3Rkfr8CNK/ffR+Aq
xW6x5GFr7D0b9CcQMi4q+A/75JNLRmC+jdmBttfeO8zOjfoK2rIFW9D3eLP3GBDjnXjQTkf8gTIx
DncU2AMXSXswW+PpXxfziwQ283cF0UXu2+JlZaXR+iOhYDMO4dDjm0VZknLiubLSEsO0XvlPmmjY
pMnAHxvJY13dbSPQHtxIQC9POPmR5EPWNznqLBdh+aZhQ80qOsHxILQxL5rWUglnCgmJuPVrcFqA
ZVuljNr6SbT4dnzG1xwghqzD85fP4CpYm9qMYKu1SrgF5J08WYJ0/cP6R740X9NAHEQXv7HYlj9W
wpj+Zm/p+RoCsv//7ha+hEcoBpkO+eGBJ83TAJ1veFugvIgACap7ouCKEwKUpA/qM6gpsKl8iExg
uLbuhuBdgCfhjhFHtTP99OmQhH7PdGYLjlAK18mh5SBNDx9fgiAZvWmyCdiPk/LzxQR9Ob6b5T80
pbohjuindw8v29yUlm+UlPUR2GCFrEhrKC+7orwxPmJxWQe/kT2VnZwCg6h27G7iAHjfhOqp8wn6
XN3L/sEdejzMEERNylAqMHfCJ/PlwhRYzK/oDmoljWLIr9Qn4IzvWECjcBV4Pdl9f21vhhyimtbP
ukgKf8XUDa97+fXY8KVhtJGOCBhSxa+OVBe/FN7P7Zdyen3z6MUCaqN8DKMWSaa20pjF9ztaeOY9
a7fMQqwW1ObZs1WdjSsbB91JGLalPEa1AJlq9diRSpj4oWX1tCBCs41nfwEeJFnyqlMDnFo9ZAFe
EcNRau0oDTaBHR9TKQ2u2lrQF9zkkUqXtQer3o7XxtcRJmJMohRmU1YkOlQi4pLObkhcFohY/9Fp
ll00wNPegQBVnghHzqRuh3Fz6MP2JSoAe7p8CMsxXE6c6dAKUHe8foT7as94v7MF7RJsbitnEccb
vsU9YjVpBSqpus0KOv3/sNYm98Jtz1zf1eaWIv5vT8AnL4kFUBfGlirju/jesT3Sfr8RVPpAHgCp
cpMg2MZhtPMwspG4Vpvy/K9HDSX+ILL0C2av0ZpBISgvAV+cLJmGdKvkeRM3300i5fPcXEecwMJ2
/+Z22GJRPsNGkyq75HqLXP9oc+NFBb02K1NmF1NDW6fuStXCymwmvIfzIJRU98i5MGFZb5n6I3Ja
CX4lp+HQnEL3wK/alq9Oceiyci2NUOpZZW8Hg4OXTftNUUrrxywzPc8WRx85sGsp+Sudh35/vCSR
uFWBTUfgn5vMG7H0jIZg+jkWGxZ5LtOGFEKuRSWRnxR1txI+I+4rRXjrrVcolg/q+daVlW4PxmUF
20v9gwio4JSBUf2Ol1bavDtdt5dyzLQ6b7E+Yo+IjGa4AF1XhLrYq92vG4BmU9Ca/pzA3xTB9Zej
5cY1PkBwMHcVLBFJrULMvfOjZJ3xE734C7N+RCN/ZgRkxViOLY6SVswiwx0LBfI4CpnBOk9jUPoJ
XePVr2hk7q2NQ7vgF96AON0HV4cIpx+T2YY+88Q2h/0U6acWmqqmkjwJtzy68gXZWSRfQDO5388b
9XUSWwV7duWQmvh1M40tp44LxDBP73AT7od7dbr1/OCRK9FyxI/RmyvnO7PKhWxJD+7tJ9+2NfrS
4Np7XBUAzGnZMPU7Il6qv+rOTQTgs9XY3aWKYpqWqpFH2VzeyExbg+G9JPXGnuZa237+67hdb1Ch
0BmvUtkjhafXMIRuQk4jX/JgcvsoIKwp8CzEuTwSrK7z+1nQqQuWZtYtdisLqliBVXDfRiVd2I6G
5tpJyvD3mBCctxBw3s0n+228Gph+8qFHe7i+38H2usglrC1CDo0hTru2qtYu5pH51GI4HhF5XE3j
SxUGejZgfvqsxTVOHHqL9QPdAejOZF1OmANk5XvRKKWLPNnfSSQ5YCKlsFzcThi0sPZjFzB2GPtS
R+Or07P7Dytxumat9k6kdnXNuGGt19ukUkXfJ+PIxs9DGdLnDHSaEHxyQq+tzxfvmJAxKWLXewz0
8/fcElilOANsruUvCIhIPSA6227figRtwQlVrV21g0fMCkOXZuiosqesgenCk6/ZNe6aMIRRHBjV
XHAw3HWS/xNOC0dITetmUQjcNu6bdsfgeroUgB0jJgd+GrsYFlT25l3H7XY/rVoWROchuMgjPFY2
rcN+Eur+c7d6SXxnIMms+4QwVXjiWwY0APcCKkp+rA==
`protect end_protected
