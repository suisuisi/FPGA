`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HemXWZ1UPU6e34YfW+rIRo8Hy2Ziurj00hpwa44wIHNePWJG450/5s4zdIVNpkH8+Z6BkUWfCalq
+P25tlG6eA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K+Z69W/c/9IEs1LL6RlQLyeeAjQGCB0EzaTfGXY1sjTDS4A2OjmoXyD7PZjLEeq1Nph9ZW5v4sBp
94l893SR1g/YV3F12/2I+2kkzNLlJV+bSMZg2ApNf6TLP0D/Vhf/ST8XWh6UYvtzyaq9rw/1QWhT
L4Iq+66ZCcse4zL3Bb0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fJbdI8aHi6K56f29tiMeNjcirC+7Ffs5gybM1f6Ufff/G06vfzN3tt7fohm/Nj/Vo6r4oEAZrajC
7cxfY3XpkRw+50NEWmzaCcO0Marql7OpcoJ6gQcXPwPAfFf4ef3oJ2930pSowb7teCNIYVx2z66a
yjBpqIaGcJ6PqSgUS3hvN1/8E8YEH8iHpDrheHG9NA5utEFQQ3RMsM0ndct0kdkY6eHKfHi6w7L3
MmIGsKLTc3aySUYuLMewnX2YA2HZ7pf0YCC+lTDcPqAtGePOSXiV/AKY9dwR0/VLoD1F1/eVEnKZ
/H9Yj5Bk8M6g6eGKyorlodmXxC9FsdDOtFbaCA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Mc2l1cncbeLMzHupYakQfs37H2gMXwgiuj+SuZBpPxyruG4Sxn2JzKUe2tt93EMvK2Z55cqQDagR
FQJVupN7Spnb/L24UFxKdzC3iUwhvq8ofYqvSDXcpBLVhmI+b8qZgt4qEdTQ/m1kGVY1uiSRB+5J
fvIz3ppsjrIl2SEDXG3C7YaNfk5Z2nxreiMy/q11R4u0EpC6TVV8oNGUlU9YGSYVMZfmaUcMHGnI
kIWxyGOudMHtgmNVvnCbBiC0GOqbrOzSYtQXkUIOU6yXal8tvmS1t7I/u/hffiibVvtjYUJtL+Xp
gEoZrfu/tajwPHPGcJrsayYVXeqnKFbWyLqTcw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vxYQLJ79gGJme4iuV9azb0wq5/+6E5ZcW5BtSEo8mnFbuO58vAJGJxdVAw8J0TtALYDxxolUVAPy
6B2kBOu25aW3152OnMvxPnRWfZmOHhaXn8Z7DwdqDi5LDrXEXKddJeKobcXoofw31DpkIl+Ezm4g
6PPmsKwOHx7rWEr6NoVOHzk49JMAZTPXjMzAgrpDrHNvbvvcio2fFlnXeIpLxnKW/MV98XfHbrzM
mzNkKfBPjY+JIIIVOffJ2+lW1jq8gmZP8Ef/Cqe+/IcXBr/TUmnMqhNo4kvZIE6R84ea4RnK2Y+P
EUjqhLNhHSwsw961ETVL0WKafm7fmmtapcHOmQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RpNfQSfnU6lBIefFRktTMg7e5TmBE2V5Au4TKrLs9W9cnqVY+VbcUeoi/jDeaF/rIuZo1QKyFHTz
7gDKl5Z3KwAm5XtW1J0lN/10zQrNx7/eSV8HO4wYyybU3Qt+laOuXQkAR2mh4zg2H2nn0kcgDEZO
um31GOe+NRLdww/6ENY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZxbnzRwGH5k/XAY8QrlGwAEqqUQ4Vb3xAhe1qc1p30qSSE293Mj9hcK8UAsREAz0h7a98iNhLuqE
y3mDaEN+PTQ9+V8uknUfb5SNhhCGYQyqyvcy0GrzoDnD659MiMH02qU2FYlEnFM77rvrksdXKz1k
rIJZfz3vNCnCPaEXnLl4cwfPm7YNCLJT3q3B1JELhtjl48G0IX449EMt/BVGZJ6wo24MaB0UIR0Q
LEfq0HwlBp+QevnEq8aMIL6eayFkTwh6+P1Y4oT/MsPl2HU89qfyPgpfH77652a3gKJxPpLBN4BY
SGGIskUrOBmb7T8oFk5ir4xaaB2tJBr6jk3gjg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175296)
`protect data_block
11+IoC/yWOtZPL0q6rHIcpYKqDxY41DSmgDGDZt8xmcyN2MvdUJsmWepLbIUcCFAZNI0aA2c7lTG
4XA7zMU5AJyO/YBLjXqWGyt1UuUHq8YE94fw0DPgq/jvY7sk+5XiuqCUEhYXcnjv7re39xipOciV
CkPmRVt209B0lARjaAkaQkI9j+9/jqdrKir/sGGRA5hFuTm/XeVUOOYjzluTdUdyA30ujXP7Fo7u
EddqZSsZuid57dqkyj6jS3miHcfq9nEfjx4xtYRrCCgaoyPtff64bQLAxGhiUhi7GvI/1obKZFfS
cvmk7YeUkIt3IZUijHPAeY+rBNhH5SIC4MP8o3C6d24SarOW8MeoPJqQSPxiSzV0ktL/gktvWUnW
XYA4yJLNF5H2vrsiXanUnma52Yj1hEXvUpKYotaazusRmdoFhKfrKAfA1I0reA+pDHLlvaVib59F
Xk7OXF43mnNyuyIc6d7mDpbDBtboAkpRuDkqVS1IOJJ0RfrPgKtpm5E+pC3xzA7EmVervd61YKJE
+H5HThgpd3a7yV7XrgkbDOc36A136QgG/jz1Cbw1tJZVIrEbbc784N3MUfZhQt/B2nzk+TcrUeuX
qGTAplV1xCg31/mWgzMp94fYl7j5fEIycgTp9iOdhwMiXHCqQkRFoPm3i9z5oyQB7gVdyGiigVXq
/P7Z1mElY0wglK+O8s5un3Z/AS+W/e54/IpXBymVcfU11NxJAjIbW3QaTVoiQE1WmdOjrh+n4jYV
wiD7BGdY6migI2pgom73/6w44CQUeRUVJ/LXiDhcesb/TlvcE5rvHuzk5ZYYbG5nrnkZ1vPb6d/u
60h3Lb5RZK+tJyRcdvOA65XjgiE/dWBSa4kWEMZ2YgMDT6pUiaqH6BGP6nz9s+mA4TZl/qJf/Jse
DDWDA03jj68njDv2rVxwzjiSy63zgP7DO34Oe3eXox+E31z3xO34BZkkKH117ab4uew1iaqffNk0
VxhvJm9wBcEIi3Bal0ZDjo7LkoXFVP3FeFzCAvjrXS/2qzazwBLrBKqGl61aPUTVhqUTiUXJEOgD
wk3h87KgJk0gIVJ7AnKB5YO2OZHP8/kRHCdrwSbubVicn++CrMq7xgiTVjxHce0c1YME36HzveUT
hXj3v67X/pKLp5SfpA6RSObdcmLmoQtB9PRC56qdStC4B/4iLtRvQr99JINyTVoGAOcGJnketduP
3MkVOmmS2dv2emn89qVRaE0Y2ABVMhoCud1FiBBVMoOOUQgLX98dK8PL8i0zFFMfPDkVin+uvu+A
2jkmOb9EV/juIfGqxkhhIQlt5CUUsl2kD1uQD62k/pIIsSP3bQ3Npe0EthbdL5AGer1GX6gsikMR
S78X3pgjDL4zurMuSk6aAckz3rhGhA0JuBws30pP46kE0pXsGcxwiw6cFNKYSI3AwciRqJxwyAKH
dTyY2SzExROt+WQkkT1pnavZfjdmGW/02ma0A/D+9Kn8TAhiUm1pWvknhCDVpYBGaMMb7/XaB1BT
vIWsBnFm4zYFxgV0EpxnUiWA/knbYGFS8zCI+7jswAgXkVpckV9nV34PUSXG5sdAdEeDaLgzh3Qt
QUOfTVdRwLomXx3puptlDOuluYHx7JLlCG3xctWWQz2hxRqsFub3+HUA6zgtIKaDay+ldKBMQEPf
YoUkvlMszgyIQUz4kN9/YPGeGhmNrVVh+XGR6u2r3D6SiMH5nKCWJGLq1bwkgN0808L+OXjjIbNw
H6WXpDILbLdDZUM3wvFWdgCpPQqxoLpMcJFT5EjpQk3/sMYAz+AV33CTgKb04UTMhL3WTwZLxVi0
pGg0vB71OrAnllRKxPDnaOjraFZFh/JHReBFUrQezp844s3Q1pKurngzPbwmghKArIt5agB6r5O7
6uNwPXTHvlrcQlae2xg307YIhobE4We4L8KAPoRX5FMabXFd06Au4jLCyvZasmblrrR6Cbfdsw1p
nIjxkSlPBO4MdDVmRXu4UQDV2tIVIRSzsa+ePWit/aee3hSnIJZ13jet1XYuKppoTGo+K6Nydq3h
4JaXWZYiL2C84tAEfGRcMWHS3GoWbS8BYBDWcZvRQ5cDc6/cl1PvAJImSanM09TP7hfujiqeQ1/a
BmwB3sy0m2ESOk++s9B//kmT0VILLFsf6Pejq9S7WkVqftRKqvlcpLAjLzH1GtEovFc/lIbhnxm7
IbsvbLjrPhHAJuac1Dt5JsDjzMhdoKI0M/e0Z9ot+tLrNy8lHVlbmXU7Q5uw4ySzDWRhtJfoq2On
6nH1W3YYDjVO29nuWhZFcnB9e0L9InfPXKMbl3paF5nPyFyrR9fCfafxYR/9sDYPBKFPFaM24MkR
XsWcUgr8Ev920Kmi6FcrFyC59vHSxkhGTjvpW25aVp7OvR8SD9eeF+Te75jmji6Hz84gzVUJf0ju
JjaqvSBea9XcFTeyamkAFd5Ryu63CZOzBzVbnk0uKlyL+U6WKNr+AkOHBUaGpCa7KHmXyCk2scUQ
7rPHLFv5dw9mOfh/pHRJF6Qk9eUecQBuNnIUnp0rJag3SHichm8a1zcddnPTYIF3raeR6VgPJu7W
MV/eAiDfEKp0WAiTopOBqm/0sa7b7WaM8V7Br8QvYwLLa/sddgt0OvwcD2An8V/PSUUbXJbHDCLc
ylEqqhZO+wJquSKydSKh7wvjj/Av0phlX/rCUoT9XKdw8APA/AylMYjC6YpHf/iabswepMPl+4o6
Wfs8YOxRPxUy44s/7lPUvfSSqtxsi3TY/T1ofzhgTsCubDrWsbqAiRQrdrfYoVHFAp9ua4FD+n2B
TKLLfU9vkn5hmDkYubum2NCoifau2q7ZH48gQRUA3Z89yuxRUVQaN9f7CqhJsI8keLjYmVPT/Wk8
o2XoSTTSSUleabvOO18mxckNO1Yu1MRWnWXqksFIdIsCz7TS4ZSuh15u0CpAQoW/+vQVY7b/9aP6
p3WjW0z9Ltciz01xWhVOQqioB5nA5UDDqcaJAZQqy9IgiJOiVLMhosQeYHX0pvLp0IbJiWjyrTA7
Gg1H8Z1EhjwWwSp282hnXGqeIFHu7kNyPtk98DZo9ZsTz2xIs1HsjX97Se+EvfbAvILkTRInIuzF
c3EwuLqjLKsRsdbGBNkqOcxSYE6gH3naK6wTZXsBmmP/0h8ICe4+PgzDXvTLCLvodQUOu8TyH1vl
oyJ96g0JHaZ4PtIGoS7AtqX5j/1XYkj6ciAhAthcyf/KsU/1TTE/2NcXN9euKWBmqq3r6B2WXaGv
0m2/Xlvxje4dKWhL75n6nnXRsMQgZTFnIvvzdBnT8CDcU23lOUYWerQgDHjsFxrEXHbKjbAG4bRv
J0AQekLbym9FbMX5e6RujVFX1MYTkRQDtC3jnd5K5jZaVzENGURlXKnf73LeqjsUy3G0aHFKZOqm
1CqpHaSoiECPPn3qATCac07WX7RMW3a+HYjeZ+JYBomSh0z9ci+Uc/OcDO44+jXdbpJ4lW5r6hXp
NyruyDwbnOoGzqO5IvOueOeJLLxcWqelIp87YHHTo7aFI/qj6eKWBdSmmQRM5z+X/8izwhY2MCqq
qjdbAIoLJqsTaXxnETzzmNXgAlaSniRBxEX/OvGSaFkSSQ8hLnRaXqifVTjObn/6/M+b5HLo8o1V
drb5LTaAdKUdab5pUio1j9Aju4BQuXjlgROAnsvAuhe5aJ4b8tic97piUamnPPpnZ5zuw5a80Ytc
rhcvdi7LsjDx3Zyg+hM75YAZZa8tMpwN7dO+MWOWVwzbB4Eovh/Wf22HGz4dg9EH7icz4hmjTFnm
WcnQcKCV77rZ//6v0ZQiBZfPVDp0EVokeryiO4UedgqcMir9pMtgwJaK5GcdO8gjo3dcKSeZBi5Y
hN5n3qZ1LAbSY9p1ZnHrjm/ru6R7zpNJmsscv/uU1I1Y/1C9KM+dRHyRGcTRWcUOp2ILdyeaWPI/
jDt9di4M2zj/1Yp8s1aJsqaKLIrqFcuTmndKH3Z0SVo+HzEQs7U5dxHGwQKteh7pARQNDDs3NUVm
ThOvbtAJ+OiH3bf6TkioNhk6g8MtOYErUv0w3sLlYEnxOmzJtmO+4vVbPYwPsimqxAMZzIyje9Yg
eP9oqU+EvuSl55XP3hAhkMv2sw4NtKftmmMflomhH4veIFGRmta3zopgYwpMvGubqXC+UWymKCrH
+KwrQXifDWH3iDhJQuM9EOMMstaUUPW4kHBk9gJKwqpBTnioZupienrPzOaT4LFRtWYMG1E4ocGa
4brE9BVTyKUNcNKaNwcBQ2E+YxZrcr6SbQp6pbEtXSAcHu+5IiZRHi5XVnXats4QlV27Breya7Z1
xfDq3ounBVH+lSETYZWfhea0+jmdYG4/9GmuFjJF4nFArqEEm6uTLgzcTDd3hZ5D9K8p+6iJ7YiR
bN7kL7I6V4uGxggbxNTltkkNi3I6h8I5CmUPdZ/pZ7JWeMeI9l06lR3IXFfXz3KegpxGUjvd7VHf
YC5FBkmdCyhCakC9MNWWGJrWE37lTLbwbXkQRc2nXImfl8MqJ733ZQ6yDxUwz405XI2oOuPK6w04
U/y9qPmv53JjeJA6LhrHDppxhQzceCRTqIYF7pIz2eGiLxA6o5m5x2MO6R6pVj4CrWssJcBzVmXS
MAYM+rrr78WZcqJND1CFtSA9Lum8K/AIOXIzT4INSPIKzIP2x1x5r9TNPtBam002b6Sen3Gbmvx4
UtXtBQhqd8SU2RewV2QrCj62JuzcJ763jXFhYVjsAuXCnnI0K9XaqYuggl+pBlfCywMBd9NMuPkQ
rApw4S1H2AbRyJrHA4FaMjc5QnjWKLsKW3OPP+DsNypBa57NLerpBCdFZZkRkQPkRRVIdt3OYkqk
t9Vtn8VXhmcENYwhPBanfAN+6PgWD7k/LQKbsh/n4SE+Jk1K2swfzsOkYz+qzdg5E1ILY+/t9JP4
t4nyqHvmyRQ2SMDDSVFF0uuDpQEv5wHzawPI68PJaQmAqQ9cecLo9KlMDQWxGGfhOtfGC/Sbefds
jGyKE+YsbTn3G7wHzOyEOkrRmRdJyHYEIsAn5z3d5kuEQGEZ1Ula8XLRlpCIuympWyV91G+UwSkA
Vm2Tr0eVXsFIkrE4QYke3FsFiUJQ57DaxPGpRBgEQo1KNAsB9+d1ePvb9cVXUysrJRq1k8CJeQHt
eeLskJcdxSoZU07sl47Lcs4l1mjve5kebnFHfBjqclvL3HqOuMoBXSrcaim8Boc0OJeCTHMcpHg8
WX9gwqR0QAzNJQtjwacGt2FULfMBd0wZLvHsQfyfYmhoibkmZ/I1zmovQot8isQehbpMs5xJEUCM
GQR/3GckIAAOOvhoC+7mXRgAuXqYf19Qg7SPV1KTTrquOnCYAdUCpQHiA+SxugxPiEdaZtOzXZSD
3M4qYr1uc9ao2Se/RVyUDRBAQXhylgXnvqeWmx9IuojtRu0n9mK85K3gheCpyFOfJPzlZOn6KAFo
duvfrfYJ8vIhWP1f+H4FrUjg3MnevU0WR6wWzYVNsLBAG9xL0GDb+aCTQvELfDAXw3nYLabKQQGy
LwRpj07b2GlNbCMdLAJVppD7JBNxkyF2abzg01iUrtPB11rO8Na05UdP1wvWnm38Jkc4B+p6ap+8
xRQ2JbmRuigB/OtgNhkaoDJmqEfUxZyOtzjRF2bZKHCpT453aN5siMe8K3xrjDJxQ1FLc4/MmFm1
uvqcB9pCedqgXRYHdqGSlQnXN0lcWEqIsztsfK/H3Ws88rdesCkFZpEI6a9MOELTUXEOBaNUfy4u
pv4oOWD4QFq5wjJNGKcjnjg5vvN7V4mVqlRby6AiPNzANg8XAQQ+ozW846JBDKp4YH42Z9gKNm6m
qZndmlGP9hBMrsOnZT7pTQfJTmWpobuaV0Ad/9Wsn+q+yMlomQDFmS+htlJlH5u1+qimvDvad2HF
pu+NkNuzSuZcC/AWFFeJTk411TpmKvHdk+gqAicsiuF7DfVkY9Mq0ikMDnQCxYMZdeEbYStiN3r5
BfyYIcWbhFY6nYRBy06sBrRMsQkyZPN9W2SssfdFAJc91LPBWo1futplYUv9c1atFX2yo2vOUFWq
SAVxBtNooN29PKk8OjbDnzFduLsMpVuD9B/OgfYcYHgvyc7WxsV0wLGfSxxRIgzaGw5RhSr20rnm
hXmkgUVzA3Zuudn8lkf8fORH91ZTOhkyzxaSaeDkgvW4KGZnFADJJuDJUrEHDyO2lj76x1hH1Ozp
PTjYbv7CLohuyHund16LvlPkNWYK0Q5yVbnYer6mpEEsbAeX2GOnbiwad3DXtR2iYNIQ9pm5Opag
HSzIQxijgw99ZWaVAXSjIDnGeUvKTuZGBnNJBosmWMIBjhPdhqzbQhbuGa0+6t9+17CI4WLCDdoZ
Z4rMjtyUT6h/7jXSr0unxEqeovupxHRKaTDxf6/5/M77VqsF3odToWUmI2F6I+CNzcCPbKIfSbG2
1YcyITk8NlIXihHK4y/Th1t+MKCwcMmonT3P5LQwwlCIP5Peril2dNVP5YsHCqPhXj8ezudv2Uek
2pewiIJLmnFeFSUdVBMyTffDWMp/71Mmi9yCRla3RpH1MVWsOKSk+EJ72jae2ruwCJtr2r5bbP1V
4PXUEWqauNNtbjmhQRlzDBHhxuo/YWLhPB8PJE5PYun4V1gmWnzG9s3daAZadn+cAPK3Uvf8EtoS
GCkgrP7FNCaP57PJT3defPXpL3pxjHO5M6DrOCo/hrN3lwVzMXwQ4GGrDbr85pFh1wvfxJ8fA+Wq
+QkGXj+MyPKJskMga+Yxg3SMxpLwcpSAnuFOFBZw6slqC/7k65SHz70r85KzdRfNva0DKI9OoLs7
3v4RIS5UxcUCwnAXEBC8L90ykFTmhLZEYVWIFjl2MnOD4QMzYdSHuJtaHN59Le9EXoF9+jEKy4UT
iApiBnvPPfNyD9RpJwDwZlj4WyeU52byaHxNjq91fm5a8zYz5Pa/2MbWMjpVCZiedueIDMhFrMhH
3lvhW5xOpRErdPSK3yIUkW/P/yLoGDtqqfFwrG7uyMYXQTU+WtLUSMV+OAOMOXuLb77rQLxd5tCR
zzpCoqqz7GTQxlzv6dT6Wfhx9VjVaxI1eT7/bS2sTbLqSoU1lSINiuZpO+/MnjXjouKTzVE3jOk/
RsBT+AS5DWR8h3+NqVmaRy01QMnAIqefqI3XeIEHlXLtHCFo4+txy5fykLzsYM5ZsDQXkjqDUFBz
kqPSaBcvzKj399xCxYBqi+k/CSJW7jeMJBCAMkeF/Hv4+oIKsKJeEqeCGcAGnWJsrLH8uizhLrLN
W3GqylLwt6m9YnmbkF4tF3C8c1RGXeJgfEafPdS/n/Q/Np67x6P3wI1wUmqt6N+U0jcPGXFK8lQi
jY9pVu+Ra9GPDKmA2YtbJtV8/gXJASxlCN6aSWSAA13tVoMbRPsh3el5+NdfHl2p0F3RZ5XYDbf/
pmFwv9DajA3FgAtCEKAC7Af4rhjM5yWTM+EyInNchqNb+Q8mKnctz1sJx+elyNMzSOvHweJbX4zw
lBpHacEKAD7e4wHxFbqgQQUU3RhtScvO8ffoSVPJqaTVowRAPCR2Wj5Pphj0sk8Sm/i9Yd5K+93M
s1ho4LSMmMcViPjDS1WcEKU5uxOLDftLwvQFh+1U/Xg3P6gtCHBdeT5/XW0l6+Nu/1BkxN8TE8w/
wIsCNbMcdAS0oJGGPK1hZtxZcvT0e2SQ0YP9aRfadJ2rKjohLLEillLUqJXNrm8ys7DEUHapLn1W
cX5YH8mqlW+HEDLCWiB2ogqKmavGKjmVgITwd7fdr6WqUx6xFemWNC/yzZ08r4SbEX+aTxgZVSYS
0bfcjYh1zzLiS7sjm3pt3TyIY9m7XvXhrr3koMC8R62dPs+JBywTqf2kzQVxaTrRPu+jn2W4TZrQ
tvz4M17l5nNjt5zlrkVAA3BX+mnXHR6NWjRI9k1tq4THZFKDo1WInGl2HZKguz7X9HxZXl+54w8F
x3dN4W8evZTz20HgqLmsp+SSYoGg6s64w9gki7tkvvTDtjzB8xQlvnok9jh/w7m1hEzRCjeFu3nQ
i43ercKMEoOEXjWcLma+oke2z+0rAigrZeBjWZO08gTAPrRs0UfaTPdmDkR2pb4BuiI+IU6nlBro
HPvUh61Y4Xw+9dnsUkVhIuf5EP+tG8tFnQjBvT/V7TAzi6rdsVos+C06vyS6ikeKWyAB/ImK+Ucm
cm9wlIVTnNHZkPqBdYSnC/B0vgs0cnMRNqlIlymNVVT1rfCu6MwkffBijO/EQmbbpol2DzkuG6Y7
hUfe4K1/tdtJBmsaKBYQvNwQYPMcm1+HwycRn6Rc6yOAnzt5USETzr+mmUY5tnxRZyuaPD3wiqjj
k4IZlFpvwZIqM7ML3SO+oYj2rNY3kbAxIxq+LfRQIGiknY4LT/gp2cgOG1pjMDZEza8z0QUqh57p
kGNobJzYTtCETjNSpzSKPjUeAtX/bctNYQIUlGDmmvc7IDpTuHxSArWlq2MFmdD9f2iM/mCPiPOm
uiZM9V9HegOkh3nYRl19SgbV1BxFuWP0816LTfaJ+Q7MKvlLbHlHy5ptWSxw8iiPsovrnjMy89pp
xovYKxbO1yVos8DEBTWvZ8ZWSpkT9Pckwm2KqWa9sPvdbaZxGC98eXzbRysQneVn8XoRid4FsPb2
ENHHc5a1Gn4uLOZczOZ7A/pOBhlcqhy+8qHk4U1piWcyqpBxszYYQRrVm/07uYEW+w4/M6fKbqSa
2ZT4h1oQnxdeL2zKOUmQx9Y4MR7ij4dS/KtofbpTU2c8gp0vYnCEuqPTBawikTlQbG/XneG3mjL2
K3nV/iQNRGvpQozARYUn/ApGRWOmPc/ivUU9aoTNvk3p9pbzuxTe8JcH+Wj1iY/Uo5zFqsNY1pcP
gOoS11F/716aEZguXw7z5yGBlB2IAqxw8tMClWqA/tIZS3AtA6i3iFFYrZHoVCHd+xLvw3ePuajB
1jdMXlhy/Tw/0TJtuA6T5NkuwVI7BgGpH9fWLvI6L97JK+2fZccyWLG53DAx/IMofkcwoVaU/8vk
Mah31ryMU6b0OC764Nnij8/46qguD65+EmSY3JTax058C/IpW9neT+BxyojcVNjEx3CUDYcyncYC
ml3/ueZeRarkM4Fo87op+8JNlywYLWc1B/ihdxwz1E6hxXC+YsabfcWoQ+11Yx1LHluHCVgiP/Hr
U6UeHfN8xPpMBZPH0f5VH0tvh411plcTXeJiLfc+s2kKGZLzkaNCbucKhVsisrooZSasuPoE5smI
QO1jJFEatycJZtzYzP0N9X9557fju68M/rttVsiaoMtN+riOcuz1ldvuqqN1FjVqbQ8UKCPQW4dD
GirMJ046ByAHyhESGcROuL56H/894RdYBWR9++BnIsiDxzqxEqaLkac4xNf0TM7ZY+XO78jKr9xp
uiCWJ+qGmUaAs0XvtFnFd9RakUJG/mmKp7hHSSe8yCVRgGLNVCLNTtVUxCSFXOViun4RGWDPVxxp
wwz59zjdVMLH1QzHyQ6LKwsWrm7k4w3+Ie41yAO2/ga+tIXODPsvo34SzTUkjty+urFrcK91X6R1
uxW0k0aC7ZHgUGcEh53pOLgXRmdYSMViGRoIiwPQr91TDKhZ3+EE/stbbaq3zQTMwBbof6PvUpOE
PrSib3XiLoGSA8Xp1/SptmFlMHyX2/ojegT/9DVBv0BWJCxQyUijwfCTTf4Tou4DyrtXYmfaAXiG
4XOben3mBCKQ2iyVBArkKtBp7dD3JBVa5ZTUZpSnPNHjBpNFv7v//JU8xmHylzvK002/OfQ+hoYS
LhrOO0g72OTIz8RAlXTk6HXx4XBW/DmnEeUMDQPIO6LheELJ9zfwkLzRmPZjtUH6K+U1/wUs7vRv
cnK8E6jNb6a+h8iZALR1iGMqYNFAfotgwrCsoeH/iwtejsDeTFAoIQMUh01UCgfJqBvjRk9Pf0Ad
lL7lHrIatY/Cn9P63/b1V76iNoVwLWX/9tlvGykXmbzbOQpsqxQiymhnDqmh+lDZyn/+5N9KL3IF
f+v7rNvb1YyFr3wHVtbj0EIL4ryACFSZxf6pVzSvCjqSPH6qzxwtl5ehub9yhKSFV0giDVWcKjJ1
L6LFutCJMAMXEO1iTeOLAHApdKkzWHjKEGKBdlYloEQctbqZcEEIg8szb1biHu0A2utjvHRQKi/o
jyTl2n7rRo75nmZbzA7z2sr133XDwWb05TOR0ugVq5L6Ggb1WnieGfUgB0x6mvcm48lWnh4bOEQW
9Jr1AGKCrt5a8ftr6/Ozxlxz6v5z5iZv/+gQF9SAy8VNq7C2BAFkBM95UoxPVF0oEtiSt3XlcbIs
e4JvZj36H35pHLKTsanWwxxzfrWyVYzIaoR9YCc5taKInWb4iK2NVHTVsvbWrndVW2Z6E+PiqAeY
rbefmf3HoT1Wk/eIEotdBsb3r8FDWTLlz5XV9NBWzqROUbTqZ59Q9OFia7yoZGL/ZqWz8iJZ6hUv
6QRsD3mEyBBuygP+osgATkbaUCpV7o6Sdszu4Ot1Zm6AjJqnSn9tZHFYxwnI2oLbNZM6q0c6/aUE
YBSkfr+Lq5JLSVR7PXVzoW4/9XLAw+5TW1nJ7P1LqXG/SN+Qtm+sbukPxHPhdoD9ME4UBYVAWHJb
8/n0A5914aeGQCUk8wIaWVR8+0bTqzT2Q2T8Vv3meM3Yyf9nqzfGmv7ybIhhaKh1OwAdq22+9VFH
wxJlb0Dol1/NXpISI7im4nwicIHCGHMOhAm78qza9i06axpTfPNtkAjgn5fKB4cKJit5gYUD+DjH
RCgWE+xq6+iaPwaP8GgCC5ahYq/+ZEOw2OujRJW4jXn1kKkii6b7tsqL5ikjsmZ3BzUyJymfh5DL
z+nTqC/BM/i4TaPcnf05FQDlD/8lsaOlp+EZ/8stHxbAe875ugbsGIO5Y6bdgmleN5tHsv1Nwgvl
YsffPfcd/WDyzzLx/+vv00xlraif8hyFvWTGqBNohxdEflRVoZUG1gXr2+4il/H83CQiAz+kY0bP
jniomzOwFiVSwfrstMQvLRWX9dIlTFtz708xyiscLj2mab71B9YsJBUT22SIgZNSQwXboAefmPYg
eIwL7BI7gjvS8q/uMhJN+nIZIPMHURjHBEVsXWuVE1joIGs+L/1sj9j9iA5ZvEqs7o6UU1iIgOu+
WAbmfEnzU46Feklxwa5Wc64Kb9Xy8s37BBiK8iKjsqCVr/4t4YXElWlYL8MefB8rJeC8cGjuqNEl
mE+5Rr3iyT6IhiRHG4tz4PK/nJayUdZWoYbgQck9SWLmDtTgNyUqZYt66jJwxLfWzCOvPpBD10O7
h9uqDt3mHjfwbolvksFcFNI/yWFXWQES3AA99DSSXP4/gg1IPBmLXbBojssntlHXnunp29qpr+Vl
+eT2hPHzwoVmJBMiRptt/pMsRbOYo3e0X5szWs/2vk5zFTQdgd5IVl6UkHdQlYdNBXRwFWJtlPBc
sj2cxuFmPDc7SJzQB0AdgfTmCkVcjAccc0HDkqmmuDIEE0bh6cDEPbDd74XnJFNZ9ThDtTyoQ10P
kSL+/v3aGo6zHOIkP6dN+4asmQyfJ6iyePD5jEbbPH/m5EN+H6mBJ4AJQrhdOfYZW1vt+SxTus9m
N+eMqLyPcQ6KflAksiEPbLslY1rCKWb/t7l8AG59jurcnTSTR7Gs01j2jAruzfF/kYKL9CALvMvB
F1bdVXUe7n9tbEHqoICelyd+22ku1/s8CflTvlvUk5iSWRggkujSjHUK3HnKMpZ3MdrEooGbID4O
YX5tWOyAluu2zhYex0zaKVKqxHadZugqHEt6TlQ/+cVJ3PpfJwDNLQ4bx75s+gb707ncLioDQC4K
L9jXKfSyhSAe+UMxmUZHKg+jaHX8OKpKZdIFIQzdyd48Wx/5Uxg9MF7MoS7p1AX/E3LskyFI1JnA
jOMmZ75utEk9UjxxzWQCI018hOC/UIUsJUUZmCIq8RPwK3xZ1YXCd3eZ+9LNSN68gfDFyYXakg3G
3OoK63EQwSUCqMsqzqlUuO/TXMcEbFGYkpGRVRm+kHN9dZ+yZ6fGE1vMi9B1TUQeGy9+bVpR70bO
MQ5uomXTcIIR81vAFx7Z39Fdb25dRY6ju4B8OKs6jXs8TFnWgEYK8rF3nYiaqUsdfCqCWK73qdWg
bnFdyGC7a0CKu1O+i5WqPL0q247dAn3RApk1NPDWw06MyYg6UL1Z3P9O3RjZ0krEcPtsNqMVGXvN
CUjZDGbDx1jRtQTQodJ3aYNT2tehG4/syuMbgPebXo+rZdEYPhwaU/XpvI5G+lv1ZdlYtedQH6Ip
kQa7uXEjnEGfHS2RKwS1fKDDaE8udCH4i7+8CMT2Cn7atfLg3Dx2apOXrQ8ENYP8oaRo02ccAr7C
NeZGceHGQ6uyS0xVjfnR1Y3rCMWEJkMG2fMY8Ff7h/cWix92T3D2/B9qHWfC7O2xLovEJC5r8WMx
xrEP1WSf33EjZpDoKvO3Ma0ycva0VqyMggPypyNO+6jndh4sdp1yvaNVim2RyqtlnzR24mlrfejS
ZdxrYtSyNDezAOJp73nECfZqkwFr8Hl41h5bBg6/r9z30yAI+ofRSxQonlWvzlB7NPL3nbqHQ+0N
ulnM6emAzGhuyQHY9qtKrI5QLZ3q7mP24yR93NK07KixYbDox3wwVT5ZubMRQFlVsTWYOkKg19dk
4ssf8F5/A/2FlkacX8u0QRvTRnIbt9c5yh1hxMkj7Kvuk1trLhIVs8jt5gmrlEfQPhyKI4rnlCQm
z3X4xAbuM++JAYpyQsKqMynVeEFHQoPPqgIhpmcRI9mZLysFyJnVynC0OHPqfkwMAn6gC9GTm3tB
RDemIF7ZLU3qgblFVLeUW1H/imIeOBEj+96UjW9DZ/3TJ5J+TyOMfMG9uPhQpwCO8fGRXK61JEFx
fFW8vReZ9arRL05AbIzlxkjmv5poI3A6+7sXk6ZZ3efN6vdE5HbtzfJmiKIo2ZnSLd9GaIPYEJqm
yaUqsU+ONq3Sa1e9mOEQY7AS/+9dXCPlTcZjCCpyh/jQEBeRSvo3DUb1HM44EnCoA8z894ryWG9U
pF8qnVpcOoeyNtUp3Ty6oixrjtHw3VZzBn540O05xoXaqdIZhpCJZtw8uhADRny4D4iYqIVQe9Oc
Wu9ugqg1un9CeEZqD82gO+F1t3AOsa8IgjHvDIycB9GekHMGWpJMzDDlHOQwFZZeD7Wd5rXkMmn/
doPlkK8aTCztoojUtY6aZUiECFYZQrAzj/W+5m0y+GawiYPTfSTL+d0Bccio9f1Cu2QtT+RDYh80
Qc9WbG9SOSrTsFGCnbfeis36UWpHO763asTfmbaC9E9UZWSooMlP0fST0KCsbebBokeZADrebmnP
+f8gze2egqblpgW7UFLZt6ww7sBwsV/O9tjO9MS6adxOa98grZC5q9q/dUfOVvmAIR003dtTpzhy
lFj75KJ4+kjV0uPP/PaaPeFHgP4HoceAsyQzMLvfcgQGnxOMjJ2vZ8V8dyG9D3bajt4mFhV6C0MC
ajQaRvvaW5RorDzcPaN9WdTpmLhejLkScXWqDgRrhuZn/fE6C/B3RBgS6Qyru8qa0KoawQk2W5NP
gPrk/TRH/OJM1v5g0gDqHpjpchxEqITDYKmcRAqtEkKInr3oHq6kqJqOMJMkVsk09bi5cymSzkii
jzubDzytdF3Lm3oItV/JFExT8rOzkBYW01bjY/oQRadHPNGcKnCTgc1MiRgp20zC9j0/mtqLCwQV
gdTjm3FI7xjbJfbu6lOy4C7DMIC4co6w8bdGc2hC0ePZ9Eg5LpnpytaoViPfBTCOY9MabMAe9tLT
ifzo2iiBb1lFpieKBw9sUXvcpeW9zUKyxU4qJ1orIkcWpFK1wBNsRu3KmclcK0XBTLcX2Te+yGNQ
9cC59iRHC1ykwzEX2l159h5UKDy/K86UOKVw1poIMPSpokBES0cCRAgEuFJNr0K12t0J6/5zXL4S
AUqyzmM8hmSeVPfgyU8zpSXT0dQyy2CLHPqz0lu6q0DS0IwYMt+C8+Ql6+DW9UpC0xmB1QKLkbg9
3rHZVVcTlQx78n4ptIZwZjCWAuCI/XlWqvPyeRfIeFqimRZwXqD+FsXJkNYMpqGSeR4pvS5jZLGh
uyWUn6VWfdQiGXrxuM8nO2RpNQMfXXJCgJhtayrBpowCCecJjU/llCxjNQHMjP4DkRC1GrPbsWlC
r49wbwLQLkGIRQvF4/uxoawig5IeVtDDbTAa+uRNg+w43uhmmHNVvxZVdOtriknHoyITKnHWjPYw
lGYVq/YZCYdZI/axXpQ5m8P56qK6N/QwpIOUvIKFreF5DHM7wFSZFBP8i6BiFTG/YLKlCmBwhQpZ
v02dm1I3neMRq/XerZ8l4ICWwWCNqk7rHdk7xQyQsDNMzHMUnDRO3ZxyFR4pKrkIhCh9X7ksBTWi
ivVlZv4BOHRiSiJOuRmmsYCx+/gYOCLJGxAd/tcdT587aBkUsTu0FynQS4vv1GiAPiGpHN/KQvmo
41qtDIZ/5fyGCC3DSLwW/Jdr4j8GJ/f+/ZPqX3FBi2wNJAeV0i7Oq+iwxGKF4mhyfR5vROSZqN27
Fczn7s8UKaPHK8okq339DzLYJdy3mlzYiTPqTUBOJhKQSkb3ey6PpJgphtMg7ym62cND10ILkOa9
XbTzw3jMnsvyKy+5/CYvEtgb//VPR7nHaiihiAXf9wEn01/aNP06pEwjOTz2UcxDQNrtSxlxBmdt
Ngyn0lfA8TWnqijMFjfJD+ToVkmVhmOTJ8mMpqKh9fpifmW3zEtGs3i3tr99CuD1EWdc8s1+pxCu
7o7ZrSBjBi2r+10qYpXN57ddxUhuVgORX1OcFj9msiFQr4GE8VDoqOGemYWUg6xh0NqJExnHX0aq
8uyI/2iFqCXgtTQ5bTjjAqvi0+5wZWcbS9YitoO090CKsF+SvYRm6pPtR4iffVeffOAF4Kh9/YQ8
VNGWO0VcDJrl7j4Ov2Eof6HV92q6d5c/AIsAMK8inP6PQ3LIc9ILKreE+MrKmKcxEwPFYBcmw9Pe
DQpqTNpnCIvhDz2SFtSQsYmSo9AjJk7F2miZbSX5C8ZPIVVbnf2FEFu32I0umIRQov1mty6Ds5cD
/jmkh+Y/vm9B3BFc9vVZYtCdCWB45z0KVXD9F9BjkGrwXsW8DJTk/YAYV9X/99ihyqp+W9AkmokI
rKksL8LT7FTlA2V1+lFuTsi3ZVLiSsJqXZoQFJ1DSz+1bY6JoQLURJe3vOYuO1nKjZekz5d4t0SJ
MEnka4jT/ERQ4S5oUttw4+FLPRGp6SKyOU70YNYDnXJL80kJGF+82JopKdUR1IGzDdzx93zqoAix
Yci9QmTRNrr5ZKWjEwqqbRVgNK88md5mSCoLW0tuD8MuvmvHrmAA1ya7M9FtsH7fCyU5teDp8Dnf
Ec4fAM0uOrETExzWV/5/ehIY184U6ENuLCuBndcH7CI9cuFflNi253VWaIgFG1YENgr0HLehNlvY
Z0RDHUIRsr3GesXD/1ndlV8SuWwFTgIIRRa4PoXKJ7bVn4vUZnMc58JY3uormsxbqIk9lUzql5Hc
5j9jVd2T/8SVdoO4O09E0DmRSXWxqeg9jQfNLrl0jwO6709AlnjwspbKCM4wQG67zBpqTRikqhdN
toOnPEP0wHOtH3hqdpcEgtFTpUdWTs64PcB/2sGcG4KJHsWzJS+OI7f3DCsF4HyblLeSmEllav15
1SDjNV5hc8aBGEjU2Q3EcTyEArtOo+GZFTtacZ4wW/pcD/wulfHBMjwqa/nr0uNzXOdrjvpBJj9Z
4exB54yNVe4+6//OLS7nF2QBxhMZgS6hDDQUhRZhtyuKYvMr5uX0jz2NDpUKyNHxdwDttIPm1bq6
EBvdOYkIG2S5ffhr+MHxOCdc7jPwCwVja7MeRVknzgbV6hnLgv8knaXIPOpFvUkUUXtAW92MWTPi
ukZHJ9KY7HZx6MPgsSRs+2jgoRmdKSDBY3JF5wlfhi26QrHCwTy8hJkrJfs5F7Sc8v9MLs/Vz4cg
itCyz72a4fjCQWbl2n274Wf/rm6z+kyJ44YinAot5fFem5kukGcl0X/C8lKiVDZpi88y++G8VfaJ
ZE3ckSaDozO3SPQEOKYD0MlHxovz9+wyAha5pKmKSrzO+i/u0KzXIzZ4No5TLdBUWXaePOSIlGOH
pFLHkav+pWn248M6BtU1jeN+946G3svlHX0P6p6u5LFxokw81tMwlZHAR20KzsDXdIQVxt6yoZks
wftCDhfhqu4CsztCTrwX7c8ScKvbc48ssHMt1DYRaQIROQwsuGgyT/Rm+LVyA0ISiWZ/27mvxwHt
S7gLqrCV1HLzdjFmnKUvUv0BmAT+/8kEOVK+mxNIpe6ctZy/e7CKAKxnC3Cjx6TJn0RH5aH+ahuz
jRNIU5X5tv6Q6T7MI4E6Ns84wwhO0rUufIy9Iz92mZ6orPovzCwuBr5DJax263cd3JryFh6146Du
8Ascq+rDQGHQmVpio1C81cDhwZaJHXYlGs1ox22POW8KHD+mek97IE0s7ewQdobkdW5Kd1BFU3FO
YKWyApwuYjXVaeA+beB4EsdTfWrSJ9UbvOG/KMYYJL6OhvDJaXxbIaw488EuqzySvKvtaQak+mNj
krabivg5ujhIXauSuyVK+Gkx0G0wQ3HZxmQZw5SCXbVQqfJiByk0498cxMa4X9pcjgUWqza/rE7v
o2AWHSv+YSUetW7SzO0LcqeDRQ5P9wcgnmqAZLKLzB4/lnbjMgP0mV7jx6U5KnTzxCNQW/DQbt16
PU1/2Fx7s94YeBCWcI5ofZMEFFsodlJdu4gL3Uk0rU0GDw+e3lCPZr9NMjVrK08PTppqLwzsHhbS
MN4IYN6Y1iCzH+rl8VxYts5rHcaij5p23k+1jsuMrOjbMX5IFAyoa3BEQVitoflbK45PcaMWxB0A
QfFtfmT6cy6szKzpLVcJN4jVSLdkzTP9NeXOCG9iohO1PRK9wrAHTclV6b59Vc3m0CnwqE8VQgVY
N2StSyVvxaK3pZM3M/XpiaZ08HD32LFDLzEbYqE0apPUtAlweReAc6BQ9BlVtub/PQT9uksMeiHW
lyiB1QEJSxMx/Tm+Muh1bZTnxepi51tFjneaLVUxfkHNNN+z5fdakFlwP2/JZS7ft+dEdeFzUADa
0FbDthUQXmQhk3tMyf2o8w+dxAmbLHgcMVCKNMG2cXwi2AqY6Qt0MnZ8MIdXQwyMWVp3p2TziEIi
viLKmG/E9ZzeoNH8WVJd8m2quSgc7BuzbabuPHs9EKWA4MeNjXdzWmr8iCG5Zlw7sKc1M5bldZtS
trkOKMQEfyWw8kToGmhN3zj9ilL1LlmsG+/9T+A0NjL0C3cdx1BG/P3PBjnn3RcnhmvAfVG64qpr
G7t8Ra24Q32EzEMTbzQJuk1pxZPQ4ikTX3Iq9SLiKaCe7Mzmpu7XF7JCT/psUXzRavKi/Oy+K35D
zkpdHY4VH5nGM8JTn3wJ70p1hVLLfuDkDcN6We4SzO9SV5Ac+DliyY19MK1uBr4BTNv6Vr6sTpnk
/vOfVCT7ohqo+MdWH7p1LjfOmZB+t/32EL3fnvy0NeyCOGy86aTVv8xssxVBjCcEKlJ7f+OFXDut
ORKKKvaC0sbz/bw/eTVE3W1/Z+6LrYEieFkVMfsb2CZgCVsARd5W4xfgJYsVBIe80bKc4Mf3P8mN
Sc1HWIAuGEyk/pVTizS4KQzmjEVcCQOKmZKGxZmX0buwbRLqAU/CH3m6rf4aw7zCJEu2TU60KKeE
SQlCzcHkFLHJIJ3qm4hDYqcG/6/Byw8z5LQG2/Ki0joIyX41+ZtPNIsZnOjv1X5UJO0htEuKsYol
kLXOmFgo783VxJAFAfoWurkCZ3qG915MYISoAyZsfuMJspJXnNRn+NoWAghX7Mv7p1FdJcErm6vp
dKsST/taWNRUWh/8dfpN2DSwvaZtcLnkl9N2kyCQoHa7QaEs5+Gfr4p3xwXht21tKrWJEKUqB2b2
RQKw6xzpTIMmwb0UpD3o6H4JFGwfdlCq2ubgCSlmA1k4hRic4CLNmJRW3jx/2J3RZ0Vxr0cPMmbP
ko2FNG+YYRYYf+qPqT09TyYc7H3fP+vufxI0duxAh+1pELH3PLAdxctdxpug66QPexFZlwJODAgH
MWlfRP6QiS7uFT6xEwta5SFFexeMObynTUP+zcU8BGJfCzV5UqCeH4qVTFgyJQMZYoFg9WhWGnGm
zK6E8gB8JemvFTDyJZ/KRmITzc4XW0y9yZpc6x0kxu+pqCIrwT85ReU4X4EtySGVZnsBgPXkE6VS
cxNO28FUVjYhrdt47LwT6I9l65sNZeP/0OaeZIxvAuiaBL7xArRzQdGSHZdSUshAqATOxSEHW3zg
oT6XJpBYp6pjv5E3fkITheHO4+5+b49i9oodFD0CFgYQagdvLqkRuMJPWlM8+byKv3n+vVC2kibQ
/ubD2m1Tb0Yo2BDLgKFBHdRRW3OSwWL41REsU7xWIO3tvOJjMjlPBAdkbSzfSyT5+eSyYQnW2Ckh
PIvMIRKVTCcB56+gOnuR7s4yLF5LtHLww1vBgYpFxMtBi4946iwudbIQgpTZXV5n3GH7dsdBNVZD
wBdwH11vqcseHJOzXPZ5YAygU1gA1wDcmJ/BJcT2hVFHSMHc0yq64J3VfF/+RboaSHnXyXsJz7iv
00z42QjWYG+CKve/zNjPV/lmMeAm575PHiijKapYiO2kZOx7fqMcWc8fOluJrYm6fjOUxHMwwX41
QR/keAQCDmMeM+pOHlzrNQtsCIyifQKxmuaHMtTwFfaGCdV3rZf16kQ49xevAYLpf3oG5aQLbMGa
v3qD5V6joXJlCa6G9de4aUI9Wrcg/8kUEXb7BPPpR2rVOyR5T1W7dyeEETw09TFLM187Wdn/uin2
Nbj880hwR7M0jaDhzK1ZNdV3M5AQmo9BW5NNBLIzIGSYBCPVOFTOuPRdR8IOSwfSZUYnyj4M1X6P
h+x8Dye59LKfIDpg5Y4nEzp3cvilahqDWpZFSTZ0nAUZqNwOa5Bc7s6aJwGlR2mYMkQazZLTr/3Y
zXnmCc0SN/G06AZurt/prvOqF/TwTBj+HJm1JgIzSpGNxK1e5V544RQIHvqru8KDfbyyuC11n8jN
Hof5pnwXPzsbQ7QK9yXOWUaUj6axtDmMGkzBx/f1Qzn0yS+wd847J4ZKE5KZyWCWOoQJ62jGM/vn
x3JI7Ch1UQ6qNWdEUACd1xEcX8wXphOjF+aagiLU14FYnd+jJ1mdcLNPAEezNg7YHOCaUdjXYfWI
oWw6mGad37W5fuvNeOl1nrRNJ2gsdcu8ZUs3HhIfY+NTQjxlRy+kPYe+WypTLuqwfQtm0xFcXsG9
bj9dP8tAYxlRG71goaK2ejCwUDS2WYEC9JX+A8tlT3GU1C76cC6C/A7/uSWlpJ0TEPudNi0Fma5V
M38ccd/xmtOtRe+Dojkeqp9XXgjPBgL5V1DZz0K+dUorS3pnsfDSUU/om3yeSvR+Y75z1g55nyTF
v8K9+GRSjyNByjJ1aOzpFXmsex5QbbF2yhbqD1Z3BiU9Vit6fRbkFneV8fTgk/ngkfIqcrGEwmj0
3z7xUReJ+tp0g3a0tKvmdnduX2WX3Xnmb63T2AK0R4m1oKDg8YQ15QdMYczu5VvdV1+46ykOmwcC
H9nnrkO1OpTmX8B4EyyCeYMM3qrRaEhG5g42Fh+BgF31MOfNmBizRXQ5Sdnyz+tZp1TmzU8GleqT
RZF5wmH2IyQx1nc/U+hNYl9rMXpmHokhLQz3cUnfgiv3ZM12gKTghiJvDnr4HKZu1Kc8RulZcSKe
Jg6apUTEprb6JWQ4rUo+/J7k5nVq1/EQAzuzPX5WL+O4dn5PzHgwGuMzbGC1Bb6kqx5NtrDtcrY/
HS7S6x73BhiBtC4JJ/dnpwioEDCJPNONc3KD5eBDhY5fTHDlXXFyM+m7+b2DQ087x0pl3z22tEq1
hxUTpiLMkqcHnGE/eXPaFxvGYEzAbZaLVRkv04rBLA7yJzoYwjJW7YUnEKQWlaDD+0yW64Y2ujdg
TAoE+4Ae9ZuZde3g5Pw8nCeEqfP2bpG6IOyh8kBV0sKrhBRVq6O02SixTNiddhl6EVxLgCTROsYf
XegYfo12Tm2utb0mIagCrFkCEm8dOVJdFGq0N+vY6B4FeX3XNXUPCZnzA91KG4hyeoscan6iBtrP
FvC/2vR/wUyfPWrGx7b3lJz8jBCEOXXWj7+HinDbLo2DH4srp7UPp1jPT/rR20uV0FGrEnOUlpW+
JK+GhKShTPcL/DNeH83/wsiE47/kiNAxOnI2ylGVxNuQV0Z8uIJ2v6U0iPAVB5VloeqgAMaRJyuQ
NBc+DvYkUrUAtf6CIhvhjInl1DEV3cK6O2a/pGDeu+xu/6dEB6kfSym8ZRtmzjt4o885S7FyinIg
JXtDqsHJeaC97109nEwQ6fA6YydD1Zg1U1gVzsq5x5wGFXqtZFLzmc4wyyH1Sr5nA6IrA8WWZLQ2
wOGQz/LKZJu8r6Xy/oJ31dJOPkqPDli3IfUAZQQzKVijozmaudBWe7Yo12mcUNxxRXNCxOxZ+aSX
pv0oKhgU9HONUyoXpv/19Y4L5w6ub3LfzGOOBujU48kgtsODpx9Y6VZHR3uj7PKpTePsh2hrWZWX
FwvTeSIi7htSCJlPbEL4bGuiQhZ0DPGr1ttJAMDjZ4llE+k9PebsyDOjn2DHL9PBHLoou4D9Xlfz
/nn6xJPAmx28r1lCZKHnZlJSegH6vvC8RisboUzMf3Lp7cM/TTFLMyLBudCCuSgux0FaE5lyK7sR
87Qax5PVapkLDhEiBtv85KqsjoHT9jOPi+dBAZbH0FSAH35FNBAWdiOywe6hMgDe3ivrEeTSJwEE
33Lxgqeekhin55EEggZcibxVi4Xe4kombgv5pllDTFidEIuXNIF0cnthpkVkVrAp2bp2jKi0X/pU
4lpudDXyXiRXhZ3mnidwmmZSB78H52iEFIvHFeeXzJykj+gdaIZniBFxu8HMdjOoGDxTE1y8Bz8/
XdUJkJlwRR61JPNGbOln404I6lCP24Fy90NSM5NNKFPfrlGYCXVjllBRv2iEB7irDIevFdtdA0ed
5/sCalPweAktJURuw3FN+bouJMrIEJdhtmO/igFP6tUECyztZGIQNyIEoE1MD1PzXTveDxqWns3M
u1VjeplfucJJX/DqVlUF2+tGRs0AVGZOGSdCPUgUKZBkpZjr7yI1X6kug8SzN1xnmPta2+pghJ7+
cidp0wj1fi25tHCy7pB2jIVEn5mPgMYqHelf3D1aJyt+z8mQ5fRLcpfJgAuzW5M9IIrQMlOXFU7/
Kxcyl1rVz/kusprw681F/KrclfNYSY18607pVEH9VSB25MA+W0QxT354HvFjVRzZ2uJdmb7V2gk0
oc78kL3dONCyuzUI6S3bQlIQFfeWMwmj1ROG4JcfUGRijIF+8I4h79l4X0fUTvc+IGXCcny/t8QU
irksR+wH+Hc4tDkO+5+kr7BbmCYZC4OXD4UGE2YpYAH+Zcsn2W05Djf535mqXwWLQowaP7mjuCCe
iI4oxHVEWxKLYua6PKnnrYnuaSwjyn4a82S59JnMWQKwSmkQzejwPUka/nWtiaraF49hdqgVyH4z
mNp2a7AguRsEkeUDcy0T32ndSm28ixppyz60H84kjM6UOuu+33u/3g4hCqq6SJmv5QzOmfIcYvJJ
O8Z+rQBIF9qBJiLwSHOe2BwbV20zqwWzCrDXO5qcXgbWGSUydMzjVXIbsSor6gFO/h8Sp9OjteVk
TW4sWYI94rD979CscKlFpoggVAZ3g24pgomLQPy9YSeZuR0H3bqcJ6khLBjJDZuUFKmn4ec2pN6x
GmYjODAJSIXGYgCFklqNTjwlYZHhxUTKp4/slo7gT9JgeHXdYeckKvz3OatqO+7S3tBM7OeIATwm
6l9toiIvWZf98nBKC/lmijKbevLncPW5H7c1mhKO4RQk0JuErEPh1B8//jQo46Ojo1xVTRa3UXrG
EGEY4+3e6riFbyeDVraN/uvzasBF9XC6JgmqcTuk0YotoeI7mvBDJOQsV6HeDzOHP4KppowGVV9I
mc17asn0fxXLo9tzeSAFv2mpV2TXGh4MhAoV6+9SSqFiruc4vrGj/SyB34VPvOCNim52AfZPzLJ0
LYMxCQZ38tCAb0u7qDDwZnwnjo0kto6SPnUV8tNZZe5z6+MdlkkA5ORhmi+/HlzJKY6T3u62qyZH
kQ/EEOuemWoD8Oqt/gYd8yJUKDkSPyHcaGFpqQ6/Du9LHu4DOKtAhzjXB7cG1ZRu1i/x4LS++3A5
5pByzeKRcDvlosvhhCR4um/b+DuIH7Kog49xQFJT8uyxvhcjLhLwtufecG5UWoWfXpmOSKtBagh5
ZUIUJrKhkYCEhgxKJ4y+Aj2liS0156Z0kXdhhNhQ4eg0a66NCMc5aC7TZ6rhVUhPBfkcNOsVDKfQ
EzbUMmyIOZ3lJH0OAKezUfATWPNFNr9bNbHZZuoyCKpoZHzD4qlqbGbopq8ojw1tadVq3cyA+RLa
Ic1dFhOIyNS15fVvaWH7xZnAkky0xUXCPQnqHMwBqKKmldNhupgU+sTO4xDn10mxPNgEG67+V7+k
gyfa9rz22UboGtZVXmjLX+8Jh99OJ4iAbKJwOATmCeEHdGp3Rge2T3ZY+KbcAAzIOG1kuJAFXfXP
zFeSYwu+TDKgHiTxw5E3yLe9fgdC4c5KSOWtfSqAAO+OCHWAnlDqyvI7atQ/+hlUEv+x7As5KolQ
SL/eb8C66dOqKeihVCey53jw4XX96HOb7MOBPN9doeBXdKmaOStDIq+fsN0E+dW5qjK1+atQLAUJ
XhWCxw8GEdFGhBw5iQoFQHqq8RKTNzkS+4Ns3DTyHPavYKMKEn4o/jKPi4kKxs209HKirWIQA1V3
CQ5Uk+hp93Vs0UI9TyKcCu5Yl1URd61KjrUvMhG7cedVdRQTuhxLeYZ+nF+NnoeGtNuOTrsFhDQI
mCr7TD+RokcymjG8pkMhwZG6r2pWTjYuEqhpZl8CkZa6oGqBBMKsDl3E18WMaUFrbzp84g6m7632
Rk4barbnn52S6pWLdbUvrXipoGRcKDCEKPUnSEDwWeS38tjszN+o5oKZ29M68YE600fo5mscx4/r
i6lrMdoG7fsQZzNUoqkrJ0/PAfoSgDqcKjkhKZw5M6+w/4TLLuOaEH8PNPXL5H5HnTDqoPBbpoah
8n/4wZK6FPjKXwPaDKtQgkPr8NUdopD79O0W0wLq1iaHbbtWhZ3BPuOhJuxLOGdiSJUMjIGx8q9m
/nNE6dqaMt7kUxVEBLikphJhLr0KupU6D/08JQWS4gdqrHqC+GJjBP2gvC7bP43PmZco1gSgJQ4c
4tv9maGxZZN+4iyONBzyx66EkVcSAUi4MnoGWggeI7BVtiAgp9IRJ48cUWuAoovWDa6Ywb88LOwN
4YlmkZCQcFeuYrZ5vuo19Uw2jxb7x3NMFpWVJZU2r7RSnMMb0NeNn96GXBksHfEDQR4QqJk4Kdlg
wlwcbUDOwOIqKutqXhzt+7N8a/D0B/WjpSG/9PgUgv7YQNm0DlVLsVwWIT8VhQDiwFeLStlptfbi
yhAXsSwRRHwJTxw/hlbQTbYVu9XNFrOpCwwqi/6YB4hil+NXaf6Niplh56nu1/xf0kp0OObxMiUk
EpLOiA+6KNPu7nZfCCw41Wn1GZshRJkfFhOtyf0LFiFVj6n9BwJX/9eCh67dRjaMyJ1J7KQLcmZv
557+I47mF1t+Wzhc9sulshpAdRCyuYSx3W3mIRUsewtU1zVF/QhdXhxcVYN5tadIoribknUT8UU1
LrRaXassOWgWANoOTxK4/gtrONysY6EBalQV0IgPMClfLkjov7SYOu8Bl4fj/CNpL8WlE+qVVCkT
cM5xuXsKpqreNQBSotFVP7SPoc99QL1rJ/9TZDHeg4qO03ZIFZB4GVed1DEMCFo7tl2qHZ26GQ+z
6nNXs8g5V9czk4hfSVE7hQfVJVKg4zQ1gaYkIvvlCgllDtVG8Iqg8EOaNIYAsUUb9kTgmvobhigG
AYIyR1DUFjw09N1vB2G+7kkV5zBo5S+ZE+G7+giQKqqqH/jZ1HjXi0lbMDDxraEwLQp505rKgUCv
+fg9H/fefsU4KbKWLn6Ggp+pgc5/iprznVWdGGTJIW31NUPcVFAxAb6vkLGXPsGwJHoAwx5D1NOA
SRflksqqt3W2Y0XDdkuQNywqFVhWHfsqGAW9AR5YWaXhlMCRrdXDY13gFlVC4/kVixIlshX7RScn
LdN7A9VZyjYkesm7WTfPAOd6i8B87pXnfhhP7usLrfl64CNin3qDenYwtWUj+VMB/2+zvMk9V1Sa
AF2HO6SPxaZBq0NY4cPtcIytXLw18T++FyBFsa4PwPC3MS0SyKR3P46u/bTDTC4OA5qtfyOo0R45
V/PV441f5Qd/wzk37n3ZRB8Bgs6KYGt2yBX+aKxEACciOk/5pwf25TM1wu9vOptYVbikaVgWo741
Esf8c3vyQfE5jgqVTk/3lWFi11XNqNkJ7aaet2pC8l7aPOLZ7XgFGm8mL+wXEm7vUGFUvxMbL1ed
54bEKPwEMYZ7K3I4BK/4D+Orjms7GAC9jTCsql616Qw5JRJfDtbp8qAUcHlgGNNJUfHAh9pVnyve
QHw+oNgyx23/NH7hGh86RRxJbBxH18CSEQGnW6xwQKfBvhduLZ9ln6hzGBBV6LNDczPDQHEiweQj
/hvYp+QMRltXCPmyAPzUYTJWZAYJr58BeyBwrokVo+6saowA5B460VYizqXvpyRY9aYQMVg/Ot/B
9Hd4UQr89iJ3da8iL/lIht2nc/7wp5dTtQwHMnsEIRjBDzBuZDau7AEXSTwWwKNUcsV+xUSy/DI6
D6LgLh24enrcKb4fUz4X8Q54gfwr4ySoK9ih6RDq7x+P7tAi2fobZ8xL9UghOsCGCthDrRHNIOpP
GtyGq6GeMGgZTcf0mjlB0COWFgxrBM20AV5MF49GxOqbTsbAIgWSJKxK18MDHBZZs0D/qWFX7K3L
lbcTN6MTwq+gmoED5229FfxRSo5G/OFpo7q25UWdpcQCMRGo19UGY1zXjlENJeTDnhcK+3m3s5YZ
GLvQlhlFp3W2YzQ/1N/D5qbn/K0ifTi5Nh29Ia1+KFxfZBbDm/USNwaPH5F0j4Om3U7hELKbKhVZ
/vMX+cByJVRVocXBF9B8A6sb3pjZHb2JFXHMis1n55b9+TMnDIet4SuIycao5z2+DtwqSazL9iya
KTUD4m2IgXd+vPoSQo64LgAt55UsKQbmjd9JxXHJ1HgeX1IGDYQrPuCwyYCnq3HRk4b8ig+zldCA
pG5J9i1YH9BxOn3OCni1Wka+B+6KNuI0euccYN+f25hGr1guf0qtuGNd71yekRwg61h3aXKpYuL/
XhiDVXvBfZAGWWjkuv9d97udzpfXOvjLhFMMArm59DYBGOGFOwKFsjt8Y7vMFngFcMXzWEsU0Rfa
ryLTuuEzJx0qFZI7/R4T+wdhA+3bPto7dCN9O+5fPJeys1ERAqQE8NS7sbTawUXq2qgQYKq5AXDb
EnU3QlntLYdloVJea1VcyUKEfltliypw+zfsybjB6U8eTUMFH9nKJyDUuORUc3taOlLpVOSKLU7g
HM9IhcACbV8UxBpcm2zV6H+ayM2dXxl8sI8zJ87M3K8guw1y7YkhXN6t9CWKJ7DqGOOIPWrHmOU8
eI49fI4y6eLyhFKr5wEGP5DJ46zl+f6GSCwBnMAjwjDTCUNEfUHEBOlKMqXXAqYmipItSGPnAVKI
UAwx48JnSNYAt0pRz+KEFGRsCYs7HokDrYbXweo59x/OSNpCzztmJ3ansXENECqyJZHosbXwabnI
htsuMCeFT/aBED3y7dOE3FEcKjDmpcpKkJp6/DxjVwo9mc6pwax2qNKz7tv5PYNs//tPq11wbibO
k0SGbPvvnADYNZfw7ZID5CtE6dLSnIMUbSvQ6zk0hIs1pOZBgIm4XJV0IxEFZoTwugaSAE7dsKMD
Mr+3uLpIqPXVl8dTf/awUpIgSz31GN3RMsmgZYW/eRlH6a0GygWfTMXOobITWTei7v45sqYc9SB4
vlV1/3araRY+/AasUrZwKxgISs5oxYysXtS4rCaYQ4Myevk+leqXO9/yUvZ9ehaQJU8XzKXtLmRj
t65dw3SbpxvuGzETpIW+MVcH4XkH8Q4krNnKYdYjYALFT/mhXa5J2hoxYLOtEV4lDT+tqfZSQtNh
tAuf48pkPgNihsrokkJjksCI8QfS+FQqw0C2WtCZqZSm1YMXnGOSRRfxPR67/NtwR/XQWbfiK2zW
T5MJdB1emIUd+yYWmRCE5IHhogoFeLcbq+DxTs+HZ8jhKMBDf5XAglj4OkctVbkFQXDBKuXfumcr
6fGvrOM3zRyiCPwCAzzv3WdnSvJzChx9S6AlUddCNu1Da+xZDd3YOarSQ/Y0IiuxqNkGYR4GPVSx
+4YQyZiXgw5D88HhNpDbhC8luFyovv++mBt42jRxDu2xmuCZGqyL/Ofz0EafupwHR2/2IDoL44fW
RJn3P9SCGZ94XHYZrpN7Pgmivyc2AIa4/KIpK1Bb65f96FiWmQdKy/+fg93NwfmSC2KmKY8fVyjw
UeYz57KKOoD4vgA0aClijuL6DzMsZGNS0LcxxApXVwJG4aeIuLr7XoCYj3l5N4luoBYVcKseDS1n
HiygI1Xy6AEOQIfs3JJWCNX6lPY2I+UZrCGbkiTCSDOoTqqcTaKbNfTomFvyRuthzsX1Yrh2S/hc
qa3YUs0bJu9KNFIhAi6UryEBnaoij53H+pYugHSs4IVx7snUiCnXr66KKV/sZuG4xlmO6oJU7sMz
dJvim03SFzMkeuQNtYZratRAUqrUYpx2rHzyyNbWNlyPNq3AkhBHRBC69YPGmZZ9/eit6EpLlbvC
7+oDF31qGaLUzyhq8+liYYZe/dMuks2+6Z13TtEVya4CeQZVZ1W4ANWRAr38l9Y8zmhw54r0RUTl
RgsXmIHXg4m5A54cQzQaED4ARF+/uaQG/M6OW/+kFWA6L9EPKcKl+MXF7n0BGrekexUEp461sgvP
D5SwmeVuWLh93MSHXNUi5zBgXUu6GsyjNfk4RA0SQtsrzSAFrU4DpHhilE4zyTe7o8cYMlUYQs5f
m/k2+6RvXxx8Puo9Dre4uQf+w1oUhHyjr2hKP1YMNM6axmvo7+0PgANPn+g4LKf6Qqgeo2SUGr9B
jHTll2Zjh3K/8m55EaAVcX0Jrl9Wn1U2ihCqNcC2okJwoyqNX6mCkMDPgEfaFOfWMOpYmvDH2RaR
+TclmI8SL3RlbAaf+AgjBCEqT23h5PUwcwMfYE/NM29VtdVBFI5X/9+/rKLaMCs2jFQGbKVwNR6b
kFM0eoHZWLXWQ0vSpK8ByLi2LiMfk5sab63CoRszbGwLs/+s/Loy+Jqftq9xz9yF9kCifZNNDsgQ
IIojP5Qraa8ndDIWBKMPXc41HZPxlh9fPmuZzCkF9jmmytpU70dSzAJmkORv81SpdV/WfnQmKTld
42JG5OZc3Y9JqfrezTPbo3wKpHLzGDhBkw7XyY1IliDjeQXUabhiGqXzd2zst4vL6QsxjvKM2ROG
8awI6d38rAeintAJwqGuKn7HNFsKbAxcVkc5UpI3Z3N4F5S8kXoAGP24tzP63H+peAy8jBMNc1OX
LqDro0FkRhB+bKScxTaoq/9VnPRammWeLLKO0SiopV6eTsujuntJoB9C80TFmo7sc7ZLQwcAOnN4
TnG8HlPrvw4NtW5DGwU/MtqnwGc5NtIxsIDthRKgFbsYVO5aOkNpvkZwiUmjqJbKalANufAvShKo
17LGxJRXpQIcdd6Hd4pnTMmxBNRRUZHs6qV8N5INOkp2DQgjJzjhYAHY/Ch8sXiwUrzU5BFD+hrg
MI7mRa+3Qbeej/oteVKCPMVmTUsUepa0Fn3z2FIWfGLakThCAzn2PB7C4uQFcZoJj94FFhGchAgc
3CoKOwM+Xd7uYa83CJr2u1T0U1f4ZxbLJpzPM5kPprkaZDGQixCMePrxeWNk5I4i0xA02ZWl2fi/
87dbg5T62khEa7gYOyHsO6C7xwXP2wt6R5KzY04Lkx4OS5mVU8p7mQ2OhuDf3zYJFaK2+qQXCkSB
nkBsOzRfo00YuSvZnIMu2aorFyJNOqjrNvDv8qsi9aCTCWCrasmoJYdMJNvlk4Y0x46UUia1XtAZ
WRc8G2cG7OiTYSraBI71wXwBhc1/su1kxeVWEeeVd/+RWkCirQrWqrjTexAZAuSz/kLXq/j+XhvQ
MDxmmK2f4fAo4fOrklAsRH1pI8AshPnxfuddzToCmfzOheeozrnqzc8BM5P0Tbw6bgke+lI10w5a
LNBF7Lb9W9DGL+Lh9orFrmnriyqbhEklwp4pfWyGa03yp9b9HUMJdwhtJWfyDmnBhvMkeVgLbuSo
6GZafr3ScNSe6lnjlpFamC77XRaU65qHjqbi0rwdfQihXgO3K28z8v8vjNeBk6Yw8UfDddQXeFUS
NZJnrVm4IKoSS8xblT8Y4g/zGJvEWZwl7jtjeXwUxbdiF+Z1T4EplcLSLBm//T8L96VodVmrO3uU
w6lK6XMlYGztd55Fxuq+U9Mtk0KVUgrVaH916V+8dHAQIv7u25I2SR2HKWYnkoBDusM4PaE4IUpM
pOuZgtcxhAHLHEGBWk78Tmf8r56n3KWWgwMhXjs6sgevLzEmyqgwG231e5OkXhzickB2H6X21xZf
y75xE06WF52TbSwge0OvhpwuyFIOrMkxJoT8F9IhLPQOlHwRSItvN32+Pe7NJdrgdfSfN7+uiiPc
Q1DVlJEpLmMBYtWx20dUHGBsjsU7Mun1iix9JYklTKnPGPNr27p5OF9Ovwaco05sbBde5tz5tPLb
Z/cgwbfLJIurTl5DTBCTxhFoleGEuE17ho1DW1DMoZFRMTxhY3ewORprOnNf3Eg503nJiBbty+Z2
GctfbB5EJ3M5OFJ38I3EF6Gaozfd6+2P/oakYN+MzkANWmS1U79TWH4P22AooN0i8wxX8D0q0Xet
p6PZ5NHn714T4MfWVWVvApd3x7SwrcfpanuhqB0VjcLdGRotLRd+5sCfUSvkyLxugLiQJcQToNGq
kqsHMNBI+wUYyp48g2osnD95GWahuVHvV+7pVjm/7hW4jHSPGuLeXbZP030Qpq1ax/nDVN5nKThZ
mhNh8peosNcKeMKh3W03Gnug+Y1AKTWP7g9n3oOk3xQ++oZyL+huKV+v5YVl0w/bwghdmhNjMbRQ
d/jfFJWUKmeZiy4G6ZcY6979gwhKEPRpH6KRwz7dqz6A0awkKsFA7Kuu09ELvMeQnUe57EHwvIBY
8S1yTnNziHPVe2OxH+4cWu2kieVjPgNUrHZuqyOrziVIGy4WQhWxmdGTnrE/u4SM/wHX3AioDGZr
ANqaRQ88NiLAqKUt1C+o9OyBVloGxE7DDvJu2TrKNO6m7SOfcfTpwvA3vA/4J7+A4nN92XJqv/YA
d6fS5t6h5p4+176NDuBX4+yCH6vfVStzf77aajipBfGMXA1tIF6bKWe2qb7P84K2YqO9hh6Z8HQC
d93qKQ0FXXi3jYbVqiuiwjWrYRDIs82PksX9hltQ0bPTFfx5S13VUdAKEC7Zu3ZhF5De1VyrD86A
CGobJo4C16AAlv5B6ZYvWbafjkuO8xVG8Bm8/E33Zo++IWvk08I40gWyGUT/T2/+bKKHH6zD0idI
aIQlovQyUF2gx8juaMOtw6MHeE6epMp6Rv6v0CjmpmdLC4BkrxARhVMPJKJQTwj3MUuBY59aSXaE
qEYMvt9iXrrhB2qvhLpKzKvLKpCFZ7CT3e/FRW4p9I5nB9tPBahS9JU+8D482Lo9/u7DsSPcJx3Y
sDcIi+gJ3LHeN35pkLuk7xowuS2yEHjsXespTsR7reIUR9t/6tnY2pcnFT6WX9nBTFUC3EJHAUEc
bkRAwTcCxAtjEdw3FFIA1xmlcqZjsvVzRZrrkPakJTiWkNF8YMMef7RBvOdEK30PjoRoQs1+U+WZ
XTsCPJq2OLZkt8EoDF/sPXX1cHiI512r8vQrnkWDXJi863abH96jNIcbzFgFoBXjuHJUkA9hUkKA
m6ufBPUdXYfQrWKSo9coqEWq9GHtmhoDU8uQoDEWrLdzRA8m/h26njLpyrZBHOCyVki882EWwq3b
IQdZ3Z9qFAUdCmTPPIe49bphcDA58m+CrQKWPoGv5C2lB+ZfFzYKBU0Mx5X2U1rz18WugbgLrKdK
ep8Qco3qy/6owhIgVwDmEu1Iv8nN5xSJ0rvRwOm0bZZUnijP9/HdgwTWCvJKPz9PXmiytEAsqKom
3zsMLVzTz65wH4BZIUOXdOIvisIZWaoDdiz+OtYqEaZ7kD8MUyyrRNPbpPUPJ4wJpqFs07fWTdzc
sR0tzt5c974gVMsQHeE0FyTn5hxaehasO5NWrMbZ3nkSz+lvIBX+UJll2o8+IbIcJS58RUoyUgJg
NYcE/i64gy2xznCbTJDzVSAhDRPWMWfXEkKmGR4nemcV7TP0grRL3DsOUuROyAOiPdZmB4E6hezg
36lHd9BkG58T1NCC1jcCuEiKqFF+038S4+CRWXHKOGnVQTRmSnvJCVTjkt1oPWR2/bqyfD7n9Kuu
1xJlmnWJ5WsWrQAj/pvJEtIh1mngjfkdTz4kkXdWtlWkHFbtL6vwZrL1aCXXFMLG8iMpdsGRsDBd
ZgN670AHVifemUps2W9mftD/c8ktRCteC6arYZnR1UO3uoeXWwTCktQQSSrSQbjTMnaI46Rxflu1
Jkqo3pvvCS9RefvvJxDxPFMnt81HaXpnMhNIvmNHju6LAnoud2XO0cgCOwAnGVpsUGJsaVzT+UfZ
Pu3OsN8jMi8yHtrzxAqlWLVKLoWzV9Zfl6+nbuIt/lLMqYjDXtw6o8iGlyoiRM1qg+7yXSiPe9EE
iwCbRwHD0sidsfEv/8ty5lKDJ9mPcJ4tAE04oCvMUGl98mY+NY4hAYu7DXfzESdyamJHn45spxQL
yJ4q+FuFH4WYcyB4K50SdSoA9KTv+l++TdoEZKGlWbmDVFA06PqNJoE5sa6NH0HSzeJyqvQFSbj5
6e4aPVsyXdT80M9nBttfVgqkcvSxhtH1a7o8URp6IlUwSJGsGigOrilYWk1s06xeiRCmmVyJ3WKx
9icW3Tdd/TqgSkYPKmu+UZtdajrqPi80Lj/zh90iTtMDqmZaPzuI4plG/Ck/iD0zYYDyIh21naSM
cFsFXzNBnuNSkK9oxtG2t5AtmQ0KBnWbrqQFP3jZGrogwmTASH6yls2h8xuXAiVxXgXnhxKHdLlx
jlDIBurRE3Wjr2M6hQ1NkZh2yCD/oM0WYN/EQgHx4ajDRHSfr9s01nJoVDKm8qWC+gJAT5Uzcnzx
xWhdYld0E10xXfwA+dRp9P1srEKVKM8I3WrXBNyyhoiY1Nkh+on5+ANs2s3L0kFm9mH7BTnTQ8OM
PDqIw9yj13MwwSoXYv7fmrptRv/LFQGm4QOzyWxtwuQMrlCo+4VBuuKnaiVyVpRxhnyXehKl9+Rm
Nbh8FAAqalquYNrMHLOBw+QbdO/S23ATFZYQYa/nB3D1qeNmgTjYl4eUvi+uIFG8hNPPuDolGMgs
yYGwmyLZdAhyZ7w/zmTx9eYoUuMbAzM0TL7D1ZUSB0WRYJ2CMafksF1j3nNAP71+/d7gk0iBFCDr
TXQxK5wy2haBHkoaLFdf5C8tpOAfO4AKmR/T7zH6wPu1urhzquT8tn/2Vs5Y+PUHw4spEudU/RFY
eZOaFsvILTK/p3ziI1ZU8Q2wlQ/yZuo9vGTqJ56XaIxpziiXDwgNagLbO2pk8sxmXziXwCF97llu
uehSWS10FlnIF1ADVBZrrD6DTUqnkfwqDDQQSmrDaKd4WeCYdVSbLl0sIluf4+Y7nhDddWtV7m6x
hUjsjG0cNpe+hcgtXjt2pTrJO1vSw89Ye3hyQnb8GVSZG6k0U5pjikElmgooSjN4/LCMhPAQxMDB
RqYAtVyIZix/MxFOIMlcZW/65REcZgWgU/qmjBnyYKxEwCy6YnCyL+5M8YsED54RqcvvGrmLtkp6
4EpJ4Lx/WnzloxqXtGON+zJsUK7F5wvcXhoGw4Luv/McBj6TzXUpQP6KVphL63cYO0zL8umIsgws
giUVgt6YFiSMsneqWAqIjNHmlkWbHr3KBSEk5U1p1GCn6MYAFtQscHTYopFeTmTEbeUDhze595oe
hVPWqhIsKZ9k4O2Khc/HQHCJ4n/OIPcpEYPk35iELLn+T47NAXSoV8qM4qNZDvxUpf6D3PH1ZEli
wGSNC9Af9Sr4ejqcazsmi2W6KLYefO0TodC4Ssx9iiap8jEQRIU3F9/xRYcUFodGnVWz8TsmChpZ
hkqhbbVoDriukDFIpTx0ZkkIf53JGAKw/apA8nRhLrFCY76yPbJDbmK/IHMzOPT1aIoh4+K2lkOp
lf7x3VGLhEkHlUf+lb+DarGKn+46uG0/qVSeeMMqAkLQhnQ2IYAm+SYyx1sjXuHPIrnxk8mo5dBe
rbVtbqXLFp787EaGY0lO6Onzaaw27DhYLB+ffFwluzGVyN+QyzDYvmJJ18JrPHx7vdedyTgQhLUR
AYQnTbbshxZB/ex49geaAdMG2Guk652XLfbwHj93uYDnaynRl08E6tCwaq3asD9+zlqitvm0BlKW
5OfQliFirWK07/+SzO7DqWCSMzN6r3jfv9tRcFHDm7Lle73JIukDYKtXEsewOpToyP+1riUIoSlD
JToGnBAuwyFk5JpIsB/ppswSaROfEyb2OOiu76w81UzoCdKzubVmlOTpizPZr1iXQwtoy4Thtbrz
OGPfmXSzyMlKBcvaF8+2phlJJiUDmq+lXef2lTYomOxXV4m/Sq+DH8nU7s+joeOYXvvz8nZ+zzH6
iPk6GLPnL5Gk5m8BXAumDJOUl8ry3zc0f9saCpc02aMwGyJ4RKcECBxIgUXWjJieuRi00qEHc3/c
J88pSMu7q4p+dTj4OX8Ovdaza+m4Ra4yZG3Jvk9dZxejncJAkXy9peff7ZRpcaeY+Vlwc03EJ43L
GRKXG7s07AMqtpYoWI2To64eWipvHO72Ngv4pJRFWdEBQynEkWgkmrOBWWmv5CvIsPEBkMa45iPj
nP1M5ARjYXcuKrb3ATwMHttvei0ujsrtX9Psls4ONkl7PKAjqf3CuGhm9tm8dRGXMxcBFu2E2R+d
ab8PI95pbfOMjJehhwdiNgvdvEUGEXBUMaDBIC4AY6TSAxK5gEVuqZ07kPs+aTkh0TMIfSQ2WBkd
cvPZUoS9foRVXH15y0PGH4W+81VUFNbJMpX2e5Y5Yis/5gr9bWjzZvqzUFh+0MtALanNWFxqELQt
NWGwDfOXBfAHXI35+SS9KFcY50iukfnc9tbBvZbfJzS3ZNwhSgeVq7w3M4bt0by40Eg7V3cA2lOT
4bBzsTG+HOZ7cjS6wURPi/Lrgqo9jLn/FOXZ9vrpBFdESd6OBLDvDzdJM2YJ1PH+6iYG9pFcp2Tb
FjO5uCCDj7PCazOPkpiq2Qyno1zT9nlSYFyKhK+izbJCfwT4v6NxYJfzBI6HVcu5/aCUdWW0A7mO
npoAOKvQN6NTsW1+f+3xx3da8ta7awNL7qaS0mN3QQHAeDQfaHA+FbT4KB3trmiLE4WRfK8W2MNW
4EdAjzV/+X5QY1Q9nPfM1akNOhBQdCwd6SxDxkbfv7LHfl3dCWeno4s9ZGs2x7k+xfTXyuA+fhNP
0GSB/ig4iupdWeo9J3p6E16YfRuS3joAxhAOxF/aD3KoYO3w+mu/bcv+5+3Cyu+MWmy/Uq1gl/4v
1CYraOKJA3C/EdJ5Fyh8K6J+JZU2dp7a1Yrj0iUdG+TxN2k2tWC9kUoHrb9phpdQiS7RSoGokvTM
nGTpqXh/JkZbvPmgEGFvNFGscr7E2hFPoXdvfby39Zcv00xQ42GjHAy73crTY3nbdmMwamF0Ukcr
QxdDFqPl/rfK4Y7bnygUg+LG26F8uzUln6bengVONlJmbxk4tmTRVF7NppMLTsruGBISqVvIblxy
72xtv/syg8RhGoKB7BVuMxPfT3IGp713/nMuHi/x5gke713y5j29TUFyBjkLxQe+gAnSZ69ptFyo
eQLqcXSBd3T/VtTFnwTJyZ4KAiyyYbeehubctmIzoQN/w/2ePMGEUckpQ4HDWIEpzNoCTKkmxFde
b3zpDA/d8KUOjYyMY5e1pKgZmnGkzsWrBPEbCHYIYoyW5tdQdU1m6x8rSL3ZtsP4puDs2mehbY84
aIGeLCHGjCBeHvLGOpqhcwvuaULDyrMaX612vPgd6t86sIV4bJLYlUu15p1nCme/phK4hjtylw3S
lKubZ6an/58b5nEtwhjIIwF2zgrfNnkQ2GVe/FnnLDZs8rANqQhVz/SzaMorl0EqpCeIC/o2HS3W
NkDbMyGT5nWCU62pg+TKnwOVp0fryCPCDqEQj6eGJIP/RWiOPjCZvigXZlY4s4U2JJveyCP0DCdO
Sd8pw2VdLWtnZYt12ckFpNclqYgSdTtBSO75GLl+Poh4cwIsoyX5WcdMxA0YQlUhl6qDB3eUE7up
1owFVx5xd7n9lj0ug4P1xhg9CtY/C1d6l96d+1ce2s+DQXtKMgP1aZ+sQgvvHwjyCq+9pkUwnCYc
Vb5tEDXQD1/zsiow/Bcf4MZnNBoKLIxc+eZ/KVveC1SWGB7G3EoIhzzU5w6TITyPOJAO4dCB+9eS
yaIYBZMq7X4Gz9jMaFBiiR+cYUJRatdbtR861nOuqHAQKCmO/qWy7jZ/ypOeun5EaODeDbl7GVgO
TJR/Mmnz0ZwNDjE/FSnMwzv02651RePckOYkuhXa3YgFD1Jo6ywJQdrjvTqJsK6qb4z7goS9g+k1
VqoTG9OF1yamuuwABoRUMUzyg8XR5/WNvdQBAxD7W2CTb5IFit+cfaynp0hMb8takHvOILqcurFs
1+kx2QMqj3Wl+yZ7JrSnuvHYwVtlNlkcEKf12nAwb+mZ3Ag4ClSKVYJvjXv6KUfJ6VsAIATS6e8k
vluhNwC9ay4P3YOyCon1b3k9ZthehBsGHecuVcVMUi78WS0IzGs29qui2G/+ZEle0hcPogmlsr8Y
JEesxWRARJ7gqPB2jM/6FkXHBFAbTOQNfI/7GW5lB7czCFTGxCcCohXVcF8qhMlgopLSRnnCKN84
wDDvj7rBXf7ixmhIhuXp3TUehzA06ekbuUhlxOa7mmmtMa+NiIWZ7MdZ8Tqv1oGNjkM5o/CzwTPZ
RVnyDS3cER1pEMgNUPUtuFdScpTohg2WEPFhqRBdaxAKX1VEhU4nbmJRYyY+U1d2eZ6jPHgrMtwm
rgpxF0tBihy02aumgTu2Dr01Dfj2gpMlb5g7LIPjBScxfb19hTJDeyopch73m29iWyE/LgsOryo3
GrYCCvdnmOxxO71R3BnkNZ5C5RJbkPeos4XOV7poj0puj1bepUDXGt/TQwk3ahy6xkGlDAdWnwcR
glnyItPBobs9ubMHfiEBd5EpiZOve8a1W6U6pCL9xm4vZJW/b8ZQ9Ab+y593ef3g2UBT6EEzwVIU
bDMCZwHRB+5G/Ic11OyoaQpdr4XVt5zuT7ws51p8UwaxoLe10fF82kVBZa1eajxqYYF8AOGS2B3z
bs0BT7ty+jingCug+L1GDyvNg+J7ZvYKPe/he4GipMxD9kNrsa//HcEH9acRs+6wzhnVZ3ZP8gEU
ADhRczSQ2gBPRuOGiGXuNpmDTgNhLOh00crRgTlUSFDe6AmAJP8lSAlPsawlJdExY66ZdpKXu1Rq
+73xnXvX5/3AWFY0wUCOqI+a/O4qaUGGEJKminlQlkb6s0GtZz9LupKy2f3tQSOyBWgwq5oI4cpv
Cl22RVsPiZ9Mjz9UO8krwgrZL246HQj+7ogstXivyLORQaLt7jjFofCnY3776ip66HI00EJdUlpZ
NEvBFuZQoWg4I5xadYJn1WdQrr3b9SZYck6pf9sYv4kU/HKOIsChCqEXUyQTg1LiLBYekzySFEMV
OLk6pEPruWSh6WFOY5M9FMJ0j9YKBLgmBDFpTZTmFsW+hjj+81YypGfy04cagE5lrcCPjk0qespO
dE3omFLVrAGxsJCn1AiC7Dx4p5XHNVNn358Rv7xWUj4xBw7Ke6vvBcNcG3MXTCpMRMMqER+hIYxe
UnirRlG2PcOy3VJ9lbysFr+6Zya9YvHcjgoVvqM4sjMxL9IC0T5/a/lO0dQarDUyEdFFo4KtsTDb
+qPkQ4heF2qdGVonEnIJUpTunbEfUyAbYWdXMVTcJzWv7TtQtKiz11nRdhFM37tp9tlAwk0iYW6m
XrTZ7iF0gtrqpA/mjnaho+XAptIJQL8cGqgKKJeKjh03aiFuOJGjGyw4s3XETipTxPnhK5bj1Pq4
wP6+wFDnWrbC/j0Y6GuazBdJlqkoXTFxiLDwTR4RpAzoh6SMOSxBD6J71Vb3pRcn9A60UYzhS2sT
Gyc1RTwfjDpMPT63iiB/HFiWzj0eB0I/nQ/QWt8ZgR6sO6fBgGzUWnxYBnEl1vNxRHC3nXUb2rpj
uNcUcBzZkoq618xJBM5OPC1FA9B+Fc7qJv1h3mmU8ubfYGW+9jZqpwnjxMoU4ddtBkdUkR4c2yS2
Iuzw9JVODUxA93CLPsV5jt64tKKanITAcjWXxv2t6GZ4bEPDYAaw/O/Zrw4C/TXuYzyYfxxOhNT1
bu04iSucNRvReRfYiReedrOdHDMT56hrZWKCVQUuVw3jR31zBaXlv5Au0waoQIjLmZ8xaEkrYdfv
Bu8xRX4DSXT39q3t1U7oiDM5aFAKI4z4BTuifN2VRRyoZUInJxsUSw/5UcjU1rGwShw8SuZPI8UB
1vUqQso8njF7P80fJlcF7zXFyVd3uqrWVlmvLk2gBrD8wihjszdQntkegOgS9zxBAgEAVBIrAviw
cQYcYJHc+Q8bjlCnhFFU/8NCtOkxBROgcZ5rFFNrlOFH+C2QUX0wDWd6YZYQlSOyqqybhCmGLEHY
BUA4ZxleEi9RpJcn5zM6wqboHrLB+iLMAq+0LdbBeOR7NKW3Yq8dWCKJStL/QjcVmI4LcimS2I7V
RACTT7fudNl1DyykJkQ1j0efxFgIjJIloor0VMxN7EtuwpoAU7Rg9KuMdGDMSKt+wK8y6NSmt0Sz
vN0vcdW+plPfwYOgeMGrw3Sy/SLpHYlU2klV8MZMo6iM9Rdi872Bes4JaytHncZvEH69QKS4fIwq
EbtyU9khyrle+MhHO9KPQf9eAMn2csZta2wqrcmZmd2bypii/JODriepdmOauRXf4tsB/PR0l21R
uSj2yjrEyqjD9JrYnntLVCiKTAeC5EdsSI7iDkE7KgwuptrFfDEuTPblh/wyYm3KBdAens46uUh3
btdmWHJrdi0xeqalZTcXcBaUbNzRD+alEswf+JbLHkl0BR7ZRRX9joUiq7Bb6tyazPZQ+VWgIhFb
DAbLbPQh/XNevLqIL2VFyvqaeMwcWyZNQpKuaYubecI1iLcjzajh31uD+WqSboY5HzqsWXElnbzN
Gf3GobpEe8+AAtzb9SoRZ3zdn8MYcdn1Emcw6GWkbAoDt5pTkwll3Pq/TnmZ0pCwQK25pA6haHi+
X06pKhbkqqfvLpbFUpclGOpRP1VVgU+38cFkjv9+8FJu6vkEO5Ghwtvo19jI6x0e+eGy4Y8HMh+h
btg+KPvL/gRSP8t/wtONiIYR7FWfELeAK6paPsCF+k3p33JyQeNYhbxCEflfieaPkqfcD6dHjnY8
zDhngSFbDwYr/bCT65cJYcvggOHcGeszZFqV6Egz1k6as7HYjH4UCWCL6846cB3+fnpVRzXOa2jJ
CFPS7dGj6yHBC8ILSWilZf1we3noVopwTVrwgf0NDrdCKRqbuNJ57eape2ZBEq8PfY6Af7lIlcEN
IhsUjylKZMo2H8lKlkYVxegXoH/19deMzsay2dNbTZS9oHliyZTBI6p8pEbqUUUBrJoA5SvFbm6j
0bb8ZF8PK6CDKgEoD+XSEe1gWvHUNBo71d2iK7dWR1hZKdLSrySbpsSdb1e3vJCZGKy2S9FuyxjS
SEie+qC1rE1+azsUgbKXH7Oo59JsJid2TUWSuGzSpcWVhP16DdbOlAglG5i65ILJ+LyaTNBjgjcO
cG8wR1rWWI8DTVlBYMwsWoVCwPhIF3EsGzaMjBvbmTk6JO5QwZNJnYHzfOpGjfD0sPZIN5Vijyjl
OIiQZr4Xqu3uSVOB/gFbGJvkSOb6vdWKDQ7PKuOZtxVg4etCcuGys2Lm3ltZ1wYWq9mOoi3aD4dF
huIqV+3Jv3Mk/qMsPDdyHuslVIUytI/0EALb/jtO1lcha0P5AqyEUjRTCCefyBu2EJO5pocjE2Nk
QDQkOTrJnXuS3fuab08mmgXI0AV5vJoJRfUfRgEO3MNnzEWG7RYA5FRfrCIM8lzajlkt8LlxmtOL
V89RwQyJGpniqmFK5SOQYPp/b/piXOfJn43s0MuHnDHf53BPfe7ZYmUEx/L3KJONVLivLakkurhZ
1V3qN9i0oarOEFtafwkLhWkRTEyw53Y0AvJs4oJMOAGMmuZvX8/hGASU0HwDXdIrRGvL+Pgw7Kj8
5XRjuhXR7tFe+Tf74qwOxVY0Y9efNvSOieiGjNiU1WWDE9vcN02zopbdgkuU2vtfrvygEZmcTSzk
7o9nO3o73dq5JIqHgR0FVY68g8GT7HqZ7+cEQcROE5DQ9PIQy4utGWWXfM5K1z+YxVUNTVDsQWfP
zQP+0TpL6PfHypKg8ft/4tunoSqMXpAXAaslXv2jhNk7ze+AR2wFOZdJezKrrZkzXaY7HYFoci5c
D+CSdI4/X2w2uVC0Z2HYDFgm8PNuPcY9oBQ0Am6h/+QGdovTCl+vqnwOIa7RBfpMh3onpiTxe1Xa
O+kc2pAm4YRMMIjJ9M4548lkCQ9T65jeJ268SwtaojJhEnMPnEXzH8j9UcglXUkWC/tyAbfN6lRA
ZDolRIiY/TGgTnAeJwM7fcH44nOh4bsN+p4lvxwccWhJHpEzcxrHMlyiyBPot6lIC4rdt7nrj9Cs
owZZokznvdvjbs5WrpF8w7hZOtgLICpydxX9IaQRpa45CdvTHy6MezIQkeIhhsgJQEoJegZFShtG
tN5lKIztDmPUWsjHlgDJwvuaozYCMcFAKPrxmSd3rFK2DKV7chUN5/iX4Sl53KXxQ/i16AQoP0W5
/3R7xD1vn6ha9Q5Zw5GXZ61/Xo9GvjOkxuO6obP1eIqIcH9EfRqIbp6sn0dL3/TPmyRaD0VnDtGC
g5IX+7fV7wzCxodpGX8GTTd2q1Dd6/A99MpFMGhsG601BJ/OEJI7iw8vrRwJciaTfsa3sjXZn7un
1M5d2XdDDxOEY6NOFYdKAGKWBXkwQBpnkKUZnXrmjDI4YHL59HwYBz+S8nxwC09TvVH1cfLF+thF
ErD/r3o0mo8daQ6zOZ/UcDGML2X7Jc6hrMAvDtJBNox0tZCS2sj3JJGNTLiSXJZ7iHowbXkL1wfJ
AWtoLEMsI3w0ynR0B5TN2CR4A9NDUdyM6zNAMY9oNd3dLa07A/fIWCdg5XNTTz6JQ0NyVfm5u4h2
jLaOamv5yDStkZHF2SZxKgioCA9iJOtZsPmKM8UxgakodJddgFNfm7ZSPW/ZvGjkCvIiHmJap8Oi
gQ7Pn8BmwcGBWm6EDDfrc+sAt1iDRitDrx7eq+h4wS4u0jjwJT3yuGYTuwTTCJdlhExcpeR3Ut+M
htChufSsgbGot93wZeHPlE6UWvftOLo03IOhQFDLD9vHhkRYpjBtKPw+w0XYO2HFTdsmb7ShRUR9
K9dtoRCCTSMwylTrl0QF85/YrdB8qyQgrsJ7wSUdYkvLLwjiflV/NaN68doLwHmTaNZLYVjA5LF+
f3rjppE5fcfL1KC19fpI3BwvelwnWtveGPQEZD8zLG1SzhiFSQ/9cKuzXepm7zCBLQl6P/hC2RXS
rO/P8HCkHtl0Z76csucZlH2JzqlmUe+0sf7DvSZM1MUty3vzbeOu8XFY77ahmTRZXI0d22ARdPtp
EyN4LcJPk2ghKUdyLKjePnzXikPTBNbFkD9wvz2ZPm5xFJBsJmjVERFVPMKllvWi5/3EWkTo/EX3
gcbc8XMrkIPf4/i/PXceA9CDjNYwJOMpzniUr9ORd43CVYWH40VNvSbsSJIzU8XkrIvwvRncAcoz
xgnEWM20OfODG7oujjoYci0RMNAwo1wS4+3G1094LMdRSfkPVcYy1UrBLqaUQynPkfGZz9Xd823n
z/Y2hC+TCIXLLtzGM5xndlTsxSVKXvDx8mlfyB6bPVZInt/9nKJ2zvsoTjGNhRHil2DaOBP3Z7PI
I/rzyySV4GUvgz+0+Z+9XGlv9+Np6fMWX5LAEBCgEk6SzBvTP9W7AIqL/M5JkrQrK4GwYrAtd8ai
rDDoKdsnGkX5bJV7lmKYqblr+Gp3uHFxXTukAW5y4ogxxVmbBLnVD5fPzWxmromzX1f60VOEd0pB
10EwTLl84Wv2nxW2Goe8Lcmsuur97Mn4UpO42janKfV1cayEqYGC7J/AawzXKqPr8Vel7poal34S
fzPbXLmXdWNaptnyYmwLWRMfaPW7QcmXgipRrF1YR8DDydp9kbztKXbaFJ5vSQgN4lVL1jtWriT3
R+Chk730dEzGnhD570lWAsSZG/gvTtgbJdZMpGZ+xopppkqA6IX/wGxGovs82xUor+yd0+S11oEE
20mlu7/nxNak9O5x4OAqfWKnq5R7O87mwK43B5xZsEzHPf7g94xJ7MqpIVQqP0ku3OUlA/S9ZFCB
k/ZglRpmkO1UPLNqyKAcrDYnBcwavEGc6Euj33Mw2cQXozp7M3M/GlpLTaXNWHl0xjU1x8lyXfK+
WQG3vXiEB93xwSea5W0tCuajfCXbpfZ0EfAfXfAznA7xDJsOfCdNWWPl9g6u1Y7z8x5k9EViQCPo
yF3j6fLxulUSFn2WQZg48kLyy95zfs6k+FwRdx9RGYRWZAu9U3c8m91HWTvS4ZNIcgjlq4tyngkd
lckE77GMFIXpebKlBZPgY7TCfpDV2yWOpx7ncjFamWtcOh1Km93eqpSVSetn6G8Y1XmaEY8xHA2x
p/hMgsgpOyppKmm+xnjrM73XYxjV51kz49H3shDF6SM6xuqbXBS2GpRY9878Dq9FL9ltVCTo8B0E
x83lhtpeqjT3WgQVM4IFH2ZmLJ2xoZQxOrmsHxwk55FLVBADL5cBNqzRUUA9sLoWlmRHYiwLd1MZ
S2axEMP9/qXzrJnatf2gFB+IX3icGtzAe08wnt/sBkbp9z8GKDG6t8dDppNY0VstJgcjW3r2crV2
CEHeoyPVR0rSTmkfr5Qw56N+lYwHR5q0zCSVVEQ5RFsSuJXqlcTu2339ynIYZP1ZroaVhlWq7Z4E
sCFuAkCVYOVByr4qQcQqXHHQKDfRl4X4FyP9e4sz/en4LqcmEI2gZKx4iZ5XvAkGjlPYZCgduqbl
tsuQ6NkWMZeatQfV1MtwS3l6mar2rnB3/iF22ecEYW+6LP/QOH+WmjSg5n4OfgKzpi6zrtaPVEA3
JahSrx8XwnvWz2VvCySW9oUpNq+zTn2maDeDRfPNSd7S57prz0KeveFieZY3KTcWTyVeXB4MiWrf
96hUydjj2lKysSdT6UGkJOQ+EHFfwviSPWPaMd6ymxHaLdOpZP0fnPQ9AuqXjcq5ynslEdFML03j
jWnHD2V/Jz8vSBRE2CAljwAZcnm6GF3mrJ3v7ewAlT+xP8Pjv0RpB+r78CiylO114+ZfhpyXI3uH
EIwJ6Br5e12kG3oeudPGafH2Q/5btDi5xAukNsEvPWRTtIbfn5+7jYR5HuziScQ8jJUNhjXOK2Ek
43h2YbUfEF6fEWgZwnRVVG/4fZ4Bd0/TaODvSFf/CpKxtExe6RW2f971eUH3pg95XoXLbQyyuMiN
/mUW3XdBNA7/fl/lkBXoXbAu9yPv6CwfOW90z/9f1WeDDLukbEXso7g3Bjy5uNHIgb8upb7MW1nt
aXEELdv6eWlOgYPt9enmfQsRIgOHl6JZTd3YDbdf0LY1bn0db1CoNoZq1x2fg6oZSWEENTFOJBtF
VuUhCqOmknPfRrtAS752k6Ozf/qyHv6n21wZ2Qi4m2ZYdsUlvWuMhv5kiCH+08kICzh3KkSiHEto
YfzE7kxuizAFYC3mf/qCMl+qOBvefFE2jBdeeZ/9riE6ruB+Dwujz/FfUGTSbRyz8++Eh/EoYg6q
B4eeEk4wRx6pCB98GAQTP3o1TKU2+TVLQYs4sbJKIYEjWa3FmtcYceUtHYTlMo9xcgBuPZohuRML
T+YuB9TxUcBozBnX/jWQfKk5aPiOR9lcxezCyG3iBJShE2s5oywdVsmhckI1cW4z1upsGOxRCz08
Dj/O6WLlWbKKnOUEVRbcI3IwWTA5ZXlNeoAbu2Lgm+yKKdb85gTgTbFSCnjvLYhsPVUSB1Dz29gr
QG5TleIs9JoXDhop5H4YmmJaZufMpxLMWKQTCSWb7hrLGr7HL6ZzdY485xYqOcyKstBC0esJswIi
csorV5f+lqaBtOrdaCXW8Oh19yjO9f7yvCSlio2kuZ4Ieea3qkFbbMDUurltj8S15cpa7Z53u10Y
ze+8LR+hu5huzd+t0xMrG5Q6ECoEuHfGsj7HL42dhAoEHnDjRvcmVIqpJ1OPn1UJL4lfz/0oGSML
EGj2XOa5z3iL+Lf/lu0imYm5EdzWSOcGe5jrMwOjNBKSrse5fWHlsP78stLNtbey89Chqjq3l+jF
Xo+ycTQfQW98OYKlAL85ytTQ/k70DucJjNQwe0HNKHHHs4jwg/mqLZSJ38IAGZm02rC5OwdHLcRm
cvuuut2t1ze+4eRijg9rwuUHzEGhPpvpNmzcVxPFkKad9R8MvggObtFBTj8pkxEOx0fvctxYUpv5
3uaiCAIA+YC4wlc9uLlfC/9EvKCJfT6DqUybrgL6r5UwhyejLiQvBJsAbD3gmkJ90eo/31cSoFU8
5j5AsQvhqChXHeWZ6/+/Plp1hwbJqJf3H/Hcyhdw6I1sz3cap/itCV1hFKLPlVdnjn6BW8LyIbNC
csUugVfDZN/oZTbq9PW1PN3eA4RzZRRG0m0JkcVbdGPoqll07PqsdoLylP3tnEN6enN1ssXQ6U1C
Qr3KxtVtyXvb3c0UJnWJ01nmdZLvSJcdcCeQOWy5cW/0MAHm8xRzkgzb83D3MS0AhGS6VFAMB1fi
JCczaVc6JQx81mz5Rsu9I3op6u5ABeaRGtc5KeLUzQL2SwuriDWDhYwcq9ohzL8RABapfiI94c6x
bvFxlo3Aw9JCMpuq+n5P54K8uf0jGA/TUpEb/nkOPPEHG3SnVs8W0vakWnVH7hS3P2yyEXBEQFea
6Sj53aU6mPRKgWW5nJcV7LeaosSvPGnlS0syDKBUSo2WF+L7KYDfg60qbGYBZmcOlYe2EKwb7xGi
eJCvUnI8QZugp04BMvLKCM0G2teicOAFgKFzBN7iOTLsCfV57lVra72dpCkQo/jgENlew9vkyhek
jNftQ6jeRStdyBy/KPn9qAX0qGTSqlZFM4dnxilwQdQMKkDpBL+UPOrtmATKNLZqFhM7hIhEfJgW
ZMPNIaSGizTx3z/iMhZNnOMmOzmln+fTXsdYum/FAeBA+ePr4Kj2Nmq15SBbRiCqfbzEoOQTRxfl
YW+xvrrPXra4QHOeJIz79A4iJ4OT3lnzvccLo6NxySW1ZpJEzCxTO+oUoD/NwgHUAAaATM9QQU8d
yUhb5HK893Wtm8vf49xWajWnpoQ3fzV5ahW3ggjNDvQQZIT7GSdZ5W8xvrNxNlkGJC5D5NSwHN3k
VYQ3QVXUKPtEoXxUIhG8rapDlf84UwpZ2hhvSA9uYpe4cR4D5K61gZMtKLhibDz9vbNMofDlQzjH
Bbg4Um2rrTugoccbVYw9u+EueNApk+xwsDGzdyr328Tmp5emYMYw6m5b5OHFB4pL5RxU1UA6CPr/
PWgmdM8p/hBJVsbpzcWQjPN9IDtPfsxeTtPy92UD64uSuBpR03+D9XVRmftu/e6LHHI7YuGd0d5d
AaJJGJRgYiolZG7Lew6UL3I1Wf46K+r43G33uyuYliEmKH47AJFQ+qrdWsimmGMY+BuVVmC3VrzU
WQja+Bg4pvPvniIGwAJmUgfLwp3XXhyxMoYCS3Mt6tgGRRfjS0L6oscLOR/ql1dPIyRb4o314uXD
uphvYe3VCDzTcHzeKg3SSDvovA0uiSVe9nqc/t3NnoPJjyr7hNXusQFYCvG3AIjX3+kZN+QJB7vb
QXERv8Uct2aIamTwuBkFt7vP0nIgc5uZep+wiNb8l7RD0bjsxsGL+4WzW6jkicjVVKG7+TFUnPmm
6BJuv95bXdy5MWi9SMQM8/Ip6PstKaSN0pDC+FaDKKO679QpwwLjOEr4e3b4ujucDf4XCtlC1F8B
xNikj1tD6mkH0dOsX2xcXaxJHzOXwX0VUcgNoxUqGPymPSBool9G/jAFtkDyv6YkAlDd8zrYVG15
ncrF9Fn3lqe+sryUU7J6dszJBwqm8nFmVWzcyoSu+OLeO8VFrkuIG+/DVGKYBzTWH2/6r9nd7pNK
Uw3ahLPxDXZpcot6ik63bAUuFiU+r+kYZUXrSM7RvxVR8Ay9o3V3PcsBuEVMmWlBTbCpzccvyZIV
upe96/dNwowKKpib1sn9Rt7g9bMBXw/mzx1BHWZtejeRXZF9NiU8f3r9i3fh1Nj5Hr5gSNjeNACe
+vCr8nD0yilwR0RZQcXynbJAqSTGXmsA9TvEqIPCUDMHuGl8JTwB9U37kt0VlzwNGbsKllQQISRb
rbmWRVHDM4bCK4aWRqq9KFjT8Vv56z/QDcfMcABsXPy+tcCanplW5b6+HIKdiDb24d203ZmUNUlg
9rGLS7bqvNK6pHTuMbNpkfxODiZh7uL7siVgqf0m3Ckey49iNqkAwFPEip36g0gzdPqj3zp/zEar
bafwRe49Su0Y49s6F2qQN5+QYsOg1s7BeGV85cwDiqykkNq80ISdaOQkJOF28ApG+Egvv1GtLblZ
A4U8GEraI3zaBCN8iPCWyhWkJQubQ+k5kn2AMFSHQVoMiU0M36of6M9Bl0ren5tyl63yg6Wyc/qA
dVf3Auwe4V0n7YEmIYYZf9KQGqZEyifDI8Ouw4eUxU1FiqyAH++kDwzjesEw5OhJr1+o01B5U9Cr
NMvHbcJZd7qJtPIZacYj/QSyYQSUI46H8dMd/BzkzSWWksoE01fl/V8GnQ2vWQzChfWVHlZ46pe7
ze68o8bTL6fsqOWGsAdy4ASfnI3nTx1J90FEY94cZBumcoFQikHVwkGQ810rgE6/TPM0awuR48ya
+TJHuyMRl8mKQ7ToMhmMkHamsGGwPvaQS+qCGZKlh+SvnfcZD9dYr+h8/mGCu0kfpl9HVIzbxjah
LSNM7jqZDp4QqR0zd4OrKz5VQY6HM4cfxWVewctaus95jWpa6i/Dh9O9vQd7nggsP9av/wsniypt
CfyY0HSKCz8uccosPgq/jmyPHvAxNuqP3hf0dbC0Kx094eJxjGLuyp0y8J5javo52vC4XWlLOYRg
Y3ppX38szL3xl+hG0Chj01OfTFiRUM4mMh1jH6unvDPrHqFM1RIG0+53vaac4FiAUAUEU7kxuHY4
Bx6PFI28vhLNyoTvNd3Jc/RsXzAnbOeNjuMPaXXWNpVG9evvmJfGqpLloi69UYi6RziKq/rOEqOH
Now/Viz6CcHa2lmfzHMLlWLP6KVyv5VNA2iB/BCMO2cTq8pnLWKcfYFNsJqsjq+W+V465vklYTYW
b9Ai8VdTHCaZz7fJ+0Dn6aFS38nmfMaUkRFZ7B4my/aquQ8j5mZ26OqyofLaeazUqFR960mXMSx1
GeQ2vFHo+B9dheJt88OP9DL1yaGvAlS2tHiuz+O+5GB3QIgePp7PL7MMdHLHIr4LAYrtJQI/CNHa
xOKAyVIdbOLDWKJlEgoEOjYXa6swbth+EV2AsZzeHns0RQpc9+SI/AshZEBZKxqYydEgI2SDrbK6
D3m64LNEjtSZpEN2sTgplPvlAIKF++hkZTU8kyZ8Z4N5/KAjFDuDK5xtijaJr/R3IFpBCdWSZB5G
dKQqzSqakkQ5g84jNYNOqkSiEsPbnX3mebZeWm4PjWJLORhYDgcDTilo0VPQXzMDMvv7LIlt79j1
3noz7UzO9wN2UbCM/xuyANd9CQx1qtYBeqPZ2vSVQTVRcVGMmEVlhVnP7ixwa9myEPOCrPGwrnKG
+x8zYYDr3vYfbA0uYoc4BiG3fKVOWu/yKa1o8j+ZIukUiPfJPEn2DTJPe1UxXbYvFHiyYGLM/Jsm
DrfJRaxjr8sAakYNnGftLdB9Ph3zDkEMzNTglc7kdP2NhPx8IhOkY9N55KZ74Hy/LnBUFYdTt7H1
FGu4OnU2M8QQjBgF2kJ81769Py+zFb5CBFaHiwontmk6lhjFe8QQ7HTMaaTpM+N1t7udeDdPeTRQ
MZtBjpLOtkWDPyImZU4KXi2IEXWocJdoi82fOGOxDpwMnBJTPiZvCTGacyjURzLOqUCnw+ylMV+s
ruC6I8k4GYfWtvUw/W2YUr75rq/Bp158HQXSlFzeA4xFIxSL6gGHYAA35ax5aVkBKA5ao/CJuDPS
8ofVNLdgQulkgJ8iLcWiZayUp7AEhy+FbwIogHNo5KScKLc5cWLXo8KHIg9KN1VKQB40A7srQ5lY
D1MPX/dcR5G0U1/HkAy2cebSO5w5u5UoRbW58ONKI633DDKBw/OKOq6D8xUaMTX1VjSHLPUZkQHV
tA7ieY2FJZ52BV/6a254YfXRpgRDCjl9al0kQoVS7/HsrWX/pSFUM7kZjz4aZsl0ew1q91z7u9R6
qx3l9zaEPC6ggp3EKM9fqr/dai03Jll/uN9v2aN3WO0hfEtjTGctPUXzjpvHnqk6d9anI+2+VHxt
PbCcv+jGUw8Y8H7rXogii/uI2g1/UZ42yYBqodiI34x9Jb3/o1oT2K5l2L/jyCRtZ/BqMghgTWj3
BqokUAKUsog9uKNLTvgu9KF1cmV+XtjsuWFcNcEQO/Ha1LnjW5CQC7Ht2FLDyqEHDsR+y7+O+3yw
Kg6D1ce0FNYlJh+OSvRO+I7OjM8dki8Y5O55cjpiP6nLkzFAC9lxuiI7BaahaDb2hj1xiXA63IHd
95SiusJbAdv/devL41Cq67BOUJcH1FUVvylucjjSrpH++qekyhL6e6wG57cX9oKVvsayK4doE0Ko
F8DkWPx7DtyA5fL0tC0/ISxQ/xCW3X0lWpmR1q7g0dzSVPB7cpInL5JTrhVKVQq8DP/Ez3cscZOz
VbXUS+KlzVzWSOne+v98990qGceD6Hsudu+IFGxszDgC/V2Zr6AQ3HOQo366Czc+5SN2sJqCuWMO
s9lv61td/xHs9qDbuSTghhtup8OeuTotUk92etZ649ExXwMR+Z2IOUMwGYWWn8RKVJ5PDzFhjpiV
JmHPn+6ZIkAA4NjE9mhgEXPNTYl6FIUupKSSOJVgt3VQXIr7x9ZF/M5zs6yvcq0AxFUdOj20pbVt
eAH0mssR7XNPt+XKkcUS02HZQMAQMB7Sqq/2l9ynrdKN8mCn6sD7Dj0YOLDGprFVLz5VXC96lrK3
nIaYIXeiWyacRxeybna5PmUrMFIgnCUdIkm0uXpVCZudTItWuhqlMdNSfCGfrajiaAlmsAiR9uQJ
XsAkkOkvIroBoJEUxpkWw3oU/zBB6/Z0daC5y4CK/VXzaZhjlXS7WazPL9G8aALOoS7C6LdpcOi9
2x//Q8E9VTattYnQVGqSnNi7HBtQwMqi8YuAAi1ka9NtlIYmO8znwsLKIyEFKNVfCbDIIQD47PWD
yme8jDx5Wb5/8Oytwp/6PI/enAXb3pXvbRC5LfBfvEW/UeImx8LaEfSlV0qK/+AFgOEBz0K7/Is9
vyhVtG4jet9xjVSrTpaCQTSjJXfHoLICCZpG6TkRV+ZDY9FPUti4eejg3Dp88RZhZewVh9eB6qwr
pfS3ejWhBpRFXfL2XOE8JuwNwDjbhjxGNJx+4lFgDRRbR5VJP28J818pNANr6GdKymFy+efR7rbF
SKxIaZLFc0c+dedixXnHduH89II7vErh7dqC3Ho75GMLR+eReiXlx5BPhd+Wvoc7wAbMVt/ZjPQe
eoEs+6f87xWROWyk8E37gcuTesAJxjpYvpLe8QviQE7MEZfNKZgvWDZxG76emdIRRqs+qKDkHOOD
54j/oc+EwfAS04DspJDjykZKqHbBOw/xKt+owAcO6oiQWcmlgOUyBi/Oakm8USfAUrnRP68U+jbO
OH3RHSzsPVzZ6ywLCbnQBsErFtUqlFjZ+nSNO3P7fx++HalDkb0Ziqr0kyyNe2wwsU/q9RLp033L
OJalJSbGCUm/Epspb4+VJOYzkZhGzFukTJnr6OUCFE3Jq9RE5BVzP0hAPwgdDN9z0TqLVJ6cG8IR
FgMwEVxHbb4Xo95RSkaAx+QgKg3HC35Sc5qdHM2lVb9exOifvy0kuTf+i5eoiBQWSwOnvASwrXYi
PuLRJX87EIhZOENm1mb8Oe0HV5359Zw8uthTHD8E07lLloUVtjWt19HX4h9F7Tku2FTiV89mqsI2
LIi93bniVScH5w5drl/iEqe8tbpNMW+BM+E4qaFoVBFGKrhPc9sCeDYMQMhPb9fkIEbm+YdN62Rl
hrYO6aSnIEp/MfZMQlXfR6EFcwngI8uI+aj0nykJ73QVlUYFQNV7NeQ/RB6ZUu0cYEHxC+9kXm4m
s4z7YGxWcz9/u3X8t+q+eLzn7/GZwKIdHhpw6HqdrqUGPaCqK0FESLp6xqTUyMMWWJEPuNJYb6Bl
zy3cN9s5TKwVmHofWb8XuiC5YIhsyRruxpC0C63M12DiaOaLXaTsqH8/Zj34vYDw9NbL7m8XSEDZ
loHMIy3XxOh0+eY1m+3pfkkfrUAT5noFlOHGpIM3tLLcEtxdqV/pORrvx9p8dFJTs/ig8X8U+6Ik
0m8G1HTdRi7w9/AWXhvEI62w6/09JiFPc+2ZCmJz5WDVhbsX36uzP1BJO+JVvLKlYZUX3qeqtseJ
cyIBdUievePcQi4vEL6a42V/cfC91+AuJoVQSwHtAAR1jQkDh6JyQzuCSgGZKYkO2eBKLvs9jhmm
ska8CtEFyn2jdhox+kjRiQOvpu75TEBaDQaceV1NT1uA+3FYPsFyBelaSWi0S8m7xPDRQ/7nFhgT
i6JAA5xZFNr9x5lvxT/SSGQrigi+8B6QvbeAW/D7gnt5ti2LsudyQy8RhDxcc0BzhobZ4DcCo9me
3EczI1nKBNkr78kIxM+d+Sk/pKTgRQjPwRAILH+MDFQHplKwszIzv77G1loSSy3l9jxsvu2Thfy6
aO7VRGlB3d1VCh9MiWTDNAuJUkgozcMJzci2xSZupfHPx32y0xxR74wQB879zke/oX6mL6OczmLl
0DifiSW+qXdYqjh9uPQ4OSi1/o4KwcYkMQHzdtYPdzw2fO94ToTI0zmHs0GpsCtRLpFN9tgDGVy5
OIArYj7Qyr1OcZ36/LBgqaYjT4h1kvJFb1s9UbK2mUFbj8KKVk8Mr2ibeGChZXeatX0zkabDj2Ca
og39TT2t4QwUVLZZpjLd/0bm53ZQaFC9KxkwiNhjY8zYOQ/g7MCsUazunHBFerUO84vfsu9Rvmdu
ih9+Bir8BrCsXIi8PuxZJ4JbbnFju9AQufOu7r2S/kY5q/yRvA14q7yo0vQ/jHLF11WMw228uTYW
QPkYinP+0WhkpGa+iby52goo6O1gwD2hbijT32RlMQuUtIOWMAgu31fg4WDRX25imMeLin1ZkDQ4
yNypZSNWBgctzUQ+PJ7wriIqKIdrMdFjqxIUbPAE+Diwi0ZeSYpkstHHGKZMBtcQG51Cl3few2KH
pNQ04ctvl6VtmG1Fxcf2sn7O+/QtUqrP0LCAN0AYMVKPB93fQMGc19BJUa9EhNd5guyUw325yx1j
fVrDlAZfIsquYKVAyN9n207E8Qhtg8uSGrmDP3XlVmKAIsb9H6IfM9ezVqcivtEn+Zkn3TUT8gio
MdYaFg4ZRqK7khD4cB2HSGWKWSJkWur2Gmh2owJlZKeyCgwDVWOsT/3DZl/um824szzpfiSWmX8A
bkU16nsnFOyTUJMyRDJ9qGVnghswKDpj24zNq6q/5Z6KGd2fqnvNWtaRBAx0KUgxH3ll2f90exLy
JGotImSb5rfrxU57QH7sJExWwFJEO5jMpx43Vk9FvqMtW3o9qp4nj0mjtCnlsoTBjPii6o2NOHV0
0OdKOlB7cUjFjlhJSl5lhABC8aIGc2MMiaQvEbm2TlZBu7uRdp9rwjVJ88uUranY3sS1GnsLzTM6
MFb/UvkXB66Nb+X91I1mK2sVB0+r/Wt8a4vFi/Y4twv+401b03+WhcofTipyACcQZ+glm6ovR/kX
zaVgryzeLtqtC6Hxm0Y2mGNB/7Le7WnP5NUyj+WKMK8coJ1cUvedhvFKmTNzIqrAMguXy/jJa3Ii
HPtkz/U1ojVlBhJculCry+FTCq/LgmrO0LAgVHXxCE3OPWvXN6C6uvsk/DKH45f2AOnvX3aVgY32
s137+V8ZL2b4nM0+DRd+DNKET3WDWr9AbdQWiw/zNtrsrkPp9p8BAOCOGkjS6qcOzWSOkGe+nbbZ
yBByFjAkf+gAAoCihV8igXMbfqBH4DYC91aBfb0QyTF3tviuZnc64ptMBGG+xkZR4ByQMPJ06p1w
Aay6AJC1MEHpYW9KcaFtuYaMif4v116dD2gsZOw2Ep6xveIfjuS2jRas7lr6+NTv2Rq8oitp5YqP
ViBHyHMi/nQdu4weyLprhISLaIXrPzY3qZbvfozKEXo1oPswzSjH6pbrBaqAjxF3zWbY60s4PXeb
nMKLv9IT+ow5gk5Sgc//QQVGJ5knaz9MOWs6Qb9uwUOCAL+eKwdbO82HLV6eJJxKay50lYvNsHsE
d8+NBHLfOvM8grdfuI0brLFilP7BBfnBzjP58SnMyER8y9unFC/7eCrWAaxsXANPgYQrEjW689a3
mihCFRbRPFebSBuwGbZqC1hNXhJ3z8asizuuJS6SipMYT/ekC9I64wczBRMppK6AflFSgR20pI6H
rJ5NZ71RREPlnH7LmCRab3VYdb7DcA6ldEwad3bLsV6O08vPr6XFX75pp3e/ki+gheCn9pkJn5fN
C2KWRKn8TDeG6I1BxJHi5zLphYfLZSAOLxIjx1fQaZ4fZMfHOmvouahxb2xbA5ZrXPXRFYMx6g2m
M7s3oKLbOMq+tM6ErHIl6EXjTihHEw09tfs4SvsnrtiHbEj0UK+n0GMi76YUo2Wyb7zryN0x91E8
xR3qBmxcljknbtbgJZupOXG7ziq++hNDQRh7tDiamuPtT0kGm/l89VWs64NQZQ/eeFasD1O7a2td
fXrBNKxCtPXAamdq1rA4ykdSgld8MkwUJLZn/QUngXAnuhxcefhfnn0rXnpaOh3lWXtUFMb+SZQV
cbH6UmOiDhjhSsnXbo0kw0faQSsaQSdRKF6pyXNUlTSb4yJefSNXvBkZN/LLuUnVICUeI6CvGxff
7xmy5/5vjVwTLasxcceX10RV5Ayo0lGu+Or/q15jb1o5t66cD76LrZM/7jKwSAhXBq1uk5PUDCJW
CIjtpj+0yZPbmpjosUlyK4+t0T27i6yBpbGb+TNudbraoTTxOKBele8aLIt8LC8/9wICz5IPsDu8
jXZili3tjgDqARiGToB+D/Lxv55oJcjWxPGQhvjXqPB/FIcAMuxr95jEIPH+ZxTweZ7uc2uXmkfH
k+VgyE9A0GaDD85cZUZ4B4P0EQt5LzbA5Mu6pR44IA3cVCuE++yCQCZbKLIIYNsK46elxGe0DAZe
aS801OeMwa9GdmQgWmJhoyQp98WpuLdyqf3/+54TsOZ4zBRpS+EznueudI1E+yC13zsH8LiV7Jze
BVpp5vYEpSoIl7JsOsVRbVmP9M8zA/4ao4/dIvZBjbjeYkCI38fJAJXkfTOdg50XVPFNNy1s7n7O
YuwtvqmtPmq/G8PwrXNKJ2OfVFflI9x1Djy1hFwzCcl7EhGfVWdQHfynPg9tUVmm5D+6MK5+f1C7
9Xb8gtO4S+TwAwuPt2G0OaFATHOyFYqySYuOaQVJ1NgWp3rponmgcO06RAYjLuzw265MVZwm5Vin
n0dL6kv7TkfGmn7g+ozSXUb/8zxaAwvfYsuCWDN1hJ9ksanSAXL5aKGkV/DKDfrN10IFqVnV4P5J
yzrudSpiw1iBFVvxYFQfBjfzDeY+x5feh8TAr9CgcQURog7WU2OxfxTmRmcYZTN+eRVF4Xccnqic
Vu823i3/+DdDqhxt85Ys8JbOPYILYNvazjZIEv/cDLMDCE1dStwtz5LOtnyzyQMaL6kt3XKz3VMt
7iEETft8NTvtZYLm1F6gfRiHocvCEqpVGu3MHN8NaIbK3OGiMyk2w5qiOQ7UjNYwozcCTUhiZTKy
xpq/1h3SjHPGsUIaWG8GpfHbT+qGooo66mdZ45w6IASTYoF3yhypxJntAm8JvizfmT+8PXyqVwZo
0khzPBodvJaetRF/95ZyCLbUlnNawhuhnVWTqDllwFH69Sccdqpyyp+ah+QlpaK9wIeSUZIkoaDu
PWNmc1725O1Vv1qWKUgj6saqYTxmswROt2FCuFKP/P2gSk+96qWNQxczWY2A+tBk2uASp0FrBuOs
xZtZx63MNgYKlGJ7I4ooyPHWLYUGooNlOnmXw8Jp5OsRIRkWVHkMLe+uf3JN8gbfDkXBC/qzAouk
ob+vH+zSfHfEuArvNGgFlam3cqSulh317OXiSKR5AKLJ7VZu404+FNesseWDKU8H9lK8uQE7wRQo
7sIET11SmJbxFNRTwUJq4qB5rpX1WJf5E+me0PSjG/wgSqrR6UOYhZNASROajgexO3VTOs1IVpOC
2PHS/QKV6a3X/sQqRfQN0cMz5udNE4rqy1XY9AVEBGrbSv3HydF7V60NCeBQ4ZWJHQb9wudohuGy
vdh9NQkBTc6jOp5fe8d4xvGKX4ShizcM6aTa/fEibI9eRm7LKDdwEBi+CqJFeoLZtwkzYwzOHpU2
WHkG3rGYY/6YvRVGCem0KERFkmNzjRvT2wpQXUySPF4tkUMl1mDDh2Dl/+UQ/XAuDGfKr+Oapvfm
liESIuF4xD2q3s58/TtJSgHZVluy+tcaInOAkAxsMUVArt44WLAklfJEL3LH8r/Zf4h3k8S41RIX
og2hj8iyTS2O7lnHmkUQQ8UKJT1czWiDXwa2JerjQtQTf7tE66BurKbUW9p+LGfLeAz92hSw2VAZ
57aZAYb98OFMQd5541jmrn6kHzIcDG3pheLH2GfjKyYI+0oUvBFXwPD/U+Z4UKInR3YxTBay8j45
8i7yRRWsDFTFCm+Ez12kcMqgaDgjLyh2fpgPjW+1h4wFvLU42uao3FsxGOGlfwNbxFEeIA1ZLzg0
GoE7arqxKqUuMPyNg+d3/wGerCothehTkUbXQHRR6gl6CUKrVu0UHTXrUA4whWYfQqcybtf4CcO/
/f74CGB0EA81w+FHMvmQwRqhIPw4aA+aXIUVKUj9xEP4pVdRi+igfuFv7AbPJNaQErveedLIF1y6
IBdiH7jABx1VyK2q2Zz6OJOoqN68RhJqNz/szmbRNT14BooLa3SZFjzpAHyBrpQjBoOosvpZ9kde
wbVuBkPMeg6JDHkbbvPWiVZ4OSgMy5knOXwc26DH1x1Zh4O2E4QhG+JlXAKfAk4DdpCaUxsjZwCd
zZlrW+FtWDBqc4SjSv4txWLkJuVBXZZto6x+HHfM9Lwa6RKX6j5VsLnr7EtKpcIrT4y88CfgkfCi
1R1S+ehWkDBetoRQvPbbShccmEYtRrlCq1jrZv0Hmh8OznOF9XyE0shj/P36bRInUAFRrFzsBY5E
IKBTL4NPcWsRM43Ac/1j6Ok1OxFQZVvnKsLyfHtKnYzWfzxkh8cXU2lsvA/vXMw/9alXRMf25KFP
u1krQDkRR4AKRfdTPpoPzeIgaWel+l5ONz4MugV0phHAT4mOpd2GlNJbw+1Vuiy1OAktFR4HP0s5
A9rHTHinKRDSK8EopfyKUYQTTuYfUpN1l6v0URmUKcivZCmqEfqQpo4nbj7NnoOiS4upxZr3NZXb
tuOwx/ufUeo+c9HDWRT0f7qDFrFFT5dpgDZ0At2d2b5fuOII+oqBMcwarnwXUrHkhtDmrhSRovy6
IW8bEihlgnW9F5U7Xsc7Vln9AzaqiouEEFEw85//NzV6rkO1C15miwcrAEhYdzc63rnATx0w1EkN
y21nI0O4bSN8q5QoVWBz4sti9w+384w9bQNAYZpFTlffVzhnOJFHXvuKN+Oe+TJ7re6S3IM9mcIj
owbaRQOWGtiF0HhSr4KT4BPQMJDajmXfzR3q1QKfAzdclV4syLECQhNZCc1p2BvoB2Fdz7BQcn5B
J3A5iV8CPRzuIv3RP+TRzhuCwE+xk6IE3PDszWxbfA9YSlfJ8N4l/8mtg8882coKxsxoQ1cXYI/U
TH5hh12wfuBFgf4lX7jMP5VX48Gl/9PsRRYDfLvVREQtt0jiFdmPhqaRA64x5AgRP++r361C6ygF
c1DZ2/5EBn1LNzTJ3BXc32jqdI1igVbaMrl8/Tx8PmeyqlvTZPlw5pTu4mI0F6DMxs5ngWyIBu60
VQJu9Jqhy8ifGCjpXR66VhLMq6QJEdsgoG19tu4epjywXWcevFFy/Y5KVgLEc2vdRPBNYMhClG4r
o7QyI8mPAvkrMdP3GLgJiIUtqQr05GapsJeYCWeHiFu0oMPVBdQNZ4kVAJ3SFH40hJ819bmoh9LN
BS0gU16e6yjQqmtpFekN08rSXzOe98XV0gET/3I4Oa13sGRrObS0njg9y+FbFgmoDzUkpJ0NVvrf
b6POpNgiKbeiQMqePqNUetKH/722j5VgpCs7ByovRHoWVioc5vzKIPGWayATudnnRucIhBpKP9Rd
2IDhEeFRN7t53L5jEIPMskohAvBMAW+bj1LKy7k5jb5MECNPbXK0oL73Jt+wvj4KjXUDDkV5nCFh
0qjBNkz/WrbiNW7K8z1I3Otsqe6pz2ugql3v3pliIeRCDazkgEtXeSbct3XOJNCTTdFEcvELkPGj
9IKM/6goHR1BTljNnB4PPpO810bJ4aY/iPtgbFESj8Gtk8xiWkDflRLxNddKxV75YWbizv3IGvE/
P3hAyyEIXTn6SnsIGL3R1o2FcjfAm2bCOwGpprCWbIB4sN7G5l6oTqedPclEq/2pzeKvkqyMpieb
kHcTraH+w4kY3oNWMIZka+RoZtHR4S8rm1aNcICbMWVVp4iAl9s1xfWUKHs2CwkJAqfyemklT7t6
gP8FxihWfJmmz61uZasiDV4GpgCBv4/ciU63McWxnTXOw+zwmeBYBefQftmDFjItyMgcOYP5RJQm
hZPW+mLcPNgs+ty+5y+9VuiY686dl2Of7jepz5SXclkV0XKm52cKE8Z4E1RcOfsG2TM0DXAfYoXd
WmyVOasCvCdcuNJSUYXt1E27lkramLYjhyCIuqjVVwHjj6vRZSzd3u6qKsnXc4rpz1Y0XdzhxQZq
Qb2RJDJ39UVsomFlquGPCBpAhZUL8TMPqU/oY5HTca0dzfAmAH5cVcg8aBd0PIjN8xfA3rY8GCss
QcXaagttbpVUuR5zDbI0bAPsui5C/LXSY/h++4UN+1opV6N2HxNfXAVBvdgYlmfhcq2UkiNawdne
5b3/lrZkbwb8KAMb0zNFisdosrDzSkpWUY3j/MgujkJ5g8u1rKIsr2q0haGC4tZ9Sj2rL2+ar/zW
N2Ub45aYW4XR1bISOSJF2FfZZH/4lx5kU5sRatFGvdfaGN2wJZD/9nKMk6Z0/N7rdzyq/nKCSwbP
KdtG75SovFehIR6OnoM4VkSOoH/YN01/e67R+MzPATdTjtf/WnZNzLADhjjYKXaK1bKg+jxwmP3C
6S1+lBR0x0/uhRE2bDiZIAwByAKjBQWjV3K2ez9U0FVAXjZaLHV+lswQkwM8S8wN7rQ0oaR92esq
lg9ZepNxhzQgMd2/bPYmnE7eoWNPpfmc0noRGsRYTqQSgx2K9CmHeDEAuz4obbg7ZpJdirRJiamI
tQrfOoXyVitRWTU1ahFCKMTsP1Rzx6pK4vMsV3+3+DbdjQyw1skhJ6t298NMFoEM/N4v3TtKSLxe
zAoouj4v47ZgqgxbGoUNYJhKkWeRGoKbBqwcvhpNypLLT44V8mPe/kjWlTWPsGR212p/HpQszEQk
CD8ECjCSesoKny9do5+5se6MkgYBfxOMZqS3Lg+GIhjJUqa1e2oj2mZz+/S4M3O19hT02aYP37Ns
nQSGNI8fcztXpZ1vCeNUxbjxJiQJvXrFH5gjN6ybmul79AmtlcZQi3Ptx8hbOlXe9hURavaINZnB
nApWFywoVE7v2N5iJlwnEdg03EJmeReevMt3yXOl35+P8odHyIOANTOScRo9ROrrl2IQnQAoFEnM
bEYQkprtB6UHrxmX0mplNfrL5CL+RQA2ArQaq1VLEUGfs1PQeZ8KYjkF5ths/Jw7+q6lGKAhNHHZ
fjnSMqWOjrFoRDD7FHK8tY2fOE8UiDgsqppXgDIqKRh9/+Fq9r5cY+5ecMzqJduJ73DMC+bIXxeE
8GGVHJSm4q3hFoKJlARNgj4MyteWxCUVLsl2EE7Q7hmAoMAjKzSWd5PlnfPn07dmL+mN3eUdtyUd
aVByhcfPFcCnBUktnvDxmdcacHpmN1DB14nMnu13MjLxedIVX4kLQCbZeJt9AtmbYdxYFN/LIGtX
bBy5qsH9t64gynaPiIgBFcBGjuvph8zc/aDWAfYnf9DqDZwzYJsctGoaKM3KnAhhqCxloepTGvlS
lPNX6Crvmjv/YdRT50aQCTHbZbQAQoZFOXSHfgRv6ElsrHzAn1pwzv+wBXyp+b30loW3fGD5IaOV
3nMS38yXqiuRtqss7k7EIZ2/G22e6FcWl4MaLEQOLOJirMyYWpSBgrN5wDAY78R1vQDDgSOLg8Cw
OibZv3uzkeM0Qa+0DGljTDVqc8fQ4xUBZSdIAEdCXYHmwB5diwog8kVKroG4lvTursHKNl++FeDk
lw8BrIY8WlwSyOXpzb2oluZnPq3Jfvzz947zXTsZwJCuWH73ifG/WhirG4gynnoxkcF/MnRcun/O
bucK/I0HItHPN9tWxofRDFkx1oWKgIedcH0Fc6UFMyTtHw/QsgcnrQZhS+b9AT3wSWoGlCB66Hc5
lxVOrx5UlNlyEps23ew2ap6v5vuEDbRZ0k0hPYPcRPwlpqvps7sdfzhLZ1VWQXMZodmSdJloLSW+
zZxRyPbQ13VbwPr4J5d5nGEH1FwsgrV7YnsD0Q4oAPybkXObhhhY7bFAVmdsKLEm1KNMAp4+j06x
dfjrx0xacnKx6iDhrQezajuKO9LE1W4tbnLftPm5k4evQwimfbHXnf5xbfpk5vtWvMI98uyUdKMw
or0qOFsvKJVQTjuXuy/idrjYyhK7JSpyquNlUqdaOmQQVXK1V+bfE/J00hoUa4AQUDWs3/Xrdsg+
X/a1TXKfBZth/QF4kkbnCUq4K28zeQRmm+1JtJcOMeMzTUbM2np2zwlIUTcV7etanvrX+Qe/TDPb
n1F3mIkwGSIp2R276nSgs8dYi+BqdVWZPLFE0TnXuM079EZDvPlbacNuV5qzNKFHr4EyBvWPxrVZ
UCO9wz32wlK5ZgN8y/Ln5EzmgyyPPL8aYm/xjJ+Wd8Pm82AYgMI6aCEF/zQPs5dki9WJwsLhqvMJ
livvX2wKE37XDoBbp7jLRkfliBeCLfgeu/l8wYjV5IWW8+iGZ4zxwYq0oqo5nZQYyOxJHm1524hf
LO0lPeScM6FiyeHjYU1zTPw6R5sULAjhreG7O58cPf8plsDlIIgG0+pH3djDBhxIi95AnLdtq9Oc
oBC4vfUvOriV0Sy9W2S9KSVnRLsnmaP0HYr93TyG1s37PQlJjdeu0Fvj+UelnmJy849YmdZ8TFVN
ZVXbLjEkrKLH5mF7WdmL/Nzw4LNmoUYqYhoz+9dd0n/oEJpJDGDDm6vr2TdrjHBLtTSmM0mkx5bE
KU15KY5M/zyTX9F3qmY9q0cRqczX8HX0nSbHlSt+5zfxjPlAGeP/mVD6ua7qNKgUOyAV4CImYSJp
uq0REqmOmlwELQkM306jh11EBqCsLt2cuzPadDAKNTZu05qv6w2M255+gMOahAbiyVsimNzF4r5n
Z+RC/IgKBpKpJrf7w8PnZFbMlKVjUBWKpZaZtwAdOd7/Cw6Yn/Soa06S7txiQT6atOHjqRLJ1sLT
wMlkoBitsexpcO0u7DdBslk57WdNafryWZi6GwVSelFGJ4i52r22l+c6J0p7fsp17K6hAAalRpZm
yDjMPcKzi6abkxDsquwP8ILyCMA/nHu5x8GiAvDitPNlPy0fyaZYPoeQBObH4kfQ7K/kel04NIey
i1KrXsLmz4a823gJZSFiDUi3XSO+VjpnT5NkRN/3NOlt3cCeLQVtGRJnv6tg32w/etXN63Nkiy/p
NSfxwHEdhQthVReSz/E49RySOz5L/iT/NMZNxtRmVHBAputUzfluZ0iayA64N7t95lMvyh7ptpts
SmMwaLOCSu5RyngfI9s9Rk0WioU8WFdXMllEDUP9F+NqIEPmAkhVlq1nznOJ33S+NQ/XyDiyRYuE
8JNvCUVen/wYGYrhwmfZYBknOPOAo+BaXfUcT/3dp7ejFZbOkdEIKO5V0tIYz6VWCHMl5zcKhfNb
P8yf/a/jrPE5cHGIcQS+2EsekSvHBjqew37iNxc/rQ2KG0Xoau2ZNdvZBb/0nvT1eyhs/hb0VORd
nuW0BYH9Eyw3PUfmODX5pxG+ei2P+jS5dhoN5ODrOveJDX7i83IiZhK6tKuqFNqPJSyTDnBbsWDn
YDB4omU44vzP0wLHhbL6awgh/pJEHc1dkC7meVRtqDy4v0OtizEoGpBf/ZBnUq8oKGNNRjYWTII0
5I7y7I7w4hZA+/w0wLUatGbceiD72xOusrnm2VZmhxdjlxt/pXEdMhlYX2FGfj+AE1GGXH1wLxpJ
bFCLfID6bY4JG797Y69+FQlNiISarY7Ly2COwXEofJs/UHpZEew7FlMNvueWpi+iM+G5xOWSc+9A
KqNJAUyMvprGN/CNSFqwWXbG30WdnVsb0A6OM5E7HvR5jbkCC3FRc5SALVN3LKXpa2NORqPNQe/6
lEIPdQBqBa8lWaQ4eg25B91XUMXZlhi+VpCjPrHsfrRQ0WT6nMrqGwCLU7jXJoqvQb0xFVnlZdfl
bF9jVPSfTvefCRAUkfnWwh+HTBeoljOuM1xZtMUxyNHHJYpHMZjE8IIyH7ixZwjC8pCw1zuyzviL
8+TfhrHpMP9w7a5CVA+HvQT6EXVWRVu00GhvzaQrvRqUQEXB0B0dCSQc7NrOePC5/OfLBypFHYit
z9crFwtusjf4Arc53z63vildGGLP843vIW1BdTbdylSC6Zgkscwk5oaZNABDJ/KV8PcWOFhTW7D6
kbXjklLwHf9og880jYatAQwqYu5LhQRP/m5wQiGmbLV5jhFKcMh6HLATdbfCCZuYTj8WnatrMNH4
YybuE21T8d+osYsWL4QqB8XMAZa+9ooYB4fAjsMYAhReo4wHe0n/Np0fTlllqMoOH4sEKzq5EOWg
wsPGLnMPrUOOLygnPBRwScjO/bgFVOw6xIRiKi95bFuxeOpyBI0e6BQ82ntRhWv2BBwcyA1+An7w
vau7GOAXMcvVbpLs2b36aBWtWHjHXFnE1AVtcR+1QB+5/0wJLwJVlHwhndlGUv+FcTed+x4CFTP4
coAGhMqApJ4ZScQwhqc/C11qUTGxWnBsR1GszN5lPJLDEaCpx+g2Dwt9ne/pVbRuxrUXSgz8OVx2
4uhQevLIiN6d05sWw0bElrmNmkAZQuHG3Mkj7cIQ6otGUh8Te+t1MlzmrPOvmiCkHaZ7x50dPtiD
J68wt9wGKozbRrQoJfq2rXrCPcECPJ3mJDjGtj8bt4OgJjWpYsKK7phMliYKfbLf3G6KCovROJqb
WqUOQXkTy5iJ2vJzlALRPCeuty65F2mkdEgcBpUC32xLwPVq3btx0/D5zV0Znza5Hglxy4uizi8M
CATEmMnGIHnCmcgwJbsbxrJSkH9H5ik8df4x3FgS1hpw02qIl0lag5kEfOWBMP+aO/Jo6PEt+G+U
HeVNoTx76+i4LQK0pMKufQp1oDP34HS6XEtOb8S+b6Aa7seTwzwWjIXu1BtT9FQ0Md0uzyGO03rn
R6X6ptgtTySPgKV+toBvmiX82Tdn9ZeB1IfDZSr/IlsVObDemByVWIGUhuFqzfmpmeARqDMir0f/
xVz8teNTKLr1jNYeUr4J9e5s8KBqp8ohoT67NEkr2LQtD8UM1//YZNxHXgDnXUNVZ0gXYozOdeHI
A/UMtBYtbDBlwLEvhx5cT9xKT5KnqIMOpOGTEF5dSx2TD73INRsodrKn2TB0fGjLqAXKmdu7ihE9
bJJ+ZGqKspsTI4W94UZQX4ed0iQUb1lXRpY4sZqBMc8ZSwKnVmGlSGMj8EXMcId67uTa4qgUmEyI
O1r8lA4siaYMHj9I/zMdWLlqw9h6fKR3LBaKd5A6XWNDNsQ4QF970s9SuMPh9xPwk5+ixHAs4J2H
BrtOkAPIRHwV9Scs6+UPW/kPTrf/WoR1e309J6ic5aQZtZ3/PqGi3C1mnGVdbeA8ieTrejAYaPte
T4vCUvNWVospCwbF11y6YvKZBas4fIqEiCVYDm1HU/7vNlF6ZTqVRSfhZ2LAvih2cRoECdnAIFUM
kURmQ6pcMSufVjk5RCBx/Lc8pgC3eKCL5jnflp3USNpU2Tv59FUNMonkl9TdpHJwEFQjtWBTHNjw
FhEZ6mpxEW5EXGzO2RxpQM9zn3fDht151eiZgPLP+6wpwss7n0lbsssaFmflSWjZd0YIiRiaRePo
x+VH8ihwyw8yEmJwY49U9kFqaqwkraBcTuiN/hhNnGAhXgOpwJl5gtv+1fGj6YLmDFNjGc6Vp/n5
IlatIdO6PBeSlbPx3XhZCpyIOL0muX1aba5kDaPnYjvYfr9zZCmY1ggCH3EaN9IHTp1QhV/OjzFe
v07oNUecU60tfelkfr6q6lTqokY2alcdJIoI2s6w6jwNXC/JWerTZ9yL8PDbF4Bo6Lkxlxtv1vl5
eal7YMmu9g+6+qSmn/7Ly2Tn3Sxj6snSB4lf4nub8EOWvnJaPdk2+I4uFY26InKzsGpIXM8kk643
drB0qNSzQtn43ULGCUm154TmJvZcLUbSBJvrbv6NFhMzH2cFWD+bjsdXW24p8fmeSb1kig+TngtG
4GOr7ftSiuKAdUi7NJXrnlG0Z4D7r05WGt23ghJZ48YLbnbzolbDLfq9MOLBtP6lP3YBwc+zAUfv
1LMcH4GCR4161bs/BjJxI/b8r6g6EyCnN+OF3bWtiWvhCdVmEoGk0wqKs00XqXn4JO2wz1Lep2Lh
hSEL1Mu+bXzBFMGhCdKnU7wCI82KJUeMVROGx9Db3oFiYUVKv1sGQ0TwXkCXCx5wTao2yKPa6pfr
qdJNyHbv+u7lrnLlv4IsuLTOnP1+slCTosGHCWHTF9Im+2aE80aO/GThzykSxyHgh6DOc0bIBRe4
82O2a+jWJu5Z1xTWv4NZz74DuZdwV/RangfN3DOSluRkvrAuLRT8Hm0nuufoF++pl5ib5L+652qA
U3kDpJhVGOGkYERCBU719kspX3EzbSPXMQbNWayHffjDBs9dAHPsiUfMqPHDQkX1oMZVuusJ9TmJ
Y0Il5feVgsK5g95ijBgd8A+EZs8gxWNRffEOSvHC+e8o90EUPa1ee2eHsGZcUN8dTBn8MfTpfq3q
1Me+YdahjW4YbREEoX8SLFGzZIznk0jx4QuugY/G+yZXv3n/0SrI+e58mqm33VuH+Dz8DJwoee3k
FlG3br3EH7Zt1TLyEg8wogat7oy8DnxtEKTbBdsaj1MMDjWOMu1Y1ZSL9aCdWW1szd50/vXEC5Bt
Ta0q8paJIg1czlU85UGhqvotm8roA1ImjYd/tDMuWthMO4RhVUpwhSGbIuXXmkFHhSV0slj3Hwqi
c2NAiG4nNI7zPGXMPeI6squLe9JTeXcnFIvoRDld1TCyPcT6XoYCVVz9VkAQFOsCo4l6pckzfbnY
YZwEKeUOyugaO9bTCYIAd6htZP8tN70FK52lM/9i58Zcb5wkVb8WUMaw6Z3sUFE8EFRUxdxp25t4
GxbUZHNNR0RF/StoulbcKJvhxzkUtgpKcAgydzUtTyVa98gDRKCxgWgdy4f5z2/f3rsJc+VbAW+h
Z12PyGm9wVAe09zmweMyoIDXOMD3J4oPVtPUKKArxqO9Z5tLfL5YnTcPSxUuLq1TEvmsLmTKFsO/
YSweZ7iC3uBIJ7VMpWGT2q17/JtB7sbrTlhhR15NK/+0zv0BgR+F41ibo5NBxWCo/cIKdv6alOiQ
91EZjeBA3qLFDZlcSkJrLc7jfiu3Um/vPe+HKguxWkipmViiLzjlc93LXJCiRYKARhza7t+LKV3T
dUhyrY0RqZL9+Sf9+7anSLapDPnuRk+uLLZVmZOGKBnk3Lfmxvh2xBGHCa2oVs2ABi/CIOYbk9m0
mK05pLFSDvLJxJPs8gN7KEy0NSqP8YnsNXCJyo2jXrSfj+380La48FWkK4afo5hpAvpBizJ98hMZ
TDTxtD3X4TmuJgmDwJF/F9BHo5Lm4Lpq5nfBsCB8td/5cOAosFXPSkKbbj5my6a/O42RT+X24Y0l
2ypWQN2HFmHsbijPuwZo+vonWrXZq9Vkm41PgS354wJZIc5oXPSq2+3SDVWCPPRYMoF+HxPZGwL8
NCGNRE2FeGTlqA3giFHfk/67yQ1UKE7EQ4LV3FWkbmDNU0IjY/ZfFSpxOX1SB0sTgE8Xd0RpxU0x
AxFPZgDHa5P4XuMhQpBD7D6CWfl6qY/YA/k8V/M4P31PntZvhg7gCJgsl0h61Gdy7qee9KSBsXrp
kDTRZP5kjGQG1zXCPOjO+8BTYKOD/peLDYevNZO5MP7WSBGbV1CkCv1PNB8b9yuqqOSOqM94AYzF
+7vZlVcuCfmuQBFO5pejbKVodchpJUOF8NORtCKMJdGwbVjOwksQSLX/qfZWIq7tb7MeqP0fZW73
O0ejzKOXCm2lfKtMIlxc5gdOv2qGxCHRt5m1H5Hwx5JajqLlRbiTqPu5xd1Cn0+axV/h9a9rrEwB
vBfHvZND8QSK4S7fh8tcEMH1Y+5qqFoHw0W4+hBjsFPeRS99UH1N+GuJDTlHboqQDNYIdYpWGnEm
qw8JFZJk1ZdceyGO9kOQWSwGw/64NY+Kk+M7WROQqx+dDJMQ2QvWHN4J9CzUIB3CN4ut0bnbJBzT
ufU2Czj9tleu1ZN5knyvjy6cThQSNGIfnklxK6E7sIx/spRShuk1/OWf0wtirzTalhtSZa8ZDlB+
QFXDzIOCmLl6jP66yrxIpWGM7Ix9oCEpMWdhSS19d6pxYdjiygulBCcSBcLGbILdmsVIIwOIM/8J
HeRN3G/HMrvR2MDFdW2CBK9wHv3OcrAHsO7tG4PoYqEorL5XFOpVN8SNX46aVj/TjCDE5J4MYY6z
gw3nlO+tMX+XntDXiehZu9qrs4aKTN0k9ovx8b5YRpBv+L0UdNGgHafcDn+eMJ68tJ8bxWw6AnvC
xN/I3NZLxi4n07DMLIzLlI8/zBkAK7J44S/gf0Z/4N6I0RetdIr7SG7RbxjD0PvBRH9Bmnp+qq/X
5OW/MhHcANJE555zEjjeQ3pUEl3gw5rPXmrCTC9b93+D/lvBYw/ridzHClyaygf/xCGAuoWbpAcn
EIHgaX0LDJJTyidyP46tUnBmv5gZHN2FBpwHpqE8ncJt2UjbisNom+5XdRIgEQb8acp1z9TSVky0
QYdqaim/7Mf8JNJAoW6/acMLfgWU000V6rcqXGlYLt+ku/cwJc6U+EMtj6CWquz7GZ2t9brMonET
/Xn2qlXqxYWq5MSR0YpdoxLzhC2+s3IAxLLgvjDhnAuEmS2uVHUyLcFiOiTMilhvwqoMbYGCHYLc
acG/wIMRGTDXZSksVMWPvCiNDMBu2sJh8WLKmFYVjKLCf+gA7TUnHNWvxM8EFKz6g/IxsBjC9LLx
YummyZRgYnXsZMEs/+LZ0G0V+0AU6eNSeDoAw7mqkWrSLhT9xAom/vXR3VWB8xyXrlHlRhD7/+tf
J9KZstwi0VAOA1j4HvSL2CC/AjXpRL2mgqCDhTJFPqKr07/O1KrjgropXc3Oh1UOGdUFBYB/x7MX
XhSDE9m4GPkPcVjkZtrG4ZpyR5gvGRzeul+S71sK2NLQCwoXCN1zVxPY3NuBP3qq60pf0Fl0sAv0
k9qX8nWZqb8ktMBrI0ttViecoH3/bLLwFrUnVhuYZJ3UqiGYD8q2tQAcwWJZbhPyJ9F2m0SXoM0t
HUsF/t2e1lQgJ7sQ4L+cDp7T7OQBvaXZf1D618cDq5ky8NwGd2yuXr5JORhwGQT8/XdDGIXo0xVS
GMBaeuchDY6OLw9W9oC74MMDKCldBqvUYFF40nRqph9lm8ow1GarduG764ZbgLxAiA693uTJ67+4
KXaRFUeTnb2ll1q3gR5DkuAMYAvL/Epq0OxxLwAtVIwCGKyCNK+ZUlItkrNhZ7MVRv4eCKRxuVek
/j8bGuUDTxSsmOS3YATR/CFwJYvoKJ/kQfrYf3M8RZjpckOMwG12nUoQX+ui0Ml+bBSS5rIvjPTn
w0barnjf23SWc0d4fP8BTsawhY/oo/OI0/m1oBQbmSxwS2wBEXXvaKJy1xVyR3hDPbms1Vp8+CTg
QXUJPvvAXDRJkr9Ui2e5qDk78/RHdq4jk47VqXQzu7CVHCSOuvDONJyRDKAPvzigJkBqplChlT2O
55vdmD0oKIBl+tjYGaqd2S7Dx0GGQjcBaLRBa1yICXNkfyaZ/kx+55GsV7l6qgWiwDt7mMOybvpu
ur/FVh3xpBy8w+mDNsCOU5yk0KhoIVimz7dCcWgQZ7LkqGxy3vDJBzOuIRV3SiQW2nNMmUdkSQrs
hwyDlLWbaJ1or/EUkxYuaB1Y6x2BNp8YGDuQDeUsHfTjfPFNXq+cniHDjmvrHZcjL5ahvys6rwHm
5LuLlgS/VA9T/zVV6Vh8I9ZV4X+SwU19638tfiIRf5ogMhWsDYCk+X/Afatz+VrkNgqB0Vy5H4fE
uYg+unvaHjhUS2HUtX7WnDcDffV5TRYgyg3tbGDkc8OwJtdJ7c9G4xO2A3W6FbRcuEoFsGB3jJcj
GsnPaaTqgWIZBCCkER4Jte4EgSNoe5Xlk5f2VTJWAhGceQ5SJyOe14tDR4SK7flV+wRmM8Wult1z
3leN4c3sWkV2X/IT1GnOMmqTicZtZqdt5Ey39CopxwfKNvFTXl2vNLZ1vRqmLNlt4Al/PRqCvAnh
RWrkwp+YKGuS8wzNtJulT9u6OdBxloq7jQkt1l0GtikPV1WZUHK0rnMOuy34XXB1o58cTDBksU0n
SgN1w9KBHIHHOM2mcPPcK2UIYG/Ogk00z93jTKf9nj0wcZ1dC23umuev7r1GFKgc3drvHQRQcHI9
ONszlkQx+GvlCbopLOeIkkJZEylemK2RTvZupkqsdohsX+45D/mQ6GzTEYJyIqELfiNCvLfELWce
rs314J3Qt72tYRAho/U7QeRZRh1T93/9+QkU3MPU6ea6l+W/J/WaoGzykwq4Sq2NyjOK5mOBg3in
yH//Hn7zsj7lKKM07oEW0EVcvETMGVDlipLjSIaYmkKBLkCMLZVQIfjOqj0QI8A4cYZ3iIWyZYtw
VsouuA3pgDNNkeTYeJQk8Ym5cKYg+yQhpdv6sLkyJBDC63ptX01thI6tQy+QseuTtjeagmv3JuQu
VkXFcWEk/cJkmBSqW8+xFt2ZZ0fycjtMRieu8tU6pMNZI7B0/EuD8BNRPWNpiykaEcN+kFpqxIaP
uYG5TrWa05BfGwKie86+cWUd9WF4ENY9zRaoRQMrfxw/A7bXS4+NjScaCqG2YolVndTSpkpEI33/
pDxReIKZMkUFEI+pQ6VvD1J+6Lq9bXJ3zNqgGzoBKMisHMISQR054cYoJcOv1iuBUKtBhIrghjj1
b5NpH5fnxifIFGLGCtjUbpA720RB8X4BBgXZNwZJDF2Nyoc9J66uDWXDtDJ7L+IyH9wVvQx4uhfd
95k6bFKuSpkJwwcwDyvQQcJ5k+pt7TLk/3UY1RxznPV7Hwb1vhE9OtWtlCDmKJESvNr3vjsOOHe6
S84v7fz6fCTA89Pl6F0KZfslgfH8F2cezJIz/evK89Uxyh49SqS9rGy1HWYrYAj6hrZqAVaptC5M
g1L/8IQ7BshJo2lghTz+1oXO/jLb50RRKgHdl0TDTH1d/BiY/cLyqRLNpqlqHCCxwUQOl/T1yAA4
vAO+GbfO2f6JStkNE32vLSIP8Fb+9b5eP1OGMCydiLZnhs/+wPLiBDkAv0pqsSXjenfIj3Ru0iNr
da387Fi3EgcmLQoBU3Gz2E6dN70ZGc7PKC6rXrQA9Tmijjccu5eN5X1CqSjTHST1S8ISELlXhepX
4za6ffsLiuIXWLoKdGiCjLiiNXBydU/ZMlaAJaN9n9zQ9jwR+LNUQfLYEWagcgb/J31IFQ+tRgeo
TUVm+pZIlB+ibWsYLs/k/0M7YGgnX30l44j+bfdFnTYHqv+rlzOlo7LLw7p+E6BJWhGENbDnz/u2
PGD1h/TltGsgWeFvDTKQ312ii1gN365tvtSuGzVJUpHVLdkWyKi8SYfq8yZ13XMiwjDgd9x8mDq4
VnUDt+mlJDXgZb/1KGwi95NWzwsy7pyGLFzKBdPN+f0EKZiejHUjErMI2cKfMi40cYu1c5moDwQ4
iWf2UMd3djSvDRWF1XufUGKkyhykaKyLhbqZq6iKaRnjvGba1uaE3KLzX4JV0LbknHcDwpdn4/5Y
quEHAv7uLqxRdUsPflYajgA/cRFwZKOtJEzc4WO/AjLKm6HiwwzRCWN55d1j5I+UqLuozUUboKIV
bVW5x28blbSdxkuOg16tFlZSCX3H3amZTnm3ypyNsI1ixUV5dMSvuz6ML4LSuQfKw1zEZyva6Bjd
yHk7EewGM2g8UsLEUzM/R4/M4JfyWc2QxM58nFhGIuVzwMh2Hwg582Q4ieFGGNlkzkJ4fOdIZ9Pu
Qn2XFHKKJWk1nAugACdAqM6mZ5zFjYOro748PljZhSbfuCFhpTscluZj7XbuUjXcbB6YMJZY7bDh
8pNP0lxJxaQSVknigirvTrlnIOI1/+TOOZzaTgOnNvncJ+NAZ8I4kC9uvIivx06GIhDoBo95OGR7
PmEt/S3P7klxVGM3Mu2D81g3guUCDJMr1n5fFGLjDiLa6aRS+OT1YFaAyAr0V5dKpSVTZA3D8BZR
2H+3nMuprzHW6MW1UkX+RsAGcOQHz4YT38k7LYzxGnm9aKetIPuVSCU7Qwjw3M+zo7xwLbZ1yAbP
UiesnhZg2VjQ5SBHd+HIVjcl9sKDMUu5yTolHQZ3b6sIiZHpzKUoOr2k84JAzQbQqiW3KANpqDN5
0imFHQt2DYnuQpXTFVyO1DEh4qx1F6yICBt5abL7YIqF/vUr6jioAXpM6SK2S8Smzq1DmrOHHbHo
YEXCImoDz0+3wg8QhX2zxZSZiP2paLEj1NlYnzX7XLinjZq52HAKlIqwmPh+lVpRzguuufSBDdRM
5YL0mTVgkPXyeX33i+Pmn7zEI2FmLkejyJs5tNhTUecwA1iYIN6u4IH5WCjMgpEfG4SwV0OoY1Fc
lL12Q2U6hD4GQNSGRGms/D0wq//Sre+LmNhD4K6HrWGwOBpu21sQQx3vCoFkBxO1ZMLWDZpV/HVt
pfE6lGr3Bdx4Tq3AkYZdYssxAOQvMT9oyyLpiWWktRZukjIxeLZL2BW3R3sA2M6BcJBDVNvLWiyw
Uuo+rhf+TeP77nkcQeExGcx3XYuu6J/F2ghv8a0NzceMEgNzr4rhMMa5ZEiFfJVh5LWeTJJpGOgg
R4/p8WQogcXHLooyxCP+dyPNl/YJB2eLrW+BE8a7mECQeuTArhj2dAHqmCJydWtTYGJf+lyjsEQR
3d11ME9aYhK2DclilBzImwH6EyvPYqazvxeFkOacF/3Rj5jQ7OtQgCHUcubPZ6VbM6tqkIwsIcy3
9Rgq1iQchjAeAu9WeCuW3lv9npB/dMpLKtVDlqG/rzEE5ESVXLVdmad18yzbJI+RfoX7z3Fju6uK
bc64GZxr85J5MVgDW5EhNL1Z82zpmO4QZ2PPIJcL4+Xey2Zb6ACBJzyONLfO0zKD43Vorg4T8pUg
TnbGOe5PfGu2ZIwYgGls6qlcqzBpz33+Io656BDcgeq9SR94KKJ5yKpEnT2bfCdC6mYkwko3XTvG
FTrMmKsOph3rDQBwLb+Ve01RWqpn/aeqHC0o8QHrrEVUSg2mFI2P2fk0YvBSI8DjbfS0vxuEEbgR
MdnyQN7kNYSqR4xN1cLdD8rEnWY5WWGw5SAa9WvYD2fXKpeg6Xaiu/E55pg0SP6Q/ryyhbaSTWzI
EkTiIVhWg38Ec8KZH0+pMK5SKPuq1pyREHs9ta41w/0D2KJjqwJkU5RDnU1Uz0wj4Ax4f213yaif
HZv814fTo3QyLosdms28MVio5h50hwoTDRC43wSGzcSPQHIZ0/ghw/Qp6EOUGskb2lrRA1ewpVJv
cwOEEWXUngXOfyPdc7SEkdPx55Zzl/T/h+dYWD09Wagy7xaLAhsyQq/kLxBm8NxVXasG515pTZv4
gkOmxsseYwKVyAj3bv855ZKPUrgaZQAAWwF8CoTPY4/E50sqy+BVFWercowvGsT/1KFdyEN1YzM2
VLJaRjoK64tdQMGztjh4LEeOEQKMkyBPgctAbyi/x+x2ze+QPuRcpLa1aGo8GSZDI7CVLRQI48yz
SraahAOWh4f+3lHHlXr+8lqc1IR/PbhBP72tWb1RiC6F0P0exDSFKOmyKoO7Jg1wRuiaM0/ngZgq
hX5jA4SioUEChO/W9lfbesskf0gPGIc2MWeWppa4mK7H1zbTIuje1OKp68FY1fgCagg+8maBeeH8
Sj77625/mpNd8U0iT8uC6PYTSMeH6c7Lnychp1IGDBTzNnNivlOcsXFouCN80Wak4Kc5YTA2o1WX
0KyaWi0qNV4r3E15o9JCkHTHCcFn60EgLlQ8uyf5QnKD86ffXoR+6z96kVgFlsJ9M2UmElO2lRxM
L7ApGjkUqFniToiY8RK5lpw02lK+jh9VcDowju9r1KaDgWgI266Sd/91dtT7RH6Z2kxvNLOIGV0M
voGj2AMWWRZBJa+/2CfmlZOiEOvmCFn+aSCaTynJnDR0CiBjsdFLHD1/G1YH83Ae8hwqAlIyn1Bk
T69UmH8t8IoCTtJlZf87jTmIg+YacqU0o7IhuaTAmBHAdL581C6yUhGwLfg3B1SoTQXkilkWyCiE
2XLjdlUN+3PpsnetGT1fxvPF4dT8/mblwdtGdGiGwi5CbmgQLueO8wsvX+leX9vFg0IQv74MDuwr
DP1a76AZkQMuCHOxvh00XdeZRZhl6S4jfHPnxdGgQ7I5Rw4HheCHqFTz5cTd8eQY3kyTRBV21J1k
3HLPF/qsZR0EOoXO4Pn/qxM5/jPOqNTOOgiFhANL82h7wQyTDUVslEieG0aPTJA5gdfTAvThHEKa
76PjRiMYAIUHRa1CBDL5OTkcD0ppwsEFX6DuBa3YogSH4on2f7bmuanj+czK7crqnqAdeZAqa+da
M6zqChFW4PP+g6pxlnHk3vAUPaRiG12Sl7McDhK2hP/PeKhfQEmMQ38QaZrukC8h9pwFtWd93jqP
jgPu+l8Tl8kaEvF+7VjQhjxD8DoFDFvN70adgnn8TlzQwdygdKmSDs1/Mj9R7zJMLPcSISbJdQq1
CUvRynJh0+alURcOU9C+ugiu/bL2UnEy2y5/c89E5NFmlcYeoIV2e7LsTX+XT8SSV/wWeUYKqgbH
GnCFPWu5KU1coEdMDrrqc/9N65f/3Xxfa5olB68G7udP4UXtTexpSFAkK7FZJ9yamiw06CValmLt
xDjKEe5+cn90F8auqfhjUt4qkf0UFzcFwMkAjn1d5APZTDK0fA1aQ2UQCra3T9OcUEc1MuS7Y7cz
1sI/+o9J9E6eE0JgaXnHvtjZwxscG8adsDF5SQcCJ7ZV0geSoNHLd+FuZf+NJmPa5dovciCAeCaA
T7Vy8l9RoeKOIezsPVf3+n5wA/hiYET8P7ZQO6y9qZ4UBovm88RIcYsOof4915N4xwSsArZn+38S
nK4aiTj+MPe4dSTrH2mkMxc2WGg8sJRj2pCWYFSoH7ZAjDV1Ijkty9ggjc5/bDkV3U67khXXquRI
9lTZ5aIcfa3gC6wm724kzyA4aD0ys4cK/3uya94KGP61i/ux+fn478tm06+gaW7cIN7Bf1JrEsdH
vVWMq7qxi54+mXBKc0KXxZ1HHzg1hOgvmNRuojgeHlJQjtXNSL1wfWMWhtmwLX5sMyJ+WXzT5Msk
828hmnAFrNJqta4v2qoMir9ncNza1K9hJvD5uJnBYbIm7vOIm/3ZxRt8Q5NulfL7QqhebOEA4JyQ
KL+jgRgykO7UWIkd96UMuCkZcNWsGdlxkUDsnZouqYVsyDOeW4R5xHDIk5nfiOTCmT00rPqfR3Vm
CGbG2NZfAj7Z+/dx9KfODVNoJdiVrzJ2WuH/kTYL0iAummRNwNmC4/DtCEJl74Sm6VVsRdG21eA0
LvABH2obs7DR2N3gQ7k1Mlsdh6DACftwQ2Vl795+JobLRbe16Ft9efcSoyYCPfN9waDgKjRSjZVd
uYCbMiOzmu5sk+umF/Lb6Kptgx7EFBHGxB6tHZwo30T1IzkGGek2cHIAOatRyGbFjPn2QvU0LEBX
SnX7Jg/qhBr3RqPlyoiGMGqWNnxLkCT0p1xSLnx/d8fJ6wJzZh/oTREZoCd7K9p/mn36c8IEbEKx
6uyt0NvCSs2So2b3D1mUx6wOYaSFqx3aHvnkMXCDmxeVLWBeCrm5o6NcJpV4bWF8CdZ5wSAP1T+B
AQm5ofPNuS0nflB+eYmS62qd7P6gLwZ/GjzG42sxCft/zmNJ0PaxRpTaafLCYYdevDG6TY250IC4
XeulVpTAdaC2fxBdaYLrUlQipevDNTm/qesZWKtqNtDv1C3BQWe7d7uw95VkKS5Nk1iXcbKp9I2R
MDVAUFG6aBeQQfXexH4QieA7g0qAyjfkxEq0DuPa4kPTa9FIAroS6c0QzN3tPefpPrUgjCpCAb+A
CO8eFrXtKo6/qNVS7+8TK1cH5RaE8OAgU0MeNf6JsfJhCyIHIb4VANWDcBO9hJv1kNgPFjTzCcYV
cCwtAmr9ANo7PJaTyiTQx7rZnE/fYLeottMjP1SVfoH0OXrDGusljIZyzylY2PEBalFhSIic/oqc
A2tQIf1d1cVgzmlKGhUkvl8UvQXdx+tpmQERINs0LK/nwextX8vCnAalEkt7z77WeWOapQT5naxO
rYFiPFLQgz163Q8SVX3OFcQ8fErXgh2saACOLzZeT3Av9eg4uFenYFO477TC7mSK21nPBqwdqeOR
IqTtsWwchdDvWMKSv962EQOj3nEKnFu4WhE/DBvchBxJ/MSL1gGuIAk1iTDBLSvpAQRiZeCoWcCC
hleit8glkwJ8ZmoqrtP4ac8a+/ni9P9vzvMl8d8sxOtkLmTVx/kQ3m/TgvGyXFKpr+QkjLDjPewC
9nVv7kyksPZEp3qWP7hmgRiL3RJ2ITuMkZaAUrGzRselm7cjgZw5SSsvwy6BhqMEPOemGasbEP1P
owu+9AJytrsWVwfPqqbPk8d8SmVxHWRbnVWLV5PN8IHbWCUIPSfUzDG6UUbVgSwuTKCwuveOy8jx
BtfYXOYekLnKVUAgWeN1CxczGzDwa3lVaFwuWCi6KI8/44iqc2JZLOVOMXNOpg6Ko0kXtaZL5Lvt
qVF0VqJ6ZXyLVZwxuv25xVlcrlfervDZHFxXq8EkH/1V/mz8C28aUdJKFSs31yg5D/IWviGaLPcV
qFXfmWxMt66lguShg12AXgY90qopc7F83NbgA5m0lhbvmfYVjcGXM9whKyhRNAVAPlCsOS81ByjE
upoZb1JKGE+l853gfddIz+X5JgFliqRqg6x5HW/+aaknn5W+9K1oPG9CmNQbooNn62dgKPiq4c5c
py2DyITkLmfpOuS+K/YKj+wEaw2SqI3kM9H/dwwZ5KNtZuKRKk5fJFSCdtK0KViYyZTytskva9Rh
WVtfHDPuF/KkOKFhFTqxXO9yaTTT0dkxryvd9Ed585NGFZUik/ELtB3reK4Fbvq2WXVfXp7qYbg4
g/mlfupizxMo1HPCfAZsdFoRGIAlv3D1CMdwbgsCVo3mAFsG8tRCNw2SJUsk7oTmdRAocjrbSxWB
XWYwWEVoLu4XBPDWz4ScKvc9AEuiv2nLMIb3aTIUlrm7YmSt3hhkOU2IrYP1BoD5rXFfasszCToq
Du0CxT3VUc0DmNwPUwei/N9bo2eNe8DbVCfgFFzGRvCKpuGhbluBBClCSnoClAmvFzFiWCGUuVpX
okjYBFeUd9n/hG1tQhwyHN7LRENWS/H5n8vqjNpZEb+lOtnXIeULIo8ozKrBRORUfyMJ8J5J7I4R
fBYeY9XWvz59vUCesgXo/hyN2gvDgqapjCxrro/ucEiuNI26VaiCxUiNeU459iJxvLw1zTJPLrhe
wNmBYmVZyvI6jbUZJFBFYrce89l0ZU31ew74PCgXDEH5VG/9QiPCNtcr2npbPiuEAgs6vJ+aQ3lS
+QE5oGewrYSu+IDdUtEnYrY8Py8FDlsCX5D8GylP9K4dj1ZLh1wyClShwS3tlxzYFCt92q1SemR+
BwfMLWP5TpWeX2TNMPbdLnOu+yc+jcFImciGDoZt6nZlt74z3E3adBvr7NuBrSXk6T5u57U726bK
rgIORDF/xZAzA57I2BgCwfY49zpHOT14SVM/LL1yq8yvEVVbLmec28o+sMIt3ove8rXN6gHbCtEY
J+v9U9dW/k367ZNWoQ7FL19HwFs2DEEXIsSoPHIRQN3O8ojkFKwdkq8I79UJ8UThxDMBgZbZJIMp
eWaSM0EFqe0x6YtD82bUh5lvg53tZOAgtqVGG6AKv9y6hNxcjrDtbRxMsbZJcNWNHcQnQRcL7NTk
h7sBGVS8rPmcRM4z1Wcmgw+yZDK6m6XsU6h8A1R/FU5mJGzIZzHq5bFsn4FvLFb3/rgaQAHX3pHa
2VfjyCywXVXN9qxfhFT/lVdi/P4UDNQmULfaUH/b+SCA5NtPz4sP/gegjl6P90ow6P2pK2lMfZ8l
bAJikWo26xWeMBzTEYAGEufV/NAUa310hNm9hWfswF8K3UTEKuJdx3DehkyP4WBNNkXIUAuMsqaU
nkPrtGHzMP38X8Sn8z8d6jAqhA3/YbD2clxECPf66xJNAIjkbbe86GIvvest4B+DDjKigEmpzfZB
bmzyaZtEt0HAjBieFS6oaitz7wSQilLqZRcIf0WHRIgGFZ5ndJ7o5IQ6YVstenvGdFFIaKB4WGzg
3/ryY9I2WBEZOCoZCTnuGFbYEjyaNRDNoFa/Ypwr5dxEHgptbHm1HrUgJQQAA/cLG9AtNsicJJ+H
nrXj0CF8Ac9Lp3uWuuwzyJQBW4IWcxN2LEmnHqvV6i+l2vKcxkbu5HOMHY/VzrCylPos64Py0Nqe
3VK9W3G/sETCKtD9ZqbKvnNV+CYaBXP1+AVCl9AV9Wr36OmAVn9MEZzULcJRCrFmMqOlFCARlCPC
9rLw6IGpd+tDbkVzVGTgiRbeWKjCZeR+xAqSZkQXIEKQjao6fKxmoSbrwwMyzyaaKlJXuzMt20WP
eZQvvSBB0ERfA/TlIeAyXHMN+hL9JmpLOd4ZZjBpA+KRYesbCDIqVk1CPNGe9DG61tqLj1Npb9DY
SiRR0F4xqp2KRn1PmmJ0kC3FkEXerivt/UrQgR5uGHqjXCyQYTqRp9PbB9ncnZYGhw6+CKWelodw
6+TYfMybfIslVWVZCbp+RzSWsnSA3CSSPF7SVq3/YJHcIjz9ETVCCWSdg0kYlRas4Qbjxppn+sHV
4wHYGY1Mnna+ln2nL9IZbw46ddpgJD84SfqTVnqFfu3E+6K+n1FH9zu6WmYQMzTroNXhsdwUWtS0
2gBCd7DXr5NGJwX5RaK7NdOs9asFk6B002SlDg8AE+d3sPLvjtse8AOaIMUppM2jqARo7GIF4+sa
0Db48ZI8ev025Vggrrj2jzje/EOAjMC0C06+C76W1FNkpgRyCUGmDrBp/8SfEI8OsVjA3dde8/UJ
e86pyA3ZobPWN4MfXZx85GK1OJ7WSQ5Fuscd3i9G+WqF+4WS4l3zwMFx5kxA+4qG6tHgiHtmiB1Y
hbdq/9+NiPaJtOP9Va6pr8khsJyL+V52kjp+0yKA77hUekW8Rg/GNNCZ/EusYo1AddCd7NtLaf+f
5dh3AAyVkfDzFE9Px6I3yYKoDvj5nX+SnuSE7RgRfBnaxjMMVQ1kbPvJgKz5JvQ6/0TZUcshC23w
Q+rpmTUZYgP6yF4DbfMviXZiOqCcH8Ifo40wAy5eJDphAQAWAUnAJbodxOVLtVc2kzsrtOwzWNq2
JZlYZZdjPoDqeVhkScDdKdGOCEozlk4sY8I+snwDHItcr4Tc34AxNFi1yb4l8IBHksoDRwekgf3Y
iRmTld84w6EQlZV0CSakqPWeCeBIyZSJCd70ollFwBj/LbgK+vSXrwcjqI+QpzcQdiUEw7uOZJK4
TQWELX9vDRFWeg8oPzlVQmO/raEs9eorORbV+ZkPpLHEmJvsaQuPpQ1OvYme2a6po0Gna0WFiMmZ
mKDUQ30rsoEz7V9g4T5z5Y6nAADcFCrUxiQPOYrX9+gdAPZ+vb4WSsUX4ajNGwNFf1vszfB6CXSO
Uh+Au0ziqAxzkwt9r3M43xj/EhE7/XnWRX6Gut6SbSnAdeNSMSh/OcL4VCiM8/Y4THUQkaLewdMc
kBJSXNDzolyiS6nNvsK8wCcBCISPTWO/yaLiBAuWMzhkhY1jHSBEHx7KVmfto9GCNuhirfATeKRq
mcEc7fCr2Z+6hXvOK+VjRxTMpz8ZHwMXlCCg9P9bk5wpY3L4FlkQDTTAqiARTB9jsy/CULsiPmhk
0fwq4UlFsevdNBB3nlKWRiv+yuQR6KUKHg2JOIcReqiXgzLBA1QZVuWu4zfPJpPBnQPt7U2BdB/G
hBA+pRz05/NT6oD+1gTHZPJpEqUJLZxZ4JNBs+cqSS6KWRkTUWax09YGwNBnXj7fE+jN9m0fdlsf
0eFIaaF7mR8nfaulXTxvVUu6IgmlsIvzvwHRlSU9DduTfTgKWizr8c0HSLNshOSWqC86123OXiLy
nG2tzs0iYu1pwfZc3eKD5ItBUcn87aZ/yqgF9Q3KwhABLcEBNDWKIbU2bixQalAD1m6YDVXvyzbi
ElDrAuigvLCKGdhSmWR1CSy3lLOPGTtWUn/y2a8Qpwn7NGdEuiltzQ0Yqqk9GxAd1c9KA5lII2s2
xrXXd2TBt8oECtBW7RDcYRXOh3ycyvm9MSNC4R9g47iRRFyvBzTmPHwiwMB6YE9qM+6HPoWkREZa
ZkgaXN4DvBUpRSZduQMzl4+MohmdHHwhl4g3MLFQ3JFY0CeNqHSpBRWPTMo5jkMI8PSv8WDtYoUN
9v6+JH1zRI/tXSewyAnQpU7JXFSZCdqgKm23kT7isxf6HBD3p3qRYnt56ts/psJhM6artsLzR0DF
6b7JB0tiEbS2UqT/jLAAzeNYfiV3/EZF881QxaojNumD3OIrMcdC2x5WXbLedRuQyP2Cfvb46UR4
T7O+FoWopakiPAK44XRHbdexmlgmtyYgZLsTgqS0zSpbydn9K7QBFwqILaBK5yIvtAFg9/1Q1KNu
JtVmzc8FgFEKf5Nfl0mnk6TDhC9AS59ovHpq3tWdCIPPZ2fDR36T0Q56wiQGgyX2vAAj36RLxO0B
GczHITLQD6UbT1UuAQnaDxUuAtR4/DqLJHzDjXgIRO9IdsERq9iALDfmXtN8r4a1aNOYsSQ00YHu
mG2XfOOWcNaYduE5ftmw0FXrYELmDkUQdIUA74L9Ltf/3BHwhIbc9ylCaP5cyHgqK2Jp9Stj2uMH
Sa95c9OBV4A6Qgi+6z/BXuIHKUNdpuQLCCHSQHQ+e0UGaJuEk0ugq1wyJfAJ1QFWgVODwXzvfUPm
x1dqkMyGrK8eRrMZj/8gfrQTG/5fCYA3NDyFPTo6j9ZIUNzu4D9AcE2Kv70DVdd+U4WH3n7QMnfl
vAEk1Y08zDiZjAzxkE2k5WPX6SB9rCm4fU/7Xn01G5rbxPOonFgZdyXKSv/0G60vq9ysBzdsc235
FaS7BIT4cksBCXqtCQHbvJPJ8Hy40u01Mx++HQt8bC1JVeYVgOTv9TBtaPkVaAhG6kLhSehAeevH
9wSns2zZzSs86X+Gv5Y+DXoVgwnWDMTIuqq7CSec4jsGsxt0+i5NniDiqPqq2Hx8v1/2G0iub9MH
euxku46y1zYt28l6GQYJM6oDMgnPsoblQq4Pww70xJAVwE9UJ6W3LVerpLIqf5/Zy3zzQtBX1sbV
hlPMFVXsW94ap8p8NTld67tlunFRZVtuEYJiB7Xbu1XJlXYlHsTRA0Q4NoJdAye7tFs6XN1RFsGc
14bE9081sFZpOTky/0rfbRHY/OxX+8XjtxZphgZIKNPXBMYhiUWpy7DwJ6X+jOuLFOUhii+i3j/r
YWhTn68CZfmsmJvyZqCsDC0lUdkvV+HPw5MSUZKC/yljeTQuqykVqsPzXURyWcSXUSEv3ZPYuNDF
PZm31riUAVTgQNERQebPv0Y1oxXV7pUp6156BuD9DjgEKWxMdHT3axx6NjiCqhauVBN/9+mC33nj
b3N+uMvKJtW6u27Kfh7M+C0RvW9k6gS1OQfMYlH2vp+if8amqCJj8QatZaljqmFttLC1vxwLMh3C
+w3eNMxO2o+yUXEylx4z6duuKtMKxEBR2sXTzNcPI9ZdG8YSMC7Usli7E15ulK5Bwgtv5xIqPLoo
+8Tj8UItt8ZXHVrQFQm2PUYE5i6Y2YPWt3cdzAcOaXgw6s0DRFxwRHIxdax0svTUZ/nXsPnPJDIh
A6apr0Wyno79C+B/gmvC9Pc+MhJypefyEB0DqzFGrcGHjPfY8Dhk6XVPCQrGJPdKdhy/aQhz50UA
9SkcwVEYwq1PHkDwW6WeLKw/Vab8DoO15TTLxRHpOxV5U81V2d6t/YXm78IwGx0Uo07+E5p8dX7s
qaW0Kj6wnpIh7ZrYBN0vNU/GytHZ6wF02p7+sYy6/rxopqxQfQLBaV8lNvkRmKzU2ThC0Hygq48B
RAErvAw86kpKXSC75uQBPNJZQG4pVW3yOHTvGgxZGLJtsUW+PIh0Djo2pU9ItqDn6ztpu+DX0PYV
rs/QbJ03h9OTQO8Kf1tei/gvyWvNud/8hzDhZEmSy4QYLFBhQOvakmDbT841IM/eA+bR8Y4lOsKh
SKPyfckhf0BFUrHYWbCRKy9AvZ9aCyufApALFAQDbOTQfzSJ2Aj8/JsyWEdOkRt/3ZW6D+uxo+kC
qQiB/+j2eQwcDlJCVes1xYJQ6sgrrRGgHbnJyBrSaLm2vJgQqy/nmBfw9WwG36h+5WiMZFod5Y2P
fOEiQ+yVE/Kot+szTcKVPKawydLKqrqfEIgFv7HyWcSpIFW77IAPxUfAYfOQYOB9vNPGv9/ebsA4
jx3hJA/0Qx1ozgzKy/F5ozVPEFDZWs+7jbV/B8xRl/qVrQJv464n2TZxcy4hEaYkz2A6z4TfKUxv
aE+UW7SeP47b3t4alOfzGeonPdQqDhQw68bQFbV/PJU1B+nBEi1m9aR60ueB5RAoWjzXaTkPKBFH
E2zC4hOHBGt/KmajX6/PuiE3nJwEyh37C6njrY6oIOMeXABnRSoO1zBNoNrYGtrb6rq6UwA8Ink7
WpJTwk6hB9gcQahWnulffhFlsXcwvGiC9tz8y4AJFec9jlkyBc5Hyi6gL4N6OLwPNVwdfkrRk08A
Pn/zEIhtsZZASuDGseezeaKsKYyylT13942vItCRbNDGqpMy5GAHaDiGZ/MvoajRdPOGxOIKbMgT
3Bp0DkSvhZi6S9JaQ4u9q99FoNL+xKobnp0VW/caFJtqKKIZdeWHDP1j1KimPw3sgz30Hc5j/GrC
NbE6ghixUoR29g2lMVufZFEesGqezXx6otKiHxepYaBJpeorto8PAylCNHbJ/G0xZDmOqW0ug6iL
UCBlP5L8QWeLz6CiXa8yMBF9I1FjJdANULYE2zZp5x9KE+W3aHMIpReN8FDeSWtfkEuLOvpKpCik
OUJYQ9E9hzOs0yFAAHbFmX1BvIXeErLkgF3dXSOFErBHIC+rf5lElaNbsRJ9T+LskE6zc4lJtZJU
ksj7RpkZoWki+R2WmUVJGGzb8qPEN3Sluhx68pSkWdDVj6NtUHzvoFo7uPi46Q6dbicDZcCUNBJL
DrqOtQm+lj9+PxtPHrf+P9oDaiMJn7HzlE5UneHysFHxH12X+Z77zyfMHxwKMbjBpcZYkAhlECxk
v0cSOLS5HDFyySG0EdHkxM+8a8xGRqDFzUxXZ/MrpH+N2pc416bN9teWJsR+EDP7VPRSH59HuhUo
krkY8ngUKPBtQYAPftGMqT9HbXmmYeoT03K8ZN0vZo1338paH97cW+9FiaEC91X/wCACTqZ7dHbO
zCaRCScWjM+2UkKIQeJNEf+07QyZQbL+8WMDj3SE7VNP9p1rPICHncbCcAWDrCLnG0Sb62IqYefQ
TREnisNkctsei6a//PSY57vYCM9Ny7ZemTLU3QpYfkmCy6C0rSbchq6Kz8SbYy1zhf9ZKn23b22J
jWSSt6n7VmlVMqdjGB4BASckb4a2MYsRPwJnSfuv7KfKccqVavkIIVm+ghH04UO92NtZfuu5Os6n
EaJ9VcaqJDqwe2s/CD/brQ2hc5jdiWZeRqp9KDn9wtEVWQU1aw3UZZQG/UjYn3yQWmkGcpWguLd2
/Ok9ygvzjCOHW8q3LjbVCezTeU2J7M/9/WU38PMr3D77qHjnR+8famMdoNRH7SjK5HMZ9piNVPFT
KTteZf/VCayJXhv+OZ0RGDLK1ptOyRCHkkjtdWXMm6YgcXOc24LfpDKo8H3aB9vuB16vjyUJ0YCc
tiO98E6VdXKHhC0tY3iSKKtYjqXiyNJ3i5a8sBjBoKqdp19XJArQ6bylB2Lupav1ZArR9eOn91fo
omX5uawuh6A3J7dHA0h1q6CKOUgDrNvvEECvJOIOy0lWA9ZDvpOVkJ/mAK5RCZCoSjAdtYf2N/Jx
hPjA3mCQIOA7xHrY2qiIOFKRhNhIL1I8W2vti6V+ZnzU6E692vi8tdUDu+Jy282UeFJNzOrzDr4+
zGv0bA7BRBsPuhOChfckHGJ5zTl4Ze7UIerX0o5YB6koe0d7OfjXTvnv83rJ1ym4MAtkBQM+8BHm
RA7v6XAPwRjriW714oE7aOOrgVit6cj6tYyfEaqta5YQ8LdQM3hXrVVx6Jim6/u5I4EX3AU11dRq
OHTbE8YXezHILUIFVgHFoi4gFIFQ4RiVwzqiCSno4L3PzqGqYPbq8POFl8DwPyEPBmfRsvUNcrED
Sk5I8QpuOcxlcr4+qxKk7DOTpBK2kpSsQL9y4rg/0UnOB3x5LzFXQj+cMnMoCp1rWGy48XFJNX8b
naXXw6wZxb/lasrD6B6wssTWUybQiJzUxnNWH+4KybTy+n+S4K0a+nY1bhcUb0+WbVDxVh+ekqV3
5gcXGVWbroIe+shWtXQZXM+9P5dhlTqPQA7PW8twOI4NBeGtRv3G02GvUjRVSmclz6AqI79C8hKl
5ysUIGrMnOIoLfFmGQGklD9y3OHdWLQwQerC7exlDX+MmyUcz22CY+uV4MMBw2XcJProt6kDkVic
X2LEHJ1VfrqTCTCvOwy/v/t6X7HGuuiYOihy9Q2lfjq6x3ckonTOstzUD97XOxJNYcH0if2n45GK
jWxK92xvqesNPHc5aeUzq3Y2QN7Gy0757PdoTol0UkJ+iRBZcFT0km7u/S2ICpgKfpeoRw2DhbAv
KqgWVXXaRh6f/xAN6SMs8YRGMOfCbMO1M+V898R/5GcDJTUDyfH20Iit47Gx47BuvJPb4fyd1nMc
8v9OYUPMyPDSY7QXzcKM295t/6y7M4dANmgAqMOOCSL5Ilu8DEre5zodxeQL08VCp3+ILxLycYAe
KIoXx4qEKB5fdtb5q9tRzOL067yx26YWAvEjM2+0VjdAWCB5k3YVA2Kq1a/o6qujY/guJE0tYuXi
ZSFCw23RhYWpiVu9F+7BPreIvWy9lo0J6Pm7ypckBeSbped3ByJk8bcCaqPjcjxReE54LFp0qjz8
5ENdh5kN9/WvygIHWi9ZeOYO9kvHJc0tyx8LOcCixL7H19amM/zE71RcYyOaT2ySasHGgnKq/Ars
dGYhI+gb7CAplVEVEgrQnFFNmmJEJgtgcRAKfbbCncnd73pbLPqfBsnt+hB5SxbGnrS2tFTzclW4
FfDY81vQ2D0IFOINgkvJAfoKUWbwtHixfiys9K8VqjKHTS2RauDUr45N5F1DyaER/xmVTP3IrHrV
8HUNMZvaOIGEY4d9dL+m72efvMq0IpTP99UQSG90I4VZnfs9IqjPzlGZyXxtv0G3lpS6rrZKjwCy
Ngvm9xB4o6enSAVlblMz1BFxhIz0kpuLnftG067WeBofYeBXXMfLlWNZ2Yj+3y8V227OS254CabA
YLopkUi7zgd61f4XtJT+y3wGpyw4QD51rEGGVzDoXn/Z8MKEPtpvOZY72rbFnBERf8hm+/GlYxFi
oY+K5tfkleeNsJenA41wfNAFvyjHusCMP3I3GO/KGcSxvE3BFu4YlD9SBQ71tHLWpracmpqxM0sK
A09DbBIoYY0SpkP98YkIL3Ol2Ohi21RdTDP0is42jp8HkZYSawzp/gJy1yrjWY40lcjmfGQKk5xQ
XpHJC50zP+95Y3a62GzlGrXUzJ5K3Jbzn4ZsCTtLyFQk53EH4+oPtbWHmZZuCUz7kRhuVD9Dqf1+
1vN9gbvzBIQfe3sDKNic2tDiKT04OnBujWNlWxfdZoNS/EVXyAiKqN7kT9XR2F+MWjrLqoOrxKfw
mcPLH3ZK8VoRz7n1nMDPTbzhgE09Fg/GXOqNoMTJ68TFqcUQPPBtp4rkhO5+g6DtZ7GLrQzXeGUK
E5DRLlW8ecn1DBNoqhM5yytZOC5wA9bdw0pQevybTKuuuoQKqbIV8TvXKDLs45t9WwMoKypXRFwV
hT4wBVsDpnTmXalbvFAQa3r7AgBsw00k8J2PHv8WJXkEsqhZDyulI/Hw0tuBUY5IqsjTDBR6wf47
wliVJ3UEgeBLDym2sQxqfanJT5NLupDaI/XWY63Glc8KeB7+xXd39GvpU2I0NAAM3RUQyUUqvabf
ZFXXVA1aRQOXu9ipAe86nMfkIK3Ao1hRUJKTw5pWGqDXA5zzI5qvjTVhLSpxsisnT/5xo5cu1OMq
hrC88i8fDRkKw7LZGcjT2bULXkLuMvv8kqtOt3r5++gdKqL+U42TxigGqSRguqODunBYMfaUveXQ
seA1be6NfUxp36Qu6Y4TrcEkS9VA2Gcj0ZB0rmzkMtw6UWspMzciStRodV6PUye8QlYoZinRM7iU
pWKTF0dMM7sW7TzdgzQtLio7icD2kxiGZUkrXCwGqEgXnKwOn7F6d1dnEL1zWj8znPb0lXsRtQV4
j1zNp3SR5TijyOtFxrpI4tycSVX65hCDVmM93pIhRfGS2TmvgMo8dxXW7HkQ5xOyu3IuVzwsi0Ix
9cDn6AaxJZ+8vz4CiIAHwlfvA69UAMJqCZteZCqbwcTbMFTXNs2VHneYhXZsTxhLRtHIsstoo238
9PU6jimFe+xm5EOm0oP/cJnZO/+dTvNW1ZG3i1LThJgU9T7eYEzvtdDzUM2rYhQmxsDRNjwNJxU7
wpzFYJVjcVZqtDNdc/iS4dUjkNrKRTmmAK22CozbnNaWz0z3pQCnjboC9hYyaDHQiXXKEx4ZpNKE
W8Zb5xCxQA4XCWTTfxf7Rhxuu9QORvHi30BGD2qXHKgYcdpA56zb5BkJFihda5HopzNFPG6K/AHP
H+KH6F27N3RrFVLtiwspvTex0KKmweIzmcO3n5s7Gda9fy/azctRERQP5noQ4Y6Bv4ModQiSSFd9
lO3/zO0DM119XTTcogjnthqURq7hppa3KzhzER2Yhlad4BBZcMz77Ix0CGg8/3QuB0X+5NA15e+G
XYdKF8SUsodIRW85BaL2Z79OfYhCiP/hmVpv6HPAEtU2zdQ8lSgX1fprWR/RDxibKzl9BBzcr4EP
iOawR+ozstNsu9nPHW4BWeDNok84BdxLPI+zXxqaE1/uJs8ULexR/ampYsGCKLFVIepxWi/g1sjh
ewVg4/w1HJmLIpQW7Tti2lmvwmEGAJeuzIwpE3pIaryPZ8w/xGpgvrcqPq6bPc6Mhy+2ok8TVV1y
425ocSpHYAHnH/9MY+Bpk8mNYxxB6gxaUIFjBqxhHwPRBLunWktanmde+2VFhCMYfIGIbGbVsLvW
DkvhjtSuLVUFdfGARcKXBUIflU3Vdd4aijBarD0RgWfDS8QuyBb2viujpWbqAZBNSKnG3whD+yFG
9aQNRnlJP/RdtwEPC0CmCcI2vzMPuCRJock8J41ImlO9vUO4Q/sQdCDhR8TI+Sz+EjzwxmZpYik3
cK2N9UnVOIuEeMDNncJVHEJ7DVUcB44ifB+ZemD4XJSLkejlGIVobBo2izbMuVtH2KW/3egy3Jwo
1i70uQk2oE6RD9wZlpyzDXRfd69rYrg9fZKZulBsVxjEydWrYYAgJr44Xf6Mv9Ne50EuHGEWQXBa
YyFl4ks19/yNvjJO0hY0VZcudWuJ68H43BmT9U7qG7cKQIZr4KGiZA+pA8ZwlGVvajmnsqi+R+nM
o4595P4O0+69iWBLgEHrdqqqLEeSYyUNKJR4X7tBLx1f26/eYiYonn6MkVOKrcQwmXuuASfmo0fX
UoV262nEA1vepuwz0E7RSKMJks6EGzhliv9kIbfcnOTeieBWFj1dL1khpS6w7IQ/ngmtd4Ig8YQm
HtgeMU55P/vCEIe4FPuhjRAxqPtGloXiY0kO6olWVTbFQAA0FyMrtAtLWCiHZoSDSjNHowr47Ta3
tmnaKynD36ZtE1gROwmTXsjBKalBpJul8Zsu9JOPi5A/cEzRePHFiCj4eESpJsljScSSGNCZ3cPh
vWXkEMCmG6kA2HDmKfyYwm9n8W0oZ78KD1C5Ij2vgeTR2gvdXv+K4uuDt0lMTrWGlNorf9ZheDry
D3/LqHHthFrncbwPblZVIyUMnR/mYu3nNKHqE6GA7gS0aeAHim8dB25zpI0/L3FW3pJVR3P44gs3
A//N2FkOUCmyWBTRn6ZQGqI9PFZpBupvJwi8g78meEvwyuUFUaF+wfRpdddXNe39va8APxkcmY6E
ZSRDVyoAehu7DpeeGHIYv4/hgsRF1+ZkP+JF1rrLkWKqVdTbC2eylvk0HGbyuCo+uwfmWBKaPR+S
i35B3bM2U7UFC29Rd2gSxcymtNvZNym6Zph8JKvQlbM0kO58/bWdmUNOlLMChmtb3dxqxBt65/+Y
9Vzt5M/mw2RbNHMgPkhthWcucNJUQp8cSXRcLfiVNE5+TDZr8ILY7V016UG0XvrUicJxoNBY4vr1
D97PPtYJ943hha5AVAwtz6hhe8FFliIZeCZ7Dre2XPrJXh0uPgkxjhozwLynhQ/sxpYSdjS0CkMr
63pwOGEiEXZKLvNP/O2Y8hX2WTXybEFv4Xf+QDY4+NWw6LGJudhacKkm5+bkPZy3Jq0WUc6aXSzs
BRHiP9GjdINyWdyYAkT4uu1l/XMZPc7FFN76AdaK1svyAQiqBiJU2g4J6RQmOStyeS4y4guE9ywo
0U9fcFJz3CYg/X+gPqm4xous3TN+3kWCufD7UBH++WF7ns6FVd2kseO59vvWEE434IRn0UTbaKVv
WJeUK9DzhPVJnklLRbCFwe4Jq6J7Vr8Ogq9i87/SBTnGNUNTXDNmJGDgB0JAcMcFjK/19fHELo66
XQbvCERyAkBTafXuoTMSbWm83TAjE0urdwlR/6b2Qbo23/PBuYcJPK7x5bvYS+bA13Z90gS3O1L2
gAPKDwwk6rGtbt9+T3hrv/5wav4mBI30DPI9XCtP+f3eaWA4aIMAvv3JizPykTqEx21x/xdBxR2J
JX4HWY7AIxwAWwmVb8wr9YnT23HB7mOoWAJflmh9CTuaHa1Abphw0djl+2bqBy3BLoTJIDXlFGPW
lQQfh5Uc/rNJ1XuH8X6rdUzu6v2nOQFJEsCXrAy6EFhmOrd4dqDjrezbxtY1rtkRgOllVBG2bOp/
dWst1oHO9l4XjX+c3HRkLmZspRZDrJ2F52qdV3JFWL8R6DAq7jRx8QcpXjjBQKh2AeX8DlSU35K5
n+xzPc51Td0D0IeoAOq5qplCAXjJ7/F5uz6LC1xPJRlaSa/gyCcYyAJOmO7KIYWPCyawchLetRN2
y/7XVudVQA9Oy/IN6vbVWJMnwrk6qzogpvcriAZZyd3KZeD0sebwqr0xbkJg4uT8quNbXoogKWtK
G2mp0nNrJyI0iZtFvA5YHHyrraPoZtEsLZXgiesM5XlDqED8aQSrF2nCiyAUwJEyWlJYWtfbFy4f
1e8KICXbi1WZ+WuIohkjLzYnPraRExLhlLA1lKBV/qfd55vP57Kyy1Tp4htuXXJyHJKmoUMFhntR
6KUykCFdb5ivVgEGOLAV9fFoMAc9NQW8nA8n2FwuKB1ZF2SwEIp8D4zOqMiBlvLCdwSD4oAhRYoV
c92oEyx4vdgIS8InCq+tVE5dF3w1SwijK5MtRuYxtYU4up6WEmBgZzvTzcxob0OsDbRl8Cor+8Lu
Ttrk86NwkW4cydjYqdBcBcQlD4BcjfJFeBM0AvInD3/EugETiIW8Nrxp/KyQf1IJBxu6EECGy+xA
thSz/3bf5+U/zUU/U2d1+5IWFmZkl+B+Knq0u0ZFUnw/glY6Esh/+Tf8d3VHnmMoHE6WyNWz4VvL
AfSZsCpfzn74KOF7j82mvgLDO4DEDCKGQHWhMI88CC2p1iV4avFdjoyCLEDHxhohMd9yXJB2FmAk
95EAb4rrZ/HaivvjH/WPCeELy3xSEkrUrooKxJBwnml7OAHlSyhe53Cfik/bpHheV46VWSYp0rW1
xTu2pvyyvu6cnSj0/S/2V5Sw+QsS+7P+7eSdJ9dW4zNWOVzMQcDrAvlW2epAf/6vRz0qgaANbLUQ
z3JNJgcOVQSHAmTS1y0RbZJ6NL470woU+kolbM/W4yw04cUYpfjeDa6bKIU+7pMZHpyV2oHp2BxE
5wIKNccxXCCHzlXjks5Ij+hjjEo2n9maXgIFVzQuzqmyxryP5KKbncWgCugDzkz4MzmE8B/mu2CC
4ymjt6NCNAcHm3B/VWfdpCRlREqX26g1ppEybfPx3z5fMFFnXv6LFN80/iIHVBDXIzp00r4UEQtk
2gqqj5+5+aeCqhwsECkxQ6jaxty7aREKhBAWxrnV2fCrjuYXrl6Duk4eDFwblkc9a5A6locCmfey
RacpPqVNNV+0u0oc4GiAI5cemfegqpO6roJT5LANDkqBiHYgOPXMJd2Ty8djb3ZoKHMJKDTYUHtg
uK4uoG11ObcFnR3YFbs2jWlA6f0WprUPK0ZUX1aiIL70Ryz0Jjdm9PoGzJvlkrjCws26URBOF3VQ
jBrdG60MfErpfA7uLfhVY9tJgT5YNNCWZK6/mA6NhX3u9MhqzgrW09eCCGJBxI6qCFls5l2JzHlR
d28kgFq5kYAoz+xAMVV5kLJzSvYatvYECJEPPPymN6a47SdKEpABvx57kHky6383kCg5zA6coioM
HdO1OKrURUpFc8zeNZ3ts+j6OdqmwBlz7zWaS2BOxCVGVwAh6UYOdelqxao6rY7w/AKcSQmlSCm6
VZshct6uUgCLonHzHWzZ5+CvX117zWovLCABOeQkhealP5DF2okbLTyDMtj6n1yqnuDGgr4y7zlr
Y/dsXOgI/befAtgn1wEFH9EdWIJ8BvLf2y7iAryQ1K55Mh2JGO9WunGIuHgZ2op1egcAKidW9uBb
B1G2BVhtZqXFNiBis4zZXB+lOfTJOTv29NLc4szwpn2743tJFw2GQLIJaMNMSD4Q5O73Ik3FTaEl
0jV95lIfq8Jo0PJf/4zDDYKAPAFV0PQFtf2LdR398rx65I5i4K7QRX6Ixayyl0drP5jdMVwpDxvM
ija/Htb/B7Kpbb2lm2SMDnhCHYZL6fyyH9S9zAu8o54uqteHBwGLqyPoyp44qrvC64P75NZbFevj
BNKBxZtMb5P7vcCS4+gE8wQPlx3gYHvMWOBbHk6cx+4TFTDqVq1Ixn9Ua1wdu/Y3j9X9h04yk10v
et6ZYVgtU0vWn2tVc1wj0NsHOU7SdVZQnB2iZnyPOV+QSHisAoTygD9mwnQ9Y7/jEW1ZuNpd2rRh
FGb4R1j1LYDcog+DeC/Qimowvxk9rq+mIbh8u5TG4V3AkXDOxgxZj4IpkSA42R9WZdX7DqXrqEpD
0X/i5Po1xB1+hrZtQWWPMT3Gmo6+EehbJeVA653F7OEY0lIq9JpofZ62FDzOP0HTyLnhx2dCYUgU
ZGPM13nCZd2+bKx+D1w8LJ1QswDmzYbyYw4s+kZwYHDmpXV83ANCEZrkLS+Ki/wl6JOUAD/gXwY/
kfCI/ioOVxyyRhqOxgFT8x2JATxeKcVQk4AWUxw6Ul1GOaFiPMs8WYKsDneO1IekWL+e7n6P2Aye
vdNjPhUvQgmHaeNAYDQlq0kDeSlvUXtZVmFjzEzsNGR9RZkc6HwcpAHm/GDxuCAftcTOJV1EotMD
tVyFvdlZL0ykXAFMme3gEvNy/hUdMh47sYKZyC/z87V71j3oNZGpVhNCb+BzI140oA2msayNp3jB
GbL58QqbL61kmthBg+5Z9ZLkEDi6E4DXFUUKvs6Mr7tgbwwNiXKKv0aDD0/oBqvqMFokUUdzQNTM
SJWUz1F3ecKLEWRCMv9YfJEInrQ52HyD3ziahCHPrYrtxme25cF4/zwNm12d0kXaj5ivyGan2axk
Reg2/rl+1nZ5tiLm4Zzl1oyzftnCFWrZdLOZM98K5bLB0IltufS+FmV/tNoVmO6X0T1k6QuxO/0X
5sAqgdrKwoDofqJzky3LDbRV33Y/8b75NVkVOgHJ1p6A50SqQo62up48N1TYzvw4BafCMYb2qo0b
m7n6PqOpbNCwozXRAGs635laRl8PpIMVKR0TLXUTXd+FSEnXURdWjFX8NMfOh7859aLKY2ESeX5J
ytfSzbX/p8uVVEb97XAgwX1jss+AiY5PUP5iQ3x7uwvsJ38K6amhUe8cLLroi0htSC9zQYkaeiF4
joHcdjDZI2Pd1CGpoux3WjsNOTeROaLS0bcCk2rY2XIa1HszQOMnmr3DFVpmoBSvLvusA82RnCeG
0q1Fo15XR0pS6ELLYVBP77wyK154RWv5xVqAcXSWllV0J1qEKbBwAsY/Yg1fB3FYeAOTtQDOeMWM
gLIIgRfuoTygEmj17fIEJqqWXQyJZB5QuPINqXT/7u3GmZ3Kp9LZATCxyJa6sOp5jsU+/Fpeb/hA
SuDucgsxJuw6UxikjixX8hTtNeLS/ob6h03a4eh5iV0buQrb3vBPgipAHx4ZyWaZkEFyiWfX7P5j
XuM/AGAFQ5g6KdwndhLzt2Q7VdHzBhenZs/4ta5YiPr98Sb+b9z8VEV9UFBuGFT4w+SlDIKMgnFp
GVPpW0S+Eum2smJaL+1v5dG0W30V6BUEkH5Vg8BlsMSKTZu5ishCoPN+X8R/gwoPA786OcVegsDu
u6TCvrz60mekcyMefaFJrv8Jl/E7dQ2OQaq0udvFZP7RAvAdEle3PIj4qxVlIrqVxvA5VPK2CuDX
OmAL7jkPxeQrp55Rs+e7Pi/nQGIM/5ySOYSYRcecqL0CMGG7Doo/Hh9z0LpJk2UucjPE9kGVxIW4
jUvgODpay1LMF6Lhd2oTapAKuIBty4Ok19inTBbaONeV+ExALkBchlTFvEgej2NbC1EuKtPAQga5
Xw0olEU+iU2kfAxlwIgilEsWh8dV9Hm7U+SFitGE3YomEavf6S9/NXy/bAfU4Z3X0hkGzB7WBRSU
zSQZ9klE/MLEFP/q0pWXJP/Fkj8aMhGzhLhHrnD/LyyYGDKTuxZHl4BWnPehbAPPOvHrEPEDdliG
Kk64tgV3z3QtxIMV3hXbcMHGm8K6ab6IiVxSg/Vq0zJZYm/b04+Zj3owtRdk2u0lYraQEQZjO/y2
EvtGvixkGDkzuJaPAoTOsiUYebvzuXtieD7AzV0Q/pbpXhdmlw/yMh8t27qrW1oNR6vil8wpsPeF
YuX49s3Q/wJHVRX+LP/P47Pss+fKC0BQlhg0wPNSTzHhg9oWN7JvjDq6hgc3tPedmnZ90kcUkX2I
TfG/K57sudJTWbuKto9b47rx1hlYYS/ZjhiB87Sn82qdrUIDjxa0EOZMYI7QXXhNczoaI74sr9Ya
nQr7znr0+4ePb/rfRqrXjIRBitC7S/DzkB74m2LGfzPSLVb9/ZWVOjInZeGR3BxSKiZYTjlt0Miy
AB3oqKNy0wpJrTQLIohXdjvjqVlQOJkPjPr0nxUmV2oufJI2U3DgpYChYrDEGBvkOEBGxQFV9Vd1
yPZh1AXHMrVQtmBPAMFnLUjZDD0NF8iq0NgnH7lAQU3SAE6RB+Ztvddr0IsEd43van5zBC2uG1p8
7vqcJHT6rQIo/78/2qiYqsKb56NYQIBx7dZ6jnDlkK8n6PvxibQkeZIy3oMzub7pVPDNdei6kAt0
q+IvxtkRnZV8wnLbkVKrjZ3Jqcc8M6zfi8Y6Nd5bssUv+O21dftRqb0V9nTTg13LxBL17+zGTM/k
LWNIi0+cXmucikgnHKX1o+4MeMdJaCE2+yf8UPHCEOErplSIu+WTQzqhHoJ2sNdHzOj/wTWHSNNN
+maLR3IGN0QzOHeIPX4rntEC4yJh4xVoK0lBsz+Y+IioyT/jUwt9RmkrE2CR/bzWq3XyaeXFAB/8
XraBNNQsRCSGQiM8PLJBEtYGBM9HX+ra2KOhx/mxplfdZ08EU3WX8oxygRZ32j5TaXlJXQQDYtML
RslLbEbBUWOWJ/NJXhWIgH+awAtbYDh7jKEI316LazLAnT/5NHOQ+JmYy/FZCi4Kdtk2zvT42eLB
xnZ+5vD5WbUSDSs9RfZ5+orVmqzCjwPpCfWh+q4z4OdfZuiibo3X5iQ+rFPUMwRD4OSYCJap4YrJ
f4AUgyB6KyH+8tHe+zcHgMCyyodAgFl/NwBJbQa9A7iEmksz+ouWZJjQFxyVIdEKvy2JFmz9ZbMh
5Yc3w498DIJNmP6mQqBamGBIlehLqudDkSV5/3RQI1cK0vl4KgnFgud5NvYZBXC3tifZ3M25p7/j
a30FIySqlx7zNYk0ofGlbDRAXeF9yFLjZ26M4W+vPZ5KFFtGYua/1QdoXxE0u4eTaMV/m31M8gln
qZpjeAV7Fc4KyrgbdXM8U1/E9XAUD+ZsjaWe+NSnk1NzPoVltNgi0fFzDkSNLuZ8V0szHopafalY
Gu/PxHPbCGb/C7bryLe/CPSX9BeOj4P3EOc9NDFTYJvZkcKkZFF1c23BiwgWoNVdNsfOGz7+MQ7N
q82oBxTJz6QV6Mpj3dOCTBvm6MYiGiHABag+uJQNwonvYvuRmKB+nxmJtt6VccaBcIva41gOM0yq
mNKqr/Ba/paRHXDCPYqeOGhSsmTn1LZHs33NzFLvfuANQePWHH+5zWuimF+NglnhPU3u4ebZGvG1
NfhfswA/Vlbmd2tkl/h4Op04zqRPvCnr/Hs+u7R8npWUwqLGKzaB7DZ0peG6ndeRHOYO/qSeMoUu
ABtdfp1PPovAE0PV67G7G+R2vmEdDmjlAGpPgTyMQrixviOXynWVa3wWzAK0vWWYwa94o3xHSSX5
oIAxKPLNzYUQ4SoNRyOQf94nguVW+aeSgdYGq3i1PVf0eHltqwTyhJuaODe9y/8PAQ+CQk/s2VMN
bVtbGjRRq84hrbFxcEg7VsHWNLXVFqFMIe2eNvxV7IayLDFQiMfJBPqRuMvdcowNbf7Pjg8ThBv4
kvzdop37ghWUcftxz8g8bBuANK5Ryks4BxUjDBj8umKUCPr5mGiVMgd4kO85A5p91PVnLQW+lJyF
csJ8FyzUQsZ3OA0a93FYH2YEXOf0Xe7w5Z+5mI+/38s3OHQNSWA7z+/3NSjurX5GGoLEFM+K/JF6
ue5pU2llm4ARhSK1t/7cR5FdT+0ZbMZTYJwk5fdAQ94T/ufCu7FYExQHNioWJ15SgjFcctSsCCgH
9IUD0YAh0fvypSw6fq4/hmSHXgbC5LBISkPjyMM+KOzr+d7EJgoZqBYVUfU6VkCoHIyLdtfF1p+P
MAylCPdaGqWaH77neRTnEWYYvCNWnUeiiwZBk6S611Ta/dFCHv4QNZSuYd16D6o/0SErDSVUo+bL
B6SVS1CvgHNENgNZYHfsWNhiL3BvcvlC8ksG1U/8JD26encteZxviO1yBTW/fC2z/2zYJw53J472
/q7YDhQvnKDkNvflCTT5NkgqC/ES6tBmW6H+M0lZxHNQUyBDMT2oUv8FzOpnSmk0nMqSwCOSysO8
MVRo6K8X5/IC+e8Iike3Zxxk+8sRBcKRrsoU3YFW/DWM7AVjnB0+IR2MvlVWFJk1OjxYQGbrA8Ba
69NaFkXPWj4osWo/jBAYfpvllRFiUmHZvY0mV+l1RhX79M/Ww6E8XoK+NiJoKijOpu9e/XDyrfKN
CO7PVjSu0yn4zvNeNv/2gDrOg5ltTOIt22Zjiqzx6donhE0UTMFWwJqYZOg2D5qzh73FUDtUs4Q0
IWOx3jPyznMYll0/ZIin+uTp2JznEn35ZrhkauG4UVqDJrEIw+cRvN5i8S9bqLWqGChMUaxlot8j
mrWFy+ixGyYHAIou31leqr3amKHTAD6tRA9Eya+6+eM7VXhjhskfJdYtUC0/SxS/KM4zMrhhtj+a
Am8I5DhLjq8Cq44hz3aT27Boj8u9IKePiYkjzXhzUlBU7o9OvK3y7l4YX/2WGWYlDIo8XUw0eY4J
ILfxjIvMCwyrh0KveV0tmVhx0YmZDDtKPZlyBeoJ814wLLI85ELm8DYUsqkSPp60acADbr+tVST7
+2P9VLn3kAFve977AVa6fbSxMfIxkCsXHFXrfgn0SI8ipgniORAtY7Eb1LqdVzOQv7rI2+SLmmVO
Vb3fYn+1b8tyenMxitcvLaJZod83wOJ39tG65/dDkIsT9MSatOOnjsbjs3+55zIHIgnMWS3LCTJ1
hXT2wkHvVXW67gYJHpEbVJuBE/xPNrZIcMQbdRZfgDcDkYnPEWewSeDNNFgF1MKz1RnGGPCQC84N
Otx+WjHcz81hHoqO+9Zv/plvPQxJrQhsoxULo5udT9vviv9zVK8I+UkQmcmEg3/iODoAeZtNZZAJ
VV7PeSv8BTFHCk5bw7QF1WS399LPISK0o2oPmRtNeAWQ2rNgYDB0ftQJyL8c0JTBReTaXikfYawe
j0lOR2qB2saFvA1mah97+XyW1A8aFm1aCw68OnE/uZYWSQm0SNiWgkOTYjT6Jvuk1MV+nkoi+0Ae
VQLBWLiOz/AnzMk8I9sYhpwin89sq5Yrijg+6XyXwscma1+4LhgW7sERm5xtyWMwrr0tHyQyhR5d
qnFV1awMLNO8DWyb5STE6kTYci6M8M+D5IgHVw0KX5K2tWk+9p2QaVcHcgsIsdbZQjUAePFABpa2
5UqyDixecdHuCkuy5Rr0SwhoC8LCZoA2I5K6vxygYrNuAoVcpe/DW8B1KcdSNQOVlJNrvQl3xRzJ
OW5I4rdjKWYvW/jFcOdId1WmFWu0QAtCmtMbRCwFB9DCezhrXCkR1N1BUXBLlBOa06XUJ3VTVl8T
oee8Jx6PYlEDZsYpzPoarJoTDWYE5aZduqPNOZaU3iqoqChehL9480fx+Nnh75w+4MNqLQAIXdny
yTPeSKIjP41bGjr89d7vfevYJeNvDUNTO1YByuAtHmhWG/b60TzAMjXRHyS1ktErXeJaT6H5le9f
4WeA/FSAaZYvM2ULBIhxHgUKrvqzTig3y78jXF9186kqc4+NFLV2viswmQnMmmGfr+zKAGd0ex9W
D60WE6P46y2yYmsPfQB22luqGstoHEGq2ToNP4Woy4r867cfpefQO2z7TrZHZz1M453dDy93dUWj
c56KMVBd6LWJSe9OP1xxfzROMT7KXSasMutcZb6+l7ZL/OEHAbjZz6Q23hWs4onc7ljECaZ6lmYX
ZO6ergKaCXYLNykOCVQa5Ewjxba6BDk+v2meJ3PovxoH437kZXF07jJDElHkmjjaCLOCGgo3FSrH
CuSvaNvVwBd1itVQ8V4R36WVzjDdqFeRJhK44bpFcqGi2rM2hXO5LaIM+keQ+bdXLqiw2+l6hvax
QBjm4D/USN7qT6F7MraKxctHRa7R+V2biJN6ABk8WDXFjfghaLQYQ7jAHVVVLJrsPk9dyyUTjaPw
/UexRFTw7GQI71Gf4FiuUWUYiWENo2CTurFPkxnz8yiVhU+d3D3Fh1IG88kcdAeTUbxxS8WcQADt
aIUKlN/9iPqBBXZlghGtjH2DJhoH/LoLFc7SpBRmbI1KMdb8hpBSCV2EZT8Pe1VdvzkGcLmAJLfX
5vQiD3JA41vybWSI2Ya6PeUNKQhXARA66+R+ER45oxzl1emiC1E46NA5rRkOR7wvrpBkCkbxtsfi
n0byRU16Ek+5MIYBYomZwqAs4EBA2K0RA1noDd3FFthRqPlmjxI4lEDbI6mVHvxaZAZ7tH6yFn09
wGDvwj6zLoj5VHRPfP4UdtbqqU3Y6KbeXRMKk1n8aZ2Pz2em09Y41O6sePya6TYBrGw56w4pWC1r
wqHB7JeEGSnoQnm8lOOio045oXLg/C7gdEBUH9ntU8x1CUu2vBqfp5Pd/Q4H4oWjIhApd67USD0O
KkIWP7065qq97avW8MP815vDQORIkSGdTuyxlYLLTv/uFNCgLJJbRKOVmr9XFgHYxbDlKikwknOA
2AYx2gPdFTCFE72jfl9BjI7dt7RwAzvZJa0Z46Zd4S7mltFJzuCWwLmBIfh+JTX4Fq6Lq6IoHIIg
xUSBtnj+y73oJDstKtLw5cKJ5FI6j9JmFAqIebuMevJLCklz4/vuRKUmKs/XNzZ9DQ9/tINRfuK0
EezWqGgRslil4lF8OsqEtSOdtuiTlCOEff9L78DTQgHUiPMwZkoiQVED73n5sZZWro2MEljwycN2
s+ofWAn96dR1Qnyfn2CyzESECp3ACZoaWDYzZQdNmHKblmLPE3HyBU474j3k7T7G6w/0VFA2z2IV
t3RJlc+MoE/kEqMq8/TTymplx1JSJ8+Wwo7YkeAHwPTbqwoUF9GIqmEW1tsp+FXZu3+sSj+sy3mu
dIXsrnrdKXJznKY5d7x4fGKJNh/oFPEtBqzfMiaOKFh+yI6zTxGokokZCHd923q86kY6bhlnzdqH
7OMgRQgEIpgTwig/zgzqkiMq4dWW73TX1LnVU87SYQVBOZqxQJctY6H/m9P/PIDSzo24STYfshze
iao2vo5ZOBLkXPXuv5K40N1olthsyRT8hihg533I5oOZwnKWqfrnY1eyS+AuLm3m1C0/ncCuFJMg
lZY6GY1abSMjxFY9M/0OtzG5MzqLy62hiXo1yF4wre/XAg+D0m+1/sbl6u1VjEIN5+GP/7RHiHc2
EH+DoQa3tl5w2MBafzf2rqcyrvVNUknE7s+rgMdASFCB9nfeWakuYQqruSxe322ZCSVJNGFL4R6S
1YJhT+nniqOZ7FQZWrPYWcDIoruk6uXXb2ERh6VSUi3TTP75lbKDppW1hhd2TtQbU4pqNLGkouB7
OzorgNKjdUUyq6KLCMHSS6DVisKFWFZABB/n86C7IMU65cP11pbtpV+oqhfehDOZVfsmRJXOJwVI
FzOh/9kHhe98ODquhulPnBth09ALKG66ZWAgVEhcPFmRHCRERMkQjL8tGHfdhnP3Bkl00maknhrj
EFuliQZgO2LE7PxDZ/XWUd2E2BsIIvP6mYwFKrkafWib+nG6rVqFLTubrljoQFYZqAmS1fPhAAqJ
6PBNuOBPxjUSk8yGQDGeXQe4V9ziVGZ4VZE2evi/trqvAnrwAgXACHNGgbJyZHTWLNaHJq/V06mi
k3nUvMiUO89HBS+B2oMhUGwOeR2rwlOLkkk2Tl1pnehUdfty5gV1AJkCNX4BYbpmw8zxC+mFUX8p
w+5SgoZiqnTmaLEc2kOw+b0/bb8bku+tXLjD0voD0CNJPrhgK/oCQYfJNk7YlX5e2tgrp9bbtTUk
ONvoS4cVZEcW/sa0LK8Itba2dccIRZ0vZ/t5y4Ar4TT1ieHcGcH5TLiStjTR/42hZQy2rGDCNYjS
diUgQ3dlVlw6z0G2Q4v7pl9tjTVKKitd78QHB1aOpLMzLqSycOOmvsfNUdybSF1hQAUSawrrtd80
L7k8QzmIaXr8km6/Ffy86GkypIZosHiqZwqC1f8RWbZeuIUH9MVkyo4L5+osxGojWYh12htN7Xj7
E008noKWv0DX+FRCHI7noovGSUPSEC5iFrkL2L47CVakHJIUlyxc8aBWn40/rfqQTDdklNeHbnmI
s2jVhULbG1CsOfmpn0cak9jDH+bhBg2D0vsK7dHxnxSmtuFfVLiCb20PLQsOWlxgVAm/FVGj3Vko
BErIYJtpnlbhWb+wBypix0FNg21ntlMDHwJxWsK3f4i+Qa6VgpSwaO/4IET2KD7BbFUOxRUG8ynE
Zol0trWR2GtSoNIhL9XpPQj7zDbn+vtsKb6PNWkXdRHvTeam7wIN3k4O3X9bLYHdgnBYTutVw6IU
9pcXhO3N73PqIcv/hLUa1vnAOlniZzNaKro78aK2vIAj2suNQO40JL3ShLRfAHklEHa++RKnsGoE
aFdDz/kgou1545VdNOgxIJE/jvkjkiMmW/CYjzKYdtgmcTYVoBzDYFMPzhwO5yQjN+Mu1FV8NQTf
mI5Y6iSKyiBH5iEIcNYjwYATd46XwGFR3aYFPCf7+zUatOg7YCQNzU8IYOoKrTbYFrzH1CJtSFfO
r33nl4kB4JbvBFfs2oQkiPrzF1aBFM+/2ss0Z3ZgmQ7XX4eaysoV9+cGazJr6PIa6D9BCHmQpKX7
KC+JdP+wAiuSLFTA3V0D4WNYvUftoPoo0p4WgygXFD/GiEy4lOR7AaVPVKGPNnP+I6/1EM4YB/cG
PQlf8iX3BiVGoq9REZDnyTQIjhYu9utf/eT3ydMs/ZY7oAZEySS7MigvceelLEz5GwgHOX6wcyg+
r87km4PIvtEqGjomo0Ml0wszshTM6OVNIw9EE3kQDjqc7iBiI01N/UHefR5sNTBom/2ryBSuhKtT
cC+hHZ6kwkpn5jMqTlorg0GsKb1pmpH9tnfZloDEAftEjMzjWaPlL6zz8PkYEzvG0RNyq8UV84ku
Kd5wjebfqnUvrWq+VByu5XP7EGEWXBQPgsqJ7dGPgoPal4O2oh7X53vsPAhKURvkoUlVBGPDGTjD
AWM6OVfhYvukZgbtR14EIf1XO5QXcDkl09P1iHFIgPlbD34oIDODJH+zumIO72De8nD7Mlm7paBS
X0nfIcpmOa6lJGbHf1Bh7W4e+2QJQog9+R60UVOtDQ2Qd7ATMcC0QvJTO/EQCfzLUjfR/LjW6/U1
6MWnJStKQTYhAolEsCrXrxLN0kuj1aTqnnquiKwNpqI9+rBaflkuExKxFpAgW85tPzBrcLtJL+om
sNsAk4XJWwG5OthY4jxdPAUpGX9PudrUPoFebzK0jOFIRGQw3/gQG9eFR3JNHQluiH86wgyF/tEm
NSItaBUGyYPSNCrFxYjQ4Bu9+ngj10FQuyCZzMHiFFmaigzGWzead/+FBbgYJveOlAQHOsgbPYgY
bZSZ/P6DLKhgUQQeoPf4mbCfiqhJ6H22Wv589ikAbCFQ0EQdplTsYOyBLZ7fnQ7jmsYCQaZmQ+6k
Cib2nFys2nZQhr4Sh2BmgjrpKbAT35EIEFLROzb+JMq2/O7woK7myr+yEeH8kG2feOuZhdiw6zvD
5Bfs+1cv44MxF0KlsFp3aZVXyfW1mvv/cNjlnk7OhPN+ZPtA2zW8K8yVZnzFE2luYKavPYHfPNrz
n8/0UYAoYWzOWitzBWVZnMnpjhB3QounoYjooZ1w9U2BU6oh3fWWZXfBPOOQYYgoRGPrHTomgQxg
wEeGFjBtU7lCGLmwFciAHTcqrDhpdJ3vQ3ALScK5WiWTwBGxBqntkHEdyBXAAbOdU72JTJBsk3yd
5ilIK3ejrgwlOWxzhyi0p+vfaztaPv7w0TNKkfZr9jXvBWaC36MS90sI41rCyBP7VN4dD0TYdfkQ
7r81uzG+4yplKY6LttYeBFJSSGr7FQeShI96EPpSlldO0FNw7aMt12QB4VpxCkTGdc+4DWdarrfg
5Tn7YMOUiGGGN3hStfdh/DZChgw1VRgyrHQ2H4lJzHQtfz5rfU9+nTV7pajTqVPyZvy6Dw10FC6P
AFcn7toAvwU/btDJZ7uQQJaeK26ieTAgC4UTPDz6ujPtenNZb9xs2i7aa9e1uvPPm9QK45/qMmzf
DsLVnwIn7beJFvuLmnQ45y1CCuK7IkcCpu4RBZnIM6lgsr4j8WowdC0wTGiDLk8Q3v4BuAuAma/C
C9nUhMRSiFoZOy7MNjHXJo4djAOphrq+PU7rqJz5vTmcr8AQoO/e3RoBYtd63XeWSRPZHlKhqVyN
TjXfLEyBgVQ6Igx06j9jBohthziwdb/QDTrGwnArz7SoeAIpc9VXHlKlhCIZhEugeST9Js+0wtLR
p4IcuuKjobtH6sYFL+lTc7vpBuiHexKJ//qLET5U2dOv/t2+UcY7NrM+RJS1CpeQC8DeIGMbdZAS
X8xGqKpXXK0/tFksJD5tlrqUG+VHIzdSfSL7SfsCaSm0SNRFGjeymgdEp/rIK4MOgY/zKpNSmqV9
dI+Tec1Z3CeKPF2LYB6SUnCOH1T+qBlcF4wBRrIuvhvN/cwd/6aNwP7oowDEf3bJfm48JXVKSLjP
fJ0GhvqoZV2OQFWVRwDIuoQ4HkJR7NANl+0Bh9ZU6LRFEjM/pfmlKnCCZ1kt9qwazT4MbObrs1sF
V/BnvYn8BRJho7jMa4oYz30TLcuXka89pZwwZPECQe9gvROErVU9XiqiTydTralbOzUY1maUcjhF
+FoTU100MVPb+JDYeImu51Oqa/laL0QRVfuCziQ/C5i4Plei7QjRuOn0jTEcJeLy5Fw2/LU4kNJq
+KI+dtOOyR4GOVZEsJBn4Y7Y3ylHPq/4P2zQWmQ+pYzxex0m1ZBEtFJPIX+0crmsBCOaNFz4z8ly
CWog25KOyD2AsNIFHZVLk6umKkLstJRafX/BeDd35/MPu6GQgtDu+LLJNesLgsH7JXnNTSQ48oLx
7bsoblkSIfODNPKreV1VwHJqMShv1bIOHyoBUanWWq1kCBM6db38kjIurb8YUqYR0rORL85V2vNL
qEojDVOqAU8jRamJxPuTJB3ciRkCu8FSuXwB4hZ3czf5c+Og68KcAW+ioKKKM1nhpWYRPRpROSl+
SrcQrwFYgqc4/KPS0FCnIov/0QbJ9l4LPbatVWMdOj3fhWnyJiAESPZ7NrFhHx51T9Bl1XmoyjvZ
z8EwDX+6Jw6G+RtCWFlTvO4eq+sEWnxpZu/S9SjB0jPFl4n0vgZ3MrPmt0k13Mnx99420kZBss3B
s6mmGBEiLxg05mRoOihaUm2O4UcPY1sMASY1qnNHw/jqIuSspdpXAIvLLXLVnrwqGxLLZT4adxrW
mac2vKT9yCcdpgSyUXgP0jKxoqnXADJTEt6zziZGda85fOBhl0yeSxYWay1qySaOoG43ChNc47yb
YerztLpQsrDUrWjDzlIswhOOagr5oeb6Rh7gh1ued+zAhA1H//Ib8LyKHCHE985XiLQ7bg/puZga
cT8ETcsyJV2YIXFUhDnK8+axKKiukp+KjQmzQF1o3Z7BrLX8Ag9mmvIPYTaMVv+mG2G0imvHbfcU
uPn+aYzM625s5mLe3kiGA7YQy00KDkXwoLYEiuMb7dpx4yZFaptta65RItQQo5iRRRx9YtztCOiI
HCgwT0tt/0qePH0JTkGLKzS5bdl4wY/nOBzujyJ4+ULEj64v0BISH28t2SOoOqLi3BylccDzx4g5
6rq0vxX6k3qUFe8arKbexCvQz2bqIqGMqxZd42Uv+4COSkPyrDrLPPqLuKeMXCESevtX+vHPa1GQ
xf+SLulYA4vXe+1xLV39sTWrt2BhPwVRX97FSBMH9r9Ud29vEL2V/r0E4RcJhVpB6Ej32V3mUwVi
Uc2QnN3NTXGfFyXWBiDk+Wpkmo7KzSOMUSci1zlzU9YvdB0FlBbAgkr4V1kQgSsLHVVNL+gC7dk5
//7cFddA2zXzEzwD7mXtzw1HqnIDCDV9xhlTVkIESJHTcOO/2NtNiDlExE+mg4uUzzN89B5XHe7S
MzAWen2cld1XhNrXDOgVQzFbGLxjOIGGRlvyAfg7eq1pEgvq4O8QPIO5jrGFJwbkXO1JbEUNrbmW
i5j56RMUCqwtW2kBi0WpIIT95w7pX7dD4Z8/atrbntwtFbDpMXqmLqYYZpLdUalJlzqM0LhjCfT5
6qW9e74G54yxS2B69H/iSFeV3h9Sdf+biphNHY63zont2OmvAAYQn9Yb9lp1wH1oCpGD+rJr4bWT
ke8OsYd2eo+vRbDFl+K8kOp+YrRXfcxO1eU2dMBeHt+fppHj9JfVcB8NNC4Wn82alQMrm1Tmrtvb
8GN3B5SP+y5spokXsqgngQhourL5ukgH0gBXkqFDe+t8R1zTB+BVHZzDnT+7czEbnlI39pB4gY9i
ThAfUtH5pi3KRc/u/+T/Tdn8+dzrDDPy0KXzqCPapSuyiOIZ6hyz7do8rWnXQ8koIBGGKoiyjnve
HHdJmhsiiwxEiQ7+0RNKZ9RjonWJS3wSrH5iY9+0q8qdE5H3PUZkcO5DBReTMhmJJxmZDQjHslgu
mDZSzuVCmIFspDeqGQh/wL38xV5FLe3s4wNQvFiTHXhJqJeHICltGkw9JU1AZ7OZgDcVEBAu7vgk
6hVlaG7ksZfQQmbIHfabPCULcJt4mMWfx/gPMuM6eQQbAnckBsgD3cJNjArnf5wx7pRitIaNidqE
iFn2VjmfxRz/EsjFhVj8UH0uo7M4jSrigz3WhbHgP1te45GkLSsVUO1wj1/BWfdmtS0uLtro7+Ev
Pc92RmkbDnZ8vMoxEBc4HDLZeNsjGOxI0UFWDNaIVZzgISLLsBYLhojpaP6Dcslc4pQbHJ08sX8q
ubcfwd3exoo8ugKmjeScIXX7zAKMRuV2mSRAI3EQW0j//8W2Se2ZKC0jKzTMWA5SIsBPIZtQTURq
lngDv7wxovWxU3QUO88anEFUnbbjDfTCatuQaZS0P+dQicN5eiNztqnGeM44VdTTETayjGR8o1Zk
ilPCOfS6w1BBxH1isFzX/5KSN1zqtbWgWzsxZJncswlVgN3Q+qpdd1ULmzxkG+pH5a/6/tlkb0rz
6YvkUVabDEjPjfP2EjS7G6CIXclLqUxqWqPa+g+cK7VuYs412pe+P+x/2cg0lQnxb4SCXE3sNgyl
Hh7jmv7Dc+YyLQv3iEpW9T2KgUXCSp4UqQ5iNIwY7iAYSdbgB4v2dR+m1Iho0IY6nh+6rUVeUU1s
Vn69zWGM1twY5E1irKv+Q+drdeTmUauvl3kcWAtmo4MIJoM621ScL2eyCAcBJ0eYosWTBjtxBv1c
ksnVf+w/ATNyouUcbsJSW1qEeM2JQg1dtANwGHQVqXH591z1jL9yoThlsg6u5fI8Nt1E2g0vMr3L
4SRzm8i3Vk08JZrkLaTHLUs8YFUrVf2bwY9V8adRMhdV+fGnet6Y2Y1j/KSgEH2bNm3l9ddfORv7
W+L3ecnoc6Y1WfAsnH2lj4DsVRBMnM4EnSSkP7K7llhkjSLvVqJNVl9u7Dd/xY3R3Q+w0EYB1FFN
a6k4ga+/Xgyxlzg874oZWBZglqLIjw/+UKvEYamdJ2EBqb5Hm+bNMH9pgKVd5j4FFo1YmdKgSirJ
zLwZkYSfyku+jyc6Iy6P8v7P8y6Kkl5gBNZ6l6BsMRTasN6G4j4DPL/7ruN7anHdgXVjoQFzaxv6
oTD94Im1pq+HpF7j6wuRFh5SEKsC6S0ZV8ZRvRudtlHmaicuneiELIZahfPXFLq3o5BmRNzVzTj7
bBYPxDTE1eC28y3QkT7xxOCj0CyWREuc/BiPraXGEDTJW9cgE9EiIySqw6bh7//yUkcBoeufLovk
NEx9eBUQKF4wvh4rQJBICDft0NRpdjaIlAyqsAACwZC5A9M4anog/JuFZpfcWzm6RkPXPRA8tu5X
+R/BTCQTLWPs2Hg7zbDBAqXHJc9Gzf6lZELWbcQFFqjViQ3vOAtqJg4njjhOOg2QiDU9TZuLUwuq
u5XTY4WRpKBT+yFrPEdonSqnlgAyjxIYCOrSWnGvMpeCz74hBFZe5ckrTnQQ0CasxfYcGUKQcaoo
IJgdp0EqhRFZjnFTzbGTn3B0u9q7CPM37fWeIE934AjwbpCntvseqv5mJzkFVq8Brtg1hVMUUBuZ
eY0sTVTin9rGTOV4VRhi9YPK6RQeJ6Kyuypy0o2+zM0nm/BIMLzKWWQvbiiwZA3TF+TWv7/i5OR4
vzeJ5V9/JKrejcd8LBcKf4bPXvIrbZ5aMy+m+p6Svt7+2Mw8/89q7zrxZkq/7KVm6M3jSwSaHL83
cgopiMh6Ny19+rgcx61pjzRRuVGEmCBJklpkPFAXGwGY+89q3qTpvtjBx7vv8lMELmjx/nk/jTNh
DjII19pae2mSrSGIQRZich5Gup3Ghw9YrEKDTZjwcBaL1/nauwHPpUIs3JCogRInyNVi1MZJkfi9
h88BigU3oKa6a40vbo5VMlrIH6pmNGMDC7p8PfkqUY75aQBPqdqFJ6WTg8J47LoTOH34s6DR4YqO
gWy6bUBE6zldVNUfE/4haSVCLTzDPX4NDT2S+dTlcRiegKMeJ9LyqPlIr2SOGz8Fy4rwBnz2Brsm
/tpwcitz+wwyisjm2Z/2ZsCSonQnnQ5NXdE1pd1L+tgACVWRhK49gFpZwN8hwucCpDM95udieCXW
KYnNRkiyiASvZZ6gmRrXVk1zikxHEZxViLbYCyRD5uUEs3J0vKfqjazGcNbZh0KJxkl9xRr8AUXP
kM72ylzexu9NX7KJ64dtlMeMYNSxMNeDpKG+d3QMcgmDp5eestNFHWpRRxJJOj3CmDvb/86/73Uf
yYiZlrJwXEM18HNpodoy4KmOGexHJRGyYPbYfewTF6l3r+TsPMtD7vFAyVYR5e2pcm2GQx3qkB6C
ftnsYZ3+xx6Kt3Hekkp3iOw0DdyffXfOfWVllm/2HCUYyTSZGv6GXZOdO8Dow786js26+i7bAvr1
klN/y477DMkbXdQpnI6WDpjI/20+a2UGZgTVYADee824X+kdM9jHpCu+BXRgC4Zl+pn5jwmECt05
B1uadVm1+O8O75FSfVuDliEvl3VR8vmETwqxsyRHI6rP97bO5JKGg3OSa6M25Dan/2Tp8OFTLIOy
l+MQoN+ZhcvII0YXg0Lf3mtwD9o2raUKwakW+T+FjT4NE3mR4KPXS8Jvp+hzW9YLVodc+DiKiNkZ
T8y0qcCevbzysYNn8UizA2Mq5oJKikasQ8jPiNmWO4NFa08MZoukrQCQT8XelciQoegA8Ue/7KfO
GdrNvHS1l1c5//WhrDmlv03ZPNiF14gZhNAC4QnE/p+hW2opqmOF8MK2YBWam58Sc/j+oFQw68X4
Ua2FARGmJXcZiQNjxS2o31k+lGzuK/tqSx1HX2hCLB+snh3q2/+zb6Ie4Drpi1WFIMtqg4CKw8mW
qtSRQ1vXvoLAF7PkmKCyuh/Z0nAIWvqQ/V2Vt4b4ylP4T/YEA5Yp6vxKjlHaNc2DUJj824tNn6wC
4AomymjMVRVV0d+raMEDpMAwglW+68+MkjUxpcx+MK6Fdl/1PiAbl3iZZFnfCjNHnqfqaEIIsUNb
QXXT0MrlXvwVQE/7PR8nRClKEu4+7juZDV4AAqHJKRvUOACRAWuf86YenCSTvqel1Lip/j8AsGVE
J13SA9J8cBH9FwPuuJOzS5W/Hr/wogT/LOsPyQj3IgSHCjkOs+POVBa4kju42YgzmYQ1wur8Ue+6
+NgwHTQ0smhL7xiIJqjqLWMdL/PwUHOgT08rJ5qtVbeYNfctHq83TkiEkU6BN2gmeVxJZDMllEH8
LYNNOA6pqr1uGvSbT3E9FGjsBDtVuZn3tXjrQBrPF3ELqtsInnJR+qNpyKX2LO+h1eAl433yRMUv
LPhgoeYrIdidogKj76xMhjXZ3dp1FMGau8HcYGztW0XvxxHcjpMInWlkRZPNMv8gllB/7x1RGnFO
5vZbDl5OWYj/BdOWa73W3ZYKXZa8a2o4HnzHeFIjPbfYDUnxxNbe5kHXngswAy0jjA0tYFyVhlaB
50mmz3VLRPVIp8a4ebPNsh6AiTAdUkKKUZoIDxfx3L05DZoOahOn9uXAbzLDW7RXp2PqxF2s6xkE
KtMaQF6p7NU57Poc+ltRp4vwjPDvq/Mknot7QxeAR18peMHwCc4tK70ch4s0VAVhBFKs/Nbllu7w
6aMSieX7cABG2KE3pcd/6/q/bBm0Vn7kVtRFj+SIkbJ+rKQCf+NcdWGrOJl4oUYQa2H5ILOdh4uP
u8GPcOIbJbHucYanFtP2Saua86BtaPGdUv5vS4atW55N35hWSKBJ7XRpnx+yWu3kZGv4DZe5FzU/
2ui3o8H5zi9X2vh72E04QoSvokkM8OGudz7VWlc3aIdk1MK8pojsTN/S6WEeCxKxI0LrQJGcVG4G
GOwRMaHt/w5+dzAon3b1uZGe4aUtOPmAE9Fga0A0ZSH2iDtY5toeCD3tsizj20JlsW+9i11GU9XV
IhMyZeu+ke6j6Or5/DMql95FsLID6O1cqWlDp7J9MeSH4abh49gWDrGSmNFS7dkWG5DbgTb0btlh
qR8IleEgRBjdcUfIXYF4Q2U7jORS/MouP4OcZmOSN1tspLFc5TT/Z5JACPIYY72ehhoPr866eETo
FPVYtA5HcPuizengePK3BHYOp8sb2ssQVaJYe3uwgd1WuR70BfdorjqQaj+YUMkkT4HSmky3Wv65
xLdFmphB+vguO2SwflSrYSQPGU4/tKnloFNGswn8Tlcr7iklqaNSbfjoRl2PHYZ/dYB9j/WYS72R
I811/vRrEdVV8EAX4lq5dwIZdsIBTT1AVB31vygTlfIRr+/x6yS/bMGuAEH0t7ypTDMjzuiWw7ZF
SRV+ucf8uMhncf9lsqtMAZ4NMptscTZkXWUvYH9ptdvXALyFSEWB+rPRLocWB3MmCE/TDSD/FDBS
TZJrX2fSJHCXMxH/zozkpuux5T0b5XrtfLRSe3SIhzVy+AO19NHwYvH/6Ic+adv/fFjfB6edTHoH
zlHrc7uw4dViedFyh/NeYI3vUmFp1v2FhRMX45WZrIqS3tuvjJuifLChgE5TsrnAeJJS1GpoKJLJ
+D6JEg91oM6kEt3qBE1hoey44l840Ytnz5WuembHnL98PZi4X3dkyJbB83t9JtFtrnLCQ8AKF5jR
504O0/0NSaUp07Q8OwIWKnUsO5M/Ujizq3auhlcFjQXi2Q6P2c7HWJRJRz2IYCaLqLuo/e2xBjBc
fUTGf/B9OFYY6GSb747EqtfWMqerwOaWJLuAm+f+KMHo0rnh/lKfnz2ezHMa7YmbxNCyZvzkw5yN
PMCmNXEP6BKxcGBwIBemvj+IyV0d4FLVQRx7DAT5V5gW69vjv9sbuuH8SbqHeLGftWCZ2uXp2Xqy
9BdkT+7lsm0/PQZgl7CFMYV+VByLD1IXYDYu97zmMlYe7B+Hy7gPNHlpbhncUWMS1p3ryVkrD+Nw
AXDyO0AY4wXzg5Yd5rIgr7nZ+Yf4yd8WmsN79GeI2qNB4jCccFAvytetu5AHsS5bVjFYTlImuUD7
9UEf0orU6FIuPAi3+hFLKe62PcrV4vPwOyIJb0/9IAnj+lfMqw99RDZWwAjzcSKvukQgCMC1OimZ
0iThr6H5uwU4xQPbk9Om5n54OhI7RE9EYrYJBLHEkFA72etvFyz4po1+WZrBLKuIew79gmWd0Lgl
NpPHJQ9TNCDAwBsTK6hfDTsEczPZId1PQoJsfEWqjuPCDMMMFVGJAo5BP0vPbJnd6bYkPkbtkvr2
a97MjXoJ8A/9nvCf7xJabM8ICyhLMY+On5yfZZNZ0T8frFlPIlLwH1YpRgk6ERfQGbyYLcUjIvIw
XY+UCZtzmETTOK5iVqGpSGlFHMsU8L4TgkUmCuqHu9OKhKHL19i7QcRv9/wC7q7AZaZeb7SlUu7j
nQqcoQpwlPGivFLySk2UyH3BBirsDrCQWA8I9Coy3FUyu2MrrNM63bFNaEXS8InrrHH33Er55SNu
PCRNBIgQCr3jL0Xp5rlBzzjRsDeB+/+Eks/IOyJLRwUthqzo7En0ccf2fJlRKjJXpa3qMHEH7wES
er4jXwyXUDJKOR/2oS2+lCQM0kN0HKfMkZeBf8hH6f5y6QsXq5K301ICdEB0gzrU0cXR7CDq7DSd
Po11biZw1GgWZG5JczfkmGdvthds0e0LuqrvpOFYCE8leLPlUNnW5MrgHAdYf/e/E4tl+f8FKlSG
q857y9SaVWgyzrOOkBTsB3voNio/6d/uBLvYaaO7JTQpMAHQoODSpxR4eIdh3zizZdp/Xfz5y5g5
cYAeazKvSMU0eGd2cA+b1+Z6/836qgt8+wy7jaAf72BIIQeQIRkhS3BdH505j/7ePyus0kVvhrt6
Dl2jQ3ot1lqLazKqNpjQrM7ncp9BkeelTJ5FTGMEReBiVMGCFhL842QsNWzS22OUHALLfHqnYzay
wScduTZliSnUzPM5T5zLBE9upsJFI+NXW+1OKAdB2ijkM9Yr6VmG93kvEr4htQBOY4HlfLbprlrs
9jb/pPMZZMhgZBmzSBEufXATBeoeIYSu7HZhuPTEHlxSClpdg6ueSWxU+F3HTuYpxumzjUw5qpzb
96jWBdlap/M8ABGTFZqWxi7i7oCs62vQxjiuMRwSqFHcAxQ9HSfEFK5NNO/PE2QT02t6KmmFmB+8
ukDMqb0ldFHbRqu33a1zEZKUJfalZJfX5KoOZrt4c0Sbim+LlB+9bpyN2aFPYO2/E+M0nskIJhxF
GIqyt/VJeVKcQ+jYPbWj2119SNisbvDtsCc616cmHW8JFWZs9HHu96Dc+EWftm9zLeqYxvaw6FV1
PxwC4+9yyo+xU5KbSCoBhWAJsj28ZHZjp8Lbizb8iruzUJD9w0SqzMjSCjSRrQqyv2+WgPbRB6E5
P3afKv0d76/Z16BvxjqVEF6S6kn1qWQANJAUMDYFkknEomwfM0bIBt/fkEgFiA2/JW3OAJd9RFTg
NOg4zUCBNXzZwRT8lr7P7lJ3MbjrxYpWTtkUgT3YKX/zZlfinFh8Fy5+k9Czv8n2/kXWsfqfz5uk
2XHk353uyUNwCkcLZGbObOGdf/s3lK38JFZmsqjGPc+9U6Hit7qQI48SR7G+1pHCpPFr3Uv8wI0E
lxgFkBMUM2/pU3EtrksQSYKAmSLlHLlr2sf2YfLjZ4TN3UD9IXBfozoDXxNOVY9rPLmOFzIO+lZd
2QNGdx0gFRnmLk9pBGeK7g71DYjcJTWEAZSB4E7/4NvWUELEI5FpTllO6r8oBFMAYW9foET3rpI/
VHc8NzyLpUEqz4I6wPW7XWHGhQVEPLIdf7fQBrwpwAS/Gxct0Bqf3ixrD7vuNlFQsB/hB3pq7Mji
62GeJwWHT+Pbmgy7OFIQ3iDy80YJY2ZdilMEpg95mpH/W0nbm/UcaYIFKeBrLcMswN2yQtWH1Mw4
8YDDX9VDUYpIySP396LzlqXX5nmBIIOfBV9Dvqp9Abi89yeZiZqKzzGQ6dP435GHI830g4UAD19P
qZsumNdgrekWmjOHKuEPV2UkCy/I1zhagJLppXDZPNeghQBngLrdKjQBABds2mDH9O9dSGvqjcMj
gZDK2+el66k6bskhNTmAMhAjS+sL9pIhW8D5I7Iiq11OtlfxSA/QnOfN00ZeFo7InvbBs3zONc3O
ODbAgtp/7xH6LQYFn+6j0lcPvQirUg4wjRoevY6+LENbq7VYTkQA63q2YPbYhbonQ3H3AuYnJF30
sixyDqqTDBDIePnI2r8bZEAKRzxkeo4on1B+MvaIfyx+62FYRkFXWClqWCea9o8I9zUIJsMEDwpk
qdFJsexA08QfBGsN51VTy2vV0LK91okyqS0ECSHe8vkqM1bpFcxpxuy6innSfXDcX7R1C5V5ATjt
Sovhfgan8Wy9e5YM3RQFDlB0Hspg+5/F/sWoTGg+eQtND+YvoQ8FkYQQZGIsC8xNOoQUAHeL8Dr8
W+EtgNGGAQh75yM8+dzZYW9lKrNGpp2tshBCcyy8TtCsjUOKwICQBpVooZ6RRbcFV8PEQKrCbu+p
wY/R68BNs1QalvQWBsKtTBH5Zk6h35jCSvebtRoqeSjITypJSAEmqJSn+5TvI1mzGnR8SxtKqFr5
wp7PCUyQxTbLPjobDfOTxIbryM9jeY7qBGuqYB9w7kkDeaPXyYHvHoO+muYPjR1k1OJfO/eEhNTm
cN2XzxR6L57NBCpt0OZ4ifcHC4PW8O16JA+SqwCcYxwBq3rhWjRgKrG6dYHVRZszCkdZXZp4EQSE
h49E5RwdA60IgXM1Ge/hKV54LJGKswgf7cv1QCX5HmyE3hVxvsInXP3S3TbkWfRujuo9NpVfOluS
g6ReBNuaA17GKoo56jnBJjAXEayjSdOWkt0p8OkrIghLBLTrWGMNLk2ZV2JTnXxsBpluF58rrApR
RcwycVoxiyJz2nk2sd2ISTBZavSX8jjNTeEcWuO8KF3oOL5FQKC/m2xeb1cUmOMkUfK1ZZXXVk5L
aJVJH4ul8uwOBtaktPz2o++YwVWTM0VXX7Dsg1pTJuAY9ecd3DT608spU6oOixmuLarBnGaEz100
Hq4kNNfjr0o7/O5YB051APHRScoM6izuIh1fw4jXfSIRQh1KHOaPwiB9IqmykDkZ3pSChm13gS3q
SyxCDhsDbdkwoScW6Ywas6v5erylnGQ1WyGAoQByXaNoeAB2efy5PBhgxNgrkvru3704X3gRytFw
sW+fJ7fSL+wl+NHFXyJikzjdrbh5Eq8cZLQzN7tQ+vblsankYhNsFB+XzjEr1nvAtXgA43EY7Xqu
cymTesrLqq09fbTE8nXjAPUaESEtI3iypekN4QiALoAR6yK7HsJzpLAb5zwfKeIdcilNzBX0CxmP
v4WAqzJ5viDI8H0hcU9jA439h/o4PhZTS7JZZMo+kyhzeqJ/CLF5XKOGjKb/eNiYkwOxF2QyvBSQ
dYd2EE2SaBOpPl7YyMm3+yhGqkItAjdodF9Hlo6gfiF+BHSvEl3Kt64qt5RnZZh+KTU1HYn50wUc
X61Z9UUsT5dQksRNasucIEQGrLg5DHqUs0bo+rR3VO3sO22RZLuwpAYQORJ7FBjZsFz9I0au4gXw
V3Ft7vlNreCCZmF/JN1bmyaPJefmRpH2qnpI0GQ4Is1NdsS4u7dVDsR3VqCtup16dYT6hKHwAFCG
tCNP+mDa4FLOls3N+OdVU1SjXsWlcDAk/1LxCEJsmm4/Q7kXFEya7zPBbSrNcEsiS/BbUKuhi2o6
iCE+DVZkQFsf4LavF9ykiSO6zWX9OtlRdj3HlaALIJPExpMJdiclwxq3pTL2GTUegfSpB8gi0fR1
KsiRVwcpBRlDBl3JvGKABBFNEIOub4roysPgTc6+j4DhOrw5iIzKH+zY+a7gxg2RM57l+ld8Vr+H
hlqEzgqey326F7FC+5QvfMHqAcSFX2CB/+Rbai4b7pMdVQPKw0CXUcBcUN6PqrWUcW1cZbuMwgBF
m50KYT2hYb4Gw7d6DxPvhTvft3JWZQUUQ8pxz8pd942wCjA0RaOFSic6P5i7RsTDkC0E7ReFdKVi
ftjIXselALc5Qhy3Cf8y2ZhuQLRhMgmucibDWJFFAARgztkkePfKjXQ3yZ6sPuNrCi6v5aG1PWem
SLK1bbQ8awxX48++IGkl4Nw3hgczQCI088uWWuLzCDGMO37TeQni90MbKANMbMwSJB/yQ5KuXqy5
8m+5eCJXfzjvvSUvRgsNNwHjypZIAnLYzJgZyrjCgWz+UNzNaW7t9OJJUOE0JXRtZUi3gZlmwgA9
j/MEK35fnhoKT18kamGqnxQ17wlSjs7x1pok9wDNDl4m7nz1VyEI//kEZ3CuBtrGW/qWno8IEGHU
jK0GfJdltnbg+4BfK5pUwr6fGR+/JqpRKsE1hcdknAxxBnH9ZMEdo8ZAHm6irhNHxj34brU15/aP
4Fm3sHzsHXi2SoX7yfORC57W/Fk2GPghB1cpvqpaDLx5yX00s4amMp+ctNZwIvowD39E9L9RJmVJ
i85U2mHLvUcGvkfVnvzx54H0Yw4iqw30d7KPDm7YtMqNl64FIrscTQfS6+4VZRo0j4abLTPs7/ns
EBS8NiVXxwlS4WhfzKEe+qXqkVT0XfYYOBVDXpgl7W8dboGoXwwcM1jeGL5hNNRl8rQ33pW3X0NT
NTkl1Fdexyot6oJpucL6A20HJdv7auJNJW5Z00YygAKBynnYBklo5OmQSCQrZ2dKpKnHG0dC1Fhj
tRgNGgZjGlBup743I+FyO9eq4Smk/ZldJwt8IVR6YUfx2EXJ7NlRf6WkHRAf+6/o/Y7W/KaTpsoS
AXP4AOAYfuu9kgM68FxZbTIUPlg9wN9CQukhqPWYYXCHBGbd8L8/tg7OAbHjiF6LMNP4wAaV6NYE
uea9rbRCFDA7UU2UmcKAgWTcODNJ9BL5w9NtUq3L7JLeLecZ+7p0MhCM6hhiGp0IxyppXGOgcQmb
9bs6Sse57Ocskvuyk+lQxRRVwd5HYWkRcryhDa5y6ADVl/S6L4hsd4x3CYh6YPk3CkdsLDkN7Sp6
mQTfYWr6hTpR88MTkqS9opvmeLbfOZ/ddY72qxc7lFUNPnZAPmqPGMU+BhvRUQbsjAb4RY1WZQGr
BxlB9uBdo/jlC08dDV14hDjIiiN5ILNZIuMA+RpFqxV/00WkFLTcURZ/4FGkp7DsN6W7PVc5mD/l
ARhXVMsRQyq11Olj0mTpiCh0hbgsWiR5OXDEErLQ4S/xhieG27KkWfCvRkIOzpYMGMry8FTnmixr
ROGeJvYFxabm0Lyxh6HPATnBg9n7IoAuGh+g9eCyLG/q7NN0hRU38QYDvemlav8OK4XMxQvpoBsJ
yB6d6xhYR+JXm/Q4g3h5oGsG+mw7MmPHDpawyQ5YCF2g7vRdHpIhwVqJHprPg18Yzhc2V3bmEcia
htE1RqmQHYQHLJ4bjJT7Noz08an8I1hLdmLk0FqXRQeZlPWz/X45m/QY5NrVW+Apx66ETpUUhF0O
H3VOs5yn5DaF3vXvK49lRQXqPQ/W4QYidAFh3SYYad7bEDVjE1TAEmzMyZUwoIZJGL2Y803686AR
QFpD8cca5TDjvemNWPs0jxD8tP1SEv+gOpurMBpEs/WjIurieFx+uAKlbb/9ZpENEZ94rWF4H/D8
/dyHXQ+oMkbzCzURiKE3PoMH2bgdo6O90CgFjzX6RXRzgcpS6XiFoTNfwNM0o2by+iaOT+UWxvIP
CmuYp4bM3ln+la2tX0T0TtFHUoRfVOGMd7s0C7rrz5OcRqk7ZuKYQTc+JCYp8jotnRbJ66ef25VC
zmxL7Vv7/yM7Xt1lGDB0eqLpijVaFbDxB07ZYZC7efwzR+H4takhPAQJIb0Y4Ei7KuH7RqesHg3Q
N4T44vQrGwz2H8l+FO34vFvy8JJ8NVgki9LLp3XC87jMtMcolvIjvgLn4t2sOBwmzNRA5isbO6rs
C2cOtsdsYWcTs/JB+Q5Fi8TYQQ0uOYiFL+v5Zyyr5hvea+78Zs4/nHuG7KIeJwiZTJMm5bBUt7hG
NWszsFeLdS/0MreC4uhYtHbsRybKAFZXNHpb2JqcPUlUJTGB4kOQdrM64ETr9Inioawy6XsX/TiQ
42OuZRRCOYTeFiuJbYdIqSGe9aweXAcVpLlfZO8D1Yyeh5pPJMD0DNo0SqSUm0fOFJ0s5nYJNmM3
PLTUquPb6YZVnsfmF45QkCgkLR8lncr6SfVMCnBcEjzBXlhe73wyzuzdPa7HqEtuqUOH5OztHsyB
STNlCd9c2dKSDQhSMgDt10rnllehr8mG0HzaS5eAYH6Vov/iumoegRE1/WvROqm2JMwnMZLPbodB
uumVSc7496SRQSoo6Mf41JdvF9sB8QmxFdEVV7gXQTYVpx3a1EFhICvUJUHmo9ypJg/QHDowFlgL
XdjZWKtcLC3Ses3yyHkY2b/Y1UfXrxs+D5UEJW7lUjMvHyqx95Zpwd4Pal1HU2JQqeIABTxT6dIB
i598tuMpqqici39rtmIq7CkDjHaS9w6DLdCsoRPxmzUaNxLgqOvNA80N9hZpF7WOapxq8+JugMdW
HVXv98mFNzZCqeouOQkViQc6I4eB9hqIkNVk9zs+xibWEZCVvq5f6UiebSs4YqIWFZwd4fSaKVhb
Qj56x/WfWW44mMueS4B8Xjfdd6pBgjMvcTGqy7nva7FFgby1dXmbT4+gFfmqCXuTBsLJrRLyOtyq
0R2bCy1XhZQ4bXg13w6K9kYChs/Ttx1lDWf619zlFg7RvVq/mbG3m0FjK/hUebQrvF0MUhD2jjm+
ujTjbF3ANtMjHF97cK1WweVTGzugYHCuApz2U5sp6clAVjt7+acMzvsRAMGahHz4AbnKLGiE9+dR
bztyna5Se5KWxUYJ93X0XZZJqv5sDfLuafpso817v0MdYrJkZSEXsZJO7T9OD4tnYp+yiGd/1oEB
Sq+Wo22qLxDrVXaMuPc8ekdKUmP9yi34L+O+kJFbysnzDItYqXvZb/m6Ul2pJ+W8y8rX2AVL3D1Q
y1Cpq5PeVMYFI18ze3+dSdPsBGxXkt5QMXUworH7/E4P6uqhUT3Ke/GUegLan0UQWs65bhZz7JGB
/sL4aVYwgHAxlQGyyD+nM0aystDd9AVrMv5tahjjC78IsUeKLlnxvYgwRJ4WPtq5S/UDiq1wlyOa
3O0kc+K9WsQFsLvEbasu5QqqemTDIyTfFygChVsjxXGh1f5xmECT79iSjLuSH7ktwjsDqqbCyxC3
qIBX4XgZuXlPCx5UOUICSRBbV4uTigcc1Dw4xnMhRmhyf30g4xEZzqd4qeHwdIUXyOCC3ECHoGKp
kZQbR4gy/KbYsPiVTTvZZAcY6T0RFPH8OYRuab0LKuT7QtuDv1+qhTp+ihArIr43Puscsx6uuveO
P7pTsJ/KGbSKUC69ZJUKjpWP6Nd7aB1VsgTzMd8OQEbr/CzSoqyoZvi3y5b7qn7XOzHZfmFVzzam
LMEfSjw7b0AyMAHaqFQ/PTt5uZbsXRUEJ/OItXdurex+xlWRc8MEvKgnInQal+k++qCdCQf1gAqh
lB/TdVRYJRJs3fSV6WPU+T0MoWXNf2guXIo0Nbfk8GkShqKYuIKkTHvt/WrBkAEKa9xSvlYxz9ZL
XW3wwrX4D8HurS5uFRLVX/aEpomeX6wWGXsKyfOWNkawV49Uy6J8uQfq0zpPphsabXepcoU/n+cX
pPby0mx6FzJ/84EBQMjWCbFrMccAnKD8gqrhv/d+OlqJHE3iznZCWxUhq5QNpw9FsDfkipdkSCG8
XR1UZ75rnRArOIh9RjbgjORV2rZ1QfeMD0g1pT/hDKCXV62QA+62DGQomZGrIiO04zlADaRMSMvl
PZZr3vj2XWvYxmjyk6yJZ0IgbYMa16/3No0naKgnkVcJsE78IrW2YSljg8t6gfRbUlrV70HVd0uM
z8Xk3WE3d+VvWFmC2iP8XGGjMq9XUmPvVul3Olm+59w4l8Tj7yQp9wAFZSux4QonUGQqBNsbOuSZ
3n6583XBgetmp7R9nhZ3R3KapKoPOCeRsXR4N+YcOMVGD/+nqtynnh69YI9hL/BEcvp5EP+iYujx
y4U26ff+LwF39YT4k3E7JTCDx+bRLZ75/JxJkk6nUHfnFErwIfuO7Y718kcbYnjvx4531F9KhWOI
No/OJQ1f/rCg0SWAP5wJx8i6ZZqL/WLjlvtZHQqtHO0URrULZnNp/0KEPfYII6DbjIaQC1/hBvRt
qzMsHqi2aEB3CSujeQahmIS2Fq+NrEpErKdyuvWllvsp+yqXGqBwHp92CemIwxJND7IV1giLRMAt
cezHat9hooWoLAjohhZyLJZRHPFSawX3klp/QkLBfJRgzJtBtQEFgfWpRkKyrKm1KxA7I87ykwLs
V4iyBv8izxqh8qi35mW8yozL328mXDEYVpggOanAkQ8K0N8N7zMKW+h6smU+eGk2iJcSGXLbH5+D
3kKiDzdL8ugGj6T/fI27VEXTGTm2xHj4W+cs5+5OXseaQgAnuUb0FQEtEGguLWW+bXwJHqfgCUvY
3KWwhc4Jb6ccYLvwdTKSExlf7Tsa+xNvg24Cxr5t4Vez7V8epM5DfgnuZjSS8WTvAiiwhkqAOyLw
VG0IJTBBqGcpLppNt32inou1YjYGS0yKFs5e6H1zJktkLTFG1monRhHYxMgBdANZRVfijYhwWmiA
dFeIZR6H7rrYFhk83/ktaSbAmm4zVKFXFlFGU0oIgSf0q/MAs1lCqHDVvuqqIwsXE80PVsRMgeC/
2rahDR208mm4g09BAjgdBakKpz6N0TuHkIDX1qjqAv1imoWC58WOJClF3aFqBMFSvM3trgok7Xxk
dQIy9q7+wAo1HEBG3LnKdBmxaTNaJxJFzKUvoNE0d44LD5ASYcPt/n+QxaDxPLo/i5Ww0WSmS/3Q
74Tbmivfi8Gs0UcHX02d15TrnaaFytMdRLYf18WQBaTm+gptjGmOfIDNbuMzQhRKBPpkVAUBPNnE
XXodYjCyRlfWbzaGWxuE0UXwl9059EvIA7HkEPbKXEZ2wfw+0OP3vHyr9nZVfjE4fksDSvSA5tSa
pKrWsyEDa79ULzErh4Vp/Ub8aUYG+9mOALJyI4Krz+Xroxy3ZXHr+TewwIbMQcs71bpYxTWPho2K
Hm4mtZJyN33PTXh1zHb/CejQn9zAMbeZYTDWT/97kz7oD1g2fkOohsLrBOeq6C6VAhi3otXj02U7
LPbyMAtmQNrZJZAkgDg/ov4hVCKaP20H8echdE5RWjHFOT0KkLMFn0TxxaA4Z6E7Av+A4gccJikq
C5h73Duig5TncMbWgCvZqmuIgKc+vLriycwde4rqJucUrumxW/eqPa3dbnwiFUCpnReEBlwcZ+uo
1/BMpu3HVpH3DOnwsJHqcz4JeEvnjicmoABxb9xOJ1oj8XxOQKQLuyI3ZWd+aj29eq9JNEi6hBxt
QyUYaEtPEHoqUMGoSrcY4Y/CowxVbrIRmdbafxaxGhZStMJ9FK9jLzNMNGQuV0kjflhi29GbPzl8
bge3XmZRE0qQf3oUpD6VqvcKHpA9pwO+GIIHyRPYwp5Ei47QH1aRybRIJVVm53D8MYNhL8R9v9Xp
lDOwwiL0cO5hXRaymH/kbepNrTCesYsopq8fdO5KXy4iH12pk+/MSZ45D0jyAwj3KmKFW74OpIIb
f97whSRXCgwUpranw3aiX+q4W16WectMTQuBUrwC9fTR1jMlxlbDy+7aDz67znDVniESFeAf8vUb
XXlXTT163TQjvwJKIew3zWKilwEja/Qe73A6sKlgGWigfWmuHLnfj7H0WaBzWlV2azZYUFGkKUhS
RfbOplqltE8y3LxpdIU/GgrhPW44LbeIC+SbHWBVfGpF0d6m/77jCXK9XGlfCtiMYNsl3yzgDekf
Mibj01Ap6fUoazG3tkMBOp9RSkusTTPTkmSVHh/5qJ4p0WOy5TgLkAl1YSsFZeLvUSP2EnxgDNMf
+5WEwSkcUf6XY5eTS3Ih3JN7sZ1NOk0G0wmBgOj3YV0o59FKsoI5rdq1Gp67u8T6NLUc0HJ1mW7V
qww/jzb3WWl8+Lqk+qQaCQ6KiwZodSkaaPE2YyHGFysoiBwG2Fg6VQ5V3Y/azbr0uezv8dDn1PMQ
LMYeeNs1lQX7YR5aPXdHVAxa2E/AaDDHxoKrCzzkzoL9UhaJXRfD67CeYxEJHx4DI7QDhXIe6pDh
BOSK5wuifZPgjWdHMDPwla34yH66e8vDIHC3iYHRdlhSfvv9m0xbsYAwzvwwAzaINTAjP1BZUa3y
fYhW2okiaIcbKgEqQf6Pxsd5rCWm+EEGAA/bVlyLeAPhg54vkHhPKBCprwszaku6NluZ7TkjLwa+
onl7SQmbgXuztnfi+ICxL7ZjA4+EzUVcJWLyl7bZ7Pgo88UJ4HZpp9xzVO1/jzzkXNiAtLEghVJM
PZC6OFZZbUkDsXarFtz3/7jkL9JnjIcECqRqT9u1fcGu7/8Qbd63UtQZj9b2ZtauDLlQYWuNL2/a
ma5otAnDknb4BRpoYXIqIRv/Wn+fLsMKZIxuD2OsZILMkoe/xalOim38ZAnDRBF4toX6CknbknR8
SILoWQHRYoENY6ycWRJL+2qIeFS/3fjq3Hc23YL66RCjwVynerEa3/dJhwIInv/qXChhnxfaKYcb
wyvfdS5hpdnXksz9ZqP+sdbpDh5u/5QdkgPsyMMcpB/td8iW0AMMrg4FH47RwDnW2p3ZQd54TwXd
MIFDOjKYNpLAoz+JkNWAlW6M+qv5yCBotl+HnXi1dBHbtjdy3nGpXHhcYhBCxVOnV/T4icZA2P+O
XO7ndn2GuCvnF7KmPZ+hclVc8/UXATeS9cfOKWJfCrqd7V44pstusniNvHXjPwE45XtU9NEVEhHs
5N0tY8g5mgv76H7UW1rfBC6kgEWo098MSbNLETV4D2zsPViBoWMxpCb/XNJ0Q0i5lGJZNVMi0POv
me3Z8iHPr2SiSGbDitW13Wk6gcbzIiWq5+wBP6xGdUNkg3apcRhp/CXnWWd7Lgp0tBfyPPUttYaR
7w2v+dd8LqefW67eenblMc+EwIZjG4EvnsGtJClAVktFgtnKpoooQ8hbU5rLlhNiVKg1y5tjzqr/
pw9jGA+9MPkGN6FvSvhQrJ+lv02iSFQMCsVlsydOypgrXuYZuR5Z1RsJZLfL65OykmQjdxYKp7Yh
gaV8/ofAvjxiyh6Pj97FWWAF+xdFGsgE8pIw0WvY+z20UBv450NvgnSRsGarJ0KMV0FvIbsTvKWe
zvUcrvVVeOd6/IIhXzsDi60ajvtal3v4Jzp+u+IFhAwes3ODTjkC8CtbIeTV+ujj+Qlg3RekF1LO
iLJigd2IUSUos4v3FTiqpYSUrnPMTvW2H+55vwA+qIHiM+HgPiH256C/71mbTfMx4ixx9/bsLXao
JbPAO8QnENLP+BmfW8qL55vlGUlVnZMJR+L8KqeBmaXwjXJObMl+QYzar3VNbW40HEyzk8BfjGAR
BHmI6HM9K9Kd8/J74hdbHL2KRGB8YGUgyg4Z/VipfdNLLHNVSxxaWyXyh6Ebqe3ReQftv6TZt1+9
dsrnu9Vo5f/cdxai9cPbDF/vMm1lgIokZ/7BKXnl2edQ8UBmDq938nf2QwpRcUGK3XaSYK20pmt3
vlKiDVX+paUz1iFg11wGcZiCiN8PlLmGpcT8ekoGF66ratfAgHuCBC1yOcs6wg0EydvnvRS2aUmg
l8lZ4qsy2rbrY7wttcTPrPsRfrJqZkIt6VXaed43PJBhHcl32phkR2w15xscjV8PXhkNc9gzrgYR
Epu6S5E9orRedVWzm9Pf08LR4087gw9bA0MtretU6c9CIYvkpuyCEkgvIUnM3fPCXPaUIySDJs09
R4HKiIga6a2rx1fj52hzKYpegpSf949RyUWOZ6xu5aQPtYr4m0uTPYExe2NdGv9BZV/SwU7B843m
QxJ6T+AKQIjpRinK2udi1tOKv1ra30ys3UJ5YpNryyoD89L/7Y7StIWIUfCOHi5nRfmX+LJRo9vx
ioSyt5EvpzlIvm4tAz5HE5Lhys7h2SJDSQJr7fkIwcdA+sxeskalDnioGWMqxH8COMuhhSpbiUuk
4hhBmzOPLSIN1vL9KmKJ6rXoQxJY4rgw4dgEpeQHkCPGpvMwWaojtgvrJSU9jU4po6+uteWVZkOx
Cd27hcqadv7JgPtM1wjtq4aMuWB0ahOg5WtNpy/OKIKdBja4fC1kKVINkWUV265TrA5Gxc+WINBg
QKF3M0BvsWqvKHc6kqSQCgNbxQkeYE5Zg2Xg+njDASWnmcjOdfa9jZtuNhDNPQ6v87zy4YF4t90A
xuWbb7Zv1AV6OJ56cnnOejVxchmjH/2Bo/v492SZhr2iA1G52yq0IDQPnQz021OUi6tAEJSqwmuG
C24Zx1DBL5sLLs0t+yMR9XIV+toQrQcaiurk4D6PxYRNOfk3h13WqBpaqaV0Ay1WyBUEzubk09Fl
ofUolT3Tg7v/NN9mcdWIj2gcLjIHL6K7AgbaL7lKHBGllPftZj5nesImH83ucBnjLHJBn8idIDt8
32uJ8A44TNqEYUyDIozkMK56dI9qnIl2oFCcomCtya+8w780ESZmjhFKcA+s5rjto6l11Kl+DuaS
wm1YoedKKsFXbAfBAH2EXrujNG4BzkQjeQ2QybWUpTKgy9lPq5BjBKWwFMaOvLEkFVwNgP1NrQ3a
Ez5RzBU6zlOl2VG0i7ij6TeH6ZneN8gxULlze5f4xlNdTtDl/Zxv1EbItF9OTjBplTh3AMqr409U
C6mV44GCq4ax4jjOI40IwzEDkfvX97KTe502jnXTFVplpGpjdttbI0kn2f+Xt0DwF9y3yCkF6sXS
KyykkUIt0y5KYMK70rV2FgwUO3YaVbb/wn8Rd7jUF6nGL8RZ43tBbwb0ktUzccIbFJ6ITh/38ZlX
1nJgOP6eAnYFsYFiSvLIG/ttzSzlQLlJoL9Ec4cwK5/zYM/3vzKLzG4cYif27pCP0PFEU7/o3kBs
XHjIoExIbcOEtLSBSASHOXPKQ/MOZ4JaichUwVz6QOqmm0JCWpGAt5q9NSq7lE5T63CAVIGXE2jS
QOYJw2zelLPUM+5qOQT/SpBDT/r4Ca8KavqAcv93FL6dIIWVFKGXSwxlFK0Oaam4KStIyXWEzUN0
xijwDF8+mUcokfahupeyhKAVngW3hrLa1UdgFpQnRu1oG5dwnBl9v5SoMvX8zRvUnpJDHMvbQt8m
84irhA4oVXBlIKw0aTjsPvkMUJii9W1UMWv/yZBNI2WOkMpg9tCFo5IVgfYAQoVXsKvBYLRHIgKC
2D3vJDpZw8/WSf9DhXZsuLyi3BOrVF1uoa1wl2vvfTip9E/h2xM1rSciMkf+bY03aMVNzWi0PRDz
id3MFKh+0fz+tkk56sUP5IvpFmqcRL5/V0aNlfrAvwncRt+YqSChftIsC5JnYckGVbkxWl97b0LV
IvACvyK2cCK0sNhswQ9DXKY6paF0zYlQbiKd2iQm0Hm/cPd8LY28ZPaeHp0uPwG8zTz0hUQQv/zx
w2hJii7hvsnoEWVMwiVYxf+X1cb0O2Gux7mvSgVbbuRZFZXRqHHaASfkTvoJVGl7Tn8j7IXdwnjQ
uxMg+k4qpsZypb8ZFDSxajyesNtCTZUMfpmPnvZn1YAuLq20f8IpAcDBoEAVpMCw7Xn8g67noYng
9Sg0wUHJfRwSRgS95PwUWGAEWS+i4cawGQsTxMFQ8T3ff9sVPHyiVUMdky3gmFnCSWcWnyG7jicu
a9csm10Pr9QtdvJk4qEbE/fQdyVcrCV80ek92s2f3mClNUrg6WgWooMSnfwTF+wUFxnVlRipMsxS
hlF/Mb1nKM3pXkI6DWU40yewfSyhp4T/s4fWv9NbsIlI3+2ALmXwF9C6NyUVb08qb8iynO45SOr2
KthUBjWfHPpVUAhBjDFAORIEqBdZl3Zlz89mzObkouagTkVFq3CEyyzMX7ESW8q8ZwS01657BDOf
SmUs/qUDBxmyUzpfL4FLqCQDdk33wWLkyockAOAVH8QfQUk7WKCRj536FWdAR1tg53QIvSnvK98v
ru8y0Yx3QjTpjRQl4Z1G1frPftMAyiC3rKZ3ifL84uIdC8IdT3A5k8nahn1WyKiFx8ouAxqpEHgO
G4zGCVu/xnOi2yYKpWVQYfYqLzbrSGxLR5+LaNBc+ykR4Gf/FE+Q/bdsLeLztZAA1hlV5f6yBR77
58Dfv9WCO+T+UK5l7MHMhHAWLzJq8sXhpQr91Xq8DPS1Ay3f//Wi7MRdvGSxEBlSz5uoi/aMsbEp
e5Pv2MK/ryf92fy0iXeXMrzONmrbIfTGJoCFzSGhx+xdpcUKp6TG5bmNGotAx12v3ASj0AnqiCUW
8RcSks018IxEKOJgCeep8glFnmfRNFjB28gPXpVRjv4GLRZRIpq1i733Ai/3aMwSGwcWRk8/lNOd
xggKxau8bK3V45UWQG/HO0luBhbXO0Eq1eph9oQujrCn3t0OCyUqQGzCF+JR3eHUi3mdeXnOgQtK
CigSNKH9on95qvPM2CItd9JaUhfyqVkPdugpPiO22G/0FAdbMUyhRZmtHBCEkGWB6eKUAb23Xo0X
w0McEoDCd5V9orbvXfFeFGlmjArj/RkqKBBKIY1m3qZCsA1E6Cxac+ArbCGEs+21fzXsZn79OdJz
n0tynD7rArJn4aT5s7Rht3jAupL1jBE1THTwj1usqmviiEFJN1Fa1LyhHDyFJa6rs6f3NK5xsung
+F3PReoeVVVIWW+eUz1Ol0OVYX4QB/gTKdwLSkNeHv3bjASRHRbb6AIAk5PBYj0rcUUs2EQmJksy
p3w2/wZD543W2wgN5DxCsExJ9fxLh7wGG8NYvEtzVsTXSwOdyOLXBP8x2YOiFRauz9mUTf35zEZi
sTAFntK7ru9uNpV8AEZmSh/4WZnGLrxO7d6m0VERPrjfoXvVDmYZml3Q2jSeWR6ROrd9uYBSlhT2
4KV31Jnjw8stu6rYEx8W2iS1MWhj0WkTT/22mfh4SQzCkU1k7GodZmy5+gCH+RyDVFIg/WMD+KBg
9Qj/nsCkREyhqk8tTGVZj/NfBbDnVSq/w3Pe8Y1QBRu/uvZD3AC1QwNEb/6Dfqa31MVJ4iI6I7sP
VXU1gquaz67mZVmD0ZZ4x+zlcNnXVH0tp0ls7JH4gbVTx1yLp3kI5GMRkUErgEXG6ZTBVa/cmNdN
cHeu7eGDtmXn90FDsT0zJKDdB+ibL0/NcBhK0Owb9oy/wGOipyMgWKK2jCscf9znVr88aSA8HriM
TcOSKy9KBLzzjh3RsMsjYp2t0cXMxXIbiUSHc2iVae/spHkZSmaryYioOIXQynnw9/yJAEgRUeSH
d1qDf2f8YfcCkhK+UYOaVAN6mIIhh2RUt18rLA7lO1SAyRaPMzA2+ridR/4CEG4oGaXyioM56Ol8
9HDcDtm43HdxMN2aiVI9RqJdA7N614TvifF3YtnRdAvfi7eaeMVXZ6YgWMiRWfLBIjiT43eNF63i
X9IPc0cEHP5QRRUEEslOSGUBZZVKq6sf4RdaUc+KJE1LMA20hPLe2E9gZO7K1nuDIdjsDLyuD6Q0
GdnNYlGVPI7oqnsWYw+/rxsW4qp9uqWZDssBxMBwgPKV91SndJWPBmQimXU/pXiHRk0xB0ympsNJ
W1HT5pkTgfVDc/3bUGbME/5JX3aW5Mli80ebhGTZGMLIwygdRt+L8/LsUWym2RLj1/R1Ygw8sp7p
qMZqi1Lt7g242Ab4b809b5ifzoCzhXmvBsGQC4AfsN799qAI6tJcLuHqw4IBHjw1A1hpiu+4sAUN
Y4iNFEb0kzUXidQCNmodwvmpkbm7YTgqx4+04qjiAeNgFRrdlJimMN3XJ5QrAGm1WUJzHHeO9l40
f5h4Nbv4UZ/K46KpJsQ36WCd5doLobQ8kHg+X+X2Uxd4SArQN6CYaUp0uWtLZKZAKRnQln+E1ho9
YgwLATXvJGBDBcA15OUeTIyDisFdAVINpjU3wWw8xQSYkdQesWd1xN7YifhM3cRW53SwDKOoRI8M
/vqQk1lG0aGqQea1aajHIxv1OXXEUMLrZzPzN4RiET+O25M+Dyw2xm3CbKLyQxr0cPX1YgZuMaAj
wff1FlUpFFkGlWyWmeblITt1YHsPFuEYZAsIx4erVjqdUUBm4xC1OYJyKBq2LOGFBcKuUXLQOE9O
sMsmEA9ynZINq/PT7tpbrAC4ljsmpnxkz8h3YXDwKioZXOJwBsEJIsXZSe7LvYQkRsgUi4Fthyba
4qkMgfgG1IAWVgt/ziTSxJBT31j4kYxVYq1CGAfk19eajEOYShuYb3vN1/9H2kue989k3e9LJ3bB
fScCYjUCHnNGxHGNAZE8anfpX/vidNRzWOdXB80pgFKEXgxYsAWxzuuPimcY1v56xv8hQAQMNrfi
oUMZXu2G722QoKJSxtxwQogsLYx7H/MCe/IWKevJrsXGNLkR9FZvKd+FX/Uyn9sK2XfJFYJyFAE0
p/D31a4GtL6xfS/VKrga71dNwv+kHblhuJ9WS3d68TztnR1Ts+SERsKGvLy/td9/xKodZxI2NlU+
qBkn/PB0o4bnPXyDgo4WmU7lOSY4ey2KaOAbHRyDAdn1OFgpDAKr0TSeXSgTIyjzMwzssrHYaiYU
rIg4u2OUwGyEtrkhR7D6wyuxQTKL903U2sxIRb2PhvLbw4/D6nqEi0J4aQQGNwAqawqPi+FzkjqJ
/dwyn7AOQZI3f5UA/K8mOZGd7U4fXECRW6Y1VHDJqWNrEXQsUGHRByVoIZUCpNlCvvhxsxqUNc8V
1SqOs0xv2Je9/ufzPl0kwNjKze1YJuJOcN+HVNzMreOBHoUE6VEpeF5J5j2ji5+G+ahvdNq1X8ZQ
2hDBBYkrDNcI3f/hvZ42HOtHPz1q3D55NxOLIIPPXXBqOFAkxMTmI3RKJEQEYWT7sYPcUy7+cKsU
x+cl6TYXcCMYf6A8WZG/M5PWkYkhTJMfTbVYpRewO9VNxvqYrsP3X7U6G3x5e8tAVCsxACddyFSg
O3MAYDeBjh6ZrdxvmzBb43B1t29xVQefvvTdQHDt625YdRShehqGdzzfrv54a44N48CRiEJy/w24
KizEPaWfEk68Z9IUwuOhNkZiFx4jN/lSl1MYLKky/28m8cGZDgbQDymfQ1ZiiT0t2k3SFO7932My
7mXxsXriw0ZGOUPVfCQfeLTvyiCiCnpsBtrvrb53pzsz9v7d1g2tqR75YjuWoMhi7EBNVcGqJ3+b
h4DPkgMXfEpihme97pCQ52q7gs40LhpTceyrFKZ8sUx740Or8HkAvnqJJ7Xp3ohqNXuNNT7prvGF
ms8lpUa6zvAwaBzcpIEFQGb9mFGAS/fWLOMMPn/Do1sNcRpeqIILHxyfL2edm3T/9r8Cb1VpA3TE
qr4zV3wG5PjKoch4f0Ye3t4EP8UElo7Jbx7YMRDygZ0uLNb0X4cp9EsJRxuIwyPyZ0b9GjVFvtqg
o50ByjdZcrddeVZfv8d1aIJLA8sEyEPCokLWQOi3U7jRQYeH9dSA5rfn2LLj0udAk1FafKY0t39u
NTwF74Pnbq37Y20j3deW8JubgDQ4HaSo5+9FyPdu2UXTQkZlOStX+yUa/mwWq1euQLP6hvDjMSmt
Ohac0LZlm0McxpMO3y4/8eRc+vlLx3kjlk4R6dODNwSopUZEi1NO/3h2lg0+XT3Y+XaZdywYLY37
m9AoZeMJ6TU80MQm+QPzhcnCFvZP3lbubG3fjMI6SF5diVqPnHtO6nqQDoBEDSXDSAs6ZeP4vwR0
lvbEWzq21bnD9uf7NWSyFRS05V63DPbpFBE5JA2adkzzHsYSlSxLAKghsu0UeLCbztqyqhH+0SF3
NU8QktS1yTwEeqsd8++CypnLYT/pdwjdHIgWYe1870/nHy9qw748CxUg/K6Sn+0/1iG9SIuDCZFH
3dm1xxXr1UHn8Z1rHv4fbR2OYC/gfTaw6Ia6h/FhWDMeiwq+W3yTqHqLPfoRewGRc29x1fa73wgF
b3XAFhy6fnFgmGD/twqa09NkHIphor+bohhzHnk0wis88vWREHOtaU8sN0fD4C+C4H/AJoI6OWY3
H+jSGVUdHRVeAq7+9uQSEDMxG/aRwje0I04tB/iBLxLWoB6hP02kFLCTsLKOACJVNJ+P2rg1uxNh
WjBt+jJ9bbUWFHx+aIMKwSJNw/ycXEJrfYpYPnyBBOZCVePF8/XqkpkGf89DU8ssljjEYP52i4rc
cBa6dQkezezw+jNm/lLd2uiKUBajgOuE0Or6o2MUxLbAqruYYsLp/44YB4ESrJ2Jcj7NUHUChits
dL2P+5xp3zYtmwWMharwmtkgYcvp9EiwIXIr5s9PRziVUslMILnbG+iS1b7sKJzU+L/Hpv4IzXJe
j+KbchTbESUKr7iABVkcZwk2PFEmz3/+kDEwqRofMZn9IpvpmS8yCRw7KtGCaHnDUxNEnSbdffy0
ygjO2ozxXxsMyi2LuEBfPfwMhYlBX9CA67Z8i8I4tYGY8fxxP5vUZxJ34PfBJcZFHJD+7ueDfhho
KQCnVsdCPJDbGMyZqU8WHvfkUV/F6SyWLFYkkggcSSiH5lXfn7uFERIAEVN86fbd/nQONgAzwA0W
Y66EMYWRAFzHbHeIs5lgX7nqIBHDk7A4Zb6vrtAa+FuO6p+L6YPwmVpZwQrFqJz09Glm98uMbBcL
Z92I2Y5mdZ9pMro2BuI/phk56dYHNMR/ygipTHgvOpnUDI5HSmaCYN8Eh+eS0JBfelfSur0C6b6u
A+r7wR43e9e/WPidTAfS8uROC9kqOVZkf8pyYF4Xx/8IUslpN+yr0Pr7UX3mDPNUEQ5xQb6NN/FQ
2W3FVyLMIRYQaM2ekXODIefEIK4KC07VJjcO/4S4udXImRf1h0XMDaLBW40sfnPjpU9jjUaMTZfV
pulfJ2FW471IYWpm/53gSet0J+Wl0EgnkuggI+r5Lue6h1A9xeJsxevv+niW8oAQpAw22vaNOP9g
Sn3a95gdXcJFBoxquZ+quFFwiHcUXLKAOUaFv0rsMTAJu31dga8FJtXEXcK/mkizLAX7hZQIMebz
SoGs7HyDNcQsRfGrDoggpMZAD0pG4EbXF3bn5YjDfBR0d9Ai1uxN2BZvgoTC61vfkqUYEVWxueZV
kfnKk9sWqOq1JOfobrv6W8ctD/ZHhLma+Pdulch1/b5uAcAc0AR+K3rdChBKrp1u3xsyM9d6Juab
U7xvd93nI3eZBOzoo2gKByoVi535FXkzoJRB4AQUPhpZdK0B/hsKVe/dZLQ3rz8u7zEpDmLi1yDM
hkqgFMpHHI5tOkEa1JDq4DJIiVj+Z5kvo9TKFA58IR2rETsE3QAu+W6Qdb1hAE9CLXZZ1NmaQH4m
wzTlcf8nOneAkB6wFPVzQUli/uQB/WCRQN//tZQbn7vEgqU2uXP7eMTxQYiLI6k8iC2w5PFWAcMx
MIuHp3u+xt6o4EOI/lw8KJwn+OgINYc9HUqQtzf3SjpDwnkjm7z741gdnCPVWECKWdZtGxXw95vy
bFDttY9R2ewEY0Z2OlMJYKWN43sG9AZcs4n+PIMYhABNxiCeZdDwblDEeW/xyGov2IyRXAIUSynQ
5H4BjI82FTemRcKikQ9tyZ8XMGNjkZYbg+vqd++kK11k7zG1NjacvpcWh68hBsgz2IwEvBND+KN3
cxjEX/1a5ENmqLGXqv6u2NAlOFm21TIDBnVy86sQHVcEtVHoMoxZtytfkyurZt2uY+9MUZi7LLmo
PFwQs5VIBYctGkPXSS9AlggvnaREE4UgAGP3qbIo3rhXxPsI4u6s2Jm6Kt5AdA2pzANf4Aec6LiY
logS+fr3/sVWZdaRXjFBcd+zO0H+JlNipOcIfjWXPx/SfcMUnAQdJDdMeiPYpae70NR9pt3GLX66
/G8abFZN/4DTrgvuXJr10cm32IoSFGoqwbtWcZCqUo+TZ87WuH6wdcFdUGtkLFz0nDKPBUFo/Ocf
g0pz6LMVKYRwMl2q2xJh+JJfZrIaRswbqhBDT02Q3CykzTgklfcaGMPpj6dWD62QOf/V0pQyINyN
MRrpeOUe1ICUKnkNoHuOSezBfSHR/F6NEkk6K2xxz6uXDzDBLrDZ5AgjNN1Xs6eiWrrF1m/WkUJ0
06ae/7uHTSg+5NlMYtk9Fs/Xf8Y6Ni88skP44e+D6Fy81Ck+f9QWCNYkEO9kU6RyUv5Rccls016a
HTutcKWNa7Ok5PiWVfb+TvrWTfQNo/VYtyHeZoBghUStqVOgJ/qY/00MDNSaknfSclP4yG2sAp23
I0utgfPnG10o3u4RGTzzfROntAyWluq7vTVDUteg7Rsy3loKnX4336xazQncq3D5J8LrPomTkl7s
vONfdCLPzB0KEAdepE8ILMcJXkINFrhBdC+pgXGpQ3RMl/ge0aFCtkVAW1exEIaCssBzoCECPgkQ
uvi+SdHKG2MqU6GjUF3tF0/9lNPdm/EMfPcJkPqE4j1R9XtjsMAgVg0UgPRegjhqt4fkud+a3pV3
a2iJzLJEHAVLvtfniOtUkOYPeDifVi1sMzOgwURJT5GSIK5UHpIhmnCb019sPky2qWaJ0m7680V5
K0ma7606DY7epciLXlXXiaa/QXpmb63OgZKlPe9w81Nc6QjndKWSjZdM2y0HOvyWNe6NZnGHxS4c
k1Rwn1RGXTbRfZozNm9i7vM0n62Kl5FBQpBi6SOdR6k2OkoDbjAsrF0F5FnZTCx4Xzut7kCdxYou
r7vSrDPTMnCnqD5u9Xmgvhvw3GpQR+xBMA7pFJow+juFUEUErgehkpb5HA9n8rxW48AGXibdKsNS
kQpQtLtCT+Jy1DDvwStMvwDQs3jnwxClL0f3fXPO2mHlqoD3tW+UPN4siP9cl2L0gRwmzjdVvSV1
wC1pTmCOTRfQTpE8FR9k3017NylvwuzeAIXOYBGp5Gl7Oh0dOpWP6cqA/AhxbnI8Mb6DoX8bQwcF
7Zm2WHYawCPgoyTcUPvuJwhx4V8FtDPX6ygnII18Ws1emnvyGHf+EaDZSwKUWKd3MaFAFC2W0E+W
0XYwM8wf29P1wkdQEqAaCusNYU1RULMl3omObzeCwoLr9Q2gn0bmZNQe96D6Oc0ZY9Q0zEwMxvo2
JdmtQA5dp2sH4goVfI5WH5ahYSWud96q60b6Ag8wK4LXOvaLJsGCb0azDK1kDIIfySgPRem7yp5l
Yxk0H+7vLwLHbXNuh/e6EjxoGWCkRwB7FeqZXRC1B1liIZbl3pxyTaeSkruI8hbKGXD84LTvKbj6
PUb2DWS1wvt6lbrI+VBX0t0rgqWN7Bym84kYPUaRK5iqggkYZRQKQRh4EwA8BM4b//3dN5hi+gcp
Hk5ckQffenaPQfKhPZ8wpElwHdIaJWgyudQpf7eGz/y4pgr76Z4pncSgEohfhlcypkMpQRLrhDDE
3+GCcRUn7gcyTBUK9zzsKMcFwsV3ZggkhU7c8BzKs4YtS4irFsL4Z+7Ux1372+JkNvTGw5jEEBag
+TskFa/X8zUFEhGyPx8pcddi9+OKfEEIfOdvqmNF4uhJPf+7XH0YVeZxwPK4EGq6fPEm7XnulBKg
XmFp/HL9XapGy6t26VcStTZOIuYTrM5U7zuBWMU9THwOp+NQK3NGAZ+d+ln1LUpBBVKxicgiq2DJ
4Z1dOBlHJ5MinRFX9YgANf0o4czm+3PMsjgXrpnleg8mKB982//JoMh3ykeIKpPvxBIVxYRjA8PT
1LiCbG1nsdi0fDmGTfnwpeiK/FO4wHCZ6bnwCQc8DsvGpfjeNBfg7dWR8z6GrorVOfGHVZJdzkki
m//sokzJFbd5Jyv6p1Y43IzxqoX9jA0E9ulMnCc4dTiimnRlhSncHRCicmkodbHA5xYnVN2FgkyQ
SMO5e1menn4ZiUrXmJjiaA/DwOrs6yYgunxr5tWfkq1ljn1gCMfTXAv/9c8rA3zMmCfH6M1E9Sn8
t51ifRlnoRddk+dR+WZhHwNP7a0pqgE7RL9+pWKke+I8YSHWoZFA2e9hiP9OxQVcVZl/bfLzBOle
Si305KoX5eunsFUE7wqrlgzPI8FIhrYN9ocC9xCvSfrOCnOIdEJJLZO+eC2RhYoO9QDzThEHkmdO
go5lnuaGsKmKRRcP4kE/D3xPipKCO0I2SEjkyaauKJ7zg5fxexysIQ+c2B6Wc/s+pBYeoAySTDbf
pV3jjBJ1AbSZ6eft7GwkJMDAS8B6GZDR5HbL9I86+fh8UGj3nit0zRoSo4qvSOs6hKyjik+b5ord
wX4qBpOqdPEoeuk13Ev2Lj5nE7NTMaxxWhd47LVoUlY8TkiHar6uLW0oQ6+V9ndYplfYt/idov4h
TWMZ6KeLE5S41JKCjdvFNoM7nk8PbGctl/yvaaZV9qed53B+kYySZI0Xm0EJ/D7I5ARDRdB1hFei
uo0fKjWHCb/8D2mX5uhuA/yzoi4qXWgAn3dJYiDF6PQa/CsO8y4MBXT4Ndrk9Plj8sMpOqYm+eKX
NLdlkcRceZIRpYIleNfFchK1EWrljnnLUcBlgYa1pSPVITm/VxF8yXyvrARxaP2mZI2mI8jRbN2W
zUY0IwwOAKfPM8zjpPJXijMXRmvm2J+64E3dFSdRielXuthpuLY3gIMXH21vM5EKRHQ4v3sv0bOC
VD9iNp0QHJy37HHMrKxUbAKc6+OXb+di1zAp9YctRSGOchhp3Bc6hXKCA1FfheZMYcQK8Of79GBn
jC4+FU8z6gfuv5SSNsmD3p1w/HuN1ROL6haMpXF4mEm6JrH+y4abCSUei8aazKIUHqPeHuShH7FI
Fa2AP6NvvoQNeqD8g07wc0o27wD6eImT9IUiujfvMGmqiBoYcQgVukZlM1ctyH1xShQMCi7KoIYx
WQnkNRMnDtDJScjhygZYHB9zlWFXoRxmFmZJBHlsLGkUmUTw98NoKPNV/mV/7bjn9c4yPUqWuljB
yqsySK+F2RtRBYKueKuOhIIqPvncFqMlKcGlVZnCES3VFPM2nFDLChE5ZSMepJEwB7W4xbGtW8F1
thlFd0p/IeVFO239HKq7tr+5VOeuO3WG9o+o6BxyPJ8OC+5aQ/I7AQrzv4nvVrNk5QgSucTvrQE0
n5tSWloeLMfIOhTt9EvvKjzreHgwbNUGei8K4tdXEHrkTL7mZvSFt12GdbWHsXYztOux0wxcXOtF
61vOXoggWD53JOFiEieJkk0KEOj933QhoKx1UU/7Ke4oiUCOCMS34xSFz9WobWyc4y+dyuo7feHx
4abt+/FLfpuqQfF1VdbV1Mnw+VbAjmLAcxI02JFYD4UA8KzCHSxJtQLALnxzhtC/qbmBVbOqDWiE
U1Zx2YtY4IrWoJQFBCjXBIf5jw2YC/yRTiLQsDvxEw0p5IyXqKWSBzBuUlT98FqkJ1FVSmQ8MwtC
Nwqn+E/2Jg3NJq/mIzBahGYjdjYlz0xrmtGvzi7mnAyzRJ7zFPblYrmzH1qFJPDA3QFs6YcJZ6LM
HJUQBisDnt1VtKF/5jPPUR7DKEwZJY/4Z9E+PK5SZ2NfHYrDF+2NFgsun6lzl4W6dAfl8KwkJyAW
d1LCfI3GplbengC0D4EHsKcraCFTW4OsayxrXrGCRnQV45B5+Pww05kCRGfoUN2N0KAfPuPRFpmM
abAYBpyuIMR3/SRQyF0FdIYSVLKpwh4bd5OpG2w6668mX29GjEs3IDIfRznhJ746lA2SP9zEoSq0
5oIHd/o4U2BgHSzjIcPDGf3rDJ2ROfHASXqfW+S7yYyx3iFcb9TkBbQ20N0HJiaWc2GjeLhU96mi
ZKpkMb4beDpGsmauwyqJgHbtqE/c6zjQkqnKX1ISYx/FF5yW+NI+uYrefNrxdMuVKUXS7qNQ4Jjo
fUHapaGEPZWLq3BvbogfO4oD357Xbo3Cut9GMziakYKXvcaysnL/tVGjwNy0S+rlIOCMLW8zQrkc
QSGhiZySs0nhwlahtQuq4cQ7ik2eXUeNPT34YAjcMZ8OxA0FNwcsT5fCaNTAE6STqw8Z7SeyT62d
afX+llzKExVUdHfFLfMLPg6Ht4X88izYLrFY0W86ze3TZwH2DUG9qoKr0PjvUFaVRgkHhhg5h+v7
2NvAHV5/DRo8YLzjaUhTpSfozUalKYaKTTeoPo7FTRT9t9Kyr7+JBzJ8xwTPYZRG+eEXzNwoHpcT
C3X+4vGSPT5Imi0aPyW+Q0sET4AvUQlQqsplmA2d2S00Cex/TuBRN3AS1CDhC48Jz06+GMoWc8SG
9WCvG19QvnVPOJDJb7daHmLKlZ6y1GHGd8ThKDpIQ10pxBZpOcn04dj16z1hcR54cvZ6G2DIZ7O5
FvB2BeRvhWNZwvldiFOkFkiVjQJkZ2P/jP+In84+MEhW2w/Yv3T+rWrL9JXrmTa5rP+P9l6AMR22
JKwvbbSrQeAt8CWZmsZPX4XdJl4b/IPxlQpw3d+X1XDJGjvDGBz4LG0gsNn0EJIxhmNuMCvlYr8r
jIIvTgZ4+g2YnOGX/dgMDDua4rIel9I3LAUniDhsFdDqM1F7d7W9wuXoJu4c4VQAErwYqPUQ765b
146MjoHd8JsS+/opTDiKvpZJq8rnKcEPJSfKbw+WKbMOLoKrvBBc6yQ5vKO1uHeRCcQwVBCJen4N
jPaA497OGgjWfSYo8suOis+hQXhiASQtAF/A7YlViI6deIyZgldw2j7Q0lX3dtUUMOkS62PuXZak
0fZCX0kOrNynghMmBRw0B8jdrOJBO0VpW4Sz2I6NpSoWuM63pqZvXNYhZ5s5xDuKyq4b1bcg6HBt
qMFAZlXvFZY7CB7uz6SDKx/r9g1cnDAs2dldUqV1lpUW0SkU4i8Kg3NlPR5+W4+yNYN63mhnC6Gw
NIEiBkCSVO3UK2rqy+OuhQD3cLth/CIYDV865aXPKymVl6DGhfhO/HLop2TnKntpyi1BP8RNfjwW
0AWAemwv2lSEKkycacymoHNprhTCeZfNRBMetCSCyAMB41g/2mlS/M8lKNcuc01hJn65Zlt2ZSb2
57yspoPRCcrvuR6k4ek52fPLyibLKWu0KBJ8KImI4MYN/PWO6vB4fDGlIfAZSvKZoK4TI8QGW9AR
FAOV3UzvMq7oOPspfVG+EB1Ie0goJ9zPWofvHS6iBSk0GW4TuvCDaEVAJICp5296jGpRZkTzUqk6
Nrxdg8VTdhxud/GlstVLy4PcLJh1iiFwwj09loYq6PHtRHAaLWTTZ6btokC9Tp8ucILjTa23ndtm
kjqwZv8XyW23fpX+PRDU0G9hM2STYeNezOqHvf2o5LCliRTuggumqC2hGSioD1Cpa5t7yR+uzpF5
rbP1pXNnSA/BoAQXq47Aep1q0hYGe6HzHPLABLqGZbGgXkVjG8zonJoZXDQckEnUmcmgWBI/XY67
hgPWZzJ1RDr8T9oEAvxGbFSw9jO5crcGEOk7IIfh0eKXHwQnPFXVRN3X2Si+WF4Q38yfbzJUgGke
+c9fgj70eRsmNZaYKEoKNVTIdB/lOetZf/W2J6q7F3IdUbG0IypppwUkkL+DcOAC/ffuz0VAU8CY
9BS/V4YJcdlv7biBLnkztijkNbT3SJiQfLcI+rYQPJg5oqVRVoCrCrrpkmrtOkkzT9DUbMwuXCWh
hzszaNRxLFbnpLiNwCr/JXUmTRSs4NS9+2FELQsol0upy1iG7Bb92jdsSCFGDzrV5j3zJo89pBLo
Un/1G324ad3KAqGCtYVMH2o2RkiCBwjK7ZJVDWExLny6nDi1KBDo6TllB9HiotW7bq1svLZGjAus
rAi2lQGXwsBWHdMDzRbilKBo8yiopXJduPJIvJot5Dr5DhjJyiqx9S3HkWVFPRrpL+7+U/QrUhs0
s3rLibPlIr6jiZxXicQGTuJE1dpbzaog9LrjE/U1hJTDT0SPD+v/CiDZnq7h47Ln8tC0dp3yxQHT
5AEcINChahrueuXIbFAZZ3oiaTrnUnz4+TMZBTwYfiH341OZOmG1bpCaOV9rURx21jXEBFFnbZaq
KuwuYfUeXf4BymSWNYoZOMevVdSDhuQqfTOkOvx7e5NU6mXkBe5u1DB9KGDLj+z6YVQQ9k3U1oVd
RmqhcnN0MdW+rTG8FCkUuiYoWeRq5xr1ijyj0s9u0QCxUbSZD9meDofgb1XHQJcVj0bw9huWdM7T
J/nF0xC+f51X+WBCdfURgGAyShkcrYlw/+sgzXjatvqET208KRueb1SFZy6PUhzcqDJ8xIghXAMj
YViodnttYhnK6YEr1pP++ITWNrS2taD+0u1RMPZxKFjvuBwf/s9OFv/r8PMSypdkoOOoGfm2Pm8u
8r6PuxFLG9DCGPS55gC+OmhAxvY1DK5zl9qHEmIpcjr0YmFXIOLH/eexHHUyF4caifEnpvWtwPlr
QZOUaOvRRSzRyTDaoEsCpZQ6VIxAyjDMNdyLt7ZjJzfHZDBsgY6uu6cafZVx6eYNcoIxudHMYy9j
DUGqPqdVNLbjXrbBkW8U+L/DoDpXCHHErp9qGNhkZQGnO+N6MtgIX8NomtnAAHZO1PXu54Z+dEKZ
jo5Ze02N28QgUA4MshEZaRzViL4KC9a+kj+wMoIRbFI7DnfRgo2DLsznmTTmcl0y76FRsDpe1lvO
0tsSeDiwJX02ObEphGjDzWvzoHPXcqWvjZNrcm8+6Qqk/0c0MMQc4zwcvgpSP9rpneruyOQeopWO
3tBNaquqXSZ0CwP3Cs+z/2UGmT7RFNnwPZvS89XN9xklaJuku74Ys7qIHQEv9QmlNKzbjJJD55RG
ZtRXsM53Y4NX+OdFiFMZVUpJ7aG84qU3q/tF4Nz+EpmEoI5b+Ktxz9LLDrLfVQeuS1YOIinyWg9O
9pXYxmWBRROTBsbfgleSaNRvqk8F/lUg6+vs3FnhDqkVpHOke9FdANfX2FIxyXuYrrqRU9w+WAy5
XuOf/1OPYHO2RD4g7jXiIqVSQhHy1sGBGvKsy1m1aCZg/HIpUSGRjrLL/tIi1NMtVwwPFYs6OSZo
zVSlfL/BhcCUCMe/k4ZNFUZeNxfYShs/AqTXZxf2OUqm+fJk89utLWqs/7AWedDEY1Gf724VQZ63
wrnGXAksUYSFz3Z9vougWQN2STdPWkTjeCvDjiNhhkd4rHu5vUJTcWEEULTUnrMGfycxv/Igr6KP
9WQycDfuyoQBfn9VqYU9c1f+Nlr3Dh2kRO5IdowEKe7zzBS1uOWbzBTBiKCJ8le8jbKf/fVKdFFm
mgLcPeKFT15xoQtnFem4dTAXaQYjMSNbYRPCFpCx+igSH7deSYKbbc4oAJgOerntLbFejmhnR030
wQutW7PzabiPyakKR7nREXPLx1I5s2+z3pwT2ORZfoECg0dQa3FU8h6b3IFmCWwgaSBmMwGLbTFy
N3QnKyGdscSPwKQjJ4OM95CRaM2+MiiWcNd+vt+XINO6raYFUk3XVi+h8ADbQSfuVyzhByE/tVVJ
5N/gERAUyvOhXPOlSFLTzv0jj+RfD5BAq1JyFXibSMsbMAnG537cUJfzYUMLmBOSTPgsq8kz0yJf
UqwkQOWn22At2j0IIomwV+GPNftiF06uKfDrnfasxVFx7LuU9zUoyegIKLebGiUqUBfRKRwqAFmR
0v/Ilh5bPdE2GB3gCK4gLYQJ1KQPCh4B4xdhDsjmuLXImh6111YDkuyNYXEw6IKkOznK+Rc8XJEu
MHpiuB2K/lJcmZM/0aOCAO+lRmIdtgUkwc89ImpeG38l6+4durD4HK0y6c63VooCjIgP733VwKt1
/Ssb/OOV+OwAX7xuI34ZudQdRWUsW2XI7aXq5RZ68G/pNrqgmnCVcQr+e4pKLPGNl5yU4YqjRjKU
0bYQY51JzQRCWWukmHh34xEIa9SO5+JMSXJuU9XcVi/FpScaTcG53Hmihbana0ZSB7uk37XOUhDS
8KdVPj1IxVOSknkN6U2R+A2JabSoL2rWM2RpRe3JjQQjMjemeb4RZjq9CuwnIKrRaZus8YQGE4Uu
Sr82bxkJiCWQN775W72eK9AY7WB2FwHtMPWevtlP4+gKI0eEWUTc3EMX0Nfoj6pj2wiWv4gQG0cb
PjnSr5jBtWN0rxkaj9zcvgj0cE0LJhGzWN+XhLSSeN9kd3Fh9dzB5i8qT0Wt2X/7gtDIYqCN3L14
QnejyDH8vQMYunOwSHxISl/pQz88EcH/7xQzGgH8ZZkM54w9XSEfbM8OFScpNDoezUVgFJ+oOLCM
CcELl3+M60xTxWy+qAPAobDrKhPFLOY7uYzqsnFp79XLiZ5RmrGKqnEY8IF89KF27SmtSpfXLyEq
g6WgnCtKMWDx/bEfxj07EeXn9+rW9KgKtbEK7FWch0qichVzFtvMzTvFHZ+Y6xHa/qoMzBRve3Fq
wv2HRdR79j9QqcoLCMWKEVwaJYnHpyw5hR0LxcEB0ZMmAYJ6DIAa35nV8UriJqBtPFZNGqOe4Jxd
sliJcvcMlvV92a+iyConq8rxHMZTItgqmRBSoY5aBnLb10+cTDGYVlEHvUv101s8B7lwqu23Bc0G
hA8RWMX+7bMTxOl+ivcJWqz4eNcD3RJAQh2AQqw/9PdBEBZGSQGgS3YDLUQZ/T+NRLpR27teSMWP
j7hS3FK7DO/u/Qgcmm5maLYOMJhLlUU71YQZOVbGQvDPR2yUaUF/9c6e2gg1tau+7I7rrxTJVJ8f
0h29Gn/1MwQnoup6SBdSJG577h5m6RWmJ2dHrMlooBBdN9eJTntLjyItFAe6rNtgJli4B/RxBDgh
49SjOrg7EMssmRvamvhqgynfY6tmgKqrHXQRPmfKJglqEDMjlz7zZofR8HAPPZnxROlcxVJ6L6PO
e2j/pUkT8cAIM4hFayIoxL4yMNXhhcMQmO3SCrd06KCyy8uy2hVXCdL2kMjalNscs4UIg2Vd5PVb
CRzVWbRRcOmxuJKSYHgY+U/hau/nS76c8K4PFpbItFEGdZEjhZRM+hM1qlRIwqZGPeGpM0QGTnaq
oyUOxeZPfZ+acLtaJ6O/EOebtdcvVHoKX7T6mpMo9H5gEh1gHHg1xtsA4AZk4NUQ62D1bQu4dBhz
09UniG0U67vBHe2p+fFoF+fqnJJnhER/loZqKcoo9SPmPh7KzEirh8Oyc7RUggt+3ZR5iow3Y+Hp
J8Pb6R8Gtl+Auh5+rwxc7wBu/iog3V9osCVc/yzP56Yr97MNzpkVU9Frl8hxRUWRUgZaSCvpIu4n
sPX4FFXvWNGq1opmaNnsBQS5G/Eo4X8c0MXP20eHIksllS3+hw29/2tZ14hXBz8cG3Ln0HXjEFXv
zxjoYYt6EVBninDDlUg97Oz9M/jacpJ9l/vhEWBs9o1UmGbir0CLspfUwIiGSzjbpotGNBz4gM+v
owogsn62+TlwP9GHpragm7VgbNYleKOwaedM4BNGoHYbaYkVVBvpNyx1Pk5UnumOzVfsYsHLgWJN
7tkkXwDeH5/Me5s2f2WzCXPpfQweYF4M5mKfnmU2nBoV+7yu3EE3npjGUmd1VzpwH0gX4/r7SOmO
0VktUu8yPT0aF3XbUgxsEOe9QlO7WeckiiFy0W+BDk0ZY7g2JfQXO+pwvIRl04TTwIEgL0x2j8gt
0+oJT7mWeizcizSDgbEOeBh4v0z91mdjlcfJ9Xe3nGwnOlZDczfooZQ7UnKuIQh57IXv/2qd3q3w
I6iFH9ahP1yqgGr4E3o9GNKh0FgV5uLIp4FeoU17juYZi+3VZzk0bexz9Yq1Gsn7Ppe0BC1z1bXC
iaG0woUL/5JJvQDieABLS7lsyeZ6wRvKWA45toPk2AS+TCS50/yWjiooSvRmcX1xzd0kt7yzw2xi
v/Z8EVsS4GNH2HjuJdyhBNcq1MrMtIVcDS9+4eIahxavchhHVFWZ2usk0IS5rs/Y+lBAqQBxp7Fl
n9W+/D0orkHO7t/OJfRj/Ht9Vl7+bmRgjDYRzcoW8UD1YK0P3Q2Ncfj5NiUe5ZavazHJcdLXueKk
fYGKeQ25g9gkaAtyOMRcOs+cXX2OXQW3kyCBVS2vTEe7ijCEEl0uijoL1zJNkxKsZgUUPdBMxsLP
MA8V8aIXBqTi1vFnf8ttsx4HFNQqtIIQltOJJNz7FbvePDdQCtYIUbr9jqoWcWx9WW2hqfT1En3b
Ujf1wqpxdvkzuBHxLuJwA2cGGLaM7LM1Cs7oM53LUn2v2+xs7lXGvqBTsO7MNmCm8U3uDaqB57uY
d0aNOqguNs+FbE8TmU3DjEPYhW2qe1UChxvHHW60Nh0UNMiMxerOV6E5dcSaCTBJT+keefBmT7xf
80UCkSje81du5BqSf+xowhBurmmO0s2jyA9jxle+6wUhYmyFtuST+idJeKPRzBknxpNG8aizHcJb
dkf5cdTDit4H1jpbWZPtreGsdu6R4krUIJyeJSTd8ASa60QsqVoPLvkRmXsRFRQ0BJnOwXumnMKB
WIn6oSd6LBOaO4PRtglfYJJ24YBAbvnoSaDn5r7v9nfPtG+bcPNIJnpuK+3fqnCfDNa3nXnc3xzS
HIRhbqIwsJIWAuR6T4nXg9bdIfMXiMmkNMXfGskkvX84V563UR2zHEjAFxDB7Z81yMRKNiZ40ivD
vRInhLO4e3R65iZfeEuiSbdgFpt+39LcPnIFumsokEV4EEQh8MFVmfp03kl+jVdTHo2dCeSxgMNU
HqHUGM765vfu3FiHJqqutPQB1BLK+JDHjbqThhU559rztQSE4dNQzoECR6Iy4IobkZHUvDslTpet
kPQ3fr3Zjawr04BUSqWXcESsX1jMcnRXFrilgFASLmGCP2Cm6mSOOEe6oWaSoqaHVusY0y/TRbBr
S9sMvUuD13y9Y0byzhWqiUOUex0ZyqQBMkiH6iTQf5l5iBoZ0rW6F/1eM3zArMVYhKsx8rPEZMDI
p7QzA+MaYW5kT5iTsZEQyuw57A1AUfLMTjGp98vduy5oK1NYfpqNFPuwHwsrnRoYY1089Aiym5sa
PYXb9c7sFbSabitHIKjXy+Wq8P1kpaACOPCoLh9Uaet01mTOr7q/4qMgOBJATmUjcPdOfutg096H
lHdCX8i74KLY35ZKzft3a4f+OSRN2s7lYGohNlnPzYQUb/+lARnV6wNldYULZPlXzhY+/ASlHVIb
M53J88B8jirvHAxFWL2go3k7/CM0u1Et7KZLNc5O5y91gnPFJo6MCYuPr0jHelrxOkojBoodoRVz
P80XYD+CXH7S14IJkVkOha8fOcF7tpxZ1wh7jVBH3i9fE/gBVJxipm9GDg9wkVKvhFT6B2pGIKia
HhqkjZyOhuuTmclwUaZDBm+QZl1Bq50l9L0Beh2KX4KbBiNh62e0cTwQDB+3iB5yS2qdF8nXdge0
fOojP+YMMmc0of5OyUbhhYEwHDW9vRS/4A5gUWnXocG9Si5R1ENbZes9YWPPO3js1lk3H4aA2FHi
jPqM/e/btrlsK1qMXK9EBDO4BtlfWQXR+ygXtwI8upbcPzXBQ1Rdqk0r3XnMhTo3VOS2BozcHaD2
0EBxf0EmOaFq17IBAgVBLZnF8qki3kEvrpqIACDHD3IW12gWE6gtS+I4xOOGwvRiAr4Iz0losQCQ
qvSCQDCljLUZc8eShWLOKUzXYiRFlN4+U8+ruwCoXrrI7en1JIdwOeYNpRGl0Dp/hqpU5POdWFFp
oTvh7pQ2rOVZ9Vz+2YCQpavIRhjwgJjKRAf7GZa89AWZ0QfjNPQf4Y+ISetTL3xkuck6g6FS8bqO
pfn2H3xDvP31txBuZnrTKuU4U+LaaNrCjowjLNDPcwX1YJ+SX63Jt0l8r+obVL11wZHtTmXdrSz4
IA4AaV5PUlQHdFyI23m2D2IhJL/F2QJw5ZUMHdJ7rCymVjZJ3Ro7LxAEAedYGAdDfeARxmhNOuag
+n4MLLoFLGWSTA0BVM/IvxLYgqG/YRKWHK4zkYkssp/8ujjzHU3CZIqSPhO4PA1t6xQ+xA3Uo+mJ
KEP09gyva/GgcoOtDki+sqjtPHiYPqLFgLCwXzT41N/PATHAoxLtVC065dDXv8E/T0jgUmDheGxK
JFW3lJL1Xz4AxPx4DXo9dQ8KRxwIUl91rNamWzAIV/7r+Qh/5jechCEWSGu6hmEYMYg45usTKnNZ
DkA2Wpc/kHVeI9JlkyzP8XBU2DKYVZKiCRXsns2+XVfzpXyWvLblC1TwFKImeEZJdD1nD59nsc72
I5P14zKdOa9SyMz9iS2TOhUb/b9iTw0hfB3OUWKNZuUlRDDjY/9ec10eMAy/wAMYK0tlT6U+b7JP
T1S8kFohS8T+cPhWXkfTZFqTZ03Qe09g9387236VYqEPLM8/AVIPJSPRXqqFi6mTX4dWxrzyNJQr
dX6I65yyQ1SG2Sv64qfezU7qQO7ewEoA+rRq9Z+1iqFua8OfAmqBrMACuBz/+5YeXVB4zkw/JC86
A/rhWGLpLxY3/8i8Bvcw9v4fZq573dY4nrtPDQC5OkRBWVX+MBeMqRfoWuZWEMnbm/UjbUq2eCAN
Q5MVU7G1visUc785K0M3y7LoyPseooUcrtJvZqK9x9I5r6GVQ3n66QRIEcU/xbdbsjAaeiXaIzJr
HwdZzaTUyZFvFeIg2LoilgrhsboRt0up6KJh+M6ENewXRxEzgvBUqHw+4GL2LA/xq1Bd+8TO4oGT
JecnQoQWyACRwagEDzyW7bzaZvHqVY6Q3+XSyfkqUFUCZYBRSree8J39gS9srTuvjo2WIMGf6251
F6NnhxZSOnKO8oR0n64wYK9ZcDE9xa9I/KD9dkOqssG1srI2VqgtCev/lN1X9gRt5eWVl7jfkeI8
bVKWhiQJCM5BNdleZRYIbhdV7XhNrEvitQWRGAX7LKRHCQxEa+3ZhJx3CtRqXSRI0sqOF0cZmjKt
FvE0FAMqIV3HSuqIaXnvZ9vbObGoP38Zxd/w/00rJ+2p09WpP6lWtAYMS1oEGRwJAughcLpkuchH
UqEVKVh3Aso/wwS4zDm4RchGzRpOmPXf5/omZepJnfnAJuTBBDmvZRPIIYbOxpC2zo3bo4RxxmaU
RuwNupXetlH+ZYgNa9YEXbMObUp6i9V1ANt7kgYasPTHDPkkY6GKD6ohkErJvMsM/4rlbGaEMsM/
lvU6OWPsAH4c3Iuz3bIkTu4Jmu/kgcjIxEmSNE3Gg5QmQbGdPZKqrvb2eh7Kho5menzytjjmGoFD
/zw5qrqj6TEYHDbt9I4HlXXjZtiYKhVW5Z4ReTHwl3HIN1IMUsNOstn8jEiDvd59hNLFLwFZVbOi
4Rim/0885UPL0m3Xm8pPfI+z2jc1YKvon3X9k+6m7SRq97nkfxq6nHqWw1itn9vwC7Gu5+mWRpVe
LabZLgo0b+ojVPWnTGWVw0psgcKj5a4A4EqD2eetVBOcqJkrsGaoNAlV/86SdghiZ2QcjInOrV9A
4nJcjoPxqhD8T9ZZJgAFdOB0v6zvVgqi0Z5FTjLK3J1SvsD2N3AYW+0lLeQ9WxxWs90qPsnBrPt+
7P0Cz46GPALF6XU+Tsyy8j3IEL79EyXQTWH9OU1ccpgyXEeYOvNbXYzj/bGSHTsr5WEOQvATShem
H7y16YH3mjS3p6Xnmg1s6XB9/fCM1QWpLTiqcfKZ8r6d/ggHbC3MI/Ae4OWOkH8jLmMBoQoohprs
KzkPkOuAqfc1/W80ILsz17+UUUzv+GDq8gMCAqScd61LL/P852F6Nwvz47KYwjOTyKp4kwkKI7Fz
g7xqGa0WwciRg+c/B8UX6Gsbu1iTk+DxmRfxYUmZAf5XO3cTwk0RD7HXVhoyYcuTcSihRz0b9LZ0
pd2ZIA/TD1sxKEjB5jUxdhYVv3utoO/1y5+BI9oGwC+V/VICZPsIhSNyg9XjtMCv6HN4Asx+yNK1
QcYzH8dl8yHv+IfKmv+Yit3GwmkqQMmaHdxZ0V+sXeiBifzJ9CAPjZPD6+rwUamoFbQFeK3IJCYM
8MDnWGEjBQWugYMxn93gU5W2J/2xFxbcvXmG55S2SDCuCUqtVvNJA4RXLeO0ExbnrCIPjpWaShr7
jU6TrlIGgbyLILos2w1J6vlEBoaySMSw4s7yonk8yLNOPkNMYHk8/OYqJ6aNPjoGo0EfbrN/q5xW
fHkOjB/Ku5B4XC6ISbJh04Rd3Wbq3ryK2ABhWJeLZ+yFbRYysIaMHkZwfRo9Qa1tpjPWa7U2JOhA
GzINcQC+wHozAwZ51Qzkj3yzegrk27wuKuAuxl6vHkGNyra+sCwCfn0npDGeSSj8Kq9ARuO/K59Z
Ai11WXLHd+qsVcX4/8e0fdnOQ/JckShBI7Y+t0BRHQLhT2vxleC6PU1RUkYP2Xpr0E5JLCmBUHmo
sVSKm6/kc+SsS9NfxEbP+D8VqHUNVuP9wRa4Zj07LKzzOgIfIbdm5N8D1lA4MdZKXyOyvHe+qEUh
TkRMcpHr458C+27e+sjPX6rgGDfOWxxBWNC+z/+hKn0Hm/orrqYvB4kWtkwbpBkD2/2mzQV7BJy8
01fDy2TC1Y2Y0TO5DPrTZgji1Q5q4NQ8MdH+uwMnUKT41efnI4xhPwFg6YT5dO1OJ3AmpJ6t68yj
6vwTTZrt8nKbZxxYqeFvyfr1Q7aSCilyR7XiAkVg+UlwhWz5YjXzvd6nMiViS7odwU9dmi62RDTi
m51KVXX+Qqb6hBytUPirO+VY6DlEyBv3ur/1fabF+k4XRWKZOb8qw+KjXjqjRGsDU3eLUSf/zWDX
zVAwg8lyrRuRAV3zubbrz+OjjsD+r7ip79Ybfnfwjo8KBZsbSkC7r3HXuHHIsCaDABL408/CR66E
Zf68y3fnQZako9IqC4qo8lFqjM47cLeRQf5HM8JNrs5D8dnt8GRTszQnh7QtPVSb0bjaE4OUwEyq
3zlJqA9rSSlG+GTcgH+0QGRNrHYp2Jb4QHCl9VhjDLV36npTC+PtLSxctbJslNCvHCokAgI23mb1
NbB5YniIkQWzaHKldcmrcKFYj36VIF8Df+AZ216bKY+pyO/dDYbUVK0S70zQgU78/WGKezppzIID
qmAYrFDRKIOZo2tnbuOpUEt7DARLLzhnJearp9nI0SvBjBYIPAhubiz5RgMvoGNDcO8KIXO9nGbU
e6DEQISroiScGI1KhkH9nX5jA2XySJiNFI2zrP+RNfjzPwjItmcHt6reth519ix+6Tp1eiak42LF
hPqhr+l3miwIBu0BD5k8PEyrNTr62249oaXoxd9ed6goIMRG6F1FACmyEH43cpl/IULdr8srY2rV
tITaBJG+49Ff8uf3FHHBNVFjvj3siOYsrc/D5iacqV788Yvb0dFJAbxHW+eofqJByDF+TudfOxcy
YCx7h8H4Qg0pYxsMSsQCrslSlzU836eVIkZbSksS4pVnVtMFNXMBe9Vj6b13zQ83mGUZ3PM9izx8
UlAX41bYms+BUtjgJ+zGd0XJ84KjorpwR7KE5QpJ5S7vw/96mQXHO4lSJtLtpK5N1TOjGKIXURK4
zvgOe2CpwxChElneUb10aUA6mpBt0dNp0nc+PuKB8cDPC3xfgnX1UncEJruI9i5L4voeCnk6U2B0
t0MwsbBjefpq+ChjHv/MIwuiA0dQhwek8rj0sW2Hk2WwKOClvMfd9IcZHIcQv8cDJVnKcnl/JWIx
U+yJBcn40F1IwrxaxoqmrO2kk3VQ2iVeYOymY//kWIcpMDEbUBQdFZCtk1ike8zbms3ciyz7Eusm
9e0TupY+/n/PUFk5lbXNI6UlWLSk4nmDik+KnzqxtgyZgpNZN8Shcf6huwI3YhhKW0/DvbaqFQNb
6hABbv8gFQpeN7iKqdip9h/TL6EX/62+lLXI7geuQRLamfiSaiwlxXJJyDrX2nPmbp1KuBhyZil1
tWkwQz/qQ+qGL1s352qyKbXlpBWswbfDsWaPYgl+oRCP3frTCX4/+yflOgXXOA2bdGcrAhhKfYUt
nxE42VuAtSTBpHIFEmxE/uSfaiBtB+VEDDljuinTX2JgM//wkrFKhq6+RvlzGt1576gI94SxNA1M
qriKTAP1gI54hqKxlnXLbl1+JaOXgXTd/OG8DdHXzaFPQQT3BLOBgp6FCv7hD7YF6usrxPmPjoUg
6Wj03hxi/eDTBNc0QqUS9KLfps+dhaQn69zlz8io/7Tt7ZE44/f1/6CVcV9vuRLGQjWhLsNskIm3
Gomonyv33MhNowGjSPllU7NsMqprMxm7C+jUDvyO1tjhhgCfgRxBiOFbz+1ij7kJCRf+shBie39Q
5Cc72z5UdBMLk4+isKznlI2M8J1VSBkGB28+7xNAoKCWa4UB5y+exx7g3mrgQJLe5uYh3WXk59Fm
bONmNsjmXHRWikPQlt3BByGiHZS51jUMIYAWiN2AQ0po4axNOhYArlt0g+ebIxoj6gzK2+SVusc1
HtYmx+FNUxCbMitZWn8Hre1Jg6AsU+zOIu/9Xoc+rf2WJb6tRuDwALYO5pUIKg2ey0fsyXnL+33p
9bD1ZARiu2lj7xZwKiwxUEPFZhKO5yJz2XneQW6CvRPNKLPGb+gqEIA36l6jplUHqupnXY3hS80e
mh3UFvNm+vSmHL7XWoGquST0esT2BF3UzsXddgCAxvl6NbE5E6tOQ7tMW5+5KWftsshWcBzRRJD4
3OZAD33qUuo33X4R/qgYXSRh6UQ6r4IQfQSQd2suDsQT7gw/eMuU2RuB0tSuToU2FFO8eA76XR9G
qSdNg8OB6Gr2wM2cK9Qbs/87rC1D4D3uWubzNA0DrQCkYYWOML6S6H3gHpFIiefiIy90Gr88gqgI
PFRdkG1OCA09fke7tEU/919j7MEhR8DBvpbMk9XFYmIL9qkpjFwU6RoPPGqhXJlZ35vd5UTfesXM
jKqLZoY1gwJIVT7wqjlGbGX/lddyZD4E6BGzJNlzJ1IBeN2umRTU6itvb7P4WFWCQBYs57VyFFiA
ArChJkiTzSBVKsFYvLatYoIXYgS5AaAR0aErs643dpzTag41SNK3yjkQTsUU2N8qRgk9+t1zkFQT
4GiaYD5ZdyOSE7g5hav0t5qgOti52UFKSx/LHZvirsfEPkyJ12pyMhxFLzotrrjq+2EaO04BlhUj
AwS9WqOWNUWmQw4UJbZPagBEafhT8tAE6S/BG69I5Ampmq9kx0g40wztjPIKHD5N5jz3UBjJUXRz
GL05eQQKb2Tq2rSnFB4nD654yoFfXPOrt0xuJ6Tlh/TkyXuVu7yVSRL6taxtZ2CC2re1faQ/ifeR
UVT/SbCpAXHCza2QrbPE8aumFhZJVQ6Y0loV5QaIbXX3nyoNAYY+FFtvjY1715AYSbsj+JNyYTjS
ZzM8UY9LGq7i+xWxYG4X1BUMsRto1TIK2Y0AUOGKddWHysoGJrLJJdaG0vZzsDRiv12fguJBcL4+
yZbuPchYQc1F5FIVb7XsJNbhcZ5e7fYzpVgw9Wra8eZjnB5/SrdEMCP0rogp2+4y+yDvgCUKq0vh
NOsg/RHe32DxXONkJJp0cj0hBKwixUBojoCFats4N9r+GnRPHUY8iCGrLWObIyQFn3B1t2V7S9g4
G8Z7Gow7yC8Xib8iyxbwXUvR6c93oXUaeewjdt6wgf+aaEy6evcIcU8k+7m/zE1iV1640fvTGg95
hu06i4uAuiGFNLgeAC7n1ZgxcfYfdOYjUzGCovPy3Zg5fqtmT2EX0r/YTo2PimpXZ+OsQtQD+B4Y
OZYvb/r+XLzZbAAD3kS6wRq+IWaLIzpkOKqfDZRgyPvmSToCWTcBSfn9bXFd7Jzp3PNQonT/JEmb
AQ/8y2Xqsx7XhhQ3VWFmR3GFQUeXCfZnZU4wQ/Tt9Vr2wSYUvTXROeMYSjWe7zDYd+bDOYBXDTmU
L5WZqb5+4nX9xqsDQn+r2rKR5rgc6EaEpl334WWNDn/0on/d3sJN2Y3xt8a9+K7/ex9QdIFqEiz5
YdxW/0qGP5YFk3Aoc0yeTh2DxrwhbamrMAlOa6vf8V7OOshtdJKntp/o4MlQkcQZBu5fLheQuPr0
IFOalRgfGnkj3MOa/q6uN1y+R3cxEhNBgPrsuooMiGNIt9GQuw9/9Pdxv/QZcAfGXljyrG4nQ2vv
xlQZqPNtT/O6NdI2VnHl7VrqAtx5pH4GHEnRlxiCGWnIzww5bhAbKbOyMfJzfXiLvi/uYK82Q2j1
ymKEPyxvewxxHH/QsTfBAscWltLHHkWXt7rkAeF9hdp+Tm2xpX4WoVGbrmjvyWhG8MIa5RJGb8QB
NrNSd6X9imU6nUgY05hrcmqt52YD8zr+5d/GYDHAA++JGaxq036V2XuwrdN6TtszcexOixgHmwAN
22MbXU1n1UoYHRt+e1vdDG0qsj/RUykH0U+kHHvXi5v+DBrohdCUNpysh+xZkCKGL2FxpUpMP86i
JRuXvB36Tcjzc2FTdcnYULRLtupIEBlDx0ael5H0nlJ5lu7vIpHlFEN3D5ZpiCT1VU3AsrOBm1Oe
6mhxWHtRZDgrNIc9I18w4k58MRZeK2vk0eMSPpBT24Rs8brCze1c5xNc9A5vu93CASE7gvuGIfwT
aK13dG/mByA2JEmz68JZ9erntecbfaAtt5mymzpJASKo8i2E23+kBjEaYDBZFDvnZgjiIKAUhBK6
WiqtmLu2Hwgcg6gnTdaiSUaWia6KOSGScrzF7PnnHEq+xhIL6oI5lyen12+RyaGI4XRqTNRPzS+H
AaEOdwYzfu5zg17sOwAS5Wy5ds3j4yiq5BwkGSkHc47LydN4uCqBnb0NOtBHKl8humY9dw6QBcVl
Zn6RFPFD1ha22/3QDqMdEFi+bjh1vO7FTr4n3KFWtdBhVDzgZtBe3h2+JfCpyugR3WbkB8Q6EEup
fyTVtAn3gHnC11yuT5XB7N9BTmcn1ORcWz6NRGkBeAn7szwNBtJeUS1O4T7XbObjgK6Ac4yVWqJA
WNN0svf7miXGGd5wUo9G1kiU/kwCysFZSMeUcHPJjDix1ZXRIAqF7B7sh/pMMK2floNW43imnjaC
XS07j7YugOLAMfDY5lSQmQQ8+ovSxKZZCFyHPnCL4P0ydtPcOs4/jVKMXi7RH/5YQSXle1rIX/Uv
1cZc2dw4ik7EJPhiIeJ335fwAjWnKv0rt72voDHI/kfSp3jM8GUmxRZp5nMqUft5CZExUo4HrhDI
xZuBP5tT2ZDMRjfVtZ1nxdqBLwTaHVgyw5OAICASjsm7lPRxJ3kzlADhsH8jaWH/C+e3cjYRF2lc
Kt4rI6bZuCfNBkrnYk0ktP0hQJ33esLslEdpXYCccVeB0s2TDWte2+njjPtJQ5guOhiHQwgPrlYk
hVkwhudhCOQA0BJ/BjZQiottkBzXY8hET6CXKOUc2y3a2YT4OczTfzezhyORQGfuB3y5bhoVCm0Z
16eyFkbrU+baGWZy60BhFZ7dwdpNp5J5e/lamvDy9kWZKTvu7lrQT64FNImC9Cm8NLmn6k4bzyVb
bghTba9waEqcsM2zj0VA6tRbbvvIhiSzGTeLmoHhxrKiPeVtDM3TpjV60rxTgT+I5yw2rsO8YDPI
meWxeB5VdMVULIlZdgHO/94SFDriNmmenFy98G3YrE/iWghT24KRnynCysypjoadTzkpAHWQXajD
DMa0HDNr3N352OLyNDUkk96r49CVoS5AtWRbTuBdQ+nzPaQwGUvtH4o9EmMpqzbYtHDBIX+IP4Gi
kbGv48XbxUqvKDDoSQizHb6XUIyPm8/McK7gCxMQSXch37ikW8LVv3idPGCrKGDcT9WIeMrPZ90V
z8rjvpYHNMAsf3pNkzr00OKw3QGNc33SPyhwL+2fERsRD+ct87X8dwzu0Bi8RndsFp0gDdWzDgSU
BaZDtBKE3GRpuFNHPwl73b1Tf6LojlHKCFO27b/I/5f+pxk/nVS1zSJJDy3wwVWOlw+BCuSaeesF
r5tXjO3GXOV3u5On9pwks5hpyUi01EpaRsLKeoPO0yOJbq1IAL2x3Jv4tyi5Z4ewCFh29bTXn1S+
JJqj8xye2Zlp37sTosSWokP0NdRX7GnzatPL5Y5tciR3b9nmVSKxIyanFI3Rj9/Jze+fj0OJcRgH
p+t+s5ny41ia6wVMjXoeIVYyoVfPRjG2MXvZr8TZMlabGFWxT0Lr2XvuZ9+MPk9Jj9CDugvlcOaj
l3+WMgE+g2uh8fFtiNslgRS0+YRH20jLMR6xG3vOjlp0CUnf4u7C/m/H/2ElH0Ml69pVXqx2j6kX
ZrZ2t1r/924O5aMG4DhgTaUBgd0R6Z/oTQcb7qFDROqe4lL2lGtuPuEyZwIHmXl6tiqL2wj6rkdv
S83YyQVK3CFwffTxB8he2ADSc59UzbhtzSY4WHLkIupYEL2OQGDagu7VNge+YhXNMRNA5jiln9/G
c1NJHHm5P+xpRVEOHrk58OT97EkBvkCTpi2Tgmw9gqS7km+woldBY8EY2oxeEx8d7s/58lP/3tkg
5joGrlg1sqUkc8T3CxuW1eLARbFt/AqA32ZMavv0FOv3ZQfvq7fwa/D9M9CULWgNL1+yBgLwHXms
C938rghFFY+Abzw1I/AIidTSbxkkpVpo4zCuumQYNhKhGCDhx5JktQVejjJkJU59zdTl/tE9NcnF
TVMD0Cprdad43jKFAl5dMiuLo34y8nL6+LUhoi8NXFy4yOkXH66juGwLKTRSsgkCv5upN2Cp2Y5z
ukLmwVD7Bc45syr5pyPfTwC4jMryQWMwPEVtfBMAYqOkI+Gg7JSehr/BiGGr2IuwFmlb6G52nL5r
/i2JO1oG7AdSyXi1Oi9bv1DIQjJ3UKx2ph85NTHxI+vYIQcPiLhlxIaNArvgG3KiycgZdxojaGmY
SV/G3N/EOK26dAgx4SkCS8RxMWmtMtoMHiTHBp4tENU40MWuTscvJUdGEQT5ji/a6HxhJYTKszk0
R1Cx4JFNbWXXSxwYq2Pt7QGys2b+chYcKanyZVbR2U6bLHETNiBGGukVQrXBXK7tlckQxWodzNA2
pyvmjPJOTeK/Ikt1h3PN8b4TxS01ZOOBXFhgzqEJrc5kljJiJXBYglTYgnD1lOpci1G7z/I05bbu
70AVAOGk5GafFU3rXWnZNfmX0WiEuTMMTL2XT4zxCE66Xu0OdoVKKiWiiYovcYoUWCppxsWX+F75
Awker6rkBUlc+5VNYFex5z8NK4FJMuWKo0lfWvSkC8qKg1BZ1MoksDM5KSeEiUqZoxAE9OxsHAaZ
2FdN2YgV4DQMD0WrLWLQxv0RYDmj4uO5eumMo3+pOEnlMCDqj+KpFc2/QYMGeJbrq4PfxZkl5VFW
AaEoby9sLNUuDPvvd/ZoVh7WsHrdpUwjFOqZ1UmB0DpVLA1kTsHrK6bcprQyw4Vzy4sStvxvLcVK
xLwoGH2rvuhKJdjC0r4ThU2gBwoWyEP3AC9CiWqMgVXcG0PnDgZiIyytOrUDsj5H9h6UnhoiaQ4R
zZKjyeXCCzL2y9T3cwzyIzrRU9FbBUPTy406H06KsQqYVF8CO2uOm8s4LaWHLiOS2WTTTGOAtK/s
/UO7GKcz9hQNDVnzi+agIBPX4N6eetuYyb+zR7uJB/wY+AWqnshqESfCkhXbCMy2lnemeY/QSGZ6
wDCzTISByGE21rqnJztSAr8pTkcWQRGSn2sD8IJ2NugviUAEuEOX7t5kkyTmpnxYEb/dFT/mZIJO
W76LR6CPsR1PSv8ry1h6ndiQcMtJbX83UhGrzNsdXeiY8o+wkt4IpKkLdCj8n/827a0ZCmIdrgnQ
7saAJUCQO+OlVVjWIopKdH9MGOCKGN2Y/4+GFe5gQCHNPc/0QdNjZ2Ok2cegT1DLIgkiUOwZUBbS
ENA/WtMjARUCW1md1l7vrIxEmOXixPVqStjkuIRhmr7zixhpyqFrkEcCbxb+Gj1AWCBp+1bdx7Se
OQTsLXDf3D74VsB1G5BvR0nZ9qX+gJvWd8D9e3IL0+7ExYhYCTjJbAelXEYNNVotNGcPOIUYk4UQ
fAf30KoqHczatEk5uRXTTlRC71UvehtR53fyN4lwHiXHkTn6YSB8bsnJOtIS82jObDPECCmCKySW
Uc8iLt1DYvnT7qpwZ/Xck1qma6B6u3kJNKwpdL+3nzLc9JTkk5e473Plm2d+DKd05JTNHADIJ0M5
iQyk+uItsh+8gsPvC77qPrRqzM/rr9QOcCjoOifQ64VytLcU3IqFzFBdHtiUG7BHgeU/rh8OtB4k
PQs2twVVBr9YhzZgE5XsIbG6qr+45mmDsNoP2YkSI3fPR7dZhGsr6VZfYu2xkiL2Qj2sTSamNHzE
Be3MICjrWp3YSFlV9ezBO2gkcIGP/OgQsuKIH0s+x7zUOLsRNFE5Lz1RRz/mop6yOPQZ49C0y42R
3OUZfLDh+8PPEVrvIyH6CSuFgWfKTOteUFUkEKftmqX+sT4iNx0GCKcaXVxZLUZ9CYTaGylcbCeX
bsa5R5uYtf61Q9AmkGWS19Z4qdV43W0UYqEfqWBTHy0h3Z9AVmjHaGhnLrikIkVBQbK8uqpKSltF
L8FUVVeL/MFE+bnZR1ibf5uqg1VhKF7I1p7ExFWtllUKr9xHwvzESZ8YMeTRb5+ZGq70LtDCy4r8
/NI/IDlmIScFjgfl349RyYWDGKNfSU1AFb4EemV9dP86YX91Xtw7bC46HfdniMt58/xOng0OvqxO
ZOCekyXpJhNIvZi4coYK3TgzEA0YjC5+6YzTD9CVx+qBO7XvsHJQzB/IM5IWUIP/jm+aVZ53MmB6
7uHPaMCroNAooHqy7l+18MwX1X9m0vhsYpbH+6L/e2R4Nseovlo6pn1qaLdFNQFFjjjDr5p+Pvkz
Zd5fO6m7DQJTsVtjgG5X7rOE+KWTPycBy5202vpENl5Ps1Ek9fs1r2ANkXlewknq2UipShe07WVI
FqzUhrfrpq1DTaN9KIUu/t8EHkO6DbPzo6PJdRwPUisk8vLB4MrETYRzfPNKKRcAzfHofWn7J/bV
S+mKQ2vl4gGfA23i7EfsPjQA/0y+w3MQyuz6QsbAPMdeODl5uVBDQZRdH2B5mrokCL4TKcrJBVZi
ZN8BBbfGgCEUXpw7ShVGElliyHy1oEsy9KGTUwmuueA/giKryIv1jVj/f/FqIzj3Bnuxv8qPu2Q9
m+6D40kINSD1p3nRwGHWgnyRrWVdhKO9yrFpw3ejg4zGWwS85+m1FUq1Kk2lYgdkClrjBDy4wlhm
X5xO/jPmYy7XaaGJHilbhliDQPc7qUbvZyFq7i2pJ8PYLW/xy45DffjkxlJ3PMUoaRUORvjz2kQp
A8qMSMUPSSoVzBErMzmDVFES+09Wq5TXSUZO3tS9gqUGmVNi4tAXNwoWSsGuwmxQg1X2cNpLPkhV
TXjIMOSRo4ppK6RkExjZXzf4um61qTPa/5G/W5GkmkbVNG+ybt+9vB0e/8ScUM3BX9cjgWzyMr4U
2g0n5qPeVv8lh8lpepH6fPfwKCKCFijb2Yz1fD8nbl3HIlFlKtZXDUhQp2uV7ZmMm97yQ2MGChPh
Wn1EvHzJaMsi3JE2AZBjrz4ICaUwo9FjiazDEec7oC77c2OEk3eP0YjJwDFILJsZqkjLfvuy3Bhe
qe8fMZgdDNd2WoYgxUJ8yFI3r/1X5AJYFyDP1harAslMNu23x+dFJlSDogiLXNe09i3MF/2nBpem
G+/xRTAZLY2H6jjLJtJD0DrBOIy42K/vC04KFOQaTsU7RpdhmO/yPLZlfnUX6aCMTeG90ED2eA9t
CZB7TtbTYqLeiasy7h4nEe2GjXIukYo/hmCUc4MMg6vQBr/vB2ndLWsJCUzKcFpwQ76zLccNnQBI
EeEQhByeCnztvhE3pb4akoCbUgptbFd9KmlshtNtypnsVkgS2kGIjB8OSaMx7T9JX7IiorxgH8fD
cdb/d6rsad9u0kv8kBl+FsCaHvmBLQDPpWtnRvqOuqYtINk4pR9GuBMjz+nQsECqobcVvhir1Yui
45OxnuuUUv5yTSEwpB74MArCuUeUvE+fkVhMADHi4kZ4SL1zPrxL401mh5RukSiMdy+j9PFMyKts
r3ZZOz8XdfjQJaJD6ueXX03qevsSHV59xRuWtGLKnIlwOAoGVuUvuAwXh0ENCAeKd21Fjq3B/Qdx
VftKNaAuS/CZJbt7skoheShFNs0sGPTB9LmfLUaUgY7gZcvJGsB+3II3ZtV+bNynME8PxQBYDcyY
H6eafQT0CcRGxIK58Cjp2VvMkajEMRaSNwp62+TQFXShb6I7aC0fFxd0bxlyU/BmrZAlSdxY9PZH
//Au9j9GKT93R2St+z//pYD8AoXjVsh3h/lVo+aUP73QDBNdY6fmy7Z7WiM5apJ4YREk05KCvujh
yNDN5PnM/bVwp/6+s+WqEMFi/kvlJdRVh38nN3BOv+0IdqORlaaIzsPRvbmcMb3Se5A2V58Z57RJ
CpFc7kwQM9Mxi2y9+PGzsmko8Okj0k407kBwDkjT+y7SbaBzzEUybbHxJvCQVNj3RTRftH2I/Qno
ORSECwx1p0+TxhtsDxvFu33UfKT1MQrAcqVTcwtnzP0VrTWQejSLCSy5RctKFgiCft8gGNmR4nSh
Lp9itT5BYRGi5jAJxOl/BtahscLdoRacgBtGUGvOflrR57AYKWZRnpu3WGWEhVD1vX8O1ORqyseW
rOLvFqQw4AbTppXqQOGh2toWamIVDckq9urK0P0RQIzvgIfZXjohStf975kH35wBTPe1CigUrijO
5CcktGrzui1z4b9zmWb69avlXDmr6cOmHADtWqQlJTNaWcXl5QG3QIOELbxlh+XCPgZL7LdBlrZH
/7LsnTJSjIExRQ3+Ql/rnv2TBeQKOyeo79QBYbS67Xa/uYtAxMqrKX1vwrpJfB+/g4lyN77Rqe5e
xQgL2kg9nU6gxyOpYckJU10kHUg231aDrbicp1aScSZj3xIS7LKQtXksUbTgTUgmsM7POWaZKBz+
g7+r26o+zC0wp+jvtMTHL0mciPYLtYjqXnbcMaeqnrKR8HyxOfrwJ4yHvbW1jw0Wk0eov+tceMNS
cbpaUChHSbuQivGCLtQVNXmYk00DRQjrin3LiYzxltHLaa1CwsIKl9yTfbPWJxdZ8yAx4fCDY7rT
z73LoJs1cfR8Le+MstFg1zWd2Brz9tj1R3UY+U7+4apxYVUzwVGG3h7bNPlJRn9RbVAsWc7tr0H5
Po9m3syZUR0aiuWGAkDGrJHtPLS7jstlJcugPHbDFqYoDPE/SK70v1XchbI/Rkb3oy6l9I2SOZEC
FV/iqyDFeYCfBBdL13IJvf2byzPgUdGIR+6mxmtitt9ztQtodHfHwKqKUxnvzdhpUNhiQqXnRw7a
Rkzc+CR6K3KwTS/+k+3YIJBZzEJ30PnqpIQbXWz6QG/CIpQVn1bsAYzaw4eO8DZfeOvTsSIWShcg
9RT+2urbZPneV16I9wELdPlp6Qlrf/xiMcyUBMawAJfEDoi8f4oixC3DEIaM5/g9lv66B0narNtc
rDJGlBRoJN5xgcm2+0dIsNveIQxf6h2r9hcX4GwF544PmrUMFGw3qmzXjVp7OioYGBTH0JgWl87/
OmeY/xGlMOKDe2tEAR8NgBh03rRkyBSBUje7MV18Ob/a5oYEE9ehohw4O31ozgNQWH6R9snkm5ZZ
rCTkNWMkTrHYpO/kTi4t96Qdkxx1U+39EhkaF7OT9X9YJNLRxixxMlXUQqyiTtVSSOAy84P/SO7E
byh0gpI6mMfw9PqGYeffLmrQVvg/rMygMi+1LzscdAe27kDEfOkbtZRqobFcVVPmdipfxaQDU0/E
viIihuIQjLnDOnejNPs8GL3sxE/xh2Pm82LRsCfcZMzLS2O91eQ9xHVbekeHU/KE3SSP8fxKoMbZ
cAl+F2lrj//F+foKpnoS1pSEVDtW8A/9yqulxWNaDZkJ0jWKBmn1JGSThviw1rAMJeNfm81oqpbj
jmoZ0RyDbxYLAnkzGUrOUsbSNAoKq/zIEKwOiEVJHAj7zygrJMhQhFViVFIDmMzESflyt3VAapoY
0TdtBrefC2OQai5uDM6b50sbB09rzOMrByx52qjtCbvqiDVBqQ1TkxdnIbzF45n7GAtxOCYRILZV
m7E/wCKrfoOF4/aqfmb0sR3SwvUY2D6ewrujBVkWSDxaxrfGoeYNO+F6QQZyu88ToB11botJvRq5
C/z+MtmclSQHHXg0ytXOm2zmuc2iOwG0vZ68XIMZL57rOnMlxD+tvDNVGMR1g2j/z3SwwD8Z0LEH
++nK45XlUd69v/3LttgwgKQAaCs4dDedENvIU8R3FFPk1gTNLT6N4cASNdWJfOam6ExRl0p2wdaY
6Kwp5bQndDMLCZGPtxJaqXGjAr2vwhPiUhUK4XNh93zSYuacPyKTyMRkGSqCIJJUHsVpW5FZwG4f
9sJycar2Hli+t1mwU5Ib1VNeMudiPh0g5A7sBFux+ElguLqgXPX3CeA/EfJnqoCr+tJr3zVR/4w6
qJoiWTz7lTkjV6eJXffXG1qn15Pr3elU/SB4VdVSB0oOKYsZ8o4dd21oi9615ooj1fBFB/CPLqPU
vhM8isoGP7Rz/n3F02DfnntSqNhILFcxk7uoU/b/WOpV6YHbdsNkB3g2eXCvDfuSV3ezdy/G94eb
RR4Ug6WAFOzI7qZhmoHN8A43nnpF1Oyvs1URrUq+shZ7Chigh8UiTRoib/977+p41DOK+OgWQrwh
gkiwQvtHK6dh3qseNznXYRdM9eUNKI9kF387rWXryFuVX08uq5NMNvFpEreThasgfO0WCf9jbBMI
dQ9FQd763Puko5jLQ+UfBvfkPQVqGiCNT2lLAUv36haybdYC0S7HP5L7LUGxaBgKllDbFsJKLvWU
eNSurcPTejm1FSvEYh9+RKK912SwXaTfsCLNiKB3g3LLOCrOCcEKlmPhjdhPzpeD0nvD4Zl+sD2I
8+6r6/cWA/MEG66I9M7XxY4eLckpysERZ+cDy5n7sekQ4bqKFXfGmpPA0kSYAL7OAnGKyD5DmLUd
BD92F7TgtX1FvcJ2xxQsMAdot1Cey3yNFJQcJHPw//AunzthP4moeGYLS8fxX8yZm2yJIJ4re4KR
8btsAX5YAH67tQ0gr/PWyjT3BTVh/vqLFigvwmb2at+6U7ErT2PtU13fx1ewW7N3pTA5ysoSutMa
jCXsQQI5ZEUAsc9qt+fntEEu3mME9dChm0gWlrKIB6b8RRrl/wBVJlQYxiA16rDK4LBxSZY6SbV/
ojSlwn7TMWcMjqSB2gDqKmC0cDB8ausyiHxy17QnnVa8/+AEKsDpqA9VMY1B4E1RGDYU0AuZ5gde
kh02GzSwYamqNCHluv1Zv1ysVnOfgwx1r30fE7F0Ypa4HEu1JwkuuGjJaz/51Odhzh9noihrlc3U
PFC8iSPBLtJ7Fk/lulT720aKnDb2kThtSI00lj6/U8v99fOqBTrdRdW1yYNMWcChoToAIY4GYBdx
bnnpFa1+OLs6pDLaHSplXPioAQ+Yw6/LE04L5gvau6xu4OalK9gkqzviKwLNzNYYmkTps/3tMbhf
xmz2XECxJb5pmRfxx/0II9/+8Y+9bCBsHq1VLYNw/YfsUTJ6oowCqqokmDRfgB1r47k3g8YCgP9V
pm+xdGXspgZR+0wVW86YYVG5Em4BMFmdhrplKwIvo0mdUcb7duLuLQbLi48Y5w6gXqMful7QQQvR
2OsrTh9HUnOCD9ukCfU0oxEubA/XPejoWPqW8FNMWgfLlgWn74Vg2jQLjPc5oHu5c/UqSjWlRBZD
IcntGKcF2EfdR2+3nQkrzldPtbq7gQEeOMxsQxmJzT7GMp8f3ik58Z2B0I05q4PI50ihiQijpyPF
hNaRav9WHnrVZB8GkaaF6AJxVt+GEdbhp9y7hkqKMWJpOpr4dDZoeBNDiH+CiBcJQKuh+g+osCyz
ZvYhxL7kfHQR4v0oRsRGwA9Zj0WY/jpOR52jpjWOI5rkvuSRwBlOloFwQrEu3OfzzHfkM3ej/9nz
1JV5ucAkxHgjO+dQESzqYn4MT2vLeb9RHfdng1U0WrIwLk2KJLCwgOrkmb9ZPOMwMHFgLMRGGRO0
4QiAJAYxE4Pra+OCk6F04nYP4Ho92S2ZCdwK1Wzr/vPgY5Q0uE1836/EH63x+lGES9BRb6pdreLz
1EBm6O8pnraxy6abEc+rztIX9rJrZb1ALUY7X9FZSWBXq8vzZv95ZsuhbTN/OL4PVtiV1JpcvsPB
ITKOC9OFW5r5GBX7FeidN3zZwU2owW2J+LVIMDs4OWgwQHc17xZKx4FUxT5QhlkqvoFzU/rk9ao7
yus4zQMxz/ti1CNXEc2WJD6oPz2Krc0i9u1a7DxJMqcgLsO79R7utOAlcHj2RHBIbc8wTGfd5FuB
Zaf4elT1ItoMWcBfA3Qg0wj2dmxtdW5rHb32uu/MkVbyu8zd5VrtU53Bd280QJCB1p/Pb+U9uadj
1C02IpdcPMuCfXLc9rSOBGSDA2Qqg6ttzwtDT1bPRp5N80uLWXo5RlNZku++r8mgy0hm6XJmBKfI
tmM9JlWgpzQI9GxPmeo77uHFGFI6DqRM4K15MlgE1uMuzAx5D0IPGU9spB3TKGSyi24l6pos1qW9
lGI7OlAoLvPLcRqHCHXA/aHds14OnHKs1bcSKUgHPRpdQJhouwvfxhokBTG3l/KegIWzoctg1Wba
9oYL5e44UOjrjcbGQ9508Etnl7agPDx9G/IW070ldbRa+OpxNmTN2HX1AQs3PyHjaGPlK0wPuZGk
9h5qV2fKBLkYAu95a0FYTr+vcUxkyZhWeBpwEExnpZ8Y2ViIacPtHWGt79I0PctZ0nLqZDbxNfPF
HB2eONftri88x8PFmnLwATBu+t+7Fr+GB82K/lAlfkLdALzwUOYRT1bYxkrsT7POn3bjQbOExrh+
ZSGCgNAFCxZlREPQD9jKndOW7MGI7p74xj06EpvPf0CAv8xjEjl84iBgMjGOgcdD8DHm9ajhKXTc
6VUBOIJSlNNsUUxNSv+cHEJyFvSXaSnsu2vaMJyrwkN3tmB8MOmKKVyOUWMdfRzALAMs3dyKuqSE
PaP3MabXEct5RUmqR0yuiXXpWekeRNXG+vU3y0WyRrRBE3khkrzAJsULT78VrRyFWbwEYxc5ex4G
Bx14a/MKu4XgcQDu3WoXm6qCpvzbAl4AW6/Su6J3fNmdnTNSyfrdROHCZ4IOcQUDkLsZjt4GBh3I
J1M3ef+M4gOxZ0JhbmkTpxfEPCvv5pciD/yy6c488v1HowCo21sJazASgSOv2isj15s65htsEtMr
4yzop49z3wxyRkPnd2RJdXiySt0T7CeL0ItRlJqjmSR/qmcAbffNTzmSEO9VryT5Goh0bFEUENMv
3O7AtDGmguX8T31c9WZrQYFzaaZExj6SUKYkyWs7BcvCxayYXxAK0zbB1ogh/j6qVCSfYCmxmKvq
+JObsIDVfklo9KQj4QJPbPdpig0XA4cD4G0X7Z5g9uNIA0cK7zPK3smFv/B41JepWvbmfax+3fs3
dmWFXiDn7KRd4ALlUcM/RMqvanQyMsWhDO4VNx2AahqgXuL3IvSuBUxBcdMd7SJEAoIpDeHMu7Cd
YNKQ82lvHQIEICULJ1jBqCTuE1sNuNEIkBp731Nn48Tgj/O5+CHuDtdYWVxJs3PHrA/oa4SkLHD6
TWCyjZQbTr89+2qx/Ah63oeWW5rUrluSuvSzl1DzU2rzM2AgI0tNrf4GWDAB1l92dY8ZX4RK1hKC
UU/y5e5sQSYKVrBffzbuRsRX3Yn7zO3bxPsz93NBLV4Q7ryvCrreeF8r4yJBNwmHLYJtVmcXOYc9
4szfEHPqzLqkp3ZwRR7IBIHt7SJtbD9X6O9tgKAw6sN7gDQrd0D6dOrAtAgfWgs3fYDXKtfMlScq
n9QjAHM4y97gtsw14cjsqdPg7zVVQc24zCADhCtTTnGe3/Hr9jkFyv+c4mwAyXZhS3DkKiV57V5r
g3RqcDXPDliLSjER5Hu7tBtMj4zSDy2dEtGANi+HcPcvlF134U1rjjdbTO5eXUw13Hq/RiNusXvY
iTN5mTE3RaYMxJFSA6auqc7pNYEBzTaLnnk8oFBLnZrbDmQKm/VkDxIkVhGugntRJj7A1ArHsmyd
bocvhbXsU3Pv7BwePiT/73obN2+aV8areUWqANUmNJusUWTRGluOCukEPIE6O5szloBnlDYUGICY
qIeFvte3ugN9eH8a0FT8wLV+njjboWQTX34Nowvw/dZ1cyH8XdDnSZp2uDq3MJIpmM3kE4K7HXdw
UkN0Z/9w8T8pD16gXwOkCu4WmyLpMKqVV6pl1d5QMKiqy6ReCjoPtp2vf0U5ILQwCL9Vh7hD9M+O
95Lsh0zySna5ZsrA74ZmjfEhS7brjpCO+bqKwE10JdLZF9LiY0G7bq5iudWY9+woDnqItyUNY14W
vBfwSU0HKFFq5Y1wRAVW9pxWUWTLWeOG47R6cmWEHvOUp6Okn1vnfhG83TVz+c/OhvhtnDq8ql7Q
zsZqf7tHtszsN6T8U05eO2HpuSgX1w2jM5g87zeOrIOsNw0SpPk3ccRsYTuQcgNBI1cRUrFR6ecv
CjAXr+f5QgHnuB+RYXqq2kqdWJduoBmuE8oCfPbCJPK5ji2LfNbmdOxJDDbAx4LX7uB6t43yEOAI
vHyYYnihAABv8CEGyN5vT3J6WWLxJyWf59r6DhyHRy7z8M8dpZk/PQNq3p4UF/4KdRc+n4M+fFfV
sHhUBx8QDichZnwFh44g2hWAqW2H07J/zXvuHrG8/fNmcH3HEzmo03HB441Ra4YnUf2BmYv8KLXw
Gp3lHubg92ltX39PvRGINP98SnLIRjWhKT5X0YvfUwOat4WRFHRafgjTA/C6n9qbb0Zj5ioi85oL
IKoH9pefaE9yYxjGSDyaAUMTqURSRF3AlffIiL9JeE+nArMhMztd/R+KEizpLM/IcvotfnnhgK2p
eyP/hLuRP5Yz6vCCS/MJgpu/xUF7IY8ijrrmDfN9bawVpWu4Ct0LJaiYAz7oLf8vK3guzW/Lu+LR
LRd/Y1sG6DzOU+TvDWrOK3+HiYOWjoSrjueAFw6wDfe86p7DNV8leo1QsKn4p4QEAnb+OqvtE7hR
XxQCGidO/YQFhtFZTpf/StZQtWt+U6GQ2IIbW6uOXWEy2nnCZF2tM2/92aSKQVmLNgricdwrT20G
XBtI5Feu5GT2FxZHUPcZ3NTIrK8K2NDkTQk87MTmP0+yMSUoqBEqFsgmJWfZxW1uHhsKSvZxuaQQ
bNmsUyz/yDoGzgRkg5fwgEAJKKsbOMiTC6Aof7bFcgvAkihErbqjqWRVoeNWEm30cQCxRn2KwivU
/4+vS/tsVzfsNzb5OP23hUoFYhtzXzK4WOmbr000pBGij4CVmOyp8bRB1D6SYpanPTFfIpI/TyWN
kqHARBntMlxCC/4w+EleBUszKHHt3DCuAiaQSNJZXS3rC0uzYPTQKN/1yZ0Eas3SwK8c6CQyW5LQ
O0tmw/EIbwwu6Ck+nSQj3d8D9oTRx5vfZ61UJzJfTZuiB+XmvGLb0l2uSIXXIRxxVvopZCmNAAnk
WcVgz3up1UUmE3c7TPWFC6+AZIZ/o6bqGicAO2OwRa9ii8d3audqvKvcausqn4LSV1ovu9DkdkXo
jvJ3qE6OiV3oGVGJp4IQu2h0sqJ+i5hZaC2KSE7Va7bWGFXAMAZvuZOhRz5hiFE2JKQRikmHEDKB
2QiMh6IXVVKUbTdkFhvAk5YiJkCjLXPW8NV8BAaIuAsyVNuQiRPX6/enguXD3CdCNyaaDdJcWc1w
kNWzg2rgJExyJAtC65XRXrDt3TlNiEz/vVb+D6ua2CbnE/PkXXg3e0IrHDM9GnxL+iJa9G3jjWb4
yjQ3j2332blg04qR2XSObEWU8wA/2JOXi/WBhCijLGqSqXnBmW+kHK9HhkorQikAz+oZPhFkRxVl
3xi1nk7bIa963iHs6xnZTPsQq5pPmCiWCGIGxaC4/bns5clNk8Vv9RbnEgvUv/wNURSRnNi/deZK
i4qb9GeIohyxgapbm4uY7w0fwMCjUfLGR4wVP+F6+W4HhdEFxnr7RLguTG6vNqWueg61tC8Yf1wl
Xq/DzXNxjGNmnbw0Y2P1AYUL20kcn4iZVx5qsuqzqRBRy2cAvYlXi8NdaTLEWuHukV5oFRQ22qJj
C1d3iEd6BYfjyAhHF86M6kBgjJPXH91OSlA8kmkgF8ZmuDufC9yUCn25/CJBCPtOKfjuT9w/+SdJ
RHAWq8z3qdcjYklD+/Vi5pJbuw62TmoEjcMG3NoFNFRxc25XyeAGa6yY+OoUMX5F4iEHmPHRevZu
A9HM0ONaVAsN3S1C5bf0emQjEyYWTWNnl8tfOrSWieKni7YGt7U/lf1SZ685BJASLst15Yv8kCar
v+b819aRHCMOso8e+eueRSaHy2SIcp7aFT4fCeq9myH7zuPG98KWnh3xhifdu/ctK/KXZ+GAnS8y
Dne52tH2+1TATmjIvaNJJztE13sEdEiq2SMB3E5L+gLzSf5Fajcfn1xnT91ra47jToTZB5KwF9sf
lJT3Xk56PsOoURU94IH0JYNqus/vFwJiAkwZ1fr5HB4WnTT5NPA8NuSdDnvZBUoKZcG/LjZxMOP1
ah4uHC0ASuhJX/zN9iwoN9LGJaSZIx+bLZ1b3cnS/UK1VgWFRAtC+xvW8xeyggBy2DidetSPqLAc
I/pNReuA6/hV+oHFJXt6iGovSxyrcZNi0gzOc+mA9mqcejF1NLIyL9ZR4IKQ7k47RJvMn+0dAZUa
jGyRqLZvdkDi1PIKVLEQug9uKTwGO4J7GzMYfjhSBnluZ3hQrpI8zNdx40moWW2TetT41cCGVrZ/
kZu1DljAmwG5p/JUxOjHtPjlEqTYFRvbHMQNrHJR8uLg0zxLgCNEAc+YJLqtXNBB0T1mY1Y4e0oQ
du00eB0sD0IC2KT6HjP0JDx1WFUPKxX/H7GojtWqYFryZtf+grrYlilAgs5poIuutApKRHxF19uN
BXyagrv0y0uxdFBkbz0F0uW7x1nNvgoMD43XLAoEhFGeJDeSH8sNbbkO2pCA5rm2i09j3dNRdQwY
wztR1VWJ1DyP/HA6yDMKnrNq4WklXBruBVOxZPY1+dZZWDhQdUGHgk02i1G6ZXC9TRV6J4k4PZuT
PuDLMXSPIVpIQLFLGabLqrcPInPZxOKgKVHPNpoZAfapgmvtqe0Y+thjn6KF4a8y2sSZBaTqC2bP
eEmT1Y8CTudJwAVumOyHUDKpXh5TK6S+mMAupuy7SJE9bQesV+DE66f3Rpr110ienyl6rLsWcQFO
UzmGiHqQn6nrDJzekVE9FXhFP08zl/jAWf/O1M/onlG/QsQcIKuMiL9saZddekLkOJhjWYO/Udhl
0fAHiLpeM1Au+gkgExUiXYI9s1LBIrlW8YZPfZsap+hc/SJGHpoctMScUN2iHVBGPf6GmXkMn0N/
dMeiiv49n98nD8Du2O284nhExKsUYpnqebQlzQQm3UfEkql4FvftSmzu0/Jn8WAxF0vFmgG/zb1l
u03swmKsQjS0189xXumTP8eiANPzQkckzmcvjGx74EqX2+ltYK+rdm4YUVjX+s2SG8HahmIZQf+j
j+Yndx7nggz6j8+ggt8XdRBNCNSdM0P1psz2+o7gX6BVtr7XXyGXI8jzDmMJLzy/+5bQpQt0eHAx
I2nwqgOtuY6bvLSwhAj5dyvFQU3MdijP6i8JG48twwpBwgnnLxAYCkGamk0tWrFRUiVJgAiANqIG
gaMq+At2n5jD+Ora6g+tHrVxSNnzCwq1Mm71LCqqxEd9foP/qPy0ouMeBEoKH/GIIiK6W894eS6B
seACbbUdA5yGRzvO1Z5+OF35b27+muAWHgDFqvxFDh4Zq4KPSyTEsqMwKbVWEy1/tY81QKKoE1Yr
e2J3tuPG6C4QKxc4lWA0vkRaxCROd5HTYi7CNKDxndNB3Uw/7eTysbmaxPoKg+02SNyVA/eC942Q
zewa1V2MIsHHnnwHDdwqgdhV2JVyVFktzBIK+Tl5dWP1aMe2kcuLNBRDA0K5yo0UozBnHv6MzLgH
qTzDw+0agdQdk+iM+EpzF5Gj4PosbMtOc7Xb3FcwmPjBrJg4qxUYqQbUJnnY522d3C1g8n04FCpz
Zj3lWj92TOwrudYNiKN8aI3U+Hwcpt1y5Sb5VtMULogk32MMy5nuZruNOml8NruNTzVlFKvwjif0
wDGO6aR33f2fkcbwL3x1fykd+3yaC8H/WHdNqpBzwdrFWiIPiR1ZAcIz/JZLeHPSsixBsuiomzEy
BxVEhYBCbgBwIKi2y+cELjR7nvko9C54Ya0eIGtkxbc/CZBlPbE/vM2DMVNNnndbs+9DkxkSsVpT
KbfclD6SKPcPgckqV+5021cFKV6HIOpIHAnEq7cUxTeeRE1q7yY5Ave2q/9xFBm1FORmVGQRyRle
zmwnlRgqMMpAEsmCHm2bklYJJEWYySfvLmtnmIY/urm18e3iWBv1ALurxbZR/mRXHx/oIF/tfYTM
uGBfkJOYPbgsWdYRROMQFquQqDoXIXQmfICOj4uG6txMxCgfzy5ZHRgOnwO9oO2uU+KCuLCNb5UF
T/cZuE4FX1d+ltO3vmE2WD6yAFnOwpaSGrMnzs1GTnhhSYY//eDBvWgJtaijjNor2WQefPMhygim
ZQTuiAyHHVFR0dk0i3xh7DP3crEdo5lBtZpjtxlAGX739y3S0vCEjdZ3S/dQTrYzrBRytLxAAvvG
AzbDqPCarHVvxarcYBkKETMQCgI9WLQ3ZVTdt/e2aDg/6Y6v7J7zU+hB7huv6eQ5HJqHurdFuXZH
u+AciHKgR5ronu4vAuNw03oOFuw6CeKb6HtpozLMv1PSxt/EEjD9aaF23cPZAfpjkUvgVImmrvBY
E1BgUiQcSeqvU2RvzC02jIuCLUR1OiKO+jwysSe70mmeeKD2+QwycnAiWlgJZm52OKvycgChnviO
uPGn+gT/rVkxjzsB74wgvKMRXFIi8LMU+x9MWcysAHBivTxK+Dz5//i0VvJHjajydHaF+ryWXY2F
PJepmwPUcaGSABhg82YEqAVDs8+mDmuiWbDy+XCkMqgm46qJN//r8e6ZA8RI/uxwrJwYCAAdS8f/
R/sg7VbKQ8DqLV0vsuU7LNEJc8LOIp5zzD2BnYAlfWE/8SLt3lF0zVc1W/xxaRrPTTsi6SNHxmmV
uezsREnNh6LF+hV3JgtpZzslkX3dKZODNOJGZLiaBlpai/I3QD6EPDHn+lg2AQ/Hnp38v9qrS1MU
lS//K5IKdEIPyVNWfQyFA3hGyjZSuDHaiuZGswImMVKGTwDJp/mWl1F2Ok04kvH9cFURNDsjtuWk
8XViHF6ZxGgAy1nALmL+3xOQ8HDUdBlMhdme8kW5lThPp7jlDrffp5ZmJQ8tguTC+Ula4dMSsRN3
Djt5yMNvyQuAO+MNmBxhkAPz/EDxw+mqLwWUHPDZz088jlcHcwYqDbAECKV4WwV1ZP9evuj8UQRj
uFT3QHn8CoXx7XypTPkNrqVDRwUFECcecymfI1GMOuvhp7/7S6uv2m2+iMRSkf78RTjDEB5jk2zZ
tjRcj2xNHHAatSfDDIldj2QW9BbsueDnF6WMc+AZw/LLcIMdtqK4vHJpdFeQndVloCHUzyuWOpA7
mtgA1t/c+e4eqQL8V2FF16DEZzgehVIUhL70i5mCQcPi8nSry7CnLkVcTkMQK7OI1E1y4DXqIZOg
xYlZF4ZEzQZPTtaodDP52AA8jjvWffr+t76zNxIKGjVDgeUI1CH/M8UCWx9XWBxgNxhhyS5lwoAr
FfdVkpWYNebKoaMZxnqoJvNy4JP3wJBgm+HVIhvaxiNyNgcJQl3TzBQnf7rS/6j/EZ3qPcmlXT7T
87ZE82PACOsAVCKwKybzI4HEI+YZ+Tkgnatnkmu3LAXjIT7itUPziXlYYDz9N1JpJC+0TT89WiM+
pziUMyFpE1XhMNQ6eV8izA75AXfVCtCUTZzg487Dmp8lDMuVvEtn9SPcTFkWT0+v8cAqyLV3nAqi
eblB2Z+sAxnGfL+u9xaDCllMIV5JgCMwBOj7Gms1MmSo2Vl+5D88KTgphcVkqpkfm4rvCqoGoMZZ
apWzlZ7oTG2f/SdVijwqAN9FFzXxp9Ki8Qujiv3zvxsb2eSfvrZIMsPEJCMe/uZEsdIqY8yWkkde
+1VT3jj3w32+yUIjqZ1xfUXpgoKChR6cLYiUBIe7fgfBMTiNbUHgn+PIW7ALBzzVU21glN/W3y31
AGxD1EcExsHBAtvvhl8+P4HXbD1adSu+2HWqY+AAFRrzCYM9UfJo8v/2fpNiIdNxyyW0Y/PxaOHX
qxW2TUjDTHMr9+QESo9iRDmWlQv4KzBma7H2o8VFrL6Gyq8NLncI6P9GxQhUSkK4QLtwvkYZ9ASi
1BSbDBhJGtrN804h8YaQqvo59Y2UA9kHcMoelk0sRjY70YnMu5lRhruiTyz9UG1mlHnx7iqwNZ3V
WZsrCC6SJRaEjYZnsTr+g3YZWVmzCpfnAR83Y1sOFJHKKiEbRU2M9K/gZHGFItXG4mvsNOqNdW8H
daSs6dMvUVTrrq6g7A3avIDV6WOrcQngJ7tFkdSsdxHwlrV7FgmN72W78Gq8qBwkj05x4rFw5eqv
wLQ4a0aVVB2ytaPdMsxNF36GsJeltRs7zY6XMRb+KSFl3/GcKGyykHUMqxMq81kWsrEZd4MUH1dK
kbJWBpUmsPNJadeiIuk1SeV1RUgz4GbvHQhoIW5tBa6hSgtSpn7E1Z+61jV2vn5dNulf3rw+Vzmi
bui/qTd+PpesI37ljhep3cIFJsu7Qm2/Hyygen8I9cw6CUq0lmzkb6ubQxe53ocVUYwqgHnRaSbP
ZDzZ8POUdemh7nPI1975D7isqf5JeBwCkAYSDfYRcLAj/r5UDy8RqE2agncfvNz3/7B+HGj5PKV9
++YqLupiQey9qguvknZCmXPKM/wm6zCAAxQsmj393H3zEjJL9WWPG3EZdZ0L7Hy6ylgJVPNSnBa0
rgXCMf8VrCk8Vo2ko8b/UuRjJcFHGnFGD0Kf/TJ25fm8GzKZmWOmm3SYMYoFPmU0eOVwePTIxLgR
Qn6OuLdzDuFjaCkiUQhE8gMAuYB2e3eHfk+1aJSOp+gG9S80YQ2CH3m56w2xmE3xlPvNm2gfhE25
gUDQ6t5Oq9vRRPfEGt8y0UUrDbC68wnpPdcf+GFn9u8yM6kmCTzzbECCurO6Hi63HW0A5v1gBiyo
6AC3uQtZaT2OXcGp/NfUey8yq9lsAJvhdfQ36qRz1sg2n25dqasqz+XZmisTVO1u1gGWvCp//+Sx
0YV53Unh5lBcqG8y1PdiBF82wIHdj2oDIwIMgbpK3UbkgQjbLLniLEoTCHF2EZVST3aotRiSQt6O
xCoYVTPHq8pyByo5BqNYgFaVdve8Zn4ji2Jq79siuzurRjLIsg6xr/hCCIpti16w6v7RAznLRq1h
j7lWX3P/1unCqDNqFF3+EOWmpCfodUvXfAuexKqr58+dz/0+nunI/CNr3TU+eeZf6OJCO0qyZZ+x
akNMtDXi8Qm56OIRjkXkqbxtD3CT4DX+eEEecf5df5PRNN2xInHuCowBUAbdQmVXaCIYWk/bW7Xz
ZuMNT+3J0zfyVp6//Iu3MqrqjXJuqmuLSKJ3tRlJLjrRQhx9DU66aNe8MirzdyySRTN3119wSuH0
AJ8aV25tRwStfmUi+UfgoPMOo6IFCmzaSZ+GQ+Vemb6v1RZj+4CQUoT9rR5kimxU2bwZQGE50R7R
ddgg5EqT55K6WWw0kCjXkpE5HmB/whvHZhmAFf5vAb2MMdTEmSzfG3yPBnGdJPkUciaq3OAKhVCb
4gc/X0dlBb3xfp3ra8XmFH4fd+jFyHWSyOGZyqtrIzzKp5EimaaZhKJ8cSbuwij1o3Oyd7lobBOc
tQlshoPcFbmdIedji252SLRBOuOkjvDHlW5wciZSZrQ/0fPQpmqZjYS6PYV0C4rHE95BdhmnnXD3
//KR/AT8oxy4HtHJsNoIdO4FaW3RvRayQchpHO2xV5AFOAgyKeqtJcit8R0ABfvjAGjYLCYUp5iX
g9loXC/WeBhbtrHz8WzXP2Kitbo9CKRojEuy9AJH9NHn1dwtCN7JOHs3omV5JxWFg01Ihlrx18Ul
53UIyDmAyI/aNkbEicPLVH0/Wm4NzY/v6jdRcTEyixOmeH5tajQF6C2NzJacpgFgXVmGLJmnA12t
yFPNrb64AgDq+lCOKhHJ10i5rOYUylLmYvXDhC9AOtEBKLL6lWBVu/GvXhkeu3IeWBCiUzVlk/tt
PC6DYXVwLYCvAwANV3I+BFHGtJ1+zG6CoqIBFnoazrGDRCNaSgZbXmKBNQvyZJwb8CNza8kUPx4T
Ctkz7z0WQweXr61Cnddm1e9NUVUohatmLPfFM2Tfka/mqJ2HMRFcsFj9wNinj8QHWAzLsWA43OVZ
VFjEFc05tJ+eTkOY0YZlf/9AjRewRqHIW6AUP/nge6uWwrr8t/amfBeVduRJZJ5V2nnCvq+RK7JJ
0n9yfXdpAptjGBwvzHDHYPIX19yWkdHjSAYIsRjPeFpbrr1+wnyoDBb+Bi3tKNGoM0khOGuyZgx4
8wY4QDRv7sem5xpdOkWnT+7+4puJxqHbAn57mGXfvqPsGGe1YsvRJtREaPeO0ih1IsTfSLsQeE/4
xv589y5TDshWNxErKE4JxA7RNUY0F1Jv3Jkp+ec9BqpTPGmwRy2AmFtAr5Uc8M+eJijty9iBo/IH
4qEqiGsjJ0bcEZZLVtqBc3pFRKbd/3wEXsu/qIl6YhRHUrljH5iHWm6p1KoZOlW6+PsRi5TIIQj0
YAlHVpDAzBHSsmYN+zJhRxu/ntDRgmXkQpU57ICmZjaWx1/brzxf4Z3983i4vgBOCktKO+WC2qVA
HeFqoj+SD+5iH/EA1v/zYzGH414Gl4XXYDDLCU6VADPIAx50rVt1D2pRFg8uz86y1JdxUFLZMG8O
eIj9YNRpEF3X64l8N1kQT3ftBKCafqdHLbOJBd3cmxXmB36CZfCNmFf6VdB2LfjK6d3kqe5AWHu/
4TQb3pJq+LA7xIH0W6Za08LI8Iv4PtzxSzknTSz+cxyCo3SPMqRMDg2hGC0ylOxDzwNrS70aRbnT
L4hfF9liThkwwrgp3gb7GYmTvzQhSXybJ8/DjN+oO0hN4w12hSpuL+ZOeYXsX7l3pBjUmfAo2rDO
yc5U/YHx/Nhehz1V5v2J0ezw90UYnq6FfUPZPjXkwBGFuf/0282MqoDJayj/jsZ8sRbI1v7AQmAk
GXVlcRNS3EAjax0irkuqiSBp1AvXQ+y36ViAjuOMBnsmCIm5ftMP/0xcpTLtldKFSwvD+E+QaLjo
p/Hhx4Yp13UpSBYTJbZiGztrdCaNe+T7HQ4ConRrDmhCYKDKeujwLM9QMyqoEnV6az2Z2QrFsqG7
FIPW3JcbqIfcTWLiHTYdCkimQlQFkyTEJ0tsh9/wOtVztOSBb39cM1D7k3V3VBAK2b66EKh2st9H
mn+7yhFGrhDETC90aBppwtQf0S633Aej1KBh8gz3jBY7gxd94jHcXFC9XzqlQYBkD7IxD/dSR4ZC
lqgMT/YC6LXJLVClAjv8m6SyNQrl2vEeH1xqREpDXtRsFy4c5ZmtMwEWHsQ8bSEkjRY7G3dBgX5S
Vs6Lx0kF4fY1Zc623H53qhzTXvPbnYvYNl36lZIlU4OlG9nBRsUq70ykZ+9ZikOyebjDvCbYcfcg
52Ne5oUEMv2RkyeopA7N1gDAMJEEIv55B5NYPD0/2RlWVUQ8+WoCTOj5620aBJsE9ajt758z3TUB
d0rv04pLrLoQWpLa20Xbo0gnvIGK1MHDoyWbRh2sy7k3BVvXr6THQMbM2Y3IeuCoVGDnIr4ZruSx
fJbXxXssqWRUCdxKY93VJJ4VULwQRANzxVaw52loJWqbPzMbMTMf0rd/E31iB3+T+cvLAl3i2UIw
KqfLPftCKjG/TVdonuF7gCOOK4mdLhYrdHjWdJRWM/TaZcNERKNSHvi4RtS6Iz1MZfxrwVqIyMR3
FjY798mdhWHk8m7wKJHQP/1Hf5pjkLj6fR3USwDiPz0WOKFPCsPFNpxRECIuxaqtR3Iltync07RG
uijMHm1krbJC38hG2J3uo27r9JXrSZ1UHngiNkx6uwxshYl3jv8Cix6LtseNmKQCEl67xm43al3g
C1QVeodUrdJSJmc201IObVtHNYowigdffRN8OlGy800T2EMFkH3NSXrSbvvE6eCNNrPYxhP0qau3
6ylENlIYgajcoMBC/tMGSYl0o8HZbv2HBoRuZDkhvaMuaK9HKMO2PBZZvWUeSl5fCm7ng978ULBX
G5OB6vfTS/g28pX4ks6vHRp+RTTmk4kCkB26Ho0/qi29bzFoBznsf/64dXXY0QqFJZH8lCdmP/uc
wj2qlI7zRmJ2N7nCe5svkk7gDqMMUUQ4IqrGG3ojYySQCTQua+/e2frynxDnvbR3opEOv3RYm7JY
LAHGdyZVDFBur5BRrh/LYhfsRXtIJnzkfTeKGsJcyme2vvuXz6jtwg79U8YbBaowGCCBlo1bwFmF
x0uvJgjZghtFcLmz++98HXVtrDhyWaUCFJ1SCl1IlT7i03r76IfJJ5Eo82uyMRZR8aWaTe5PiJ89
BQCF1PhkBRtcIdIiWRJlaT6oPTCIHK6qi6LPKtPClyGX2EsAkexd7UwPcIkt+vQE5K/GQT3H29dN
TFRdGjGWVnxCEOzUqknxdNbjs4osEtw+jaZLtFHuld0m/JaCq6cH1EeVgvUVSuvhCBuDJ6x5Hqxj
5vWE65CBC6plQ+tKtQCqdIGQHRWzDbGgtkhVixHJCxCURSHiPwZ/iVNHEtdRgoX8Z0byhRz83q/A
jl/+Hin2BoJIAb0pOhErS34tE43vQrci8ottd8jLnzvwqpuP+vunJ7zkpziq+li1BnV+PaFwW0Eb
Vpr/SD9c38oAjSc3MmKJ2atvLka6HY6WD0cyShHjAN0WebRI606ZYVssPEUPJ5Yc8vKI5JWUOqun
n8NR9I0iUZB1huMPXsPC0FqIFvcl0vYKYALgy626ysZ+19w9vS6w1pxfwvd4523ueroqdcjFsJ4J
hlCltue2KA8c361Z8vhgjf81ZM8VrDxrW9akgKvcTyYomiBx2+NEIJZwpJF2lt6pNpGMyslQsr+U
qenuxYBxDlOhlLJWilCZ5UUhYiLVuK+5dH8G7rKQ/SL2mQf/Ui1cdJtGOX6ukh5VWaBaJp2cIl7q
/T9HVa1XgECVl7zNi+3O9Cy/9HK6FJz40/qWVbaAiMihtp28eNd+NzPTI8gg1k6Y3PKylnUtECOz
NNOGdw3MQMv5ZOLG4cZsltpyuiVMdf7ykc4hYBKjS5BuxpwQnB1llynJ7ducanzt62DZ9KOT0/2e
/UH8FH8+2rrTzGO7vtoKp5bIyicXXIMZPl469D4XERsuOgxcEN3qm8BjtJySL/E8FFKtg+dXWJp4
vB0SKPu9CWJy8Y9UtJONBT5nKQDVWNt8GafnSJD64dbwpT03dRLCkqrciugYRkgAP7HVLe2p0HZO
MkaDTFP6SFhE2E2mRxHAWku9Gobv7V0j9NTORePsbxo/ldFe8ZAdurObHnoA4jRWWxNm2tGOGxNo
sqv0prrNsi2Qubg7jnv9qinlAGljyiioUN3Qp1GTtjm5aS9C3hzhNkiPDzfjS3CgljM9RqGXh7xi
nEn7T7kRByINGhzL95wxYjU8evQsuGGE56ncV25eUlEezmRaiGzpBzV5KXQ8hMQN4kFb1x82sIP/
sjXc0vG9wn+Lc/2D6V+N5v8GGHBhgOJVY+L9ug+mED7aBwPbVH4dx3twNgfqcydBGb78W9tMOWEC
DPURLsfsVlHARo4Jd9ovtuhdec4Z+JUmb7Ahyv3GCbzA99UrYUCIw7bybG6htscug9tb8t2r6LB+
2QWgtPra3gZibmGUCWfGLoykTUuJxAFJk9hWYbfM5zz7Jr+7yX34vTEen1pLjSCuob4mDzsZDQ6t
hauyTIj4IohhGxFHn6v+q+XGiNGamKd1cfn1wRahYXXTzXESFRyESEs3nBgMcp52FUneMzb4DG0E
ak6aM7b81QuzIJEhHNjEX3eCVCRd4F0cZt6nLrNtSvOQ0rnhM+Yype/J4OlQWUmaPAZvBjCpvzNe
jPt8R4Qxu3YMaSpgSflViF+6orIu38avONl44GZewfzdPHo1YHJga3qO7UkGfLvLKTdPwaJk8xn0
30OS9z/fKAWg2qUgAYmIjUeFqePv7XbIMbJZXuuvi9NkHGaSZywC4inF90DvkXIG9uuWvcxA1baA
RxA5+OWQRMeUysoW9kRGi8NTEl2D9XJRtPw5y31iwzGYI+k1YeIQhaK0SWpfnkP5rGo3Dzo1kC1R
5SujWjVBSrs8Ob9Y6qlAhCbD5fb6awL4PKakdgmal7dTFFkswxM+isoVniJdAtgQ3+T37Dk3AntA
FRraA0YaHkKLR3DM2RN6WXk4U2VnztJVhEUw+BjxS1z6t/GciHhpJEse6Lc3wWl6xrZoiXKSQOp/
il+jwXVnfBrMH+fxuF8ih07RcGI20JGuTGVUgXuS4BuRttK6ffUUKx2nZCNJD+lPya2uCam0ES2L
fz2dbihS+32GUePza9V8JqTRdF+oUri1mckN+SJOvM1An8C9iQJcZHiLJBn6mEoc9pV0N6Njcdl6
2JezS0uvQuRsea5lEodLVH+1fD5w8C/TdshQP9G+X7cRR9ugBZhpQXjinFagfBI6vt5OuFkSiD2f
qew4amiDiT2aegU7g7BO7bUA1bj90d72LlNpa+d2ehx1KXvi8l6KlYar8tuv8copGmhc7XhWzUif
cVNJXzBKAu8nWnREEAU+YxPTHlf/t3j5er+MVEBZ6xv2fFbXazs1diit/00TIZ86M3Hn0nWIMpmi
m2ON3oD9p9aR3TbXoQhPL+e2c31DIwBy1c0CNTWI1AAzmt1CHoC1KHQGu907i+y+OIt3nt/Cj3X8
VtzmdwDe8fV4ZFsDiIRJqYXrhRicyVIWOyhjxn9Qmbpmx2ixWZAl3DDQKPyvXv3CC7wisMNJ1tLT
ggMZJCPgbath+3F0HrlPLYq+oc8V1JE7+mnF7by9hOPApbBsf3QQbbMEi3obqDd2ruSWoGzZZ1tB
CnTr/tmxKsXkpAUCy23c42IzVDzIRPxYqigFKeLaNC/bDjGRMRHhq7ov79S3RdwneuUug+MrVOuZ
SJP4hJm0LKclCcWqnDzM50BSdoJj4WSWw/MNrDVZRERjIvYuLC74a9GuPJ0NDC45zO1N9mXdWnU2
6myk4eyUosjgTlbX+vST1Jq5OqRLvdEQTGdaQSvOdyBx10/KzAD2jkBAr2wFBAW23DAORMq8pTHx
D4xVY7j2bP0LingRHL4FYIAUMAbvedcmFbiCeYQ8p6CYEgnCsUD63m9Q0cXT0vpxFNW88r2PhpZq
fah4CEK//G9oweBoelaqeK/lrl8kbQsmJiKc/m/IYSazHAlW6aAnFylW2W16bH+JdzKPF7Yn7hqE
35cBojC9hITWmNrYK8YIzac8+sF1oYxvueX+69zybEPjLpJb5XIjLQqi9x0VD9QELTUnnQcVkvZ+
NBg5AZH8+mnCkuc07/S37YgSEnZGcpM2uOBIM8BGa5k6wKlD26IY59AfjqVFmGFgqmjxcVm87Yv/
00hExg7JApJobpJkYbiJahQZhl4rKKhwlRL4eStBIC/UOxKPVoDQF6KKxSzZtu/16MP5DS8XAjMj
WDCR3L/B0KHrHpKUSk6h70sgGJvRjyNAMhUI4rOCIzLnqLlV45POPS83hhnGsGyTPyF+lTJBXvXd
tZ2LZxTWVVV0Nx4V1zBjCzY33xpLRN/XR03Iy8kaBwzhd7udKe5oAYQ83fgSEZyMW6QIMoo+PNMC
gqacKyrxvQgFGt1EcdOTmRV968ZjPUamF+wuEW3J4KdM393WVs5ZWFZYCCDcrLUsrp1/z1yFided
cI0YNQ3AmxLTJVqK4ZjLqJACc7a3l720J66Px6x8Y260aKYy9W1CReBq/DshWIMcHMNbhpicdfT4
5GqL2/VrBIz1TwKuAuDqe0XIznVjOYc5E1g/JC5mHgA3RsPYKWswfsnvvZg+zFwWAu28MXkY6pYq
PUJ5bRhX5touU7K42phVpympY0C2HaR/xo1DCcJnTmichPwTO9RctAM9iXQQgMD6/gjmBe9Wx4hS
UGwHvJNNrW4L9LfL+0qultecnVZTBC+Po/CZiPFv40+hhUbN+KBAGF7RiTdmTnsVFDtvyJsWHjNk
FIj+Rgks1Hey4p7GvPBEU14ekg8dZ/CEy9pJmeuaup6kmod4Em2J3LHMkMpntuArO/P/wfkNDJjg
94O85Bxs4nYEFPWhIPujcOX9wKrwsE0WwtOeeo2WXRlKO6p21ScTlW+esFcILLG4OIHyGb+TF5Ik
+pX/VAsqqYQjbqNq98AXz2YMMLO+GEkboImZ0Aapsqktv0/0BiT7sU2UteHatOzK8hEk8aZX5AFq
szOUl0OCPu+p3NKVb+I65yELrisN8s56K5sQSo7A5HhtjP1Vsba6yybM77D30F5Y5me6+kSmDWOk
WwPEPXqWtD4I2O0hI7bYUQtTO8k4VuoS6gocshp4zzZXzs1jLQmRNUfYjmQM4+j80aemxasXjG8B
X40LfwiPOmDyudvCzkyTd4o81LU6sBBYwO1jbh4mxUaZ6vWjNaZhudPJmW2ZyEMxiL1Fnh4zKs0o
uWsiJNF+PfsyBx3rlWbpSl4BUP8CkfbSvp2CBbJmJpmMo/VUDl8+O9gOH80DBrcD7HTd36golNPU
mbcD0CznT/+sXIrZbP4anIZUhtZ5wK5B7oA/4r3RXgRC08A+l/P+LuG3/tYdhW27OnEecEtj0hcV
Y+i6lemqNAyfD0nURHc/0li71AJ2GW1ucyYXcaxR5ZQ4b2tb69Q8r2/gl7O93prwBPddsfvieCbJ
8wdR3gaEwRuFYQeu9jLlQjOtqKqYhU2JpQzPNNPwM3LaGWsOoX+cv5buj7TWZNvuaDA02E6SCm4d
YFJeGe7cStm5RonCTLeLcOWz86QKkxZDwsXB3w/kxLoX57F0uT+dMDusjyV4LLP8VVBuCSaIFcdI
GW9aKg5XCAqpN1QGIHHVAYHQ02DPoD16aedVYPJL/KwvCLM/CA4/XPxbFqk0OqACAct7+d9FdG3a
zh4554wxg/kMObBQbglYMPaV3Yy5yWatc6xs+V04K9y9Z3uTTtQoUaHYVg1RQGA45umXwxx7sm3i
sAHTYD8MFWY7+a10oadhKcwX6QHaZs8kxNKff0BKv/pSm7zS8YuFFDYRF7fR2AwEqRbMCmRgx0pc
YBvpWwVoPPFeeKRBZNLbjoCYYjQRrBWn3Hnnqsc0X4WRhnL3Qpyastnng1wldeFYxEhQ0HDAlOBC
DIdKIgC+uj6P+bgAkmNlrm+plJfer8ROH8j4es9LR62XPLPBExQQanB5csKYLRI2JdJdSYnEF9fX
pMMXrEujbkBEfp3gmznBct9d/z5Q75PXDt47N54Y48dT1B8efWE6LH9vwlkT58HnMJPE6CjG7Wr9
xcyWEQYh+PWDmRK3zXGsBRDkqtL3FxJ0a9wiDlmmo0m1Cd1E5fS5DI4DS0Tc/GNnnOAo0YxspvMo
krm/UZxHjXXTAlUR97c79tZC73Z/8jgkVApfUI/GYgb5MTExvLHcoZOjW4Hr5QcNwAKXLOKzeAS7
cJ1g1c7nniQtL+RbuEeyiwZOgLbooRyvWYj5NaMj7u44oqEAPxJyT5njIKLSjWRh0fqovND2ne3A
AeegWvMTaoaMisQssFPnqUfjl3lS3Ra3xxsT/Ey44ycUyGBNUu2XtXpZ7sqFOHcitxJ1aJ1cny6J
Iz1i3VnEmoFEXghUF+7S7ISxy2p+8WGkbbfNvUbmJ/J+r5slx0PtGHghwbgRwRZ1cCWqWZTziHrB
/6NDzVSa6dkfFWA2uwm8Y3sa1GA7wAEquc96rnHu4qoVadSQnCqSHqQf03SWCz8F4z4es2vW3Szr
eYJsTHTG0OXjygR4b9v04Wn3DtKJs8DUj0FxumgYNy/VXm8n03CZF+8UJbYxs9Q5ZuW7I/9kwbDf
jQzwRW6R1RUAmzTK4eHOkL28Tkz1sBmcde4cRiDD5nhNr8DH7Cu4Cv8dhfQF8Jkxqwx+oxe4OsdZ
JSeCDGv6T3M3J3yXJc0HCX9GjXdRK2YXN92olTt/402b+nSlA+mONQV+Su6DzDZLMSge2tAlcEpc
izzozOTL2SQoE6afqERwTzNOqGpLTCanIXQ3QC8JsLzWR7+edMlSMbIdFvXJu5SUqFlfyhzqv4ln
SAcNfZ2NFiXLRgVJNTX6niBJrdbEMIQYUhLjyLUATnUCqveZGSmP8tCYQTx3v8oUTkP5wxwbTgTP
zYf5kb8AXQTY60yOXwLrEdFFHs0zWxR4ScilWqIGKf93QDxyoZ+2nKpvWeUYJx+lfPhp9YwFDvTo
wXNvv8C4Sb4kbrGIAQAc6fSgQwCI3Q1Bx4jATB1FH7lEgBvvGUSKpwLhzxeMTYDmQRsNwq989IP3
12WGWh+/B2+R0wL2BXBCIg2OhOUdQv/xOhnyhifGahuQPJG0pixGtKVPJX3VLGe71ZoCSndnc349
GDdByUAPc34ZPHtz3ztOh4fDxB0idQUmDz0EtIVqtgfAzBXWxGHA+MhDBoKTg+4Ns0G7ASlEpy4x
+SPg3MDhUr5vxgjYLWFwxA9jSAAGyQRi6SMEvdi7SXymmLUxYRXqfiaqYevRhJ26+Wmjgt1GbnzE
ugT6YOj+Hd5YUM+gOLTiGtXOQ4/pCg+ceErqAFYH3qL/Dh1lqPyiwVhWf0aNK0KCiE7pxDaE+YQX
BrKc8+cnWDyLMxtx0Sj/dt+TMR9EJrLOmudw42yM534XQiyxqCInWrf+mseIrnxdlH5oTrSO9oKY
/xoX2CLh6p9vGI4eIBgN44qLporwKaGtrufGHjvTtVt0zfmJvCYDUMvThbytevK4PmWROuB9Crt4
CbeY893x9NzkwTi3epjUUivd9iPXfEbi4V6czyJStwRFXwSK5cO9jh3+E1Mn1i1WW+catY7GQMXt
AocR6s3eGG/b0ZeB7cEtgEgWXNBlCr3yEebwMAWEpbKsCZyqFAheOmMijP7hZGbZcTllpGtBh5BJ
k4FdivEOA3krlXS+Lzvtw83SBhZqdj7tfEPgYnKu3VgoagNBqk8amn6dN+REfHXwMxl2YR3I4Tej
2dmSY2R7LGFAVBxsIh0QcF/BS13Xu1MchobW0GGNBtwRf7PzgTNjsWJmsokbOf8f+Ou4L3A9b+Q0
fyBfRgkbLmou8oGPt3Vrs/QLGqj57b6do2l7UBvAk50TfKkX1ibIv6XqqcNWO3jR4LOhlO96v+v5
wzJXXH47rFvrhrfJ1F26YNmkLbBi41y8nPl1O0JZXacuKF6Og4wLsM/Lh0VbUCe4Z0xzbqEISQS2
4Fbdb1x+qRh/f7BXgHTyWoLiy8PjgVoKDeo1hM2lPbyGZcZAWi+sW5pmuc9s2nhgejFJ7xlJRfpK
0w1SecU5q+G4BOKGTTFhbuJ5IUc46S28LwG3VytykC+nFd24SC7vtqogOdraef8d4AWAYeleX30b
U+DvUdCYAETfzBcinkKaFoZ3zjzBytxeraCue5XTpZB2LYOCYQ9Vw0qIkgTnQTWdfEZVoZmgwtW5
VG1n9YVqS9/sBH8l9axIeFgQ8ft3fPwo714omLw+453PP9JQKNZ5xvVuqHSzIikj3LoKiSJqUdyI
dOzyNy65V9YLwC+B7naOpTdaJfVHpgPQ8k+f8YefNvIr+Ofzds9IiWR5npVlS34bDUaEfvfMb+rl
1hhBY4spEu4bOd8mc8RYX2hj9xeEobI2vww0S+uSVmoCL0TseYkOPOadvJMutcKdR4ICktX6hslo
cn5H0qE5nxwphYqqReE4pWP2WLL2Ji34FWGvrnN8djCoZrKNvg5eIWYiU1B8N6ojd2W00vNQeFbn
9UtgBB3uY5WIgvkMgoZcq2TiagHO4jPaizZwkp22HvuOKj0oEdQ1/jgFlJ6rcFKOmA7I/KSaRymV
1Em2T3S671/ruTmmzLxjKgh8plLbdfMH1dcjNlhtVZJNksSX8Z0aRr64Y2Nq9OaD3kbP3wDyxk0O
8PPlCBc2gWqKt/Ty05en5jN5DrqPQXZIzwrXAu6MzwZAuXGR8rSiK4ATuxftlAgMt4J9hY7PWB7B
RA+E4aISGZWOSKSYHvZ0ftB2F3JxY3R3vmpJOlwlgpD9GQITZjfx7oPiNu0mr5CyaZFnw6K+0NCg
ho5HioOdmF1eLYK0uAokFwM0AN9l75Tu+3elACbhpef8c8JjMELrvWQi4c6yCkG2ptUQ7pnUSn8M
j578Bfm92zYVMI8UUM5Itx2L5nAURk2V1ndYdEd3fyseM1d9IpTqCg/9jS25xfluBaZLOpVyvNU1
m1rbh5n+/zjUto+c0VvexrUpfn7ZZsfx945dcO5ALo+fM1kJl206rUR2pO+Boy/RbICAwlNoFTxx
3TAafsIPjPLiY2HzPACKaWuHStODLd3dT/KndGSkYG+u8o5TOOYf/FKc3mYp+igz5VQUBJEkt84N
e1x4JZuLgw/VLRQdX8wMrVw5cnqUEUMNC1wgWyiVVWBUpFzUQcKHIAOaPFTsbDzHUaQ53sdUhW/+
gw9uDNW3cRaVOOidf864HLYa29Rurijz3L2TINEZXjTBiR7dy4T3Liw1CfZocsAghoOtbtRjT3VA
u4ZYP1HGjg9xd2EXxB4rxFiHZgXGnt+DhwFhoCrDUg+F7gSHMT/Nda0am2N+9K0un1A+kcEJ8NH2
OkeTkglLG+4fHOIJfnLLFhxLrKXLQXmBegJD55e+70WHakLqSAv2WKNM5B32lkjXrFgGBMNYPPzp
PiQseAJ30HObxympjF0UL1CdisfY53cttBJ8pA/+EXJBayYpfBa3Axx2pSuiwr6z2Gr+/Ezzza5r
eKxYvqz071RPw+xj7Am9N8Pw5Ff7yRPenfCccBMM5eym0vyCCTb0Dm/PvBoDs1aNXbPv+63THMRK
ZlAjHH2a6lAvXQM5+UwHxUHWTt7rdU9PX5lfhKbtDmRgkizyNDIQ87FpfgVFJ9NyWr5WIfJb5xAI
nTUvOtEjfO84FzbRwM51qDM7/OF+rTmU5tyCQctTPSLLZ/X+QDAYG8OJ1LooNkLxNCd+62OFkIKE
dUP3mGCQPFa4wpNrs61owTX0P+K54P005nQ6YXAsv8TdgunApS1Rmj8ERHUTt5Vc7z+mf9Qwrk9t
t/TmtCvVBo8IllnQ/7394fDgtC52PFj9EPlSZw4vpFgToPTKddpKCWp/2A7A3yXK+11Oq5sqLdb8
fZJ/2x8WNn6DyQzDXaL2w28cu6c9M5gePGXrb7Q1kYBvJilLP2votn3FnyXUU6IzhnnXeybF9yNY
A3Sfp1vEHJFMswKEEy0pZR4fAQxLUJc9Qb9rd15wyUUawEHf22BpwW0csc2plc9JZCEfAJ9STS7a
lnkVP/uOfOlnr36uJRS47zpH89RPiaLCO/feiRskutWBpGB3ZuX11qJLP2Ud5XV+b6SKkfhLvr4d
0j8ZXbvbfR0VCXp9YmVUJ0gYsoMdu+PgS25x3K3mWBr+vNRK9zSTXl12aj3IaDbT23WY4uUhothp
fET91ZPMoDp+8leGu9g9A96pqtZZh5W927cwrOGx08alf9hYT0R4+AYbcfDKA2NFimrL10k6O/wy
oPw5ygr7Uw7e6AhyjhfscRiK39PkzYQcG7IXF/L19hmAE5cd+zxtJp4mtnPEuzAlNL4vAgB4FZcm
Ap2TnRXhnWLJqxuZMEGvTUiiwRerOydoSvzTcwkdiTpIzxu2fd4dYTBiyXBxTSdnCDETemmqk3tY
nDuOM/K39cf6IYzPRZBaY8+1grUT75Tnb1RZCC5glM/+7sDT1nVD/PM/Nc35h4Adc1GaOdxajkOH
8sp4pWEZFpynlpfi3lKvXQxvwt4PSm7o8O6yNY2eyAiK8uBm6TvmCT4JExUCRpj7+aBMLRRfL008
Xl7bpov2sGapikVp69i/6zSdHaXtBKYRLCjLwoN7b33nYCard8FlJFgglM5tKy4Ej4+lCeWvgzgr
h7O2yzPaaWxqECSpQ1i/rbFYOEsor0mXYKhKPdbYIqjMJCixqbejzjQl/BuTOIywA9oORZ1pHEs5
FjUIiQ1sWglhHuMGQ9mMeEwdRc9LUk8Lfw/FmYhRdJmDgicb9YI0K77sNA0zn0fsbUyewA3B0je7
J2lwXtB0JIJhcRkTsI0rW+2PRT8SQurxLcW8JVgY4TEJ8bstDu4+9+OqyKPqn99RIjjB+XLCudbF
SSUASZ0wC5b0H0ALEqB/06n//cs6DJwtWqxFa5THkPNkSKrVWvI0XednsRa++JAluR9V+hlVFQGz
FnV7a9oGF2D5EudM1krWclSToEdGIpGurH35pb89o5bP+NJH//sRMsVIYZFVv0jRDy51Ab3/jUYU
65Q5KLufReLXM+A4jkd1D9WN0E9IP/3+LmOEWH5WUoWLrsin9TESsb95x3fokEBPSXV3GK1kMXPM
CXPAWJxEFe+WyQF8zo9Ti6QhzNDkhHcX69tSM8GLaudFVr5bhhHI8XN+6exoPcRZ1x72BOTp7ydA
WFn0tscfbbGHGrFWniLS88us2FkZaxmk+9gvEaYXoLTwnHdkB4Y4jJ4AmsqR+LFsF3+Uzkudafng
0qRJHHo4hBZoUMr6bM0vAbNWgMhVy4hIvXlWDzySK/0Z/Ya/ixjRjTFPO+02u0/ONLRbt2a3QcKC
uZ23m/RJ7OkRV3E5de/BhvsE7xTmKEo2F89kKXrObtsiae1u1z5eKL+0VrZHDE1BbI+pe0Bfgv0f
ZRN4zEAtappaN0c1P84JBWb50a6BKnY/tZpO64AcQjgMiWhptv6XYXo4DmpYHTOcuv2wXkjbQA6s
SLFwyiJephJn678kHxyTQuN1X7bccAVgU3uGLwb/nSzFxdOd2u2g/cDq2Eslvf6JD516wgbfStml
X2BYnGqkDHax5sV1+Gb8rnQ486Fi5e9VRNJLypcIwNP8MAqZimYKzsdLBlufqjTkt3MUFvoeNAID
tdtIGEaWhh+QYArPZHDA1cYmBnyF4d3snLGMwgbZNG1yRK/OxB6zDPw0ejM8TPGp8oatak9vBKwv
06lQkObC8nHflh0s2MG+rHjHJJXDYqutb+ZB7UbPl6eje0svaOJeNnQn2qBDOwvAYeqLQ2n2Tqs0
XBAiPsF9IxDDejZOKdOl4/8OsW3edkf8QGcYyq5oUTqGgG765u8Lo2sgyB6go0BZ4nlGxrUs1HaH
GmzxhbR71joiHe9w4MrqiO+EeO/P+B7AMbeRBfywllTypkbo4WnO96c5I2aEmRM9s3ZGH9kF0MN1
nCtaiBeJCtC4gCAbklN9Y1rweeEFHTbqdWGwEkdVBLHVw6MELDaM/saiMBcUX4G8JhmVa/m07TeQ
Gddgvb+y7ZvcwS5bDR1O9D1FEcwjTfwxSUVgHKzC3zNDAMkKljiIsXUTVqkFNz6G9QExbucYwhf+
bcSeBos7e8BbwIpNZ3KjdaXdtp/QscuKrFZ7oe3M9uYlpzf9xLGL/+kRSoY9d3LT/qTXstX1khll
9VNzMgQMD2MOIFMEk4E2rXNANUvDC9J6WIA9RntZgQU+zLbRB9eR4nVScb5udrhTeONMHB6O3wSN
Mi3UIStN1KBGbckC5NHpNlSmsKg4hIck/tp6AR8Hs9C0lXYgsn4rY8PpMEdXYtdumjgefS869KeB
Nx/I7WHrA3KP0y/OK2sWLS4a6nfZi6urd6XLg2GMlELQ054uq+0P5CODLVh7QWHXrc1SBvDNVgfe
BWYZRqglE+cVrnD8pDJntqGa5rngXwDgNfozq4wsvUXnPiJzZ7BRq64XZQLo7+5KnMcp9ublKr5N
nkjJQK0eMXfawH/p9fM4mTWWUF3vAqEe6nrRF2Bb/DtCrrUibljZIAojMQ8RQLIIHzktGHyXMxAW
VFw8oFuALq8BNYxYgRpA9QXfHWcjHKO8VwRkh5bZlxAUDFjxhLxRFM1h0h5m9QZR8XDFMCM4vSz+
RsVTeT4vtWPMtxGjnYeHQQBxuH5qf5xxlGVeljNiLwGr+SdTOb3xd4Ze+2SBVXdgcDnOCeDZRGQs
P1aJRfkVWaO4vvm7i3I/3K4E5O5jSZIeNm86SNGgzVMCsH1Cpinjy/JwnKWovMExYYmwNem4njRP
VsFYs0LsTC1w5LPs56oTrjt2O5wsmAate2GrvpXLmgb5F1m3MsEZ/PzyRuilk4sYmrUPxIS5P/6N
MsJKLlVTbFA69eY28aW26AcQvp4x3LnfzyaBugNur4SWUyZBXfxO3P81ofa+z/diTxnZ2Xryy4yt
jx7A65dwCw9ixILkku/p2U1A+muftAQL+337WH98kpoke9ZLj5TECaqu00qbj4dT82ODOKvcXb/r
qfM6RDssFzJfpQKUccIDfByIyhNB4VHBVMgjkTJt804BP95T18N3basRTthgC/uCAWANnv0dfARa
j2ecDt20uSQ/qnFqOFRHUPOTYCWBwZDsmxcBQA4lwjtMmrNoResOqa7YKdwNqCLX69RbX153yLJr
CgVLu5bkk8bZ3piHFcpMJTBWZsEr0zeluKTeMxD5p1gfZpUcRqwkSF/xiTQmVMenlNJc7N3otIZB
TA09Oqq/FxSVTHo21NpADSPtgMbqDXjqZ33DZvFoIeE50whPYsLrHyrl0a45Fhnmmsk38uj6PSm4
fg+WGD2nXo0FyeRZr28xBklFCrqOThQv492dqC73Ykz+yno3tYpN2TBAh4KxowdQEZ1k4uuaRE4N
etS0TieMAIQENJvmp018i2ONSrFQ/c7c35oCrhUGqoDKMqtoOVn8klwKy/Lll9ep7riBP0eCMT+u
eJZGjREWrrWGdKae8soQ2ZWBnHXs8TItUCvZkBbAS7JYKCmEROPBMcUTNqYBgvXcoh0VEZwwAtWY
/a5dtHlUSoLZi0G5ObCrSMfc0oJ3G0xQJIecQpHu+oEZhtHN1RF1X23UbRBR1TuH9nW9Z4z6iKo4
PDa7o20dRFp+owym6nN1EBIRRzNf9vxCbe63VXos6QziOhVK7gPBMjks1FhDQ2vwnqgk6CE00wS7
xFnx5aBL9RH8BLg1r3X9DxebY5g5pK+QkmLWXd7A+q+WykxjDBqOet+v3KSZTvcjH5Cax24OveTw
8wEtZIGU9fkVMaz429II29ZuN2Ns2AVY8TNhyUju5QRVkmVuRfJ0v4KTHj6FR/aXhNowL28Evjfh
h26nryFI00ZEdM/YsGt18mAmnhZZgsUNLpMIckvUhDMLdKIIa2BoUbQN3ZsphzcgxCMY2CwnmEAO
QLeIZk89S1xBB5lR1Cy3twKXaBnmMg9KgE3/oz6KPxmp65jlmKXAYApDBec0A/ue004lK3PGV8AA
Y/qtTpd9onF5mf4KtdtuLiuSTEbZeBtB6DeynUgONHlNukNTIvoSHG49uqP7LIBBx92DxI6GTmSs
mrbMuw81GCJVQg/hQYp/flKH+/Pvet0/HJP+l1buqwmU1dHeav0PGGriJiKYQxHIkACe0ZccaocU
zEQFGxNnF4x4c9bS7FUDy0GbYWGcCzd6TKGVrcbypVdTnrELfJ6i1V1ucv5E+yjI8W7QdH8sZYF3
DMoxPLRABNreSdtNrOBvmojK3FCVG6dwu/xe8iNdmsI9tiAVuxA97bGaHQ+VRM0SbZX7rUqDY0dl
eo/R14eY+6vsqLzjMVZiqbn0uN51VlkojhHA+/K3YuzPuCkasXckpNuV3r7UTlEh5Why2m3O5Era
nNFF5ipAGRv3ryw3gxtVYSTnQAJdm6EJtlTK1ewYYARqVkFUkvp4FI1ayW3ettEUv6gsc9TWFhE+
aPRfQoXreD1rjOPKt+xjGRMhGaWZQMWgZn1/ZcA8EJlD2fWtVnfs9GPkDZzsqQZHkVkWR6pQYEiC
Cl4XPGG0an2g+fklzHF565JwIYZPLcbRJfoyvvqdI0vKQFsczNf/w93Shh51nCnuPeqXxFuLOTCE
DtLBVI+b7D0kROFuLOS9Sblw2FWeblIZo3kiaixMQ34vnOOh9jM5iPlJrZWfNQMWLREgmwQzkj81
ps6J9duKR9oUhQUOmOZEYpgIk4qWnXBLYNsqeCaaJ0tQwg7UeOLmBhVANuYmkqXANNQ8S8/p7xVH
FWQA9CM/VLeLZW0kifKs5YKgTIi/PnFaLuuEO8vZ5UENB18bSFq368wOMXBhpuSA4F+vBUkYyaVh
YV+eR2FxCKbvu0n3HF2vS3JTkeBGYwNn4k3pcKaj3cKHnPQX9I6Bi/kbeQhffzkaV3CvKbuZMnVe
PfQFQLZy4WHqRbx+OfEqIhDzlGYDELevGtZkGW9jdU+w28fTqy4A/WrzPnD4skOuECDi9jIN2O8Q
QlcIVTDdrUxp1zJLOJ9RgogPd7zjytAMNmNmMXo1ap9QPzmIA7HyapBhyElKU9qdNPtktFsF+4pM
sKppFV2EkPPMbTIS5OZXwo8m3KpiiJNDoXtimDhxMChOCY5pfotxfj+474nvFgJ1ESYpAs2lDBcy
Jcg+fCspnLjRm6x5iLtGO7LcfKXH6k6kkyCbBLjkcTKOKrnU4WKaJ4Id3kRkGTRD/dLi6sVbiCko
DsrluBPFQhBAtY9vp1+Kcv+6p0caYNvYX0S4w8yA9JjmECWQXXPISTsfapoTYbY/vh+mjHYYBsf9
ELx5xkw6bek8LNL16LuxqiJONIkOa0PAIVUBP7+5mr8HZOwavUe9XKCP4grZMy6YZzotM8exTDZj
aJZiF9CNUTVMbmVtVVxmQeYzE45tPWy2uZGKe/srZKOvIcYfeeyKjwUOkxboikfBKUz8cnarwxvF
CU8E4A7Joyl9UTa1/qJ8+oln+HpYuTx2q4cSAvUgEarC+FaOPZ3B3wqt50e49X4ir/94iLUFRfOU
qlArjJyg02HQymunOdmzApJLKuqPJOVy+E1UesWkSFxDvy4F7Jy5Rc5yeBWESkFgiOhbUqmXD/hL
qmM71qtV2HEABr4qVHBo0fPN8bT2YnRMRBWEL/lU86IZWqzkUoRMAgCaK5TMJObWs5z9yyDiQacF
VDoJeAyJGPUFCQ4z7CiCA8efdadtPf27sJbP/w3JE9L9y2TXutalPATaPTVhuN0EUIRSk8Er48ch
1C1MT7U23aOYeKv1WRYzIjNXffq9QQQw/U2gFYEaL1UFoHpH+uAA3he5+jDwr0llAFGQwAmC+sC0
n3KV+XDrP6nacrYZU8jDK18z0Fq4k5JLCSvgRpB8BvQ5KU7gStLwtuKp+nCu0u4L0JJeC2GbAZy4
AHg+JCWfs503h/tx4y/ZL9Tqu3fNR89wjHzOAQ+03qTjtKaCgZWQby1Tsb77htW2+pSNqoEAkUOq
zjxcr/qvpXryTN00BC4qIfMW6lv7wZKVKjANWGjreHuoZM4qvC19b2ppHvZvY6R+R/HNy9EeFF3y
5Ec8tIaSkHDAKxnq3PP5mkfV6hby7fcW1aYkc24DDSeh7RG6UlqMFJ2W3g/yxkVGePw8o8XEHsS1
aOSYPYDcByVjKfa7CZ35z80OnBTWDkoP9xtUWU2VKNpCU8AB8gAJdYm5U54XD3BD4ft58txb/kSP
l0LGDbIqLpmkxpjjp6LrmwELJtbpwTMphhWI8tgZ5ODnUOBP1rYrBHd5QIjfjXO6s65v6iFEc8VA
r65QTWuXTfRCF4x2/3kj6S2xc6SC4b9CuRIR1QvjBEqhnVKt6TwNY/gJ4/qmeyxAmXpste03c6QK
JvfSCFroDiS7/Q8edWwXFcJagr3hK4jHd2H5oiKnNQWW06XO0OSL930AQ9mYi+GJYCXozc+XQ0Yk
4b7xGPkscd1a1Zdoq07VGL6KZNixg1HPR2HtiQzs+1rCUJKI5pSJPReXExkKkBjPNN8UTN+D/SaZ
zyxE7flVw1Sslh7NIrgqGop3sZauXTCpk6aFO8kaOyU9OtDz9Mv4purLsITyTLIPs89Nqg8PtOYo
7xFP5VNWjQLQjHscR+VyA66F0XXuvAmArf7F4SRshJp9Rxb2S6i8jNqWeSIi8614eyHfTPkt44kK
kw98zmEylNyiatSFrmtrlknEMRyhn+Er0DfvCO+Eaz9QrAivVUpedoLgXL9XERL6wTGVa9b33MKC
6bus4wSpXRr/pS5PlObVauPP8EOiOVMXujLJ/FuVVd8m/Stpd4C7Dg66jCfEAm6gd339+rt5MK8g
gNNlpilY7zUdJ2oyj6ajT0hvcC75x/7+0C+oiqWHkXGbOwn5PXtwoceHR+Ew5a2GJX6XqsSy4ksb
9kx/doRJzQeaFSTPhfI7FSsBWvk8/YBImyjh1LOiF4D+cw2nV7+ZIMm1tBxB1XPW0vALJPwl+RPW
lp4DSj9ij7GdC/eeNAcIqwra/NErgRpNIxu1Lf7csqmsJIWCSPx3pTNvy5UfOC4Jc61EQdV5v5A/
GM5wq6ruudMWVq/dONX+tGUhg6fZSuYO+09lmQKL1sS0/VcxqoIeprrenPp5XQDZvBwU0GvEu6K0
mkT3oMl5TSdc+Kb7G+lbr6tPabgm0Xz5zgKjFkNZW/c7xABxaSeiLeat4JR4sgcl91ZMKhIFM2v0
WYeG9cWboOlUPT0GNLH+aMqU2U7UBzqjL8h05hqNE1ISEX7dNhKsXRKku60T83Ze7ocmwApx26eb
GlTI6RjjA/zBgw7PBctzn2E1fdoKgUvr/wuCb8MJqNuPXP7vw0hfHfnCqm/wBOLEENyjGRZfEW3v
8BErK05kooWN6f0rtMtqnZW41j0KzZvRYZcYvaFaVuj+Csp6LO6ObFxkbgVLkQTFdXq5TOSbKD11
dTcIg2Q8wQiX4ZIwEn9yM/ljNAsbNcltd2sbsPIe7Gutxp8uFm/f1IHAwOLSPypwzSX2YeF6JCMO
lL+YcddPHehtZaJRYUq26W+eCrggP9mO5tV9mneDntmXs75cp3bw/p4JYaJxu6a1ysemEsyJFRFq
hN0ZSRGqvzy4nqFh/NCIsQ9Dm+D7yxfM+qEUNCMcyfOjC9E+tGOC07c12dzsxKu9y6kTBb6MGbYu
UgQlMwgq2jozpZME+7CKvrrFm8P9T37Ed2VpmNtLA29+l5xNzAnu1a6Vf7srloK/085nxbqMsN/e
HiOSEmCR3YEB5ax1v0eXpRpJ7r0jgajlb3ANeZW/4VbPlr0upmzbsJHwNuBYjkjH+s0C7CGjfoNE
7BLVBA+xHMZ2j4955lid9JkwAd3EKS666rGdsmDq1hGfvLMja861fd4T2y8ltEUu3DqC1B0szAXv
qA+FTleLIKCakCOyfJ0vgVFANFTOpJ3r7E7NWPzC8cRLALbogJhBnhGLM7r32klHD+Ai6OUOjw/U
YYTgZNBxoQDRK8z/2nL7zsENyWiVsxAL3wgYjfpS86quMMRyO/NVIWLIjzrcvFmk+2OltR/2Qxj7
kRd3+YeNC4McLXd4qmGjNvRqzNzERvs76C6+/P8M+25I6V/Z/2PbctfSSBUhVt6RqprOaeyyIhYW
NHYt1RLhAZ0jQ/Vqn/fw5Xhwze7AYi+bG7FuN/h5j/HPrxxAB2zZIJlxA/yyXtjr4vq9I7m9AUqc
Yr/ZwIy2Z9pFMBT5K19zTdurKr2utWfiyxDhfiAN+SD85epAm2zGL5qvi+hsMUgCRb5ErBGHcBDl
6jAfchForPUZEQ2xMDnzO61SZ1Sr9a19aOxiuEr+XwqzvzsnqPlPLVZvacV2cVQX0csh2IZOtpa7
PFgwi4jj9fcjPIyo79t610sGfIJJiMUP8WKJQ7II9ia4AEFrxZ+eYzUqZi1AYUrKK28v7QrEsGdb
lMV/Ac2RFlCTklEchZDtwe1d6xTVGwosUSpEgrQ2YsGGX86nBIMHdYSUuIDsn3c60n7g1F0MJNEX
xQ+er3CMMwe+gqg6PNgviS9PCKmjTh/rhuSsH1+KqEgo6ElAdP5FnuO1xVACZA0NTa3YQbGVWocD
ZfH8+lJghW/vp4pQYhTWg80G5NDe6OzOwpJ2mOeJaqQQM+P1b4DO2pPW1yMaI12TobuWOpD/4c3x
1uEsjBO4l8FU1RKg7zp1aQrPMqxT7W/BJnQ36fCCSqb2elkIqMEH/TxaJe1BsZXgCmLc9+Oy0ksd
g1D73znTfgNs/KoKF3AUwX9gFLXOYmkpH9mVHG6VcOFaf/RnIbsp2C1K4r6cvUMUJXpaxk0wuYU7
dHcFKo8gbePYECVPNnasr6EXGjzLTEzYvs9NK4hpLyAtdBqlhapKG53X1y88c+KxCo+0NLriiY0m
bTBNnFNcIlS6Iu6gL7Mn1tduOV2VBrHNbqf/iIWgIVyNjCcb5H1uoyttxwnLXnpmTyQHfYxr7IkU
NEhsYYTlpDrjDxw940YMJT8KimPFGkOK2ZRy3sqeHT+jSd/nNVxzvg3uioe8w33dCF0phlq6NzbC
kMNn3+RkSI2V2DjPLtbunRDVtyNARl5H6qsfuB7mZxreMjXyPI34V/Doq6PqCCt5kVy6kgfjg2Kv
Sope9bFH1XLtabdrSclLPyXiidLEcW9sMJ55KMRbPnaEm006oNzeLBdsi7OSWWLxl0qRU6499sre
CCFLGCAaZNLfNf38xSS5/OGpNlhKXouwdM7Nv9hgfHfHA7qidNgXBBWPLTFVmX1KI0Zt6f8jBd8A
APFunRZF+GSeXoZ91o2joEj3dYPp9JgWYWjBC0HF4/PvQMt0JQHvAm/YJNQz09yKIKZ2EuabdL4t
oTzUSaKPmF8bQbM3l+NzOWdf9zwwxoo6obw71gPuEwLpeXM+zBZXzB4RuSTGhYiGEEto+XKGVgCG
A7sNa0a3ISinuvsK3JWVkKUXrFkYadbEFNMIm37F6ETGGRvalUIF4lx74zeMqC1howsV9hwcaZTS
j+Mv0VRyfymBLWYkVX5HZ+xICbDxsaSO0yc/oQwYHCP/7aiRhKKopWcNKKIporxLA/5DGdQlyPse
bp2BkxVfKATw1fPty67CS31x1tMIQklo9fEmuA6B/HYtj/JixBqBL3P5hAUMrgJnZQOGcf6c4VJV
ymqN6NtFf9wYtTBq5MMnZZC/udOHyqLa5w1nBSbiVgeby5JDVv4wKVJYl7BrftBRtndFvZQJpaIo
a9lvMMAjBKlx0qfFZ5LyVNgQPNjMkvxhR7oruJmPcyAb9OgVIBzJTpF9s70sqBAD3ScAf60FhGQO
pjOVWj4r2FO0IfomWiVqk85sgyEbkjBxQ8pxc2rBxRw5EdmwDtghMN0dpGmtn9gJKkPs3XeobzzK
jJbGn0glnLw/GZK2zREHxx+nkiFbrzBqVYnU9RRqU6lYxD4HmYGltA3fB19JxEGLJq7zsNpme4/u
+M3ylFf7ERyY9G5t7783cBQDO112LBzaXySMW+RgFAeYviFrUgS2OfaB1I7iDVyz9DCKQ8hUqots
oN4o+EzXL9p+jl1L8tKA9HOiYn251gM+FawWinXu9DnelSNlfeFk5v2Y8OeBttKHwsT3BV72evnu
xmN33p2d1u6SaCB3g9K6ejz3lNgezdQ4Wt3IZXQx4ouYX7m/f1HQ457VQbdcQIPFxs1hxU6RlY4A
mtQILyrMMaMQua8hbsme5hZjbCqWljlzGjUsMvdEoKaOVIggOlKx1LhQQbXwj9v5bd8BU56B+vph
3Lsli7BiGeKXedctsu4CV/A688OSvjoVaHz8U39H6NMWNfTmjNW5Kj0rgwzdV0JIZA9wJ4wesw2w
VQhgDyXvSkXgu761Wl2tZ5ZpEZXZnIQJLr3PtoBiZf1VnrFp6k4prL2RvOgorGRF4bxTOxu2E2Mz
WEMQ8M+sga7VfirN7GEbodufPo+XTuZPml1qKA6Et1OIk8j+jAtt8e/Eo7EpyjTtPZOP0ndrW0JD
RyGCxG8uonsChkwHtYu6VH2vxTXZ3GkdZg7bbHHDsp3fOHGAKHS4M/p0dhaye5/wHyo/pzzOFm9W
U6uKrKRh+J5aMDvRNSw7ovBet50+rI6c8UdYBNRQN/EXRmyDpiUFtRqexh8YNfXzt8p+h7PPTHRx
wqWDjrXGHmqNB8EDEx/Kf09KENNJOEvDjOwuY7XEGwWlI/qNo0J53eOVgk9DQt8QnnLaxFQ6IT+Z
7N4wXYvHeW4ydwvi9SRxlvcGm1O4gvHacuScgpYbr8CayaJuS7kQKGoX5xVu1UkMM8dLJBr0AJgm
YKtkId6StxyXd6Nd+U3FkEuTcWuH3o9qZ0S77XqnYninB+YytCEpV6sHXsquM3QgtyANR+EICi+E
zDwh0SP6GdMdA1pr9iMFUAJzoM1COz1hYG+nIS8F5YLvgiF3evLaZreMZqy74qCOQAFQXIvK9015
qREeJsWJe8fxeXn4r5vy95RZion7rOo5tPn4is1bfzQBF+xpdvS74YVlnlA5wSCjllF4re/+OOIo
A5vCstx8KtNm/Ic9SulAYB0dhVaCOQ5syPZdfHiMkxGuPGaGER8wI53lqJNeuFwJDiMrCo9r1U0m
ENkjYDreUWpPnGWJeRiE1EjbtlMxTqP0LZLjO1/pClizXJe5zWGJpHEawYQ0b4MhgQqsw44gPKkX
S6hJYq/Yyfk/9hbJCUuz31fbQAn+4AeZJ+NmR26zPUGd9bELJZ8K5wi6Uoae0rniLAhGIpp9yZAH
13U7XmQUsHH7o8X1YFeCGRM+358yykaCEQg3d9+1509LlHsvTN4kGDWcIv8T1XiuWolLj7KpYRBp
EKGEvVlFWXLCqkubo6nATJ/Zf3p+wqvXOi7JOmQhYFCQYMMVOgsv56OuoZP/iqfjHBwMb7qo38E1
MrXJq48YyH660LtaYkwDkNdqfZYgZAxo0NZaWl1REPoNBucM/TJ3FgqRr/mNRpjqU6lA1y8TlMPQ
En5Q+sYnLO1ZfmwUIIt0dCrYaaCaM67g917ssYzBmzJSjHV5/pPntKYKb0hcQkah9+NFyS0G68cU
77G58QbH2pq5fkPlHWDSzyx2RBU8U1zfQNlVr1M/YXsKQuG7X3rko2YnEsV+FV9eOMFfbUdho1D4
zzs1bLmg6oKNNkA7d3XkXsBMorLns5YpiUGhu/81zXPR/6X4byMEoGSi20jbKftW49u6jlpDrv9Z
CZhZFUKCts9wWw1NRtkSHrHnEbuVO9cxjFDK7hZKMhdVcyng49W1O0mySTZEl9tdXVPv19M6gK22
fBXl1K3Fc0pZ7A/Gqd4xKNvPlM4Mu9Oqbrjo+mnYFrWg10pKfZ/9xlAaja5hCatMDmTuea4Ad1E5
THzWBZJlCD97Dd/yCYVLVoQgu+6FE6CH/wFEpmDBTuair1+M9n9U54ur0z48TwklI7jATmWVzvcm
44XkTbfVgT0DwWbvlv0D9Xjn7uy5GwRSe7rkaSnreZz3UU28SD+LRP2zmpX0mfuXEomKGplUm7f2
o25PCFuwiFie9ndc19n+yIZkgSL3gSfB2jLF5Z2NQ9hjtJIkKAiTfZYp38nLC3hejOcP+gk5CliF
44csfJbvdHonrDgp4OdBGe3Iho3VDzRAdooYqNRVllHeJUw8d1uIo3UFQrGlOoAkVQBi4rf4Jw5Y
VaFC0rhtuPUbQpbinpDZSYVkzfNneUy9scA/UCJ54EqJRLyfXkfVstOcT257zB+G73T6L+YgOcEs
OqJ95H5j8cLJpwvXxgxPnIvQ25MxMpyziDGdgIbU5tIwRrGdB9KBheVpo0BAR2Ea8wymIXVRfHJm
fmMPyHfjaRxGW4V7ALrViFWsuK7VBOi6UU9Pmogki/F46U1Ohhpvr3WeT/T22V3d7Z09n7lVTfXp
7IAVrB6HidFlMQrKZ1YYKRJ/x4CDl98x2uwGu9Y022JJfZHHWxIqAUljUWCR2EXBC3YSAtAs9T3b
d328dGCunf94YlF/Yk89aTdf8CAOw57+iad3ob3aa3Ago5iV0MoRbpEmnwkqR9lZpdCNEmu0sHQG
/EkcC6QK3x8bBr8GZclI01aAdxdNc1izBSYEx/3fNwxEg07fEZFEr7nYP6YLpAijj3M18ucz8cEf
n5xtrTHgOofd7a6dVyILygfwXHi/Cn7CsrC41jZCOhRxaYrPgQvWX0qH9nuOOoTCbZZq/yMth1vY
PmuzZAZO+nYuXDzWBzpN3c/YDf2aB1oybUZE5avvfS+xKwfUqifmyzIaMPyZJ/a9cHMo6ZoQ5X02
vgUxnFZly73phfvyiozXei0XhEph48AZxfY41lnx8nezAesEeQ7qfGfqXvP+AmjVm1vzdVTTP85d
30eJ1RzjLXveB13xFoh7TmuhTDtJqsLeUVzrAId8azBEz07fhlIulj7xgp9LfKWW/4mlMnXi5Nq/
/PYfmnsSh4nfA+q8tRSGFYmi10kM91dQBj6/VHWUYLLLbHLbZffOiaKpLYV5+zkr3spY+7j76nye
04FXwpPoENoKUK6TH2gAjoCpdgNVXbA4PkzQ02VDnLodLW8/DT5apEm+dtm/tb++6O7qHja8+tuq
lHv2wgsBB77KJCNHykZjl2bRdEteFf/cLi4RPJMcZ061F6L/9m6u0HXfczh6HEavFXYnIuuShYM+
3Wozp76ieaRIP4llmjSy06DeDOl4A2R8hnNWG8TRZLfE5Qph2GMA1KZHu4fDzjpPImrNjWgGndQ5
iHj1uEeQv3tEzy8FB9rAKk6Zu0Ng2Xc2yIDAol4tIj3cVEkm3S/GwuK7EmuPHXmyvhvyf2vSW+MR
JmqOLlv2tY/lDATEL53VmgYXNGdNDZhk75fiGYXwghd6J/PdCoJUFmi9N+Lp7O0cDlDpdUpW4lWl
dkL3cwUX1Mw6YYRe/SCkFPJGIoDue2MlyETzCWIlU2acUGRmykLrk8Kizurcqh18fi0PcLdKcFhg
O0Rtllhbs5jxkxpVF80lgkGMXLy/4gwBFF6Bb31WYxv1gEUSRPC/ty7GayqY6ps4CjYsuzbQE17m
mjn0H0gys8KEAvys8xF7/Yy3EcjgO0lbteJdFykQ+8u1VR0JpS49vmfsyDwVOYhfYFoZdjaNwW+U
XqGqYy+BHVUcPrf9cMjO+roDzDXiOXpIRXPXlFUFCXKyEBWi/hA/hYsNap5TdO/7ThH8T+N+NrMc
J1FdQJzI3U2f6Py0/0t5XDl+7TLL03jPrJdpmeFv0CSe0mVPHOfmx3ttTMOPVMUskjvehZuotHCS
JuZB4nd4cFElbE5w0Qq7+yvJ3H3VFmLkVhY19bedhXOhk0qdYqLHE8r3ZhFXxNrwyglu5GF7l3KI
4a1olfOOlOjS2Om1OOOZoqAOx5e00HRQDcN0PvuRQunIYZbhJLUVpl3y/RloXQsYKLhnyQosNkML
UHL/NMfgw4zFkDrD2hVbo+iji+gPI4QWbXl9QMV+yVtWoadfDF4zbhUSX0m2fmUbfpWp9mmtq8kI
OjzTc/Q6mbjteAq087adqSpNxJx2hBWwwXPkn5/bqHTqZ4s0PbtwdkDN52sSWAVUv5r5nWjVRppy
9v5TiCUUL4vDLkMU3JaeKG1GhfpWmPWMFJND+rJepiyOcTK4cpVZ+XUi8HUx0mVRZy0SdwMwfJiU
29FkdNJkqZL+WELPxbGG9F7IzZfhIkxBJOcgQ3RKumG7v/f5bgdMYADEka8f44nUxWl9s7n6Ic1g
jSADn1RrA8jpstZzh5YyPIAMKw7xVJ9f4pVc7p5/DJ8deMgkrp5NJEvPsgRWv3X/13NS099OSL0C
fatXJE38vqHdeEsrM1HalyzGXVVpixlCTAFkDmkaAtJnHQp/KoRGdnNO2JHE0c5swJuSYKAb2eFY
mVMEyLpAQcfpkFABlBqH0D3t7R9X6CSo5WmN4W4n939mZb8Ra5mN0zJ42w72k+EhOuzuy48SGxzJ
iafXt78PLrqlIXZiiI+5BuuNyi+ody9aorrOJiysSTcDQenVYMq3bTL0ce75mxA27tfueZ7OmbZ3
wjF6NDM+o4hwCPkuI3K/z/8uf2pgG5SbACQ6OvhhXZApzyS+NDsAVh51vpibj3fvW2D2n9rjpFSR
Ez1fu84DHEFJuW489OmjQr7ziwcAZ+eogUqys9wX2Bpj122FXmvg5XzTi6hzgi6G8LD5oieQqPMb
zVeMmrpXN25FsMH5C9YG0VWYxke7mbfGzp3tlPL4WMFggkXdYREWKAmo4wsnwwWxj6PtD9cSyTqJ
yJokYpF13tFE5d6GPw7NHJgmU4JP9b80XofrZBvXBg8Y8JzXvmgURnZzVaY+aw7HDOaZ6rA+/oBP
pQkn/izQEc2mGaH3gbO8hr4e/iYTIebzPhY2JQKEIEHQeVj1sJaV7FlGnu+NeiE6FneG4NrkmKac
2u/GsVu0XafekwgpTcjNmjZzmN1zTLQTFn9GjX4hrFZRjcc0v58rmi9wmAgB9svKiw/K4EnPHp79
EAZWWizbpTHqmvuDUf89DDvkSgIiKGY+zhw1XCrZn6dym6bGFvVb32XsQyP5O8QtbU8h8BQC6dpi
2CpaSfo/ByJ8tCxuD3DdyEuT0myHc2sibjHoGSqwWpGAisUw1oZOfW6H7fGBdBku/ud8lu6p8PgD
E5ublFLZN9WGeTYXOOi5hiGf3nBfMxDf0YYdW8ytMawSH2wPmrjhrMcQ965Kh0d1lpXIywtr/SvM
JH4B0VykPnD/vZ3i1dfJaadIpKzpGc5AoD6Y6knffUDZ+UKXfdUVah+u87SbD7lxczY359d5OoD/
1aujzxCtEeCxYiPkDWBks7W40BuLP/aiGsqKRzgVSmzquY/a4hBbunFgZjmIwh2+uxcgNMdvQH/U
JOxmKnmniEIYkAXlnLtuCGPCVAth6X/7Yqkm7/q2Wdpwi4s+8iLibA3B5/G24CfXn+UvnoMZVGrw
Fe5vZBsrohkKwWssw4zcpTwztWEer3YFJbcVSIpAy5FBUv6g8qn65qzf7Y8S0iM8CAnjKkOri5MW
VuVM7x6bgcVk0YgqFDhcer6LduYFM/rQUyLmzxupS33Dn7irqF8B914cqZIyTbd0WpAZay95sODL
hPX9eBd+1HBazkLaEyn4U3o6R0goULrJ3xe1WIcwENm1FlTyh5UJozvkSvfg3y5grF4zmfP8FtJP
Cb5L5+0FQBRbcioFmb3cLGQkANKdOsS1rGAAbt7a86HdVv8UZfqzKWYjkc2MBkxOo/kuyxKVi6bG
Kxc6uIcR1uI1KfWG4z+shsFUM2CgIv5snJINUlbnk5PPOMA3Z8PR591WVGBzkRd66Sb+N+oMHU+S
/219MNPja+AKqANXSwtVzc7Aqw7SZRprjRqFhQYD9XkBfV/f1uzVz9vaOaYe3wu0kseZwTpt5Kpf
LYXLLkt9cHpjHlK3U8aOgCklWvDN/X8U6ose9p/GjpL5RpWEq9ckVI2jwQeOnU/Ixry8Rzd9+I+l
KuoP7TqVoJpbXQM8iC+SoVVSfL7Al1F4xOs3kGgIcl8/dy4qt2blymCxQ2eMV374u7AZ6YSrBdwC
IRcCrjcf5NlZXGgyCZC9um9gR2JkEooKdStzyADz/JyArL/8ziwWiBdS1ZVh4S2oRq+3Q1RrjN1f
igSIVe6JP2jiV3lIojHViD0hs4IoZko/u7iR3CFA/V2wKeWyWjlKBn/+OkQC/BlzSuR2V1xgNlmW
YuUovOV+x2Kj9vQZ8BWCEJ0YkhiGA2ZhNqFX3KFtvZiIF+sKuydzQ8fDuRhS2pONHKi4AAn8KVWl
vFN0KZg19x+MZgWJ/iUySVYNJPWGjKYcaaAGhM0Q5OJnMFtBSd/4WtA5OLKpMM5mhJH2UUhWqQTC
ygvRD/W0DHHCDfwho5BXQSmBVp4833eBszTSDxzxQMJxq9Z/r3guzljnqkKHkdppOI9ZYl7xAMaj
4nQtR/RZlMSgU5RwC1QutTJEie3OFt6kssp+uuK4FZR+xIbUBj4x8QsVfFe4EWnNUyQQJ/acULOZ
NNHkXpk+H1YLl52O9kF4xbZg+6V0Npcl6blHQ8HcvALtJagGe64fpMeZygVb+l9clow7sniO3zEn
OVVboOIZnf3E50UIWgRV0ZLC1S06tdeVWtxnRx9LNO2FtHlNVsPpNBtuOc+mB91UNvMYUU4G255V
UYtrCaeYPwxE+RuLdhPJyl815f+58QuOVJ0mGeqZdIm7XNS9xB4RuX3JXT3EJHim9emMTidfv0LQ
vBORXGsEeiYDzVkbkjS/Jv9MDpfthtiB8PsKpSWvVTSIluKK3YOTiALTvbJCIY4+zB/fuXqmSnQ/
mYtNWyOVpzL7YafEkti3uwxLqMYpgVn5f3u1ycrGp7ie0jzQa2j05AC0GlFevofMrge88pGN/vpT
C7itUys4aNbs8VVoDknPmQRg7BsORz+FGzjGpGD1Mkx6Yexj3m6vFHL1pe1fssTNi4fglLIrJapz
FrzWFkh0yu18YOyZ2o5waQkx0EZpFAZOLl2mHO9AMDDWBKcTcSIG3B8Tchux5Gcp83VY0OEMgq9I
9gTvrJUGMJsciDO+QWxndWdDnhmLABy8AJQGHNQel29s86x/NhzUHfmdCl3i/zydWPUY0Zd8Afev
1NVmV9oV09AuDAFA9Rmr+rQS+UAjtlxsj4ImBBkL9PUvGJ7AAJIqdmIaoRKDROrf8DFKD2KbGNPE
E5RXBPssUxDo2zJg/LRivnS/yM4mvxRC3vxHG7fcp9S0uqnxfuo1MwoGFeA8jiBgkdB2FfqufGXj
hC4Ke4T+MHd+P2XvPr62pkcCj2GrjUzPgiNzDx8qmfPQljyYoj//F0LJZ/BQl0BGDIB8kwdRmjhK
1nTiGfcRz1eS79OKssEXY7jgTfteCEQ9UxxxmTU+5cIMAHrHRGP9kwsTXVarfkFkusycEvDoQr0l
cXq5pXmdjoVFEhavaxXjh35J24zNCJ0UnFJWQnJXU4Rq9xz/5Jk1CufsBJMtS8lCr81xV+j7NvGk
UfPLpCdVSTAMR8hUNdehVaZlY2OAdcxJwNkRiZyxSpCX1s4VTVUx7ObWGtGloJlZIr1VeMt39Eq4
SRFo0WvsHSY7ujC9IXIq8pUGEc6EMPCBo/KWPEtxZt/me3H4XHuGJNKdo6Gxe6PjI00kr/200K92
azXPyemtwjQFbk2EeH8xnSjJ52hewOUDf31f14s1/Vi8dHoeW8Z4oLUiueqHfLdA3tab2KLa8bTS
ARKdNjTkhDbNEk2QpKyd6CjSK04r7t66GtNQiqlS3JtI0m07ELq74fcRo7la6APTgr1At6GBvUQ9
ze1dA6YvuCv8dIH/VjxhmHOguiJelzwnzfPTCMAlEr5t6p2Pt1JvE1aLB2mvOggbdhHlcczH3TvP
I7xubbQKIyViNTb8Evkr8XeeQCpYBpFQNRWrzqAy1j5ksIOw/K0l+tz+C1pRw6PQ/32y76dq2SRO
nc1YHcmt7ImczIavqJ33OIz4XC9ywzAji6al7nk5OMd+0VAnRWi4UP+a55iHnuavtfhPwtm1CJDH
gpLtF/OxVVNaUXLEOKIKLDoxjwQF2Py2DlUwnvPM5eSdcIA/4yIAl0Hc1GMVqaVBXwbzlng9R/TR
1CmdM2Xk/DFHbBdlXo9WabEez3AbwyjMBjUbIEaFk5VUC8H45qJarDYNqUCVq7nXimM/rYdof0+e
AmW65krp/HjwCAl5gPKnahYkQKyllTe8amLE+JM2fwBwvM4RhJparuR/tSn/Z/Xw65HK7bnhEibh
QQ8AphEvkBThR1eDSrQAlUwTjPYvNT5FkI7vRe0wUmcDhM+PtCaMubu7AySbJfu7R+KNKVq9FtAG
pAIqZSiTm1Qc7EQOp5wUYEIUmzrOYGvwgsUdJeH/H2rarwMXtaiSf3WRvXns5y7g2q9QsqZewVfA
bXS5aqSE3sTD222QzAZptIFT5V8XkTBh+MKdgeM5DVZwc3JUQXwWOb1BpEIvfm23mG61NiH44LJr
EDZUryg93TybeXTI/mjwNkI1fiZS64KOHS99Dcg72la6nHBZMEcoj/RWsDyJfmaBgpx2gaozvVny
/RSKkpRMX6qUNn4tfVh0IfRSBDQBWgvz6BDZKVW9pXvqGzOXWefarkV8Yzylju7Fz384kYUBC4in
7qHrUDzpOYBPXB78hafyVdF7yeMZeeRG2V73RCoEvfMXc/8Uzfn2ZXaBuR8dajhDjwrJqO+pSy0A
wNKA0OHeHQ2WujE8rC0r28UFrmQsTysBrIfpdqMiyGSTApMcBVjoe1wQ6vZP8OKNjaKmbkMqKDTV
MOsQdFP1IUyvUNvjquQ85lN5xamJyQ2grWTKcxgGF0ZGMX5mmGyXTzsgRn06YTMoG7qSTcxm51Pj
4dxDDL3z0Ztg6CHWK+pO8N1YOB6ocwO1TE1dzNGzXgPs+Dp/HH5YQIWBVjZKGDAwNWc2V/DzGrv1
SqyZJXEBT4uez/0KPyNBALSJSUwS4RYgVALVcuswywRQ9Xh8zbDvuipcyDcRu9F63UpJvcx1KwIU
zxvMXK2y0MwVC96nYvDhaNwbsku/tnVkCPA9E1RYqijGlMO68EQ6Ex6/va0nQGHm3cQIfFKJtKW2
GD0Bhd9iKGWqSElPln1PaT8yR8J3GMxrSV4CkTaq2g2PevuHaMlcvlg0IlLZYrfMCLwDf+jnpkM3
6r2aAKHqiX7C/5dffuKPVHe9FI0hHP/rz4vw5L0WwT7CBI21kgi66fMiwoxoEp/t7jKX4HB3xJl3
h6hxQPnNgqM/IQMOQFi+fxQY7LNJ0dtsaoP5B1SNGM5LvgRKXu5VEbILL5/gioF7IeymbKbDoXzv
WnrmgWbvZDYd4j6ylSNYriXmgwSZsvkRQ1g0tIq770SR5yioi4YxWoEaYFWL2PUnxQc9bn+hmue9
OhjBZurGx3Gi6IGU/V0JJJ9LSLgWplVsmL+L8PVVK1K2hc3A6HkTtaRgSvhp9Y8s3jbRTWwW7WcV
kpv0CT9yCMnYv3zOvLOQcrtDFwQbQH4vA7x/iUbVGFN/sQ4Hr9FGBRfH0xDnfjJwiPH05NqE7YQe
76ik5TaT++pwObwUEBQUNUEUjOGUtphaDTRUeqIm9IekB+7ValYHXLa/NWDGpHnX8xmiSVZik7Zg
PUK+l4liwV+gk/IXa17wTVqkymfuDfvJMEQDm8ksxQoSEL9c4tjMt8GXWGs0YdGpR7bVcGmUC5F6
ED7LtMJdjPddpP4piJuzGL+x+Wp0RSpkwOWv+khItWE8hxs6MFTYBo2TUimdS8JILVdT8ZeRUfqr
g23cTpgjZWpg9d14PIg7U2BDUvincodAFwePI7tbMhjB1o5mt/QoEqnfpidL7Y2cYn6h3wJ8IF4D
t+XszMPGTWkLSGNHH6mWC6iKai1vBxxdSKyg3EOYXqiJQjNctO9BmoJJ+e/vq0263CVf3ViN5EtE
UeN1S217B/zFYZcrd3cZzsCaq3hjbMOUprdBxUMgg3VpmD+G/D37LX6N9/7ffzUDniYXbnShv7o4
ziAbW1esrJtKoVUo7I6DRnFVk+UaB6gHnYh4X/PFz/gqraXk+2fEaFm96a3JwQEGcLa+52yyh7ij
2o78hvSthIcCFfuZadu4/FgGGBIFmPW3okIdiXb2gWGPnuOh5Uq611uyRPrv2owlhbajgcqeEJWU
Ub1yutQZCTdz27jodrYsftAYKDn0QKQ8x9amNlC9USW7im9/Fn6LDRqpGhZ6SK5MHger3EUb/O8s
uuslBDF7apJUYt/lcBFQzuwdPVKCbKN/1+ZltRlUx0cAVXgXyBga2jDIp4AHc7h4WEp5E784C+hh
sjQBuUHM+VqkwjqM3Zx19OR8pOUJxZBVSuH03rLCkP0YDtSeASSfxpPXdtoMmSz0cojifcXBZf8G
X+eerq6dkGpZaJfpg0vIyCgTZloNxnelWNHnjudgcffx/ktvxcPdSgfwTtEhhogreYceDK6QLIh0
0Vm/hxsgLyYJwQsg1oH/Ttf28Ja4zFB6p9bztw+8GQ4fAcWNmFa1dEclanq4u7+PGgPXb2BMPIcp
0JY54y8YE1G5Twsh5VedS3fcXnP0Wf3k74Uv8oFHE5igVI35E/c3Lkt+ucO5DC1pImgy5zXTLM9V
0Im0/VCwLwcv3o0yEYMMJhY8WfjNlJ/xNpvtLYA/RQ1akuwcqHOuZtIhimiqGsHUmA7rxricCeic
yoYdXPu5sIWyLjgt6EcLVCHf/FxbPPKfbZx6omX6MobwNxFkH+xRkK3FsDPECuID1cbLdTSWLgrb
rb0Fteg1JIdIqLAOei4wM1MrG9+lX9X2vwlUrgFdVueRkC68Z+lh1MdrKRNfkT2tHdZRw7qi1svh
BDKN22W7zvsg94kxtD9R2tjlznW1UXc14M/Q+k3CzGSFsH1F1vTKg6ekxPTUEbZigB+lBbhTMV6+
9ll52/Nv+TJ2rAgogSYtb+xgch7THqSXYYDAgFHpbSBlHK3XsaavKvMz0KNBWMQSkbwK6XChnz3r
go+rsUE9I2FjuYmkgJXNavbR4AFOP1wn/Qql1Sd/1xZ4CwEpZG2bKdiEvYQQKe0PdJgcDfNl45kY
lfEamJgOPgs/WUmJMTh3vfspAGILHf/P1wo/3Yu27VExTQNz/n7xKtMu6LMtERMwpKEEJBM09Kj8
UnBxD7euZtOolPcc/TQ+NFMK2gdCbM4MQeJ53PpG15fALhYWAxRkw/IO1kV0K60JyKfAJrLV8CjA
wjMiWoeXxXKt0oth9nCwCwLT5ggMEzCuUbZZk1nItbbdhyBYRXeuONGSH2dFfjR2ZZ7hEYwMrQi8
kcrOazAueov1DwQCadZBvM8XuBSVSoV3JX164LkGrA6/Wfa9pM1o+hwSNKAe1RNOmbGq+kCADAnt
QnZnH3tIFeSdKTwH8LpcdLZx7IwIrQjUynsGzhxiAyREv/4STmH7w4Abp52rOKjWnorS2heNk8Tq
Vy87B25Fi/bHk0VSJH0shRValVi/ZFm3W28JlZ2T10e/MNzc/7L9ByKQEa453j/WWRNeTbjtTwZK
88MRvzpGkaNtRSubdEQkcx1+CV7dqN+w+PDKJJoWbAfVKVxG0SCTkJgiA4C17gkSSp7pYVITLdEq
gU60WQrOwAvTXlybnl/k1tZ/kiK1PEqaJoUBUN4m8wO2MPUhlq81qliOgrrq1x0ihXykxPolK8xR
mLKHk3FVa6JCVrrR7ngImxIe2LmdoDN2vwXW5d+t2hrkcXE9iLmfeVgWi1GK0STPsxSSc3Y3dy5+
C8c1R7vAp3DgO9Opd03pHWZ2yepMgKq8ovnW7cmu6o05lnk1Joy7rBiLxPIWPKJ1PTZLtDkj2ju4
3t8DOYqSWGD4L+VV7JZV3rTqYzfxLh6NqjMHlKV17i7rQlKI3jOZeQXDv/51oNaVzurDpI2FqvXj
BAEp7IYnC9WWrMFeLWB4aiM1laEs6Z8yX4ThKxIJ1ipaNRbAnS8JfYaKBwvSLO1eFbG2TGfD+dJw
l0jSYyMzT53QxNBUanwdUi0xtoyCe/xTXsH8nS+zSP9uW6UvLRvivgpulWrZjO0IMonwwdGwJ7XN
q/qEZFYQFETYj86gmUK9+lAF3fZbn9Za+rLY3HTxF/Cy1Hr7hZqqKWeTymz8kq3EY2p/jo2UcUl1
gW4PWP4MsYNBYeilSWs5T093qgrJqSGboeyqv5qUU02Fl3It2Zt+3IBUG21U9BHsKPc9quj/pQZT
Hh94v82pq+JaOH/cjU6RhadJiMpI3XVBvFRWdlOO/izH3S9weUNRF53Xzkafqnoh9UyCJtwMN1ui
FtfqNh09uYBHTRN1r8WtzOJCLGQDgru7FnQrp0V/X2J/DTph2NWPwqv0K+3Hr1SkAzswvSMrkJou
yQFz4RJEM3Kx5r/JGQI3llU/WflxvP/4ZFOfUNlY3DNJRKjOlEqp9BPMrE2yuFhdeJZu7iOmx5VZ
kpY96t5geg8uyOTHHtwVZxo1GqwW76RfXu2aLq3LWPuezhr2HvTHQ3qcc3Tz+z5NCGLpe821USop
rchSC9ULk05BqfFBK51EHCk1g1pBZrxlvI1iYFWomacnMsoJtgw5qEO2xcl/sqY4sXocXjAPuB1O
Ql2qwLL5l4lKhHpFE9bNcNyIzJ8TAIws6/RarLgmLhHdr9znLyb3Pja0+9gWwWS5C7UbPNG5l45W
WXg6cIAHKtzx84pWE0M31inOFTjc16RTOv/J6GeNwdiJEFTf60T6guY6iERjKQcgv40x5hCC/nHk
OAQ6Hkhll+xt2MjjwYRTwXcl3u4SvCC467gAKKO+6c3JCAlbvG/uy8GNY37jEeCHbaKE5qK8DpRl
M/gwlKymOz0ohm93WV9waLdFNS/sYBPakVFOtxROeWx1gUZz721rWXLZXJxHzKeNsVHSSzvJigsZ
fBnmdqErB2iKwDz4iOWGK4gslClmiN6RRkMk33HiA+ndQXBq4Hzyeq2MK4AHKdXuZj1hX4RAqcPP
v7iiQf7o7xzAn1MFzff/oCKqukebmwbtew8FR5rda74SC6aiayXZoKrsNx1EZen7/+o2WxDGnDdp
D5a1PwMvQtkxmOCR5fu2e8Cfn5LPKmSXzvv0vh7kyefoU8HYfnAQmyEFw3KxvLTKKmNKblqNCW7E
vDPIjZ8in3X2iUq+VjoO/N2laPNb6fVtvnPUpikr1szNOwX5EoJ3zEfIlUZWfUv0e26C5DzEqaBp
w2Z65XHm/Dk94CkiTPN2t/i6FHpJCfJXrFb6F3oLgMRFhsPoYfCpmtmFb7QirZ3x80252MhK036f
77UxwP0W340v4VnotQAX1HSdVvgz/hc8sbIaj2+fTtaTuSfGlMp0fFBIme0RcQu8QB9lu8Vu+xPC
aIO2A0dQ2NgM2vZ0E0vbbFUk55Tm93Kgkxc5Jt6GsXYVnEemZiiPyGJ1PK4Io0/jEjNPWOFq9EUH
WdqXmm9ESgKOQO/Q/DzR7wNgXE+ryOiSkkWRh5T6F4GVkcOij1C7+HcrulsyqFLY2FjKcoRUmsar
rxY7TaU7XMycLdBH8D2DtFo/ZoQrqtuUmltV/b6jDFid4zpxqbvsrKlFbibKgwYoLreFXlvLAh5I
Q0i1fFC60ttTOi3FTrCXddebF1S9DxZ6BfcVeESBaitBbrefSdWZB5IHeTliTlfC8gkc+etoAlCn
8NrK+Gvk9AvyZN3i4jt+735f3qA8oHJjZyZcaN4SewJCmITqrq2tfZXXgO0osoNkCwApp8OdvpO3
YV9YuFer43JuUkJiwsiFTORpKkGH/SV45CB9u3noQzN3j8+V7YOYVYb8bCHxUeYqbvgNFvvja6ZM
/0GA+616qLaKWA3iq4jiuvPKZZIfZttZoYmxZcq5jKeaRPNCEJ5AMa+TjKOWLZNtvWFZpFz8iTPv
G/wKSdtVDMD7GohfJor/aZSM0+Srn6yf6Ys5q0Jyof3p+jiHHFIyWVYeJSxXp72mtgTjbbg0ythf
RmCyKQFiWw88gi/d19fj/h2q5Fip9ccI4n4LfRhctq2CZtkHeZZjxIyCN//E3TOsk7BE18qGILvJ
5CaGhhlOeRy/+Bg3wIBL5P/rKqwTsVP6tXOsQvsZMOdEHA5WKEp4xvQDEQIv6G6EW0OdLom6w8O2
y/uU/NtjsJaze+eJjjkKwxTvoCH1OHI8o/j2nSZfXMYxtCgvv7tP71U3zXNoN3lL7Tq3ri6PCGUY
z+7oWuyYrm52bc/4Iyq+NSoomTjkKDUkHAgEAFlQ1QPROumT/J564gZsR0rf7jr24xIHGlZrKH9a
hWsTlsAGelyTRAqVJlQkJx9CzpYbrZv5oR1/6RVczk1vDTkQXAK0zk63My3Ms+wfvDaIFMuKeYYh
e6fzgH+kt4FuDqXIJdD0AhuLwY5Xx2RfHVWunt3nLhegqNTZz+GJQwMlBaicItdIL2oxEWIvNrhc
HDuVpEWpge5L9gabsTJMx0UorcdI8TRiKLWfJ9pmf/pDMIvty6sIZCfW6xI59U5W8SgOTdp/YGs9
TSVop+2CIqsOP+S/GIauHI+7Y+y9xb3k1q57F/P+l9jlpKDp2mMnNi3Sk7kDIbWhkOxFHM7LzdAf
KW6+694j3ESlrOrmpGRyhWlGp+zlXVhlBQ9/YY407uhvqUJhjO5x9hHAZFMHYo3lnV8rqT97xY+J
dnXZkkxGe2ozS4kYyOtwa56Qfb5OXzqTlkh5+ToN7OtFD4ZWg8DsDNoIZ3SwvC6rnAUcxGLBoOeB
kKgPZ13xephGjywVYPFdudvaaL0f7qIZ3HeeNJ5hieKCIP24bYdZbbpSEEgepsOvOhBLDFqlgbGf
Fj/cWIM7ifuI0vvHroaHgcwn/FGaFmPEqKmQd8SQENf5uazg+yq20d6GfsCCB97nYv1WEnkcrLE9
OrN9IiZ3nNmIanLmCOfGfoSZP3+o9+lXO0hY17hF/mA+AcOn6bCqH21mwtyYBpkgYRlENuUOHvZM
ArYGqebdeif/CRUclg+O1FsFUotNUEGspVrhwg9nFXlBt3Mf3QqbqgxtafEOPPOA/6ZGYv9mICvL
uRw0Z54wCEf4K0tJzzm4+ZlSyWk3cE1+nRBgrlYs3qwxf0Jel4p73V+ug/f2yuK1ZyrqBiQAzUuq
GG0zGuGnEk2hebRDAzTqlh3i1XYBDchs9ffYTKM7ceN6bIX56TQqIpjsEsaxsEmQ1iiPqekUQaKF
SUHCn2aA36ZinNifjJ1IzYro3/N+faWyyGASy5f6khcmt7jaMn8rtDAblXUR6UY5O5Qa9XSBzDq8
I/3BZmxd99rTro07QNMtpbpHN6vVct4PP4b3TF6xKu+rD+RDgDhlPptBX5ZFboSsP8V5N/R4KHR9
aCtciBn1XxRMt1I5k/j+msBouOetkJIPzfCnY66RSELPWdFibCCFE12UcBI0r17TOyCYWPn1AAcG
ngqMdi1kZMJYnblWHZIOwa8p7RIitfJBLlj+8YPZIY5Enyb5MoUGNRNba7AtUQABwflT2egu/9tk
wl8/zK9e6leL7E4gOjhBkGlfpNfwX42kAa58KL3CiUFvBPtmyqs943ndAA8GVpmJO/9v8AkIInMp
LVYm0dcbsD5SdLbOsZshXgvsVolpzI4NfTYjdwM18b/jdfySkTVa3jGt068Dn162jhuVH2FZKgwR
3S+wCI5talQ4qyiJKRy5tY6wFjwwJz1Idbhte2RbbeCDCj0EHP2EqF/4zsMtqNzC3Lx3Chng0Jto
aqBKI9TKvrVb5G87O5lzRmlgQBnqCN3gDZygeq25QTb8NNoj2SwDEj670FAFuOt1H31gUyWTNftV
AA1+v2ynYKdZLz20DLGk/RyvX+PomNFqbzFgoN8uJ1MEklgK0npnDWzDydlkwx8FpCQrl0jd1VqK
AyBxa8ZqrF5hU3ijPxYWcclYh9v4vwPxDL5SYV2dRtAZ+QnzEXIzA7mdbjuuyRp+i/CxNGA8nyXk
od73WC0RUkK1Zico9gc2IIvPs3wVt5/8HiF2o9yL9qeNR03B/foUb+pbtpRWyBZDYDEs01nEA2xF
FEnB0zAFYVRniq2EL3bAJpuVUpDHztzm9pWvBoYQXizwrkWQDfmQ23I5iLZb61Vuf7evx0NzA7rF
XiYp4CUjLmvu08Dam7HPYJv3iApEfHaQE31ZsrpfDBX5N8342fd1CYc3uypEgVr+LJvfvSsnBtsw
3HT8zOwzT1i5mBmEQUo4OUuRIdn9m+G5gca1QAh7UpWWvsqIxAu6Wuecp2yuiWK9pzXlLwSzkC8D
E2YtpPF7de2Y5PkLBW3CHyiq5enqQxYWfUlefkiSSR7gHviVhcfVBVXazMoSuNZCZ03m6rYqFZZ0
MSi7yMdQIau/5bh1G9WGwYe/U8HyBl8E1s9iP/d0cF6+eAgqzRuQAcShsdVHEgGZY672OFxfIy+M
j5WE+6LFXzQIW648viG9iEbTL7007oc/pnEEXayIy7Ht6LcuQy8YFVvj/U7a0C+ah2jwfstQyOR4
8NykRsRIMDoGOpyQomi9tLPJf5Xq6Mvk5u7iKivfap+J13iDnYIHkcntq03Z3Q8Xe4+0Tos+zT+L
KKpYeZk3KldjqMYwS/oegPLhCjT+gWTDwJXbyzmDr/hbEQGc+9flZUqFFyZkHSyyrQIBgV86WXuh
D7Iej/I7mKOFks2zNr4KiuwaZaFkFnxkcmeJS5xyuASRu8pplx+LRvnIrgbkaiOMhPxhZvfHrGC/
tLGXivU/JaTPsOqPA/QlLwNMMiq6C6i9j/dTROVHGu1Ee5/mEkDqxvknNm6G0qjHoxhcxVygPwmo
bF3+r54izzuRJ0KlNs4ohjQ31rjWwJ+zVoMqEEEubqB6m+3uyfs89M2Fz1g8gI566KIV0LNx7GYd
IuKPV38/nL69kDrxtQL/OFK7ATHx678N7AOWZc6hgiJepHyhH8AFVb0fOe6SDYzXaYYY5qjYi8Ef
tfIqMseItDTfSCSE2JxebL3zpCDeaOmcU5yibRavnlCxLpMoC9CCFYVaAFTBEDEZVnUMsJ84I311
63xTSMfLHSWRvwMvvCWmi71C6wKGBwFfurfTMx9sLcATdaYUhDiZdbTtS/pm48WHgJatVG0rQjON
fugelZWAP58KguTv5P46r++nHbQaW7xdGlHTN652PkTdIFOSsGP8JkUAiIsjmi0FqjdamtGNz7KY
WLELHLF/3FLOWjhxv9xTGdH0SoK/40hXVwGM2sREA8Sx+C+zbSc/LOAlbE4ry/1f7cWwOgOws+OI
YG46DGhHF6NiVXC+fQpha9KJQv88gSAxRTT936p8HJWSuvL0Jcf96PAuSOGJ1oO39HRaHzdqpNuh
fpRqd0KTgt8DqTd4Wx96DEnbjsQQH5cBQ/+/lqfX7spFP0fCxyWegiZV3vxGnSv+uELaRn5Up2Vz
rmBLTXZEiaKtx3UZQA2jBi2TCdQDraLxbt2+OwmApgJxz+UErh//ShsbTlYP5rN2DhydYFmjd+q6
aRBY4dD7D7IYYQKmL00Xo9zokmIpNZtabmQ7TCzWN3fHHC7WFkTu/ZA1tosRfcGiyPT3xdp5E8OC
yeQXghu9C4p2wO4l5ERAdwY4sAg6gJmdE1+YmFwHNA2F/fBgyltJLSB4TBwsSt8TDBPd4bkZ4B/U
jEw1FawK8QC8/aY/yopMf68EWUj3rFfKGa4U4b+5TIa95PFeNu5HFmqy6oajePk9qONkE0syHrA9
3oXZit1CXxYYmGsQLVqOUB8S9x+M54xv7K0dBSXY8gEWD8Ok67RJMLRuNWDcpSd7uI2kBKQDG2sq
30/hEgivkOZvW/Y17LU8MClyP8b7wVlO8Ng5BjPLPkT1quAEZtOZ6qs89PgNEvSYDOaODu1qu84G
eYyog0WgWFCVhAagU7c2r2yFoewqIujJ2v1RCrUb7jm125Rug/G7v0cQNkadJq1iyyy9pGObk4fX
/IGp5iftdjqLBIKqJcYwfltliPcM1Cl94W5RJ3pzdZAyyWAMjEDoRL5PnPteywMH13WGvZbe5XXs
eRBdTW/VcEaOtAHcplJ0SdzNIVobE73y2H9qOGXHPMYtw6PTqXPcwFFhjlDoM9MlpZhzes5Vq1RC
YGSRrWnn+ABNyhQlzOD7U+Mb+UyqMvM8ZOP0BLV2apMKjpSzxmU98ppRqUgwARVTRsniVo93CVyV
hK16aYP8KJ4rUNHPUc0PXYq8+Iz4G0u+zbcHcSbFs/vnnF1px9j4lIGW0mk8tt3rtwHNiXXLWEqE
8rxk21jxGnc+PoB3RHhQi2QbgucyNKYJ4hyGmRVtTboAoer0oBHnFjbWW0ijlrB6WOfzeM0ZwMSF
E0hSEVEClwiD7ImH+1aQOumFj2OIMFZ7chdHfPagyRumei7hJ/mpWYYkCTsw82XuJNHch1O59x0m
9bxpwc4nP/W1RIc0KTfpbznpduVJse45SHDmEy67A80tzPmnsErUP6g0acJxE2rG+JPJOE6fbbiN
r4d15izsgzuHdEqjX2r4OBMizNqCEK/p3tkyjCjZy1y9vpeBrXoLPLAkaO2KHgd6HSIQ85UvDdQZ
2z9O3q4kpjY0V75p2cwk1SjyGs8DNHQkoEOYE8weKZdwuAsw6VsypMyMG51uA6byF1k1l1hELDpy
ur+noFQPuz5P/YGCxLIF333/zIaPW3TeVVHZyla6MItNKMj33TpRiWifARBfF9TrepdLqBZ9Gvbc
XF6xynnUcsrsKLoojGX54UHVG54PZQjQ8D5iVsPNkPJcCDbOcGMt+rml8mSF1nJQLWglguKZ6ux8
hcDTsMDhLufGfosg+pOLbgVAKbapSiVIFrcBACpL6ExIh5qffgCnolrRw6JmnZkIbYtl/7D1osjh
Z3BWpbHKtnI2dRf1TJQSpXV+D17P9aSyNI0ndxdPDfHNtkT6SZoZj/Nngpbj5fF+eygVI1CwIe3/
Hmpz70N5WKsw+K2Y3gDotsU+uIxOthBoUsqW94E/wr1DkQQ6bhz9hd4SKk/6wYTNOuJiJQq0xevE
nTSBpissUKfbXzMP55PC9MokgKXNiu5awMHqpLm8xUquvGUFRsWLfaJsQx1Tn8wliLYIPDHlaIz1
2UJTt81AMkgoZT2+33B0uKPieX+IT6FLROeVxJ+v6qREK8p2Z3Nh8aS+23MffatTY1fNxtNsCAAq
DbEE187iKKIidUMnZossDIfDN7nE2dPuLpGHf+yEyhX+UK3EoMcxGWDFWZhRvrz7IQsEppjM91By
lN+4luDvf6vGBVHhLZsmK2vf01X5M8GnZY2P0so5Xs/A9aIXVmiyFkI4wetCyetcsjA7MCHEsChU
E2MOZ+e9birhHS0KaJXv7vVXnWRz2zVEQJDnDLnc8a/EDiKK8Ag5cuu5pIkD1kMweVvp3gbUYJfn
+ZJpu/GE+Eu8CLB/8UyXDvwX2kAbkkfCJN5FH4tdDoVvQq0rEivGVpWGeIAG7KqkTPdWOuW31y8s
34wnli0l/P7u00H/GcVUxYwqHDnT8oQHbnIi4Z8++cTDwqYEBKkjJn3NhsNpeR8tY7Z4PF5B/FSS
oWXDo/jTBhPsMS3ayED0fux/v3dfmODKdaeHo0heowErEyOgdl1skKCrAX+b1U0CTJGxotpQW9xd
NQhoNK1Iu6Uxy61Rq+U2N5xAmCnzw6WQNB21jvV4nMMgXeZS6ZbGko6E4wPZqG1slmPYcpgZQYyC
FPEn/jQFeuFKDGMfySOOV7c353LI/YKJUEoXIUAREoOOgFhT8rTz1zHo0bYUvnDL3o2uTyP2+PBP
g50XTIedmnTwZD18HZPfkw0v2gJ52hsTxg4fD8Qb/FZK5CLShQTrqQqj+VPuF6bgyHrrtOx3vxkl
glqbL2aG4pf+zbKoCx2vgvjwCWlXixnGqQZntusbmP4uUpV/iJO6KUb9e3VkDoNw/2kAmlmOhFm5
d3CME5tohVBK6+oV2M4dZNOxYOa0Z9W/K/v7bP2incfx75KZlNxD7c9Qi4j5tkm56T5qSCWjW6Lq
R0mTI9ux0sA2jPgs9pOd8MeplUidEZ4o+N7oDxTKyWY8QVeKMoZR3TzwmNkSlBc+P3kiV/Ndi8gH
rA2Z+SZ1CrE0wv/1erLsteABIpnB2c3gieTt8FxHDrdhwu9hUm2gMzmMiwJ7zdxfMCYk+kre9n8H
9Ui6k2/fKogVYuZtEhmSyYiXditlMWoBRwZMHV8tA8/bhWily951POv3Lf9XW8Lzuqr8Rigw9gbB
YeM7u4Qb+4rB3pbw2u5JZGmX7TsXvCDRKptZXtyuuikldzQoHwJyCPPPGOnenZxZHqgRUGUvTowm
+jn6zZ2IB+EhgIC4ROy1mNqHtUrXeMqucs/Kw5Iy6sqI6iYuatk0+57NKK2QHicYURvsgmyVA5jn
pWe8xBjz6VNf2GhPd0EQUrJWVWwWcCg2ViKUfI+jRVUsytbhtRDgUjYghoYNmTn5ctgDHONjAbUE
FijO5VoNrMU8rFPZvwpQSxHb1KnJHwQLALmRCuVW3ijcsVUW5DY4tgkyW7STaTqn3YLBmFPWOJif
2I9D7L5LuWngUynYDfGWlsReQ20JJt78LYQ8ZknhejWJwZZmTYtysKADjGvBTRn6JJXHlgfDGWO4
Yq0+S+ZXhI6EylaPu/N1xpAgqffNhOD7WCkp2uhqeS1xv8N2S33ukeUEpYQzTMdxmCMtUs8HAG+e
UT14GWaQdKEN6z1UZRv4gpBFZWGARNzM/xEToEJXCGXCOLuBlmPFOqHKBXxZw5lcLHhij/tFLJrb
t7DzW0VQIGUvx6rF1xnk60ZFNVhZ8G95WE2susrUuh4pOfLAC5if6vlrbzfe+FykcgXyRoiZUdUp
eTtQzPzL1MTW8g99G+S6iBKRoTWwgR7YISwePVUu0e5hviGCk8yFyerFX2Yd7mlgcWGPd5SqnWbk
AH6GiO8BdwD6U93vnLBdQgbEdTl7j/wXEYfvKjWYnXTTWP8VnyIQXdxdP4Q336BXaeps5JuCHJRf
aDpgYaf7kgt1ejx22DEEmAa8ilixAUop6vBkxXdl8NUUzNnBHToed4Vggf3aMh5nwIyZdi+hm/Xa
MQXjcNsYr+xSRdStzeYpJaxyvpmktAobkWgIHo7jDzqYPgPOh6EccLKF7TY8w7KdZ8myH55X5U77
6UMGXUGGMjxJo+00xQYNn7r3uBSgRtecr4LvepiXqStPIfRNeorDdX5HShY04kClv7d5PktqFEbN
bp4JuntQPW5Fsa9Ymiwd+4UuM2xZp+P6AGDsfGUFVMMyoR3WbLWKkaz6UO/ypxNKrLTrzf8jayq2
ny3eIUPQnTP+wQyPt1g7cNn/Ke5DMibh6lEJNvDanhNKivTGrVtPM7i3GqZsds+Vle5LmuYc9pqj
3C+kdKHzS3hglqOhlDNR8fMD/o7mK+PKXXnlhz1ZLKGrlZ+f8cZyeY8VI6eVQekPiUAlUOfTX8Pq
Q3Ti7jE4jm2YjFtu3dn6UZkkT+mH231zL+klcP3Qfck6od+mNoIDPyeQ9kddiHfK0bXBvEswWN2B
TI66pjMxeotrvJU66KekpSi/sUWcWHLkvbp+8V8UFbJ/XChEr3YOTmWrCdI7d4MUWK+GMCQ71Vdc
62r1Ke7OnXaGur+4nQLGp7kioXNxnU0F5WJ5axJPH8qmdhhiSiw/vjonmiqhL1MmeFsXYUaDXiXZ
I7WwmvH7RjsXQsAlX4UXS52mjRxFRjDxhS1BSDizzhvX0/j+0aqzsDTS7SOlbvdRsWjBmQdfyeyp
0R9k8Ym7FNzEFO/9xAUt2Wg4ARo/m/NJ+gRuRCb3K2iVYl6miSlGRgwMxcAljcrbejQNLNuU6iH/
VAmzuPk9ob/bSg1biYNWy4lfMn1aIMx17TG/K3iSDf4LLrHx8nh5nxy/9gB3DMAzaASbxLhDTS1r
E6FonJHDIxOPPcpXH8hFCA/ujoZu4zLQetTz9pSsVgEFhbEMhP1LOWpbcnfdThpWjAcfvIwLtdZG
EmtWGDw9n+JN6AFplrTx0CacAgsx8h+ex0b6XZWtLidyvtEZKEGsnYCokJaGdBsKtryOwi54DXp8
rVD3IMSs7O6taENXUuME60On4XkEeVLVmdoAWxiQ6FjVrDicoVSHxF9yItsgNgEgGI/kx0mABlqV
oSnANgoW2CL9KYzFSgdbeotLeY/xM7TEmUUVPgJeBFxw1bB5yHrfmW5C+C1CMLWaThJg3dIPKZ9b
6DvqqH8+UxoF/y5Cn7bXt0uNdSakfl4+8dZRw0QK9j4HfjgvZxxToid3YRYuGwf6U1HNuah0Putr
lXZJCoxouAYAve35fCRdtNSXHf8TH16MXkC8fMf4unCLQii5EwSwD09ovgOgps7piHGESHSV3npy
zx5MdYkffscpWFTo2jeVxbyVlSVIz8JeVnmUwZoj2YttgYYmQFRpLs9+aqqsNEIixNcEsyuJ5q48
2fHx1EZWZciU3RxEILUw8KFQrDjCZIvsfDfwiOQLKFM2KQszakI3pNZF3vT8ENdLXDTSTjXo5vUU
OKwtWpHN2ehcSBb9SVO7r6XyWDLrwimBwLDnZTKlXzlA1TyEby096jG0r6Y3mlsPzajZOMPl00G6
5WnxLLPcr4p+vIOSAxPc+SttaW+aguk5IPCtsE8xPaBFsmhfSIxqxezSteVCMChdgBkBa90obTsx
Dvs20KebNAuZBaEy/NVSCfSIVYMm48Fob08kNQmnmihQrNk0WvGr5Uv6H40n13HTmZY4+Cnx/VTY
A2CIKcP4uG6Vo9s0US4D7pYRoM6JNGVN2qeTu62b4s9mT/E/SJhaBWT2Jc38YSKSl/pDMmtZ134m
mKwGgbSVKajN+/IsaWxpCYGwFguZZnSyyLsRTrW6H+9edg6mPPNO0G+WZv7BPjlw0kW+9JpW8oye
rQx14Nr4OXxfETaWt7cHN2Deq0S34iBCGh0itYdSYwTfEB5swuL6FXH1MAuuz2fhOm5Wk/rVR2iQ
7KyTe/OGGV+TMDpBzZj7WQPEod7ygD+gDEl9QjVcT55or5YRMTahnJgC2ulafkxf0mIxcr+3rakX
jdeiIzjesBE5btaTYMz1uD7MJIyGPOZf6UUIAZvc678YMJwyj0F+G+dolv8v0kFNBw8ez0FIEQsf
dFU/1xHw8uIPDGE+f+PDdJ4K7vw6weVqWcq4uTcwYYD6gGzMtH4UXDBNTSMiI38Ig60NBu6KHquw
0W/L9Fzvu10XT8kh2ZDvTiHksJbcEGrc9hIO4RV53j6HqfkEpRVr4NFe+6li+0gCEnS7qaXGOUPS
qGb9c6IrVzV3/4TGzQHoyIMhTfiIdSzCb/5qFbqqM4fx5dOUNr3iSWuOzmX3GKvAF/23vxuOucPV
f1iNIEzn38XLUfoWAgyAWvZmtiApI6z05jtsLnqITMSXqEMTdsEqw6px00zfv36YDV4f5GbmoPpD
6RR8VR8YjJISOHIkbvnt2wGEanMQPQ7jmZdLG/xdOfjPycm9/J55qrqPpEfU5gQdcifogXasbSzy
h35bb2//D6qOxnz4ceYLE9T5rlMzci0OFkyLmOmUt6Z5XO9G823wLLLjcStfCaeyfQm1KHHAM2xB
cEF9x+0UuOvsO+mRkl0p6gEy7OSDW2ddptha15yGLCLQVi1kZZxGqQ+kTYLmHyMTVpRdVWNjL3i2
5i4pm4Ev0dhfEORqJOExrVMEqWM2NHfFaqZUoP+DTbLLwye3iW+sxo3IrSvbuh4m2ejIM/8qOfEM
6vmL1MI0B/EYtZ74R7tXZRbSaTHSGxMMBQZ3Y3Y/etNJcFxlRQo/QMpzs0KIkKcH+P0OvZiWhW1N
NJGCmTgu4Vs028yCq3wzDqfsQfDMdeRuTqfUSNKo7bjK5Y873PxgbdYEvxIwlFxSNQnjQwBIwIKb
wa4hcU58xJ5OTd8e/iXiW6BAN8b54sta9uqTw5iQreYCVDnoFsPLiKc8c2YLsmM58+K1X9g0n9Ji
DrdXuIPqVrXxK0xfrU2U9ZIK5MR6mcGUPUtxh0O0M5oVUmucdss5NlmkhyqjGwty4En4QcfYjpCZ
fJduw7GKLrO9/vUQGZOw+DP3G6PcnrHsyWIWNrvNqIjnviFUsnXoKzBtiWIxyKYtiSNyYzvM6/4e
/mPR7culDm25y1/1C1tvbYCaL/d0s193rljgKUoVXqTdHbZcZ7LOl8g197bHr9ja38bmIHa7IyBE
hKeo87Rj+5+gXzSrpAdzvckrBdZmvWZTgV1/4176+0LV5K+mNFYvgFdzUlCrmtIRLUfJaorpm8qq
hspAbQpzB70nJkvqBJbHnJN4BR2O7/BAirNS7XFhEdTSvZ4C932gXotEq1HegsXMO05vgXhhy20F
H4VGcTFzlWgcUkPQTf+r10CeA66MLp40OMo7U83DH2voRg43xe0jsHKr2OWQ5mBNb5GwiW5Rvq97
nMGuU2wtKrUco7/FfYKjLk76JIZagtsJkCH504HA1fudwxgnGRc9fTWy6Q4TsPhBAxXETJkw6pBv
cjMd6k5lYbRUkZFSTRrEtKzJr4OErEv3uUUojnSDnyLQhWKrI4HFEAFkPcYrB0esHqiYd+NAaaQ7
I30YaAgLUXqUnxP2cS//7eMt4C2RpIBglvTepDEacBKGGS46I5KjSEPFs2gpWDZpq4SWk9Xl5rzw
KsARk4FmABl9vJ7WEVha8/JkIyjG41lslubTEDk0cTdAtlcFSAZzJTrJV1QKh5Z3jUNNSVDaItYx
g8vxvlM6IX3TICuo7Ue5tDtgOh8liI1aiB2619PDEALbc4ehme4S4doHFXMwlyrqDu2m38yK6IEL
pt7EdVvQ4Ld8mLvo6EbFi07LxfYKedodzm5HdKQD7LeG0HhlkJ1CIh0dSvhSLXht6MQhaWWv/UOO
8odl2St+UjU7vhMdNocC0gRRqls3tr/z21lIeR28c9TTkAP2gQYBvH3RX7PI+DRSmq1trU9XpCj5
Vhwlp093kqVevdOpkk3b5YkXJoTSdiMUjOeQ9cLK7aYjHuUnrEaqjTTYqD7MDc5rwBJbshH9ngEF
5zdbAyNK3Yhh1hWkNiPjZorA/k4CNuMJj0EKcqDWAwrzKfLkDgqh2B4O++IE4lkfVwiqE22Y4ejB
tI7Y5R8Mue2nyg+gfDE8dMMgAZX+xL+qMiUChw0vN5up6TvyPW20x6HoCsm1GySnGE7idecJKM+w
7laQtZsL7lXnukD4HrvW2NRgIbd+yHvqor1I+Mf9GqYCa/DS70JzkdyGK9oJOBKQknfoenf2luE+
Tr4N82kU1VlQNydaZXLQT7VbuOduNKqnaf7ohP9Foo36gbJxPbUiygo4b6tH/6gaAm0iDizwd6sn
z35yDSymnXmGt68sJJiam8bVixBWsDxRoIx2NipjyQISPhZX/2K/zbcykP8QRXnPR93A5bM8t1N/
fDRpeeVm/CsfrKWGKkzVckP9QVKgvkzGPnSNHGKzkkcm4oPLj6NJrYz59Kaphvy8F+6Jj8S4YbQm
vFBMkwPclfqahxuNmlewveMpxy5yTzz3ns92Y46X1N/G5bN7LL5RBgBw2dtFVdV+8WPk4IPJg/5w
Z2LfPhe+JT/4D7xAGS19ya6p6dPczkjG8E9V6jv/ecGDrHSJQ1hobuMFnt46DSw5dHzg9dUUspjc
9PuPMU6ktNAG1wwqrofpfMqr3ZDwvm12y3G+JIZBhdEMQDhtWceylBvExOYrphScTtS8NIWcP0eb
rODWw+3DPqy3Ug7iFCQXeR2Nc45PZrYnS+Mi5yD0BsDc1yGbHLqSmnuxWDrx0Lpwkp995EvOqYR4
cjhakS4yA1+iSGIY4wLvPNQMRPlcSOOiLp4orynv+vH/TZOLo1Vs8Bee5ypTRdJRdUBo8RqP+XSh
ENxfB+33iJELIwKIrwn+BEE3/yiNfspE6G8NxyNG7dGexAqGZJXM7boY/O+a/9DgQD8O4FFv2UVq
csdLOYEiDF3zSuUCVwqqLHYhMmEZWJFwGYQWpkHdTLYJmD1K0Fjii4jjbKJBxFPr5uD+9CqNher1
guTasRP2BTI9eEqN5qMlwjy3+uJtKckDJGj6tXfWSSHDMwiyf8NM0k9tQez5rzFZnGUfPTgJpXMT
JdoJCymZ0U6uQCvyvj64718cleAzHax8/wTVIp4oGBThJhdZCHXxsL3KXxosYN18BmIyXuXEF4v9
av2up2tSKDgvNmteuTG+Rr9gzB7vS/3TKj3J392Cgan3b0LrmtDW/Dorsd5LUXWQvs425Gf5nzUK
R00lWvUu2MtPbXBVL7mcu4Znw8vrb//gpHdEURcKKlakni1gFxrPOydEma94UdWlqxk1Fs1TSBvc
W0XK1KlPrvrGKbw1QXpzg5ZZwkFgVhnYGTb2Z4FLs5lQuNC2mtnGbagpfd5bdYb9UdSZE7KdmA2l
d3bTaaeZiNwRsCVH/DH2bryZ4epBqG8TNaXsxZBytfV59cYS0kbQs4M8rFS2GI9v+SVYcv5+Q1IX
88wR/HN4WWdWWYmYbfFLCwVqKnUxgk0Z7unvKuYLvV9EEosZf72M4V/8SPncQG02GoGGFWXdlU8e
0D5psLPwC1fWdDBGsfVqCusmXLKJL5O7geUU+6DwJoqW8t6Ftxtg2NlotZ47Pp/dflQIoZBXM7gA
Fchsm23du5pAoEpjo4pyWnVaSfI5bvI49CWWad1EBQcqIaRNPz218TbUXO0C4s8sRPXCG9yLbdPB
1YyXTr5o0+JnaPU5CyLHUPV7NuKdR7CufrQStg+oiMwcQW10/LPTeKnqkfbefc20QP5Qs0Way2Sr
1KGGECRQZZn9tcSo2/EFbbTSbD1vAc/kdzh8mkMBwNbnerr5zfC0j0BLIYqH6xfHobAKUkrLC/Zz
b5Hwn7iBMnB+ik444WtOpmoklqejJgrhBx+vYwQ+Jd/GeabghgPqJ37mDqxZFe2D4uMJxDQiOKWr
UkWH/F43V7xucLCxoPaEE9QxmIxt5sgFGdey2pOMl8h5fn6VVyyFZ7n2ez0194kd95QLp9zv+iRW
7gphntMpetE9JVnsTaLFrOlVgkWBKO8T/twkk+LNxW+AG98HH2SwCP9nq5GkzVcpdZIMbbdHrM7v
muOunIeBPZbxz8mo7++ZpI3zgK2vtI9YXSux2miEc+wXhbXA4RZ+WB0cKC1Q26gnFa4TIb2kuhK1
4pFxwwwjG4gDzIxwgh8PtGjmJbNppwfdq8LXHsg/h2pl0zTlHa4zlcKcp8aGHBFfW+Y7f/lsPe3c
+5Umf37vn9KcF+4Zm1Q5fgPoPAu5FTblwSCzfPxX0cXFSJSUolrKIXlcYzkomCusCEQr2BY0Z14P
zxd8ItqiFWN532L8b5lO24nQtTTfVYREyUL2tUk+Ji6nGG/tXH4+cgnu+XEklFCa1oFwQ1WGImvw
mUU/keny3GAkajL7NLjiIVSUi1ScpGSVf3DNxa7PnEJDyur+8xTlYvvTfOx/qMzocR688+HY0yn4
lyO8XsaMAQ9OKwLFH0KXhgXGw9OI/CvPqX39VUqU8zt7TFt/HH+aLHPvfxuyvdcjyfJocgi7jbt7
TDNyfTKG1lQXcjn3+CIMfc8GERXFDqEgp3qV9vmA17nt0g6Z6Se7Iz23ynCc++ieD1piszjZlhXc
kWpSIrytw+vqwOGw5g86Mu14vejBAeT7TZlBwmFz2s0qRn0KfM2wLiJGDzJNjuffJmrtVmPB+X3r
rclqWFRqtjD7DgAfu53eKq5pdTZp0NPjkeeZRx6/PWl7vhWwzrKAkt2aKO3FxD1CTOuzET7tN2Nb
xqS07N5brTBGLNMhsB3BOYrb3hHQxG51Xh87KcvPH2FU0hr0l7eJcSA+BzIOoasDbWcIYGaUudWs
DjA/2xf1tuxjfYiVuaaIn+jIUcxPEjVVTB70SmU6RN8Z5ArEAX4aB/kdk1Rg3RBjGnw7Aajg54rZ
nvJqW5zVVtJqPxogVt79a0SY9/8N0kltmiRy4QJXn1rR5fpzvCAMkujbKrlAr8XlpUNGtqGZgL+T
fKFL+dvLYK3iuSvhlwBjNBQY7Y9D+fFF2dyHt14TAsDAaA9/JCl5vklh1GYlq/8xrL9oFhoLpGar
Ao3x81cG3WIvhsFpFOfBlHhGZn0Vi/P5iY/WkYxJnYv2XTdW6bqRMRi1MagibbUnKJaBpZWHzaj0
ZI9FBsql81AqJc/GMHV77WRiGOzeceagrioaC4xyT34rlDNGn5wSRwsxFHguhqHh4Zy49Rb0FJ6X
EDmDSaqiO74Q6lI8hnkqrvRyn11FUoa4xcKDREEw97d7YxJ9jVAJSrYzwfwmNC52VhOL39in9HjW
0oDiwA6Pfm1ORp5dWldJ+QNi+JbohpWeZt21nFpRv84o4Ned4Fv7ZHYj5eHz1lQNKYCoFedPGQy1
dNYSqK6YvuH6yTRDXwJiERrsCSALVC6fO/7Ijdnv0wR+2Grzemn9IrnE6//7qFGAel7dG015581d
C9iSmkoRTNMbeqMDVc60YObTbnEax42RbloNWqpL1KncFJUHJkCwEtC1PzO7F07mgJWLuxfHUVjy
nBJjmCm1Q2G8PEhG2LNq0l7JgqgVrKA5S3lxN+P4R6tE6LrbEHeVu+eO7NgwbJ0Up9NZvuQ/py/I
YgcMVsuNOmKPseEs75KFVK8poEXsYRJZ74MXNvS905ROnKVAjv+0uA1ZE1NWOyX+CxvzDddzLvnj
huh+btIhQ/jfX/ihU/0CabELJhRZro9FMnIujwIzVXp7Anxgj0tULZ5Hl02y8dw5yx6mIOEuP25H
JG971h5VnQs5RkZVSi7sfDSPedTIkE9Ex4kFVnpxNsXR4C4brFtDID2Kimle9+0jqhKTv+hThMi1
7W8IFd72rYhWLWERct3CS2sJaEXd0LZmCD0gYLci5ADpNbiRq9G+ynDJEICDtsnu6BNDXJd82IGd
Os3+Mg6lbEkomCjv6Tdjb8IFakkGnR1OVpilg6oyOT2vvboIrEgUGxqfohfY+TCF304orcrhsdrQ
vSeGHIyWb1zjOtjZ5U1xqKpWQHu43xUl8v0z3ojGpnMOGrKsFWcLSXGiOxL/eB2oQegixmjz/a+j
h7jVwDLQ9HCuX8hZjuEPO/AlcTJ4KnCeTV3sUP5bsRrpULY6mxphEdc364m9s7Tn2hl0W5uLfPB6
I36JQLDtuADEH+rWept5vDqSW7d9Fq/4+2jn6mUJkCzVH4gzu6fGi8oNbzA74E2L3CxokAn5keVH
SsExTeX1JuZMh2STGw1ZKiDe0dB7ifyZ02ZJbgKkSpXDxUJTySsH5PD84Kt+KK4ab1rxI0ssYo8b
IQSiychs1DYtIDO6qMpC2qBURLGRR0PMpb9+0F5rnJCDXhN2iJQW8zmwHm2GOelcjyPX5KwKDfsn
RE7VTKUd9Udu3Mzrr24g3yuKW/bMFOtATXHIcZiUm3NtAT5vt1bWu4mQ71xmnXUVPbX+8aBSwseA
Thn1n2wAs0aDr2ElsI1wiSzzmQBkKVCug6SJ7vlu8E7uCJuGIGxgyjsaMIDtCHxXk4LHwuT8uhvZ
bIg4O7nCiqtOqgbPZYVmEMzOJC9RaEsviNQBnpOGMpYWk+2wjhDVhQ3nuNkg4Ezz7J0mXqaYPUyI
Fn/hvlqVILb8UY8lnhSeh8QE4TK+1tHdWMtqGtDG3i6sVVVRjVRt2s6IUys1XdW29ILcS8TNsh0g
dy56s2dqubUT92XvLprIskdrwr1tb2iq1VFg35Ce0t7d7Wi/s6eb8q9yTwwKhK0cz5pMpmtu/Lcv
+La+vwutN0vXZS18J0CMm2DwxJKBLyL6d7a7FnhgXEi88h7EOj/J0RCLz5MjV0qSK425/MLK1s7M
HzzW4IH2xtgKexgfPSSndZpB5B2zVI5Rp/4/fGyyXLGhW4fLzz/GIYGfQDCz7sIMNFNqetm0/iSW
skiBpAv5xqjzggV1YxD/otL67krDO5fCZWRDHk5T2ROXKkh+uL2R9zdN3McSezIjwODuq0trxWIJ
a47YX/CR9Xid8nhYeMCyuHa+dvpY7XRykZ9ATTxmg0NxgnBVjKUr1LH/VLbU4+/0HZE/jprud259
foywcVp1OGxLhaWdDLuqg84+IacZ3o+jyNlSOHmYecZ4bvhYZDUlnqiHrHfVtZP2ntI/1kBLNhqe
8sRGQmvyB+JTbSroUxNFTriFtl7yGUK1CldNs6W/JD0bwdVfJ0unjyp2104NzznzM/viP77vcSBs
RKHtPCrztG0rQxoew/2kMnd+22V038EU0Bcwcu+uW/ZRSSbsmivp9YY657qHYEjT/xtoMBAdHPuO
430H/aho4JZ2rKXi/xrZAXPHNquGyGpj8F2m+yOQZfgRBY9GnP7VjEnXqY4OZ97Ygz+WCEbwZqC9
mk50uHhI+f8sb7lLUBfwfDQq4fWtpfUH+I7KHN69T5/8vHcimELVh8aNcjTgL43jVbRajfUtGeFq
A/QG5pP1/WPspsz45IVIBz+fw9T+vb/lafUr59zTIqHn5Q9PtB0WWJa4pX+yW/hXRhnZrat+UQ2o
cQ9sUq5C2vk/EV6El3vhfYYpvNYTMuYY9/JFuNWEm8CsLmRPW3Y0Shgw/gs0aZpslPQ/rzz/enb8
BzfSs1d7md+++qQ8iLpy4+sc4hjHeabKrk+ZHhQWdX/DTF6riJu+4rzdoPXz/MNzIFqktArP6sO+
FhJQQUI/6ZAFLo9WUXeHAmHZkoDWDSlaZnHs+C7HW93gtGQl8VxoD+sKgVRVEDBxpenRZLVKXRgV
ZtNqp0Hb0hmPIJ9qDFLyq/f4kyqHDRYBJMuG8cXU4n0TH30dDToXbTta2K5kNuMS2cUX5OlyRhtB
JxMfe/gHw1NL283jrBVelHToSgANO/bA4vmCnQv3JCeRJ6TS4mEZYbAHy07gP6dbhLLu/sOEzslH
SHw2lxwtSt3yGe0PCKA22ytZztiWgDFkQIhJ5btiFiTzI9l9z1XSczjLozTXcbZfm3Q+J8i5svTt
QjkaNYovzQcNfErT0shyLtMPLX3ZOeJq2TQZUe+OsAQNglJQKAHkZBDe8QBSP5mkF6QXXthW7IIK
/TF2+91WhDErHE2IgZ4iLrZlcOej6XXfy1d5+3oFN30Q2XP4Ehavu3CqXGLQFbMnK/BgegP+pKfM
kj9AVFQeV1khdwIZCYvcmNGfckBLQ8tZFDqEB4lq0lHFtYcfkJB7zBVRgSbPoCH3x4QAg0GgimEv
nMeOICUgKtWss0nAvB649DGoyHBE8JJaoEQ1GDh595x21h4BQXoAzg6zuPYI48ib37iiWH27nLXC
OfZw3poBXgSP7rKQOLYYv3SUbs20d9ZMLIedbP89uXBjVkkFtPpWITNuU5Bh0svtFFtBbrdtDAbu
sfniSOHNGjcDctKg7TT96eM4q2+Qb6td+Y44960zixw+OYxtoykIL1mbKUxYTRnURmrUU/XjC/rJ
y0s627lrzSOGwA9Fu/xLbQxbDhdWv/p+UE3bp2KmfKG5rI39faxYnOezECWlTcWVwKUszTX5fDWw
fYyRdFc3OSYwdySe4dayI3hgbHP9FtoFm2P357hsPJbF28KZq9mpBLikbSQtqKsKCLHkJcg8tVtl
vU/RXwMeZy/XOY7MmzcXZWKLEGB5FG4SBPId53j18dUV9/it8EsxhF0rF7GLMRcTPHlufhXhhNnk
4apw72YkZuwun1UggLl4liqKfat17dGWGJGhXGbY3L5RUYdcMe3nooQ1VpMFudRnWZKLn0ulD1Wm
Bv1tBkkW/rG6irh8MvRAZle6QfBj+fMJ72S/TMGqFc/PBKCPyFhwZ3fJvesOUkaxQp3hb2yJ/yv4
nXokOx3F3GdLLzMjIbF2/3SGNlxcWvIdHvGWDA9GZUmpYzGSJF9EOr6yDo7GI2/8aJ6j4vIkcCMk
xAPcAakQFO709iBACOZIEi0U1FUfKz/+MAjiryJAo9MevzErWuGZ7x4w8rZooLD6VVIN24y/R7p4
QelcKDr+nHwSityvsJ2mItIvrgQItoWg/fqKS1NO4ygz4m7Uhf6q47/ZBmu/DUuoDkUtiu3AdFvP
2ZVBKJiMxuhr/qbsvYP20akYLgdaa4XnKsHu2mbnh/+HeKOBX5POzj85yLNkvtEhHyzTlAbtmz5M
6ML7AeIDL+nQ6pojoagzjiVu4pbEl445CiKJGAF4rIhkhH7i8ZILLSGQAGudvN9m+V/6qOIqSzgB
JWSGc3jrEZXaR06GZlqrZKeqN2gc5DPaMfE3c5pOmwg67NDA+/O9JXX5jGqkcLCGSV9l2DEDVFhK
K4G7ifeFDFefub9XoEucg3GFtbbtZm1TA55ABAqjc966tYEAcW3gzWTeWEHNUxmnHAzs9viI+j5x
NcN68UCaf1QgU5gL8+7SQ8TDR6uMHWkunNIV050wpvJ80Cz9zsJBltP8bb0orf87bj8WG/htPIkc
DRkCMfNuaOOUhnabkdwS/B0KKV6pvYjR+DOQ24BOysypcTFsbp45ChaXA2ylsRwRaJ9iiqrBNHzd
tSYDHwTGl2BBm7kOcSjwiZsMQJtkGNyiiGkP/wpEG70RP7RBRKZRcQHiwRIF06LC5rCsjqwx7Aat
FiN+OGM+qle8W7aYWKV19sm7zKbzt0VsUiCs2VfO/yFL4fRpyT19o8TSoMM+04zoqDLIuhT/SRA9
Z3qjFo3MO/1seunrPiB13wItnHD6TURZIOZ9c0eTWqpmHN4MB8BQ2M6Te/d8uWqWEt4+9e6NLnYf
xRKQwxolZ0iLiMz8ypugxbRdm4c2MQrWzd/X09jRNYwqPTapoWo7po5krdCxmtURypgHhy+Y8JpX
6buhA1Va1nf7e9VsfnRQZ52VKSYACL3HgeXJpuERF2pUSAszSM/+zNP+953ENpiPpXQsPST6t2BG
QTuIwUOepgeB5pNV4JgMfd696zrHiIZ7njXwKnbdyOqwlxDJd2I9yTOet1loA8o7PDoaCtahcrnx
Z7li4ljPVt7dlu82Am0HT+Fvs/g8S7P1tqTFSK+rI96uhOWODakimwL9rhp96TB//XBM0lM2kH9Q
2Y2nLLm1KVhya4elwtdw23QqYyDFVWvjZ6bMEiTH99K19DCYaJNGG3MhxP5cHld0EYhMj6bHG23A
8m9m7J7yxYomiIVvYDH0jwdKGt8JZrFbgzAGEMVaEO1UHJ9qFNM+1eX13gtBk8e1mKus4Gi80o/d
yC6U46rUqRH17CtXUko9JHUx684tsAb2Ns261RWA8dZ8rZHjynLzXnLnhFfr2DNNWj9XG7NxZipd
otPmgiyT9dmj3ygrxtcu8SK1CZiLgDVlf/J0RKq80E9d+Z8RR+D5xsSjcUMaU0JqOYSb8g5M+01N
YEFEGjMuj6gRb0D/7MYBLBJIVpu+1NtM8X9t0kgZRaVu8Z/dAY1jNlXFOSVKlLvKVMHkX+pMukrr
1ighcxOwsXDKcwqjdjT/edVQacmqJk0h8tkPmjzxEdNXIhzATBmoMxxAoB6eJs8D6pkXIlieoUKp
UuliNXHXes1+MZxtwIYj/jMqXq//HLx9yS8aPmQtVq/ge9FMarc3LVxV7HDi0p+D8YO1ukptwyyD
3HwpdCyWGOytPZ6T4pvGQoih2nK9IcY3/8buHJ27/onkofeq5/Otu9Sk3ptFgFCjVdWFPKLUVoNj
kpZzy84v6LjtKBoZwnnoPHofM6kzXfRRftyVqi+e1WwUkxFNkBXTIZ0aSY8NpPN6O78ReDJN9aLO
D4n2YHCLbXsII8eVGpBW8i5CYmfGW1gYftZ2lU6btRmPBBi8hFmOuKZ0fanBGYitxWewnadF0El9
9qbZqk23qwrLDyRLiZ1+jQzHnaQ1O4UiEsE/9GQDqFxD/7kQH3+8Slo+ZQx+46q7hNGYRxM+OCrk
uUdKtwXW1wI41Byk1KxCxnRfcGED8Epw8xGaYoM2gFdemOqA4Rj0mQbrMPPUAToH83ZAXXBBil9n
g0ke1B/8Tp73L6hXIFOi/VSfG5N/6HtGoY3vqeTxVnq15L6p3T85Huk1Dr8B5KySVAlxapIvAh4R
cZ2NA4KuQjqgGGe1/48jIZ0j6aSKs617hTxvK5pPEa0p0HWvCA+uXFHT7VCiTJzcRJoU1U9VMiMP
1C2BQm3ZtJPexkKNzHcQUKnHzC6A4kNh6lgGc0BNUX1l0Prz9mB/WponOiUb7kjk2fltwF50DKUP
ieNYIedIko5do9edUXRL0DHtpSnXwFYvzCtXdGiiXRYoX/6H2SCl6gZuk4Qlt3QoorYxdv0cRf/B
vSEEVCCMIUdvPz6a3c0b/MwXtMXNQhlR6PXohrRJPMamtK3/gk2t5qkvPYTps3F/t55GtC9ZwU0B
13o+RD30wlkYJsIFW42A61YineHJ4nGYwXAMUQ0Y6i4tNGcrI2X649iG/ciXFvOlaF/tA61qkxwd
gr1u9byc74evgf3ceJ2jiTR++j8t9s3S9pzJkugebnBa3ypM+XL4KK9R6W7pvz6xIgqcs6XxQPkp
/onLds3AcPAWVXn+T0gBqFiwcX1KpBYgWSGh1Q0rHwlUymoYPAzlt6G02fj4mr+pzjfRaWElCZ90
ODJXUbK120raXJqotn73+tPLPOKsJuEQYpzgihcL/sj7qRUrjVlmULoWRKL1686gjKsYCeF7kBk/
sSLLoaBwv4qLFdfDOHZ7DHGSH8kIcV3PAE+9D1285hdASpV0d943VSCzS8KCj3Zkh0PZXT3sDt7O
MX52LIJrJvn4susvLaKrJyxgap9/KbTa+Ze+1Zf5iBylBeyqUCHh/pVBiC88mAFDLXn1vRgaFzV6
oatHjZI7eDBNBEYJV6lMni4DZth8fb9SEsdXTQsvPivNWxm0vcNjlG1GmW64yqv/Ss87HPR3f0Ka
YnI3C90EgWVKwBgQySmpnbpJsWrNpRyjYtEg/7oqwSmJF0wU8hpM6+Q+uxw/CylhMNqnqLSH5nt/
psx5nTVCUlxRYZKfcmRUaY+0tE4f7Ie3c+5XGrDISud1c3CzkcXtAv1M2DN+NcG2JLbL09w3ddGm
v8XMGIXo68yILtVTgnUbdvJSRHfdSOqYFGBNIXHw0PK25t+jFkTvrleM4fre6R8r1bJoL8yW8o11
FrFXhkY8iBq9+vOyu8qCTHPwowxfdD1itfrxMBmLS+NrlGzAF4gQ7BZS2Dd1Bv3+8S/ybQyfcnSY
MO5KVKRlwosR80jr8YHr1oTloifaw1btFvm4+TDyA0YUCi7DpUyPFY/Y/6GLIFsZQhly67fIQeiz
lu2VxIrmmhpJGdvmpUaOmemaUooRdWJvb8EXGfUZYOuoFomGcnkyrJuJcT4cBkrIZ9VUZHa+OJbH
6KtjKsU/tqy/i0f4OuYqoDcSzC7DFD/DTQUWAY46zx2VJk4AE0+CQ9HKwMTKB4pL9K9GlDJV/Aha
JKE+4/NhY4adCpYl8ERWzRSsfWf+hzZIfmy03ZYOpNaRBw7kPNHsIZ3tAmNANaDvu99QhIp8vhxi
BqJAjMlEU/wnKJiUjHsLGA3chM5gd9rvcOcWvoqmuxxKVeZy3Sz89BZDou6tMg1BjPFFHY/drK0p
TT6rKE9EeUyCvFMw+Cd/uXk2TG9qKHMW1XNuEku6iF3B+j3g3+CJyOk3ni1wxdj84uLlQ2SkeFuY
OfmRNd8liYhlLpiWpxpVpvbp3ntU0PGfvRmxVsEu8tP93uSREhUuwguyKdT2i2h2mZERkjnG3RI1
RAut2IeboqbW4cxJEtEEOp5vVyWOkTsmtNpNsazM9VK0MUoVu04JnaOCgIvqxfew/2wcWCb05ltX
a++XcixnJpnr2/jTS+bvTYGCG4LEsMYUUqXU9a9841jgpXVqD1E2vgDjRfo2kiC2ITlRb4sMCnMr
kw/wmpJK78Tk+4KWV5ZYA2EpjcCsPgViFPbNMYmWTioNsis27Agnuyfb0piCMdO2/HjHDHWcqdOi
vPE9AZYMAhGnpJTWymj/fe6RMqXu+esmVSonPU7e+8SNX3rkr+ViPyb1l9HuZRml467TomU1865B
FHmDM13CzM6raDZp42W0lxrIW9O2ddYFFKiJMniq/7C67x/msn+xfBu41yqf4n0VEjKnD0TvHAVZ
S0duhSHiT9kY4gMKNwo+k1MUBco+Xdiahufk5mt6DTpqmb9+k0U3e3JvsPWqeQRjvE6DpQegVgkc
bZm5W6FHt9Br84UcGTcEUOzFRM3cX4gd9d1a6H8SMJbjU/OhgkECPPxW82bkS6U0LR6ok2gBJfmP
GBBMXM7kwgel70CFpcgbKvaQxUhuOk1OnO8L1zS0i0wkg3+LHucOZFnGHaC1HzlZU0l347Ogejmb
ZvxWF17eD2NQT3rWTEME6DvSwSZsYlE3tnPGqDAlTlEvAKh7fE1cFZH7bh5RRdtGBVwIHuPOLJDq
AEqg+slbUubrcsL7UrpjnK2VFG46isyNKekVopaCY4tz9ayOrF6O0bh6A1OX01XlkbjQrIYlZ6cD
QfwI2os6xn3F5W6bpW2CD+2clWvGtIQpn7v4+Tw76UN+OAE0mhEOfB/dpFu1SPr7/AqY7Wf2qDSj
+dDCxX2FQ5qAmqJNBcUCxNwaY7P+N89vhBZ97PozoxSah8iaTFiA3OpjPMNGx+ZzKsSoi5/kSSR6
s+TVfL9ykmaPb4g7Qu37LXJrjg48YfSQ+e0mp1MuDVPgrayfwWurRDg9FyIeCt49rJ2uQ2p5WADT
tznFDEbY8JeIMhvvFRZKDVtZkme2phrpabrHxaXF3CUHCfC+T2Me0m8kKs+vtCbDPLactXy17cU5
zexa18T4RrL0zcOKWThHzVqWZTXQdjgw2Yqe+PbiJipDSfU8jUtsigbET/LAb5/ArnC+wzj37YPB
S31QUPL2qSUPJMw/+/W/DlHq4zdIKEaLmTxSv+lk+zbQBKhqnh8dpZadNc16EgJpHTUlMarJnOfE
ZWXwtDjQpRNIhiRhSZZGtyU07kEAvdDu1rCImQCTk/prho09ASkETenFhSKY6gm8kvFOlwKwT3ai
uKPs8mqeK4sQSk4etkYp3R0m1eYYr9wHZomduj/ijgMyr8bSq4LkmPyNIqJf4gEw7x3ZeuoAIh+z
rSXZTERBdZRIL3nlH5qZO34+zg+UYVaCrO4kt1DTrx8wfrSerUmQ/0fDSJsLJoauXwlf8XtijCOR
xwX3687fnMdPjLAX3mx4m7Ku61AF0PFS7xOaBk+9tkmPa2KdguS+1+CMrOXVzHngPngHqxgFvXK0
0EdyfeujTor6lSE+l643ljJWhG1Eikmr6pQ4xI85enb81tSuEeTUCT26cMZnDcJ3q1YxRQVTQtCR
ZKc/APQmdc6uthXvTlIg9fe5eZOKN2XWp0GVZCEJaM7AqErTJAH++1tHx6OBjcg9StETHoLn0cKQ
1uQ/p74v8LKTT74n/uRfZX8AbQpYqcx8JFmBQZLhHBcw2VJIEa/ERGvHE1ET1umSIUSHZgMA//tO
9ECeaK62jQYoxSDvX+ZIX6QfN8SxCEh8Shy9RLsf+PYgsNDs11RSXg42bBUOVkmv8w6APKHGY+ND
C8YzKOjU9R7nv+D5RvuuMLPGHlSCIe6OCGxTZrkRcx43r5BudNdZwVeaIe0Wc6j4SbYPPDI4YgqX
cBH/L0hvHDTqNtgGlogk3O5EkQFYE8dA7AKAOixmE1Zi3yKNEzpepvhgUBNYX5rvjcWK1qQPF0Zw
JBKG2X+GW+JqS+ubt4ngndZdfi/Wqktt33oSXU8Ve44P++JVrYrwckFfO26keiYYszlekosHPgqK
ov21ypGDeEiQc9HQ9EtyKZe7OeXcnjyahg5gYghIZwlt3cBqbd18g6Cc3pf/Ykm4B52itlvGE23n
gxBgDQz5uUthObxzrVpjcMGDrIYGrq8osyfVwMiVkbhwKcC5pI7PBLrx2+FzndDEYjOAMfKt/K8f
7x/1sTCl8OUk3VSRzmFyL8BTDD8VqtSSLQyIP0Jv/JaT/WkxIDzpFkebgZLJQiPcyet8TKQMwlV3
bOpkRD5I1HZ26UO82gFQDANrgrhfADgEQSe8fBaSEXZKwc7T+nHP6z1aFUKsDxn8qVeV41UEwkf7
3RrVbJS1XIr+4vD21fdIh65PvXjIUS00bYpqUUyoUrVI3WdEJSEVBu3HkbOpgkbeZcf6Zjq9IHwY
gxDCuORqLH1d7cSW9SQNhdrTyuP8NTgqMuqk/uM4RjD+PsfR155QTyxxQoTQQDfbN913gn9jsis0
jAF/EwLFfPofWln7YTr6pnuM/ytUjYt987P9QqtQ9EHTpVMOSAGOL0Dcdv/O+xBlVZw9LZbQii2N
odsRKOBGkqoZexso9kVG9JEpEyKlmKfdd65rhFSIOC5jEdILZtrI+4jfioIczsI/4J+hC6Qtw9QW
bz6e0ZSw8e56GiLo+0WxsbP1GrmQV4chvTpciAL6w1uw/Xo4/W7aPi7hD2hIB2rIyF2GR7wZEW3O
AFWocsUZYFxoBYp8zydnossWgJaRGUSo2w7OahNHWxzHKwM9Bk3MpVrGgjhbX6RlrAEW+4Ggyul1
/mkTXEL1PmjEycynz9OzJV7BJnAUzarh6F0j2TxKpBE1rHpVBU7XIB8wNCdCiGTlZ1WaQCY6vdPk
z3zlS7uWNU13yWooOuRP+LoP2IIEefHXkW4hwSWRYr9xu7T7MQaw8grJmPuN1gw9FUdIEmtk5u95
KxNmv/zH3pfxbtvJDtKRBj87vAgBPXWnACxfBjXbHZnj0xduV/iVZA3QJz6Yb8VAgfoWfjfCHqRW
X8BA22x++XYBaS5Qb/xcukOnxIw7bEshzuGugBMhItGxmF46jWAxGR8zEH8FnsGUWeunW8FIZmRn
bJLREybpdNZYfKYkas+OgvE0g31inmTlU76LO+epwq501zMPgkcRMFcE8BmbXv+YUAOUQPm1R8Xd
5OXZ9PQEzk2k327ZIci2KIs403RALzKZnyjsITeAhbfrBK0ei2DMiyvuVd6qp9H/p+Mdaf7Z2DUf
ntYvAsFUdix6BuR5TUK0Uowx1U/BsQR3HslTSoXeTtvbzJKYhD/2vK1fLQRREn+6JDyRe54pjqNY
ROv/HsGhs6VNZ2dTWSFq0/odAMu1wnAIYXi0iMSn0NRfQ4l6M7e/K40nTn6Jw3FyXb0sPfE5mo55
VhrXvZLBXg+x4rXtFstlWhHmYR7adJJKyKRL0s3ccVx/xFePcMqjzodWVjnV9JKSwq77TmAgVpnN
GPaK6RQZsRxYTyciuV9ST1jUKy5Qmk3lyavGEuQN7f/q8ZTew5PxYRZP4QV45w7qeLa6nqtReeFm
T8akxDJaW2SpFIzGrhbyij4KVMCR0FwJHqWvDP8JOgnVkhC9gwa3/BnzeL+LZRUHgaBm6Qimys2C
/rEIpxhn5SnIw9aKnLJPI8W/PKPVuK6mRewoVMYWwyfGl8zdgsEJcu1xpeS75Pr318oRp37E613m
/7ROPMMW/PgaE/IZZphFk7R1KRtdPCW2pOQvar0sIyqzNAgPFeqoR54XYP0ZIr+Z7dC4SeR/w+TK
KEpjOtKIxFAmQJR942sHZWh3dEwPVivg0wQCUj3Est86/WLMOjZ1TbnTilr+ada/hW+QlDZKWvZC
7F9vgNIrnc62mJV90Rg2Mgs1dk1mMgC3Kh2VkN/TEsCc1eLdWLMLoMveIyZjkaj63RheF9cbQUVG
H1Ic4RC33aOdK1ZKDAFm2VTWQJS8CPq/iA+APdUG/+upocq7Mbg1e4JIT0SCFiH0jIQEgXaW2MP9
5GW3pAaj/velS1uVbaQACF1AgwX1Nxy3SY68TkPv59hiJRzcFCXduBXDSsrdr7y7WXiztIEKqbx9
QM0umlInOswYmULZ6HaPUJsbSn5J0sDH42kz39c8x0NTUkTud/qoagloNotVanrKfV/Q/ev05Mk/
Km4WE0sC4U1alWQzrABV2SvThbUVGXpP2CCfxxnm/tkD82RoSFbQhyo4RPcFWgX/XB4Nxk7P9etB
cB7tIdhx6pGkVFVLGUMdQI0qwypK5JN3Hz4N21BKxjjp1Qwsx+KvSGwZGRHy1oBkgq58lFGwwaic
VgTqLVdQ95BVFRdb1NAg0p/It51rnLebW5FL55mF3DNccQUmoOfL4MtYo3wqFOpcyBeUxZQzJEQF
wZsqhp1i1G84k/dIRsSwmbOfRI/Tq1/PtIi0ud/uuukNwdTlHQdQfausGcn0IVQ7tVD2RtM+bfAq
3EnWvIkpnsrZSxG2VN8njiNib+fPAmcVeX7FEyW8BgzvJhFRc7gEywbStbuIe9FwDWYv7P+S7Hoy
d5Vz0lhyIudSUNZid9RNvbKx/Jtg9kEpUJXJ4RIquSVN11gdAucuEkQvbpz7cGSEGiXA3Lo+Stq7
M3TCgoqo3tcGTchi2kKUM6OIba7WGZwKx++4nu8Yeph7DzF0nehFAeoxyU+Lup9lo13jCIVSrMXX
0rQ0Vm8P838ZmjA5D56Zx954rPT/F0OkWzG+iYWv/hITr4jzicsDAv5CNH9vxFqqeu1cl2T4eLPa
2eptznharmyYgUhavxhK3/UnuetM6nlN//oWhKBnjQxJMfsV7Rj22jlQxT2kwDsC+Bs+uFFY1E2E
ID6COe1bMDRGVJH9e1Y9Ok7c3WlE47XKjXFgJx1Ln+QXfnmx/MKBOkguZBv/KqY04gD07jWEWNIr
ep0wdlfpjZdCSUZIruHltmxCFT0TUw2nDwQtrgASBjh8tcxw6c0R3phXCQToaQV9GuOrTS/6c373
v+LhWcZBOzAmOyBrjcMlIfkZunFKkJ2wA0t6SQq9C27/+A1oaM9jvjrBuXnSp+GoZtU8G40vda53
zkkMAvmqJFZ2IRzyj9z6BjCzXYiR04Zbhg3MK4TOpxUmlLpeIsHkNevestW8dzAUlE24hJno8AuH
oc/O57U+6LV8qVj64I9k/6ThjA0K4oIE1nIaJ+7PLwrGvfKd1BeJJBni11Mfr9K13eExDhmHUVDz
59OSu5REjMAT+jwmbGM5NRsiR918nb67CjglnAWMYyWnCCndqcXOmfpD5SGFvOADDjTUpOzGiN9I
LozS7b+Hgce93535mJCSxF+VZzeIaRzT8soZWg2AVJc4lyeJAeS6INPECfV/U7D/gobWhjHkTYOE
BLsxnBMk23nMKkcqB7JIwg0lHCyQm+OLYh1nuINKZVjniq0OlGenQzue7IcNCj5GlZ5cTWIaq075
SzBWdyPQr8qw88g/1lJk5nEZRe10ouHX6AOGhCjGoLsREOwMNrVcCAdfJhbJar0KoeAZAmE3szde
ETRe66NGGW1R9SnRvicSMTgg9IfV07z2AOTiMo7/5bHr9nV2zhz7UlTjtT29D1mskR8waaPaMnZb
Z8b8ScDqfSLq7zJEYt8UCEAU3flbRcLUMYUfx4Bmf9JzjQAwGZ2AOlPP1bbw2ffStxRS7PNK6vQm
fS4kSE/lMutugBHDSFakud7gc4tCv8poqsJjG6vXUjojc0X4s7f73t2ikKKBNvJuIAveNPJ5YJ0Q
EPdd8asvheKkmc/w8DAOoAHTx2iTf+9BApLaVhal0bv+GaIuH/SRZeIkJOo2B5BVIhYFrk4emCXv
+ftO6XSdH0rMw5cOEEPnzAi0hDxFlLC1FioWZ11uQxLS/+y8l+SMuRiCvlrC3nZpF4K04oLOqsQe
tZiXJnyhKgeicNDwclR+NZhyNH2Ac33RquHa2eGPOKcbq0OVNluoQvFiDA6bQ4MFHKWg0g9LM8t6
9ylJuYoEBLMydMnJ6z5rDqNAyp/hrwBOn8W8tcwwMflb6Igk3iifXCJAuYW1qfevYchjEv9apF1t
UAEmMyuaLDeNGzOUCB2evtifC5xkGkbTJwO0NU7eQOlTTD4Ih6IdyzrGFhEevRwFpsZr3+Ie8Csi
MgRkUenYNLVhqQd5MhdKds0TcnAwUKSnrsKYEr4yAp4siipS7AjtiRTcmw+NifJOYCRJUBMXT2Mo
2ZX+oKgwPchKzDBGpQ5DB+2YM+9xLl16klk2N40SuXNIGwKskdNs0f6bXsrfl/VI04Yg2fbD6oNh
vTYjUbBAn90wdSdTWE4XIqapa7bxx8Un7Y50pYu79JXRsDP0ltW/U44ljkKM5/DH6KC+AsVAwZdq
kWOPpzQ4LcaBXzpo6u1WlZDD1fV4ZjDNw06YAEu/Y7s2PfqsfBUqbkN88NrdIh4aEP+4lrjZ+6Jk
ajZbonanhEqKbNCdkCPdvj59ibpp+2m/GxJapOjevA6wp0jyZxsYYHGjdkmBDYEUkprt3ltg5d8A
k7qKCadJVYmmh7ZF1dyVFy4xO+HbrGtUAFWRZlPmUdsmGwzrlZS03MB+JIIWDWYWPNHdGGaFTGAW
NniTsDzV3Zny4qI+wg6Fe9pzQDDjVF/7Mnt0i3SxDElRuNjLH5H0cMlkAcuaY3YRrCTnxEHGzkjF
Sxu5DG3x+RzWNQN6BRcqeDOY5AQnTp2Ju+qoxKKm463Ok7ePitysJmwjDnCZVu0mrdB/bUDaatPx
sc2RI/u+CjZasQ5+EBs9nLERkVV5gL/dyQdwmItuM6Dys784qiiudWbkhbqLTxaCPgv43tlPjVTn
IEmvWZa9OVXdmtcHu04MnnneP0C0sLuoTY3doR3kPGHHmZPBSMIVTLy/lwfndAdh3gLM4Gn3OEL/
7vV44uj5fTEPrfI091ns+42OIz7H2sOv7qdotJC2mul/OorvuCEkQjeFX+QqY7rQj7oY9DvbMwNV
j66DwrH5FjDEnPFmT21PTB+zOHOoYKqjOgV3GQFk5q+TU+a/Phx9mcMU33COA0UhIZrgiecOK5Q3
puJx0SKdOIW9hz2lt34qdjkq53BusD9B3Ru/wAEAaTPPlq/yGG3HQNWM5yNlU7xSb+mDtP0ZsLh3
jJE0w93ENjCdkalwHObEh4r89+g/omnY5FA9rvJ6dcorlxMkfGNRhWkaHLBGlxBHUMUHVa8OzuXl
NmIX83oYflfbC2DNaYDygTf+fu6z1Du1gbCmmKOvq8tUN46r96bentfpng4pjlNd6+sB6yHXQFTX
EDBYsqYI5gtgcPO1HjPqdEJ7l6qSIh+JOET4nAH5LYoR2sdAuAlpObQ72oHFMO9pzzTt52IuLFcz
EeiEOWTUMXnOYSyg2m1gUXcSdP9r6039bBPfx8/6/gOuULCP30yxRa5aNSXwQLsLgWaR/pxRkTRH
j60V61TzFQXrCHNSF0+IgqpNEVua60J2mt7d8xdp5rbUeQ4k28fXgLqswIWqEtnjOjBZw77tUuXG
Z1q6a8nuCULVEv7rZieQhSLhaBNLNPyYk0hc0lE/N/g0KTNVi7RQUgFQxHhYQXB+oHLfOyCqnb3v
/zf8R+Ljm3eJxpwuprInN7S+YIxpbMmKy1dt2ON8Mjeo75G/OHGN78wu9AFdbj0Ify0/Txmss2X8
uEhzonsCLEiCHSspc3ykowO0ZuF7H3nLtYMO+DIcn8LCIZb1Nqva4h2BxdAku6r+4dL5Czyd8p0X
nFpwHDMVv9tpiC6XdHsOq8nvD/GTV+wOEeiKvXQJrpc/C0+G0vrQA+KNo7FCseCJC0T/PAOy7VPT
+FoIetvWMbm9NsZ4RS7pjC2Ma3wkd0KM2q8fhdLeVgo3CfZ6K3e0lP1LFpDDtORNaGvN+mZvkn3U
qaUk4+fcf499fUpHQaS6tjoyPqVgoStwP5OTvgaRCdbtpokdNf2PyPSvDcDD65KEJXtUZ+ayLup7
oUMr56abGGP6xqnfVCrORN1FOKKOk1YRrwGUWpMXyWyPS+EGcpOKFOTMgR0/sThdO/UtHFAOqmVX
ohjy6OFmOitCO4xDBTpZaqzqzjdSPOvtUw/oqMp0eReGESJoriAYIpsfrsY7T1ARv9cmyk2g6QiO
dMRIPrzWcn7JAmEwWWrK1c8doNLnrub5BKw2mtBb+hAAke8dNvlIXt+OEEcFZalgYBJcmYRcL2Tb
L+KXk1n7QwWf2QpOflh7dAuHxItFDFf0vlaYuu6dTJWtHn2KhqzGqasxL4PqD7jJwFMF0IYtgISY
8rHb/gVMPCzD35bhsCW7u/pimUutfa3lRPgnOjOZ2ILpY96WN6OUYVToHqntqpSohHaJCw1p22dm
qftgSkaYj/OtFXMx4U/NmoW6zWcn6dCQvGNLoq1WHnZfy+R34CdfSdVgJWEaBI4G6eK2lgL7mdCF
6ZCYlxQUTG3G8oOqQ8Wyt2ITVmB48j+lAyz4zWkq4FTD3P/+HDM8vYmRTR4TxanZmKK5USfX3XJM
f/cJ2e52IwSMicF2j9URFtk7Lm4XYxfXIsfg+ErID6n9hXgAVvz20Md9cUhSXUOaRcQy2iR1qJg9
XzHfvNh2LNVd+GDiAdYQFk1zBB7CaNNWyp+HUxCKrx0Aa5bX8cat9TKZkKr4T5OANdTRWlIGqj1l
n7/vDkIWu2idJqRE6VLCSJd3GUEIfRHGbsJlHAtgf1z/HA03aTsXudtKnIyWoYuXwPbJiWDq1+Hh
b16XEezb1zxIonrWPNrxTx+Ylv1LLxilP8R5RNEyj0QQwSr+u6SouNpBgpyQBa8cY2+Fm+IYeppm
rpckZVlrWFJeObMbIerqnxnvuigETPUxUWMIFsw+xdNppxcp1nd5eKwEx7jSjOMaBeBD+ks92aGs
njhTNmZWdCFodq0xVBSCIkCdqa1xEPe7eGw7h021tpkMtSalpobO4/1NxZYaJkw9w62pNYp5Jt26
up0f0HZfUcIDlSeknSTwv+C3nxbHuZwhQySTSAFld3M9z4QQknSn25wSlfE0JCbpYOSQRvbWDZRV
wyugsyVhTFUfwh4hrUOjvR2F/2I7uT3bkv65p0NSUbh7c61Ci+JjLXAQaCO3Lg+dk/0pDCtkIHQr
IWp6wb8AimNTQWNe9QRhlLCb19A834pMp1vRTNBa7B88qqcZbK1MhvgdQBxQTitFeupGoAppC9Q4
AOIHK4ZOKL/YlUsF18IEn0C+Xo+EMPc4WIJn0VQY/9rS/1XLLx+8QA4a9PMUqsdXh0fHn6EIrv9I
EERWbtZ1Vwgblu3uYNE/RWoF3WkTqRlvihSDeCcxF0TwWBLBuI1C6WFimIKUrwe+S39txM0RbOvH
lFQVvQFDx+ng2SjUy1rcGDWviRngFvB7+se10HNkbBewg4JMwkOb8fQSM8O2DVhHx1VIOLtESIjI
Sqo+J/5RF/2NxF6HZFjaD/dFuF9myJEUFM+r+adR2uS1C8DYYfuhmK49pXlJGTqJLcPCY1A1ISM2
aohIKRcrrEo2bejeIte9XPMZC7aHUq8xCNWSgLvTsCsVzmLTHeyM4Pj1n+ZLNZbpbSP1STq6ASdf
ysx614d2s7kSjhPz9gQMWOu0dSyN19ydpde5SABJfivGrY5ELAud6E3r6CFT+ASKIPgADT/q7VyL
+wuHoTjZejjZ1+4fxw6sF4VKYXGXPGPJUoGkE03Y4n3ZFVI5+FyUYlgTM+KizLP+qqxPPE4pDdYj
WCJVvDhRabAjx8+jsOjViGHi6BLxr5M1lkKbGILAhVU3zM66Y2Hq70wuHcQwe6fekae6Ouh20Vgy
gDhMhaeM4B7uhEuIMi/T+iRgzPnLXOOnfKB0oOURcpx1OFohVSdLbwvTvSS2q4AaduvGUc+iBBQi
kBd1WgBq3MwSdsrXcTan1pTNF0uZSSgs1ah0gtvng0E8SwjLrHa19bEF30mBz7FtIwP2ocJ6Q6ty
owyo0mi4x+G/gca0VXF4doxnxxOadfB5Q2tUsn9sFZk0om3mBOyWrysw/qiepeAP2LMudXjo6zpv
lAtNvWWW9c/jMeBCK9w+iUGoTYc3L2RUbNWPRHGs1CV0R5FgV/oIoAYp5eW85qBfrmYJ9uwRMz3Q
dM9p8yTL+pXFcVVd+x8ou/Mg8oppLNFhSdku2fYgoatIcwvVjsIgGKe5lufLoDG2d5jzVsQtuY3g
F+Pk5RaYzRPNN2ijlnUxu+n1m8znEu+NM6ZT8X3xTh3+bwoERlbVw99FGfbpIe8s2s5ZQGsmWgBt
iH/3hQbW/VJtRG/jvNjw12xSngvJUpa1CWIXJbTaA3IIZMVrRW/lgVBBhTf87ZWPRsQrTN/AbNMP
c1tsLcLTLCxactejAq4nua+xMc8Tc4rYmod8YJR6gzAnKnUQKDQShWRfm/FXaWepTHHo7Y3rtNbR
ITACGSwgg4T581206cDOQslX5zEpkBf9Sf3LZym8r2w2lINzBZRM1QVOHtyLoH0FzGUj0Xkc4MU5
7WuPsdDZTaUAxc+lV+gIJCq23bbgVKSvf8oEeIsXTsjx2Sg4/5x4LXowGLhoAbAGFXPp77qxBAY4
jFq2pijAnB2E32qMixF0MnTaXljU2IChJzULZJ47v+5VrghUpJYixa75XXrTtyOK0qrdDCESRDFW
SkbO824kl1u/TIcAzFDsS54sC8+kq6+U6UaiHNXEfbaJ8CrNIYLrczL4AssR7BnRcDypUtd+n/wF
nSzmULyAjCfkEzeqqN8ZgPO3bTh8vZBdYxDPkbr3xtM1YY4yl3FzAv/NBNosq17Pty9yDMYUHFAj
M8LdaZS0aU/83slJ0xC7u2sbZbniL4H4eQq8yYBkKuDpCEZCOWxNs9HMphJ5kiyq36eg4RotYSRb
Wlz9vhkuY5fo07r+tjIzztRcq+VOJDdmm4db+3tBQsFVYDUDw8pSo9h7IFPBXOx3LEY1Xbv4ROWj
BpZSMr1P2jOKyUkrleDynV7w6C8FSlJx0Ital9QEzYFQ7vlyNg3qXlt0JsiTEmAQ2y7f7GTUhwWU
wGOyn7+poHfa6ODi+zGY09J/ITNUbDTsM3ILabOJXS6eZ823JmGqfeEnkOYcDts2OBCLl4KqhnaT
zCjANN3+XTlao4IG2v1uu+qJTJsIYy6kVbIOouqUiDh+Gvn6rMriXWiJLJxI31bmpxDXJ3/mWgE9
N2C/4ClxqMZaPM5LDk0sBeaYLhokoRJxMUy1YoA7pieSNm80pGCmTSKBe2cmKwKiitK+bQ+1XiF2
bGb/TKTFmP6QqWcaYq4I0xCLhs5ohkd0Nf1ImTiXBSOeBfJRUA4qgugoryJKxz4RcLJ/v93qpEFv
LZrKQnMQj5VTAAYFX3NwBU97d89kmw9okHOz1zjkOBgKNUddSb1RRETUNsa6R+REAdYU6k3IZkPo
sjsKUdRhNdMjym1c5PYdSejlC5ggZYXrF7WPbEQLZror6QgWSqfmjmSdLhizN8MiOqWX33yDzG1m
Z97jmtb+WX5awiAjMGEy9yAH1pPeTM6fcNRI8I2VRBbr+KeEEWfsco4UYB5IDzkIuSt+d0q8lG6u
Etjij+O9DQoGTp0wxFiJ2nKryRd8K6eubQC0c+Mi1TxHWV6bq84+cXd+zThBDsoyFt4WvKO/sOEj
OWkAXZBsO8ww906fT2BjVRL/amKLLKcBmJIfA4HF+JrandEZL+fHMtBT2D7xmxlBPGQeh8/K3LX/
ZGOBPqWKcwAGRl2jfYAzJqIpBS5UzkY8rwSyKH5Uk5wibNBzxNx90QK8yQtbbWan4NQHrGcRBlgr
1hPt50m2gxaxC3qfiPtA3I5+YYw/UfkMK3RKXNNlZzyzNqydemzP5vZydWqIsXV4y/rydOLRYiZd
adcWeMFwPZAAiNs4TIOWkC/zO9XRrsLvqD66nK6NhnB8eS2R2YJSkmQIDHK0D0S2wDzKhyx/PLXI
Bt5zaAg4V+9I0Dcl9venilQO57IpK+UyHupz1QM/Ny/e6cJ8oHpoFMZytic/hmb7RR9l+imijhvo
NYa1WnEnnDYMWz4dpc2NLo9KHbiGzjeI5AzNKSimn2HiUHvHG7lJ0U9cP4P5zSmjCi+H1+hcA9fX
OacgrADsKQcSqGJjM3TRtPJr+ZN5tlCyM/lQZ+n7qPKfl86ESMrtVyv9U1XRrRj7sV0ofk+P9K8J
9iAvSdu+GEJBK93Sb3d0ZPwNkKWbnuVHbXFDncpWBI0O3CzZGKTyUZmtf2CnA/5PCQ+tPsdKKSkq
vDeZE6uT1f0gbtvUlzm7vjYgCPcE7XZi7le0oQAjCHuuvlDA5XeA4U5I92WZOXy6VMc/DGq1b2qq
e5lWqGhYhLl9JSDTWko6ANP7mh5V7wptLN9WZt7b7+Rnky+wr6Pybp2Y1u+PF1u7IeoQMv8mihpo
wzyOOSqVBkZ8r4mKyqGNXlO3VQulCpU3ZpmdlTSg/VN66184msY4QomFBGzb4kafsJmqX3gvDtc/
UYS803irQMdpdXSoWyJ/LKuGzgofdqqPkBMtw3URjGLx3Uu7owDfJ6rC2D3xjn/mSzUS9BKs5bvs
iBwytS4JKKTy0SKw2id9A6vpWbR2WI2WkEqVauisx7Xp5eB6dhi6e83FGY9BV/KBZ0hr39vrsyHj
d3mMDzotCjLQ2sxwL6+MTyw9UWjI7DRE/5AyHPIetVREhvuXPBZoE6rnmwbFzpDJrVGGDa9GVKm5
JQE3AoKDBM5aUN/+f3cSfTa/Q8C/GiRYRk3MBhpwf3QrVaSlYW3E8erm+bqDjW3cnJyVemSH3SdQ
9HkythILPcaZwGqOb0JAJcHgMwOordK+2qZWGNwg9X2f83qK0vt/Euw05h7Wd87Iq7XzkT6xdj73
w42CV34qR3+umkQJNHfGRbwf0Ich2Ghx1XE2AYlnTXzp/QngEi0VZR0Fy6rUw9jyRnjrqmgDZGLN
nV7JCgZuT+2Q2tRWPg47FcOvVdMfMr5gTcGOc39etL70zKV5Ur+0K7dKeDDf5+0NFEON2gkvbiW/
y+lQaxtlbLDDc5Tk2Sl27wfxRp/nGyisJJUKVM+Z53cTsik/YQSO9ZU1H0KGfGf15G4Rw0OstObC
UeNUr9ozvgcx1LPSiSSG8qZzn0ngZcB7/L2AhBLoof0WqvXGtjPQjl6mFa9Qm40qJ1GlBwh1k5HK
3uGyUDJC0z+lEr2Z+hhFLYjAQj73EhHLOqWbuIdEnN1+qFzII1Fv1WXjYS5esOprqsQj4a+8z2cC
035Y5c+jyT8tQiK430HST4crnJgrmc7XvjqHBO/NWmV//leOY0IOqmDHMsyzYbF415j4oT8cGcdv
2JS+JpnyAYKNe03sjlH44jFvW8w2i1f+OSvBarPfwTuId9KYrLmheJEOG6dowBo9q2FTCAgqHp7o
l5hapFIdP1u1EtmQytif/4cEH5IRzvNWeNwX6JaMUxPINuSONtA0HzIkgo1AbCk16UtlFtRHbYpq
HVWhLQmnguf2qTXeDawypFSNf0hTDo2wsJFFm7mOz1N6nyKvdyn8zBN9lhD/GwthvRUFaucPiXiP
h4wkuaR6Aufr7YyX+aGI0/LuwAN3o4Gt2WE4o9s9DTa2CPIPzhIfxYz9TAkQay/BlRKHUcEvmfT7
suWC3R7p2i1urYY06oXO9ev/C0D7TVDM6V/pCFsqEdjLbjjg/6se3w51zsccHM191LjEo9oCAghL
dGk8CcmnbNYPKhvuS02cam4W9HMYVcz6HQweQV0Cy5bQhAbT7d4ywg4iTMUu1K/tmTB9mfTWkw7e
aoDnGN73AmN1rq2908Ct1N45+dE32Es2Aowoo3496I7kGZbgDKDDVypLpU9qYLzhbMe1cbrrsHa+
nd0t5VuVydg6bQ4RnY2yd1zIg+6iOOfWc8diN4JzBHFLi31bSc98KD9oFYLpRD4EUUHTBLFf+mwO
hs/eRt4MZq5cdsPaqDenXurSs/sUHZUOmdL+zzsgDFJYQ+N9cvHPZW5RVmeGwFs/sepuM2+t082l
SwGZTkd/mJ/f5+fy+j11GgAikJ2Wa0sLZOk4R4ITu2Mv331wn9grNM9GmDauRkml/fdcXl/tfYdN
RqqQZ13/eJsDTQ6NgqWqCWsRrSuS3nTln/L0Nq7LQqbAu8uwZIbtLfO/DVVHChfDSJd8yrE23xPt
JMORm1MNWXZtTLIokqKcGqYuiL0CDgfMhYVll5we3naFgZk5bhPBYaPr14rEVYZjhO4MR70hhqqf
aSXpZmocveApZb62rB3DVDH+nqOW6v6hPVGhZhlByxuskXsExLz4ZoT3tAC0uJnNchZPY7nJJD8f
WVJ+jJwIlosc84p7d85d45c2Ii7cApeyjoiMpNh94bwWPNzF5MEikSLwQkHlH5d5jNk5iKx0mXUx
wZsN9jF8RTXgHGx06Yvw8ykn57mX
`protect end_protected
