`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kv0N+ODrJQAnD45jVEsSEPytnysm3pvAbJ05V2JaqTdEQNJrijqrY29nJXOyqQOIioMFCyAehxdh
SS8dEy2RvQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wl26nrMFXa6fm7UAkMFkRbwMiWczBO907OqYX8JeRapSfb54ShwQXeaNsbVvqp4GNYQWgD8fiWsc
Rg1ZH/ALNgmzzsXH1hqu9qf40O6LpbgjO9M5gvRZkEo/Tsa2oqZnRuXHxvGdfSUWwgm16QfnXWFD
HONMKYo+TnX1BbyoHuA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cF9G3LQheZJrMO7arGfYkxyoON6brspPywtxFKpTvNhoNGqsA1QaxZgfesvqKSR6jIrBuWrdpeSm
PoQl517JxEpEF310dys+9f254GuonHdyipWsWNgWjbTCuw6rYLvLG1y7lYwgHlSqKUNrBaGYERTL
bx0Arf8JZijWzxoSQ9FVJxjXj/PfvGzrh6e0n/oHLpafMxMPZcDI+yx5HuAhNXSr705mAXB8bgRf
GS+N50n6SUyWqcyUqw3kHjqQ2U4vJW+j5ZC3mQaQb3xJkZgzHfCaBKMstoXIjqY6XkB5Su6aeqKF
tsdYwq2h1uyBfljsOFo3IsRsUpNIiryBaM1j5w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fN4hvSzwAQXVTyvBcSPI9qSFGq1b0QWYvne9odu5QkpUwhn44DFKeJSRI90o/blLQLnT5fdJ1IVC
mwqzRlL7DmT25nQgDxB1mM1knf9aPQaDbovHFOWTzAPBPJqGcsU8B7iu5g++kkRlIJA/0D9NUZP/
zdeXDuR/f3RpGDQ9X3WIBcSwde7JdAaZPxu8gycDj+eAg//eJ+Ch+IApwl6KjZF7Lov59CHOoVNR
udrlY4+R4MFUEO48SwDCDlqVGTYZykUVxSqzXifsrNKc0qKvKF4GbqbVHDidoVCoh7f7Jnj0snvM
x3DFGPDnokqNpDBX7xF9L6+GYPELuxQwMV3Yog==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MECPOWJAU4w/UvBGQeSeElgdlWQuUK1on5QTAzUF7zMKC1Dzhpw/yWAmwgERdTOHF4jFwSXDGCYX
dcq7yoSgrYHNe1Z9FD7/4uOTgF7lUDYslV5k/HR/cVW9QWbwl5jLUaoa4U/BsWl+xPk3gCXBhT1o
1qrFxMGkr18FyvER+gYFNuGtJOdwhkp3EWSeT0uUZpww9gD8GQxRUyHQJxyLO7OrJ+p6c8iZL8us
t83ykRj64BZ4A7H8a4gi13wX2JOPHaLBMG6QaY9NxFK4P+cAlJ5tz1UR5CiOSua4Nbo8RZAnEv5U
qSe9Ctk2cb+fZHyT1Jbe89K38c/68dSDrW+q0Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JGQumRp5idVwKA3zzoqht/27epSOGyhvfg4tXP+tPHgo6OfP/FU3H6/X1Nd4Y66ilN9i+iugj0ng
ehLY04ISDe8fLdY/NaZ+qOkmAGDYirT/RxSo79rIeXhylLKnHv9FphaO49Z/wGAPNVJcMj7acDAt
BmSxt3Wb7gOV2zsovZM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FGXHNsFzSGXjbxp7bvoF47vhF8reHgBm6BrifhO2QcSTwMmIfvC72GA44UQ8v8jHIWHgPlay/nGH
qq6loQoHzagZ/voRdMzWla+HchA2la644cxBm8f8Fq9WGjAfrRKdp+ka7tSEmDbdQiKs1i43XT8z
Q9z55GPf5g5GdS4wXPj3ZM9TkEPcyM6MWas1txHsPj+r/l+N/OJNLRx9g9A23yQcrqoY/ibZoyFW
/7no0S9W9Nh+BPh8OXy4CwqtsvPd0/Zl0/JDLnm5d0hcEAn+3TkTvrZq0NgpjAEEOfrxtp+HqvpD
SE2gPjJVpUBZWou1zkZKYyakXZCQodq+NDtzNw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
/b+hsXv7QB5NXIuqN/9PIi9mnXtntkBUS9iBqRCDb9/noHCR5PxTmmQy6IsRYRIEQvPmiBmiKup9
7WDDxzxVYRuTIDXtOLptAWLHL+Fjr7p4iiUq3Q2fxru5nMBQnboWN/hFdi/446J6MQgnq3YQRBf/
e1fTJqDOxrT4l2FjEf+E0c4R5H3XYnjjoGIwVwJ+tYejDxewD+9eLjOgKNKboZ0GNp0DCcLMxE+A
1+OX9r+L21gOad76mSNJbWxzmlmv0maK4iaFHCmrKpno4i5wsiYIZKpsyeENJu1DvMH2WRIFXGEr
5y6E3ABQIBdJ0d5h7MinqpunikgwxDXUSOYiIBPmBDBrm7bLcsFgwPTwP8trsbOgkEXnEWn0EisR
zRRPMCCk1Zl9uv97Q1xWppSR9vndG8MP2Oc/H/00FtxYwZ2jHU+XErnkT8LlfkwbKp2/fWOo2gWr
eJClU4/NIiOdgMtteC3XkB6imu2pAtYtBiPG+/mG9ucMI7aZAp/cQ8az8JEOZBKbKjR00K9s9uge
O7LDv3gpDzNv2EyZckxJm345qCZwp4OcCT+ldqwWm01Y/v90s0K8MvD4UI+VVPtBxv1NdrwGdVLx
Lpzk2krrodEPeYdmjP6OwBTzyIc/uL2VFxxguu4CZ4suZnfX9+qKUWhwcdE2Aw6VQSlb2I6C2xdl
vmpP1Y9KgpjLCBoiMSvRKaYpsAHgX5ysVTVnXDejNs+C0hsUXfX3calcJbHrxKe5/iDVg016ost0
UhLiEzVw2RStx+uiQOuES5IUJ3U6dIAjW4YfS/dZZ9vlBdxULkmKc3FLbPJnCObIwz5SlUOF3+0f
PL15lwz7mp7oGVhufJ15P3ZhYdW9c7J9uvjfswiMjubf4JKbmaIxJ5ZDwgDQgzspJJhD19ryN1KF
r+kdZDaYXMz2TCNNQHXvn/Ru7Pi05CaFsCLezT3fjcHy62b5+ukJl6joTXcN4QHedUrZ9Fzbm3On
IFaomI0sNSbl+PLEpvQO8/7mtVgOsgf3AeONxmRtaTCwK+RBdOX9G49LkURs8AuX92BgaLokG8oU
tjgoDYAyHTnnJv1RWh2+BSDCMjRAbl5eTQU/0I1KovzJKLY/KOu9H/kpVxlythmLHYRQLgo9pycr
ijACazQD13I1haOZ9s4T0ZwzN8rTa1biH3JDyZxNwLoeq39GkwtLY1fUSLRIPdaUh3MA9X1wO2jr
ybNAwDhc6vtSoC61+ue8NsRD8WurbSUVuZnEG2pIqE9qm/tmvY6AB62Se3bWV+q2KqT2w8/2qBho
3nnB4ACG1vedW1l3hTSWhuNWkmzGDNOoqiymPwsKLcPTamLHd3gFyaC0lNYMdkBLjYuzmnWWO7Ic
KjrXYZ/8BkgGqsGy5OFNLFkezvgwme1pKkjKvBZkcfZ6p1gpplVGC4AXq5665bVtK0zP5JxJvKZx
lBZRrC88kZkDNftZHdDDqTnwRud+SZ5GMWI5HROvkPoH7beE/r6a7YMeoGJRxh4EggmlqALvEatn
o2xNB59e+izmYXAlAPXH4MaWiajtO3kCDJewz5mAwBVNn+Qvf9IR5oMuIM2k7vtiqqQAVTd4Ii0q
zYp1xdgO+1BPN2b0sNeGGA0mjeyfFriQxTVKaV9Kk+N3rQ/xqN2qevIDylBcBK8+y/iJnMcpdG+6
jhKWmOISyV+eRRMeOL0oDTT/pLV9fOszuhb2E8adX41DWmv7rPF0A3N177S+J1vjbXShvTI7fZk3
6hf6Jy6SxQ4acSLBGzcx0qd4+D0of3PRaVr4BS4ftGNVK6Q4xb9X+u6hzd33KaN7XAlpsyzH8mU3
a0x8L5HSSReHIlC3BCZcBCo0/6V1ZeT31nKIG89Ypsd6P1pqq7AecwvE2AeqM5WLswm0LJ9b8yOV
rFEQRom11ORTNIyfO3rg0ttBnyRzPS2O0bgy+blyZ/4X3O4SU66fHdRRtW99Wmz7LSkDv9YLcj/9
t/W3bpG+o/FmR+PTpmKQUovyZigDDSc09OX4n9SD26ZB1gspdhkEwIU2N0xWb+J8+Z3z+fG1Ih2f
K9LuJn9MbBWzzShXkhfFg/mKoq+jUcU92NxdZ885b1zptaaEjARVsvKCRI84tAOsUVzfqFrcgfDc
97C4UGG6MNuwQucV3VdpU/QXdezB7Vu3AViIMgGePs2AUr9Bze+vnTL/+eHn1Q1v2x2bd5unw+WI
/GuRrUfdyQOe3duBaQO/0wXd/Wvp2NUAcoNZB1Kd0ePhUM6Hpe3Ilt2doK+OvKMqk1s+A2+HY1st
e/wvHxXVrb6AqBc3Yn74PPR2FnsSByJN3G0dXqAPMRX2Z3bOAvzw1Ig5zJLOwDxBfk0WfjgWeTq2
bGflZEALrk1Flal0F5u0yPx57egvb5xYwzJlvy+IzICGDHTr7LSR2hSqr6tUAB7rlDK1RC5sFqiB
90z+jmWpdccbNiFiIAnj4+HC2hUOqmy1A+9hTJOgaCrRSkCzb3nG0r16p5DobG7Pp/LoPraDRgcT
n8mfIBTDexTR8gQxw18mrvaX9L79pVykIhIjmaGGvv9EmHP5Q8Z5q23zKPRiI0G7wY1YtdeQEFks
i0H4IEsJoymxR1iimr1DGJoPjs9CdZdG+qDdIA99UGgpJ1I9WR6eXHFLZSSLDGYA4Xx16RHzt2mE
7Rjvxxkt4iDx6Eb293FCBpT1jn9eWQityUz/y73h00jjNJWT4//pp5DydpPy1MnJiFsrAAuRSsYA
HEzndjJKjZSnRr91/PtnUy1hjIi34i9a9NMR+fqtFpozcaMyLHqYZC7cgLIuheJEFpARChLfYyoQ
Jw8u7dt9LneNSIf6hTPyb4JAkGaqNxzSrCa9G3/UPkgMdwfwVvPpEw+YtVseV6saoTKeRU3WthKc
V6NEmK2W5xdXCJplhHztuPi56M2rHN6vJPUxUtEW3MnLVggnC/2GinA0CJHRPIppCJ083l8aRQG0
HOMuzuuh5WAVLioMzi8LZ3SASKunqcAA7irHH13zC569xbJovIq95+wcTfp4WpAGcRRbcm+gWwXv
waKKUc8hJGSCsEaz/xOxUhVnLKDpvspbTAYtwllLEs5xFZ7cLz7wO+vpnsC5oYnTJ7gB+Ev+5k1+
9R+fAlqgN1AuKJmBjN15TPE08O2ALbeMT1pQ48V2fuhGHwzSAH3CZBDPqIoF8oSHpLF4lJEpx+tN
CKQRl9ZXRDeMyecbgB9Bct05gXB/HcGXVwV+dOOSC3YXmNjk8a1W/Ttv+fb4Zs+rxbHMEqS24qwi
CBOUq2mx32Gt1CcK+92tmB1T/KKhs/d5s9NZagerZmROdQcQFGPqnAZg6Le3koZ8qxib/aBC6p0M
A/UselyQwQHe/Zqo7NzNHxi3husTGS5U1pHKmst4oS9ZF8a7OKOV5lDpwnBPAe19rg+vbRaSk1WR
b5nzhstR8zPyDUVYssIFXBrNrU2Zv4yZygOfr5NEp1jv/e7HpbGvZS3D/4ZLoraufBuPSyv3vpa9
wA6cqOYxWGqqYU/DBpNj2xSJpUdm2hPNxiPtBkFCxzBR4QQ0nkc9i0V0cETon0Vq/Wtj3HCGrIwW
mdq14rCAZSCg/neQOrd8fdNZ1uFkdBQm2WJiMkiVwbVN/X+uEjp1NebRWZVNV0yAi86BEE/CmS/u
Inm3pvnlb6ttLZqCSLD68QcQSUxc+ty0o58hnh9WEvxTfbn+ngLZWIBRUJT/oB7oFx8RKTyhc7UZ
6yxEqf3xek0GE+Hde75VoaigCT0sRTzKuG46z+Cx/DRhJnvKF3ZehUPJo7JovpIqOzQqnmpQVcfH
PwK+lWAT9ExfBjTKSu/U8TQw89bQkuANk7jsfMEEEJfuPObS71ooCe5yvF5ynhpbSM9iT1V19C/U
VQvR5wesmUweM7AlPKf/zQuJy6UiXG+thXo8M7iSTGdRn7dBumwMTw5g1mcnMXFaXNEga0kpg7cD
5cXk4HD7u5cV5dehJHgAZkmHUSWE8Z2ENFPYkWMoLgnLEYOuFz4r6LsTy5CTiKVZOoYcDqoPOkrW
MJHfZ2VKo9xVOaSo3lCwh5FeNuunZQyAdysYVvf5bMaEpgqiCYboooOifS9P328Kq2HjE5X1c0SJ
6SpUPtZB+mB1M0aLcnrE1fxDH7y868LH0MQ5a6i09jAVUMTGAehRv5jEv18spm8sxJxzzt+UkTdZ
OatTk2wUVwozWuJraJW28teBwuR0c/c5nLA5tInAK2Qv+L4Rw5mU9tBgtakeHf2Pp0Y41rdkHdol
eXbu7q0hpp4enW6FuQXXbsIDWDGWLsTcGJ+SA4vCk6y3CxaGDRqvW1Zl2WnY7EbH3GbBbnGhG+zd
M3oXb89Tl5dU/vaFdLqlSAoBsiH4qI+AuH4nqCg9fpZzgz/jQa7Bd3j/UqCtEKJFXIMFQq4kgHLF
6qDZHnB6VdOOJTSXluaLPTvL490qoPr2THoQrjIsm69liDOPg/r8cnMPodOFLEtBZ3Du9ZjUwYMd
G6XZUykZG3Ej0xfMlNOX+nbZO/tAz0v5v4ljF2ur9p5na88hmZKstRwGBc4gJmYTYCac10Aae9+r
8z4XneSZ22IbG0YXy8mwJ5SqpgJRwNtcc/ihxOfWVNcpqFctruArF3mOEqbDeOqnUwrgkX1Fd01A
Ds7qISWgO/iiVF4WYb9ay9Lzry/XyMbeoeQpDs8qxiwky3bhzTBoDrHvchaGSB5k7fjA/2Zsn6zu
DheXJM1f7g3u/VfJEIEZ9fBC6TBD6GfAkSxCQMJbcTTySvbKl7NrenjvxEw3YxhZrMmP6XY6NY8D
Gwj4JMMjLYpT8n/E/tuH1a65LN/CeZKIXKLi1GgvaQo7LbpWmR6O8YgSWfX4JT48XtsPlKEoFpkd
v/YABd9Vj7HdBHFbt5WvgkgZaP1W7AFnC1P2lhjvqGF0AKYTQifgVpY58Y9up6tmZum3tG8eK/N9
fiSizk9iEEGtCnAcUGpjqh2pylIrs/GJ6B5hfMspTjLR3Tut6jp7QiAlphDAAMQslsP3umPBCuLW
rEKcMZNvXrw0c+Zxv3FgeD9pth0lNf60W/Lz80TDDUSTD5eEhZgAKVP7ihGiDqmy4w3D92VdINfP
NUWIsO/oA/ApaXpEFo1m+iBgzd5iI2Vyx8O3ScnNm74MIlhav8TDRxujn3gtV+YkMkJdWvC9P2g7
pixQNm2DS1wxrVMNGyG0bENzReitCLB+hLJK6xdm7PqhidXoKn47nlVhgSydle9zjeHZC4wjIeEs
CQuj+Y63xV6eCS7AtDdHt29MOmx8FEChodxtOT8m6ooyNrfn1OwFHij/1m+6t7kWdWfkeRnLgCaZ
0vp+OB5xQpAqoRxamouDZMv0D1MZtHYe5yiNAKe5Lc+TXuO1K960utVe3XHp0k4AWh4rJCL9ryRq
lbgnappEaLqkhlJX1HAXH/rFLm38i7enawYnTYg+Z7MDdEowvMnfpBOkM20NY12Zcqp2vin8l32M
uldrr8ShdE/KXKCjvDMmaZ93PN+MBM4t35csn2YH7IwLNXXxXl0SzFu/XjH2yPBH64cMDa3/Z4yg
sJ8uMw6H7VpDRwR0U1r/2h2PWQNopTSPFsUn7hzNsIbEG/KgEAgTZeQhmdYLF2XBZ9lk0Dk5SpK1
1A1uSBC/8L308/lajaJ26Xk52IAC48pRpI0KitdHIYExSHd/Ww8b0Rv/byVRKNSio4WdrCbqbijk
UhE4OL1J9AopVldcBLVp51r2W/6svIEFxCc3CLgLiE2UJSPOsZFLb5Emmt7v25LFbgD98Tv/BRoF
ELw+N4jL6ykUDknl9kclmzh55aeY7R0eYr96YBSXDkIFfOvzYBZVC3V3NyTVvCuXF5lEzzkevnJn
ZibexO0HEVEmFjoxYaUO2++XeL/qeifOwvfGG2mXJHAI0BNm5RmVSwfRHqsBF91eaW9bFeYAIR9W
KfCrfV+lKj41W5bBnB7+Q+vQMlukOoj2IjTldZVOCm/7JUvw14Q3i8Qpgd0a3n72y7z6UwBgofGT
WmldIllicc54CQtG6Q6Ss8xRb4SuzBDBe2Ozj4okiLzKqzYK6KtooNBEHSj4SZtkwwFr6IUOC58I
f07AsIaz4Qyx1TjQblZ0p8db6geaGAcGD68st7fTiacz7NxUbJSSqsRCsaJZz4JKDv+qiTx5tTlP
aowyrNVL1xC1hFXw4OtVfZGG12/O9TGjf6Zf+Hj6uwQCUcZVv+dWeR2VK7ZmhDA3KwofOlBXvnN2
lJUQVPFA5aVQ2xS0HFL8dG8mwzy/M9ildTyQY7NkrvlbgAugzMaB/hQCoBN9I9NKswWMixJSKbBX
B6qYmbVM66ciOhBuuY7fRDCiLoxdAc2l6BQKHZyI/u9s4ClG+kP9KG5TdHA6Y/1+bhLnhkxtC0k9
QAkh078UQ5kEFjus+hRRQaVDcqcCC+/fa8ZKRnbSU6ztBk/T8p4wh6Dpak0EXlZEEYbjPupzkFTc
5R2CqFmPE5vBezIB48mtGGqRz24wAzIn3faMP/bReKONtGYznklF8n1TRrh7woAagNNapjHVZ3Qf
fz8CXdbaf2nA/fxofSvbpHKUiYFO0QozaYt6Hny0g3GidPatbYVTfYuiJzqpiIcSCQN7EILhIJg5
oNv4isxjLtuDinNehI66BjyuM9ea7ghSZac9q+HtNdkMJy33J8bZoZRAY0ZeNIcb6jCIiuoOndN3
NzrK4EBnt9WKZP7OPugT9oqAvwCKaKaKoirEPY5Umu6Z39xnERRF3b6B2377TVoGqaou5ncTwK7V
lYghYPTb4kGQEY67mVCz5IbPKFp8Gtim+5YFkBih0ilBN+e2kDuMqoylZsDsbRA+zE00tX5RPUuL
PII7oS9VZ8bpnE5hHoFXN3rMHYd7AN1wetE/6vtIGO4atyA7AMD4YEu2OfvnmKpswtVg5bC4BSSW
H2TpzKBpeKs72bG7ppx2vvyZLhx1PTiEE1nipUL5P4s/KBlV9/HamxNMJYl6oTEM7YwuBhkTXIyg
sRTVavpLOelMG5grAqbTybK67AEqykRq5bQQVqpAM4csvlcIxU7Ytp9kxDk2foEZLd4F09Xw7a3j
sQXHcSLhJxE+AdjfbZxO+eQ+EQ93IaVvr2YDj0cDXjFHCACmO+SMyaXB429IRJKFEz0p7syIO8Y1
lcP0ODV6NBXnudopwDoTV+LRoAYKr8UN0YYNCeHzhC+IU5lITcVtLFnwOwftR56Sd9QSPwnF5H+l
BKrekombol1o7iDvw/uiDaYvE+uYcErtFvE5p0dDtJQg7KralHtj8lxM3qFzXMzY/Rfu5yZhjzrx
Si6GI5W8ZbGNB8YvWi/zNgaDkhf3DoNJyljyGJirxezarBN2XkMJNNmHq4ft2PNOwktAN3TFtS8F
Kw3JG7JC2jWAz297lOsM6zrrcflMtZHph4LqQ6EcrEYBw3c9w08MrDKW+VRQ97eqT4VmAX7TtKJy
JodBRF7ti2Nad5yiRAu1HPjtg5ynuIH2okliCLmjho+C70FdvCNbfWP5gbfPWDjBKft0/2Eqil3K
w+ZOQ2vfvOrI7vPN9cr/iyaWL44WrlAoLDnSos8gFraanmcmDyPIGBk6NEJCl6PaZPFVm+S1/LS7
U9mwhLpx2cfNf2nV2pBwkBfgSmI1DAki4OGRe1lTk6kqAACq/Moet4fsz9mGgJenayyIRKHhHk7r
O12bzHpdMtyiC1ZwF+HmWKqNpHNl8W88zGGfjLUjc5tF6fdv7eMkIrbHR+MCnkRERE9vxbIY2bEY
6kodxyzR7j2BUQFhmH923Qz28GS7kpQczvoo2uqPx7jGE4511sysqROHPi2/Mk2bhI+jGA32z9jb
iBgV3qPqj32wTmRC+KaT588Lu8gBFHStNvzN3eGD6wePEzmTLWXjNfVg5CfZ1ZH7P4lYAc1AJXcX
O28c7uSJi+4iNLoSXLqOodTcwTjCqPCTs3RE+etv7JCnTN81VtrUPOyJE3JHyg/8UyLAsG1C24Es
e9aAD4CO/olWjjjqmwqb5vf1udfuIWKKJ7ooClIQL9ISVhkOhxBi+xG3tlk/KA3MIIm7/qRtZrBB
aM4OCPOtgpmKsvz8gs1RPUII/1dcxiHuucAmDsE5eG+i89cDUzAjXWNhLAmtsiE10bv3zrKg+N74
C/M+FSY3KfQjp8joijAwXlC9hSlsNB0szQd+4kHU4XAmz0FU8t0TIuUB1aQkRSBsE5UclQJwv4Ma
MPhjHFds+Cmp7IHPdKwFavhNkod/2bXaKZRtaPM2Q81k+LJKnQAsL1QGZRFpeoZwkTaC97P2Kkmm
BOVHBclyoUxvR6/mqGBDg48zl5F2giiN2fhbDvftZf4CwibpTt0j9rniDUoDvdoeX9ma59CkhNu5
1hi4YI8Bvg3rfgAjIuMVSkfG06DJOFBc3oxd6bfx2q2cfHKYi9D3fOpZYiEZM2EVM+nFg7jPOZcn
6Pts7JMgB1vlS0SaHOOoywr884gYXFBUBmzjjwLA7kexFBJppI3DxhTLK3NPYrmwv7PnCm2KrPb+
4F+dY/NRgzLu7pWZyo853HWo6ZfSV9nEmaBR08SUOzGlcD6G+g54On348ssYWoUBQFOJ33qCrqD4
37axpREyd3kKE14ItiGfczK1+9Xt7s15ulldLn45jazY93ayl1RBgrorlFUD+qm79378cXooUKpM
GImUmehZloZwYtbXjj2reefwAWgipUbqOKOMFN7ZgDn6eBpH71JpQcU4J59zf/61pfB6wo4CVk8s
Absz+pek+EaB64g7AHEgXvYiTvXgorUY9A6FWGCobkg2OKs330RlklGDH+b8kq8FLbH+jFO52tnk
St4YwCx+nZlp5nPdUs72k1Ort42ieanZhR3NNYyQ4EUuCF37RC8priFjP1pgpwqkBjuakg2W86hN
bRhgeyv7qyVhp6zA377AoyqzbnOQSiRRgBTDJlMbEz9jYPWB5dU+m4vD6SFmUFeemoLBoFn+j6dh
JnVRWuphs81O68VhAbTa80YNxO3LWrGIHS9SxMGS4HRKiROm0bIAEbLAMAHzPm/aQ/w0fmdAXUlK
WBq1GvnJbZsYP+AsO95E9TxzOhgW49Fr29YNfPi3bT8+6ut6VRE2nIHaUhY1JfPO5dEn6R55ibXV
ozKvSdlfAbdCV7zc3eUX0/mz7MDG4xNbwHbaEHW+YlUj1azCPn1UAovwOXgZElXmoVur4WhdGw6u
X8qlLgy8rdnLqx67gMgqLlZTrUjQh6V5QljKKbMhdM0ro0NYOxGbHc9V6VCQ3fVHs2Kl5U6S/8XS
CbTdf87HRI4HNKj4+NX2lZLfWUoFMxfS5Ee/K44nZJbNEo/GX2mt/h/bBxQCQp9/xSpkqR67pzuY
z2P3vdBx3GBIYLo0XoV/+RjEqVMDb6eThW0GJdhVRqM99EhKhWMF9/jQE6iopuAfLpy+jkahYqk+
fvgEE3QDEJgqsaq4SMux0ZF+0ipXcrus68iYl7Ajn4VDtL4hFaAhuUJK4+jVjkdsIDG4/vlqZDFP
xAXhVNTUrfG1XWyf75i7hUpZkpRwumlWzg75mWWgdzg+n+vz2bmojaNru9uddh+BoG9nMjEp+iON
bMar2LPTy7wP5YwYMtnbaVq4KyYUHMF/qWrozaKP1SaIHIK/qnJLCcHmdWUiWlrKEiSpx/8CGQXh
cO+au2Wbzs3Y8f/G0MhiKrm5hZbBCq83Uul9yyShVg0+f6CbHe4KIC82ZM5rcI8eI4H9QpcPTLHk
CaOqysYRaTj/AeRaZAlHCG2maYOvEG53t1YnD22uT4SHJJHEqaJ+6r7fS8hQX2+uD+ffIcfdPTD5
Y8LkwolBYQz1YIitDFAB83ZJRmKzXN5yaQIcisAmkYpZId37DmNR+14DYTyP4exa7nN64HXDJycn
iSWB5QxYns1QtvBfSUwgRD3R38l1QMCzPmFDTc2xF0wv8F4hzsXcSZx3BhybK6fu4OCaD/yufs+a
kmNNsdtHWdUZd0djVPJsiUlpEmzNKI70dnyA5WkvhmaDbtVPx41znPMQb62rDVs6qaDpaAA8j6NG
P0tnPStuwDEiTPgcbSRTBEF2XMnLlWouOYuxmBffjx5HLLy+c5nUwuQ7zLu+1rbbqELm9DE4cdbf
v8tjkI8yBz+qM4uzfeHZ1aWNHzwoUNGmoR8USYF1s0B/ADWQ8h85hSKuyp+ZVi8r4JS4SbvmJr52
BxCVP9jhaZA6VfJRQJtKIGuEvz/A6uV1RZGdKSdZjj67LEmzN9rsSsHJ890Rp5Sz19PfYI/dlLfg
g+AWk4VXblRLqEhSDVyCpvlNw+r7hW+F0aItLT9hEVXPA4IEa9DGSGG1wVRXcVZjcLVOOW5963ie
6t37ziUlZGrw1EjyjgscUNEJoFo/rHj20rlhzQi6IwUzXp1iFOCqV0b3MkQWmus1iCkVr+AivTIC
Kvo1tA6buqQHFyYBVnZvrAc5UToh/S0olzlWhuu4SuoEWh1/9udQXCrdfKHh86VPOUiJUG0CjiKO
1EGcm/7mPXXEFukaxLTC4FCJvbihHSXU4Knx7HJCbtg2zouksWjZ0lpZbyQlPI0cuiOVO4zNE4sY
raLYjfpvPUafB5it4njZipp5THIEBGP3NolrEDnirPv6uYTPTaLWccw/wEOcZ1OB9uwxU0A+H4uP
PBf/iqnMyY5lb5u1IQmxOzMmfB/DG6sC9bwalyuH7HkHQoP+LGLc2u9XBxvQwroqsVSG+U/GWOLt
lAo0dnM4+hD765z1R9NJTq0/B9G6JWu+mmJgKEg0+amMn/WE5G6FlZ9HQdoInKBUhlmn1G1d3fOj
pZdjNTfC7YXzs884TsdT7zss84kR1qN936FPYtIo28L52xTuKftUIYn/LBxuyyPFzyYYIGkVEkwg
b/bQlOJ7wmyniinmNds8xxJREYA8X+fEhIFlfPwPGG5iAc6TfKKCp1aqdO+s24KYlPK3LJcBbHCH
GIGuZgCx493dP8vP896SlKbfX7PKcnylfM4kusmW/R5a/eM45LYO7tHqM4rshiAo1i+wWNqOjqAN
5gOKN7p0rlbI/sqBnF9lVh+oHqSxeIege1/r/usfRED5GlbYpwCgdVQhM4wAMdXcn+L4mIF8XmB3
gnOPUblKxK7vLbuEFAZaH0OAP0VYV5+rpn3Kb937jRMyFJ6f4BzJocvZEZVCNShwvN6KAP2ZZTpF
O0zKQMgYcEML2NxtCaWmkRW6P7RS1S54O7jdcQhJlHneXiLyCXenXmJLAecxB67MR60r6tb7hDCu
mj3ZS6gZVzLG5EceRIFED1qBLS8vsVsG2Lj5O8wStjqY8s3HXPrVd0RNtbcuFXvCCl68HEmSZzAE
F3rN98QV2gDKWPFVs5riL44HFExpDpYzE/m2USRkQKbzv55+HuN4yZrhou7Wl/wUKEaLpYm5zX/r
EHSgg7oBmGBpSEMgBkMzdY9hkOmoJwahKkrS4PljM6w4JZU0Z8mE0aKDb97NlrppK6Dl0GnSFuIc
pka4/UgxjzTfFgfbGJN7x7ubj9vnPFTiuk//kcmnW6+tQ1ZrJP/ZfF6jI8qMAAYI/xa+FW2Zxijq
JauzluMnaSBM+H5voINmp4TiEMlAPpXqrQCVc5qqU8QQFxUxTK/Eo0dHpv5bzA5j7G13WF7PQT7b
AvREYS9AKwK7WZICnq8auTTBKI9/Qx+06aRTCUn+t4MSDlMtv/h5eeA+VN7XROCXqhaYmDvQFVsu
Wja1i/xpCYXfWFUSZCbkJnqfBJ7dX3B7hLTd4mVe7EGSstDFLCsdhZd0fHMa6EpvLrA2tpkQNFvA
LKceWPYd1wtZpTLTvCUDgPjISeFctoaY+nvpgd1LHBbypS9kQKl3NfGnEM4Ao3QTFXd3ev7qaA+I
0h0qav0rPuli1RpC9CNuMKl+MG5e9sa5WQRqdHArq8/Bp9EQj6atLwOFEek2VJGLtN9j/fcYFCWH
scbcEluN8TtHjdroKPkdYruDjrM9ulBJRYukHvlFnyexEFtAEUeWbvsGB5ew26NLsc1Hrea7UDCB
0DpkCSj2Eqt+TwrlS+0lRQwHvZLApLRVWoTX2sPsYTyxgz057mSYuRQXqel6evSmND0rY4+/895j
fHv3Nts9nd8mZ8weC/sMOAdvePjxQMlZLwuARt8Ai9Idll5LYj2rJ6+z6HcQKJMoqkT8JC/1HEgH
q70HfnB2QM5mPXiwmNBwSUeSoRXvT1xHnoUt6gLNrKmYk43sYj9wRKUft1lbSsv7t+w9iQFYT1ZI
mBaN2KFOCh4KfmC+TzOLIJGV+Y0iVvzYQmTzT/mWASrj7ppPtjObNkaIkLEhmFWc5rwuDRk4BjyT
AMy+0T2OxsiS5XRsO27QhcE20qF6+lT0TeLz9FOCVuvfXD2DAXJEQolmUuAqwhqxz9v0r3i8ICrv
w3cUKy2K/WpjMFPxJMfqE64P4/ajYf64CsdiPnrvWNvbEFg+vI6G1K5H+Av87vkHHB3VBSZTZqjU
ZGqW7hbnsUPYwtgRe7UFLh6kMdbuqSG9w35FZctCcX7pMvMO+4H1gezcy99YQ+IYvdbn5e57Jo96
t1DyguN8mUdri/9LQ63v3PqRXMHMLrzdaSg1b1O8TtVd48JVpmPNWoqILv/BZSGgNm6T16MVPtPe
7sQyj12HwHSIwKOj0htRX818dxhb8OG3Dw75gdQJ4YSHCY+3JSwd36+baWUK2NbO+oLeT6FkMl16
6WMpPD+NOD0e/JDgaDePHVZoEwnynzNDi+QBGZX6+E9btzTGibvcV/h1hagQtblgVXgLNzGVkAg+
WoD4JsicPGRNzlxHZPDghRAHqLx9uDbxDwpIK2yqEsR0aiIKnfqojAOjji4tK+j1a3XzSVkHSvTG
JVyYKdoRSPGoxSsLUWPypnifCR4NnC014xjBqSfSlVZ1NX9xjNYcAfyUokp+SYLsirOXAFrrZSDT
kdgWhGH/SDOlRcwRjKNQ33IxAaBVuE0rWSmTcgBe+zDWy7rYpnBCSw1G53rWOoubfNfHdgr9HPbn
ovXSHMApbioxKHxW3BAZ5De7dHtf4ty10Vo2DBsFD6kwsWlVuNJ+g0R0arqlFGMKjQFeVwn864um
VmeGKYnmzEwcAPKXZO8NXwOHiwAofk+bnDu0hkXKjg/L35m4o1Kp43zjBM8B+iLXswwFfNK7zJT6
iRDvm0P8wGihSfiP32tnErSldiVJYYnr5xMOaqq11xDLDMxShCO++TQV1eMZXsgJTfhjiGvz8aja
U/TPUtv49rlZYcMCuBRptsLUGchJqEAtUEJR7VnBy8X6MZL3VfTDyn9ztSXbaIs1XB2MTlsHzf+z
edPXDBD1p3kJtZfnDD1h8Aq5iai4zIpSLIBrd5suIFf6iIHRU731LN7txRqy9BAACXdrACuQMDk/
dffNOrrLNf7YpkDfm47n21IQbKFZQJNkbU+GJBGw1qS/cnTmcL1NadwgqDclbagU6Oqe06/AJoxB
pIEPulqgHB7S3x9YMgbYtf9lupuwyub6YASp2Dcb2mWYLXvAHzdoxWADEOV7lQtv/9rU10+Wt1VP
dbKbsblaAudZ6onpULBJSWq7feApd1X95IObAbZA7/ndIy/Y0E6AW7GyvBwHEwt6YnGsigD14kl5
oyuRvDyfW84EvCywCfb5PjhRp4nCqA1VWUTH2P7mKSzEK//OwGEDiLPvpFRoBcjkMuGPuKXV0rSo
2mB8HP3ugP1kgZatEc543huijYOcnldcApKw6YWUeqlYco7BBBB5EcATNYCeKroIsFEq6FJHvUmP
cgonvqlWduF6WRr/xLyTjlp0IQ1+DI3E8D0u0/fwQ3Q4Q90wRcLeg+VxxNwZUEep/LjBqZ3FtVDy
bTsasdyltzIjeIh1hN0DdFrYITFgFxn9IvrBwNgwNZIx+3RuvjqsQkqlPPREIBhSEqNyUHxTbh9k
j+iLkSGyp69Fg0qF3H16PDQ2gKb9uDj/YcKGrYGWopnl3LgCglN8Ocrtj6mSmRV/W3Cnpb9uVCx7
RNe0d0/0kfUWS/WFoHesS+8hnx0b/znyjczOPBX4YFSUL+BqZaI1SXdG0/EKLH6Qye0Aa/YYsVlO
m7hMCJqtNkP15dohYyc13KlyttvCyI+fqnKTU7G+PqbRKglXJveBnnfgjD+sLx6Duz4Fx4nx6Lrd
ghUTJmRKk5R75+deVka0Vqt009AbiUFKaJuMUXeDufiMbgTx3TzU7ANsE6MudqzTFL9BkBpIvPiW
02mFDO+3AdOpD/1BKa99uH9rqyTvTuAPslFrho7VSJph4eCR7MsIcwhqovj9E6BQmY3WiUbb3VKH
RgvgLn7H+hQsR1ZlyDeYraUTlv/3jNG8/57DgoaSXnRskBObc098Xl5RCWkuUGSt19xw0ekLT6wO
DGyTMJfsRS/DJOTItqb4hAkJfGDDamJUScKZ563K02BuIDGQGWYnTQi+uQUiDIEkHYqrrZwhkZWC
JzIQP3JGy6EkSLoYP0ArhceYbqduK0fYT4KYhslmxdW++NE112Ul7+966h0FzXyhfwDInXdtQC9m
84sF2Op8Ly5FnhwNHXjNz9vJg5e0WHcbstvh90bz4YjAXztW2hFPNO84WXXyTdGRSQW4+COTLvv9
RTq0+2vgd5wm34KjnEKb9z1aaVZTgzW4imBBGH1Je/uwCPVHtCd4vF2/fqxvtjikH94x/wpJ0fca
s4Cx+y5jNYR2Lx9UuLbSl80fRsrZje2OzjT/IJO0jt2mk9I7FPpjYOO8wS6aD3WhTrAyHx6uTii0
tNP/k49vODy1p0u3w9T5kwwME2ysmOVvSlU8cfsjlXPEt00CcaAYDqWTmhH7wsREqAI0XOZGSU2h
j7gdwAuX2ZnjfCu1BFclBYollzdylAn4P8u9/0NQLoavsKRgwRJdUkONvTKotHPD6FlT8XWP+xOW
LgEqObBAmw1LRZQyxu1g8zzyxZ48ZsrWOkZYylSS+2hITU+nJkLk1JroR83JwLJ/C98n1Ia5QVRr
m8W1MRpANceak+o4WbbNzhsef7/iPzNkJYmIWjzKyoSDKepnDZ00M6lwaGv70BxC3AGJj9+agVe1
ul4hGGGom8pyMs93ZeK0ebW1lJKAKMUfSPaVq30qBXQOQLoqeGT5H3AcD3MGuDAW7S9cXHZjIPZL
CEHcjZI0N59tjtGK/eJbXEKHZDtdH6Iu93f2qulDWclPDpZC0tbRfBexbmC7gdRR2pAuPMwGjiyh
sugQbm255J79jbgVL3ZQaZTUI24OYeTjlxgk1Wudx3YJEPN7x5L8dAxD+HQiqq6A3iJTELzOSRAC
P8YTyqO0bRVSN//jUVJIKNTzDSNic90SjPmyK1mQeWF0fYI6ODDAU2/kn/mrtes3WwguRGhbh2AN
FC6uHqC+W9lu+XBHH0RXrgL1Kcl2YyIH5UcgfTo+T114Fh+TFJGiGRsRIaGrhJFScYtFSmt8hwIM
ht5ba6nRkwHvWb+vtkUraVgDD0sXNkjhGCgz9Hp2pcnuUnfFsp7ghQbRrumW1Jot7XkptdyzXZ3Z
gm5IZ5fdduXmo0sZrQ9zMSGJs5YhyEAkwKsQbZDVXgd441QJ5gGhUR6tzk3Fs+kSWE/4HnwAOzEW
p8JicrzAYD7kIo9xgJf/DMD2NQBaitEnvxtpWR2y1SZdS34f8lL7EEY+g2RRucvnmy9/wnUku/i0
bz4qdlBB/HK/8Vrqy4eQDTZoosPjIAQBMw0+OtLuzGETOeiLPA7hl7ckviQraL5dXwGEVWdOyUZf
tvaZ7B6uoCNFPPbNenAHMbdn+d7OSvx/J/JTpPcfCO9JDpFca0bWXkSNrlHSx5zg1UOh4az1uPa2
zxrMUqSRfCwl4HPvdmKpNb+z92QTRwtQ5iVakUiH01NQQL5PjVe1RUQNKhr4awVyz6DuC7CetfLd
pIfwEcx2X/EwyLGcOn2qEc6vUexgdBzaGqXE6hB/7vDK1ObZNn5CouWIcBY4wF31fSqyTERJE1i9
+3OrM52dQ831eU5lHro/g/X0lBf9KtjuYqFqOUbIQZwXHEaUegv1WTVqXdsUAq5Jofb9mNtZQB7i
GbSkYyLAhbxcV/vZL6RoUnHfayGxMYQEeLZbpf3aScufW38VCfYZLusEfFC27mAODi6EibEgbvfQ
iGM8dxQ/B7eY6Qzc1vXa08cBsQOEVTqJP0cQ9448Ti0JvcU0/nEHzmcxsWxUwPQA90Oux1WlOrbA
lZh2opL3CWgLjTz5QUfWy0vv/gHEMU9Jv03HjsvYos+YxTeIL5r3cttBTL7tvjlrT3RA8fY3JXja
dpPIJas0UiiNwk6Ssp5qYGPwICWDnMcaWjn8NTxy4Wf8fDEiqoOXkM/BxaBaTIJalMfRHr60hjJ3
7cX3NNKNHoOS5RDDmx84RLzX+DHuWKiuhQMXm7eRnQAMeAPUHrCMlFYCDoJc4RVHm5XL9dS07mya
s5ClCW/PZsBjUrHHAgOi8AFWdsGKRwaDOU+Db2bWP1gwnFW4wvPlkzsCCdhidUHlMtbB2FIgB9vB
Ht3Xp/0h7BGGyP1YaB2rRUL57Ktf2bCS+YRQ21FBNM3FE0UKDCljpcUcEkB62OEzeeCrbtH9frct
HO5627YWvuj6BRurmklvaGqsM2YBRdeW14pKEKR2ZPnKx7qYTZXeQyj0A33yWaXhcbT/wkU2KAHo
hUb/7MOok/q/H6vhkRlxaKYrUqOOanR85gCRadFtJrdiwwSnWdTvZWsnzZoxwKbDTdXRNdNe4uu2
BRSLTulVhA5nEuOwkng5hUk6kFuvQ+Edv4YKZG8QRQc5BYr9xGJ3GjRcyJMq5M14xXURNAXyBJFz
FHeAIMZC/Ku/6jmyfiklOGCQ9WCKF2I2W6XjveBLujUueZYkubPDSB5gtiIwBr6TQDP9nHb23VDd
kZv/urwOQZAuWmE9sG6Am/2ObmB6WuWDFPtIdsyS34m/iRNx80e3/k1jjyrri+WKzs+M7LPsHGOi
fN0i9C5PHH32ysVQG8pXncKSoZ0hu6DO54/W+jl7QgxdVISeS9JWVpVzOdFvKWCxDFExIBFyhPSF
Df7wd7IU+wPgumaDtI0v9WC7agvFyCv7xJ/WfPPxDohKRJuy94QixHWVTrrn4wgqsoUPhRpKam0t
shNwMr5QispAb6GyiotN3bl+1RtJuEBtwIAKBFk/owZaRVNOAt510tTvxoRH9MqAwvAZLkU5SJOd
7D6RmHgQR/Em77n2bGcgW4E6DOTq31xupWfeXpMQFBazqLN7z6VruGLWkOM4E09r3Jvzey5foI7C
FgcT/3PoOT7iv+4x5skCJuyVeJip72LiYo8ptr9fIsQjqBToaBhSVIAqyDa2rQFcBf6aAJedcZu6
sUgoFjzomlq9+ezL+zEaL/aqkh7P8gP14Ywc5tkLviCi6C4RlnKylvkr/Qy2XgOSkYjHKTjSely8
r/4XaAvqVwFumerrgdvoyMPKAIF9kSWVm3nqpmGXDqKscTQXe6vl4KbvlIfwKYsF79mzf8l5M+tg
ncUyUb3A7URSMl+aoU/k5NSc4eqnbTIwo5q1gRMpz7R856xxcIIp79UpD13MvizUX9jx/ElXlfKR
bHBY+ZW8jP8kPtAauGpFTxiS2yXVqlZ2fQuG0sjr2apPKe5vMFrhMqfjCY+PWuYbbnog3GauUuyx
VDH4jLq5SAtfFOOXBxB18QekFB40s49BqjGEPjFUo5r7u+jmj37ezoff4jfoTabDoiIMfzY5QION
bYL6frXsL7E9E3r0qaMgYO9wp8X7pE9oIEGp9X9aSai/359xVwky+56Q+aHzpVxm0x70U1vdHC9h
ofLBLR5tpuiOwUsosu6r2+h/2Qezsal5u0jAvztwFVub3+UFjba0GRrqQ6dy66ZjDqwYAn9dhJLQ
Kk6LJglEFWWMlJunBymVywV0OEgZDA+od/ZMs61rmoW+wFJHhju2mQR6keAT41yB2OQ/7wkplibX
Y3SAL0sKLwkVyJWfpyuKXth2HnxgMgqO/biT9ahcyV7bu4YqPdPfGdL38SDoPbdQSwiV0QBKQj10
0K/utRKBVabJfmsmo3wIFobwzQJ/NtrNyxx1o62ES09tnA67rElXkr5JP802+RDOeVUWlCKxHvCn
yDtKasd4ZEfmw4Nd9eOwvbQhkQf9Vw/Tcrj4/zodqfy+41cSjjIf7COlXpJsGVRteBYUpWQkf8me
2EZN2sLTHiMr6MIJVnnVZq05FV20eFG468HILWo2TAvjSpo2NJNXrp0XXqpXYeByKfkUNNQr3xzO
ONK+oAI+Eq18urewmOGGHKrewRZl+ulRvt7W0f9aBmun5FX6ar8gX5Sha6r+qGT5JKihhjmujsrg
OQliXWVc75aRpWA4f/UOkDVKaoBBZmG9MBG7J2K1vnfoxHKTLxj1oGR4gaxi/h3uQqY67tYQJAw2
veirxj4AfjVJdfUHGxNBQXfuI7CCE50LnpfFBzOe+GWtgngzYzCqdc3SLTM0OJlyo5F95OIuCsYJ
oSsspAYlTPOemACcFkFzbMk7WKCCz/HF4NbjWh6W8LPi7SWUl3f2lgqECZmzDtiqR6PacLY5a3jY
0HTfftE/arAW+74szwHeSjFdry1KTBr4AVy7EiIZ0SJYz/i1i4GY+tANu6F3wJd3vm7ea/nShI0r
Fb435Hv5S1RyyTGGcZg7/Qkl+i/AnBW4Ul8AfDZ3MbJOE2uiS2PQU+VOOevmeu36pvN7Fi2Eps5U
UrX8IdXqlqFJ5dJdXAconwi50BNjIBX8VRu//68nyaxz9puPCsXbpDzSh3eZ7lka+YO4cseHeadk
RXj5YKAS238P2Rd0oQTs2TlwaI6JOMFtVLpOY9Cq2GrN45xoGcRLWhhJZwsM58tgBMsLEeM0wbr5
rb73mEDquylHFHQ4NcmMA3fPk/1dPaVNNfnBklTe16QfwMKAQh17pTYHUnRGdPAe96T9ArBFHZXP
mMeen7Ic1GKDphombrGhSDnULqMU/LejbPpHB/F/7BjKMl1xbtlu5INOD4EX9YaWAOXkTyW1Dx1g
D3UgXCK0Hb4Wl2rq0iEQdvScoUu4tOHHFqONPPUrZs09v1mMbYjSKOsix84fpd5RkpTaf2zQsjs6
ZfmgL3TFsBXoEtoC3l8vQjfi+MvWTxqzL/TLjaGN6DAeZSExb2j/ZvGKZGXnR4tPf6Q5osz6iNLg
Yp7aw3BziHf/Pb+8/5Mcn+hY+QqzW18LBKANAKbEUkw9dt1uh/sGU9hNfD79rhgG4vGsbtixPORN
u4243MrhT3tEpYRanMxLBQaYWotbPAoG02uth3+8m0DAKC9qZhAtULqVOreyFOuKsq+ppwlrh5Ww
spr/P4IZDt+TsB2P6gC0uVfaIxoFbI3q1cMbL+bpGechii8gEyibueoH9HdAJF3vwcmj6N/ffiRN
pHa2pjEstR3v0p3qWcn+OnZSYIY1TM/Luamz4waiHFsAW77b25J5M4/pmBFuzbkm5JoW+S6bue3H
Kh4F0DFSci0dHxEblUE+BDdpCp6N3k0yXjRaQ/+DY7iWVxepuRGf96lYi9QaY4cnIxUNT5iDNZ5f
C7RBahblMxwkJthDiokFBabQ8DQdzxlJwa1ZuGFiwQvgMgmJZFNGeQX6zpGacRIZ9Xw6K2kfQHni
iCjYhjnb3SpoFycOLc4hbjyLSVA9QksIW8XuKSe2KOrM6QGqnVhus2T9xq20nnoycPMgzDgCUH88
cD1WuQIC8XuV3rI+aWRNmnyuucyTlxRo1kHuwsSbm0vN80jiIJdcj8KV9cnvCpEAkT1N+1N7PlVk
AkmdPUimxXzG6wpIhS+HiFEzR5x7kGuxeHUsuq8XOcWHMrUcTyzoQ4LzTYVZFclhX/IUzJC9zDwH
dNY3mOcSYYxKi42fOjYDW54hAM3zgO/ChjSXCm9g94Qf0ET16j4dkknRoDq6DgRBNr03vU8EPPO1
rs3szaZPQdKqN4KlKE7r8QQsj5RtjsgVOFZahOROjXtMt+p+zNgRpy0DlUvIrnQx4ggmYMZtbqBO
3g3VeD8fXGuvFp/C2gNTn9TrMHFdwz24Uoo0UP7Wntbhp1TQjF2t013hYEiMtvCvckt9zjzPfQ8+
7b5lac8OMULzOw32J1YSjlVKzxUO51px6bjthhHoyNL7kCCXOKlstddyrebfPnLeoQRWYAxILo1K
E2gLrWyRjK4806SyqySxb1324QLQkIRt6chYS2DT2iWtHsVmm21K6CPZm1HTj17D22jezebdssSZ
vAUnOkhMC4/QBy42s18GPtVeEJwrafjkqtWYPqQFqAGF8ykLSN+8AMqqMYfDDn36MO7vLHPNnUvx
91sLPLQUM4FWOhrE7yI4jJGS0sxFNsrc3oUROVPOiondEzfbMyENE64rmaM60SzEIIqHkmxj5iEE
fja4fna7kfMwK30vOGqpsN2U4+Q3oBuUoFz2O2vzSeJgqmID73w1GlB3RLEDttPW2aNHeHpdv69k
rF8HIdjeJgSD6lqKMChU9T1nb/T2zSYrpezKC0udDJ+MSt1tkm1y/kPI/m0zsSCL5HKAJF48keX6
Swmymd77id0gQ9fdGNyN6Yq4ZNveXj3WOY9HiVor9crOUJnGTa5LOxQHaJkXCspe1yIqw2pwSVNc
JKkkLu5JJEZ+qoUeVXiNHW8Ft8RFSJxp6bTZaglC9OyrM5s3BFDTS6tgWDgXR/HhDM7m+nB5eWHO
0mQ5rPcwKMhTvtT8jEXYvywsMNnOZEGQpg2eOYvc+bF49En+it245Pzu5L9zPh8JQ82Kf/456rvr
lVsM9gFDr0nEeAJ3P7lyNqrbTXfhTmfLXqYg1Eef9+giK2sCZF5Qgo0RNrN4qocFAGT+E/GHu/Iu
8Inrib7RweuUbtMqH5cS7yxQ8QITe4iHHBQ8AI0Cp1xbHZhMhwuBbQ5n0eyKNl+PVznCWxZHMnT0
kFeqIIGZn/oNzqOj9p7kgm8CyZmoZRij99l3553iuR392mBabV/lUfTWyzuHYHgl2eVLCumdroe9
359JUnwNZR+n5hmMmhT6zwSHv1aTQR5i0O1rXOuomCOkGgPoN1t3yF00INjKBQ3YqrLf//dYBKGN
xo7mzm1PieHCgKG0FPCL0IzuQPu0UEMDiAG3rgvwSLB9sHHAFrOg4rJepr2xpiO71lVOP0rxHkAw
EMtUt695PJ2/3LQZ8VvX7J3ftDB2FcmBHYHB94X3yonfOdBQ0fzCiHaKq1ouZZIl8A6eJFNGNBZA
mNmWzoC5IQZRq74JecxdD5T5NRYtgepv+Y92sdA70FQCPH2ZfY6OGfOLhEyN9e/iNnET3bPCAm3E
XugvQImrYYtbsNKn+XOtIr8eOrVW03BglrNmOemXwsSOhwpzlzus/qIHeLnPbOz2yz9ILPq8ekuQ
BjogGUq9zImwbfPV3FgDRp/i23JVnTa027cHo77ASTb/cJMBBiW9C5Kw5rp9rP0aEFWgelwIF433
7uDiInpPF++I89nN5tEjShWzAj6cCvy2UcxWpjmOXH8mYfQu+SjycWA/jOf7QqxvAN5wML4ww5dk
+crOzaJwtPui8jXBTgtvy3RnljJPTaejK2Q8/T0ziz8+8KUtp3JYY9AAAxen0r9OAdw6mbQZSjXD
5YjPkQnCLcLqkIrSrGulHk+v5csT2tfN4TXMwPwmhLli5nrfMQjCviDhPQ6ApkhKOd4O9p7caq0H
CyW63d9f7483l2hGcZDqnXnBzSq4RJPTnRRdcaxxKdMNzUXJdN213PtS/JNBE0/J8hLVNnyyb0nh
g5bIvSmTlWk0M2j/5XbUqKKUQSQG71CvSuNT9FtXEnrflG/yCCkeuMXf30fbiqMpx71XNebrx210
0Vx8jq8yqPZRISn12OZrAkxgEpB/7M5JwZzF3olF4P7n3aKqPyTpUgjFQbQXskpB8HYLK9HZs2d4
qTBUc7nEG69D+ALHm49Fjf8Ipdz2hkQyJ+XMplhpWPkXvZmwdw7BNRoi/56qswR9E2z675H3yOnc
jePX9YrsQCW9prL/GqTMhsWbyM8PpCtJXJH8w/4zNa/AaDuKcCPqeEE5cueCzHqHtvuEmkAKotRB
0xcKyasjIWddDVSlbgh20c0LXk07oSNH2uKpIy3A9i47Qc/Xzvf3CROlibh7jdcZnMlWxwf7qD4w
mtCKKzYG8FbECnDwYpiWN1gPVKcSQe3zLlNbreYOMob5xhYRsNc8RRZnjjJlCaOuGOtXlfaZaPIQ
dnaLb05qJE3+mKawDXjoIeR9aK9gMUE5AHyMTSMb0F6dhlLURlEjfl2Ftt/OCpOCHltkdVOD+m7q
6QXfCHa42jyk1cPnOxLt55DUDGs8gVH3ncJpdXizZ9e9iHqr2c77ujT0kd94o4OOkqiMy9rLZvhE
OPBmS2AsRSpXWHGIbTvVGT3VqZ2XVXc4FJzn92acRK+eYCro2b9Q1erlBj3gIKB5yZntXI5Px2Zq
grlfNCduR2wrpumWd7FXDmexjPJQH6TgZT0/QKlvZ+c6IovDgBWhPFu2+b9OwcqC/ML5mnuq2KOB
nE+bj5fR1E4Zb9kLdDmo8Vx6NrSyR0R5ND/cBNw1sbO+nZvAqiv9gbXEFXD2qT1eywGNOLb9ApBA
IBo8jXs59eS+1bqAl8MrC6athGCy7tsX+TL+eMn2UI4wtsJP8QQR//4aXFXf86Ad4VLLl3NwEp9E
GLlq8x5K8OXHiM2D/SdnIZLCyxdjcQHrsQDvVSWJMYwhlc/A8pVAFoOqQhNJI4s1xTYNjbGTP67x
O2dabSaLIUKZcTm2lQyUlwoaHv/rvVqyU/8c+l450kBvctGCZxXQteY5nrmRqrd+2PACo02t63aA
SNLZOjaI2zsKUKUx73by3psEGLHa9NyJC5AJgaytFzo7qkJR2I5xeOf85le+tML/ixZ2eX3ozANv
R8RzyUBJaS6BAwOfIFPuzsSYkItygJZZl1gJztwYKJOgRp/UhT7ftMupdrFc+jsrkiTHCQaw1mWQ
VYBrU6JX3Xq6d+sv86hATgezyPsRdiLvbZqW+jQqF4OO9QxKCOR/hbI3TUT7XI8XqaIWcCxd68mQ
gIsm1TcSrhjIi/iZirNtkjOIH0cHD5JP6/JoN+KDLkGXKr3cimrE5OOVvOxo/5WIZyFZIGQnj3f6
O+k0nZHvehibtyteuSU7WRULQ4RnTWJAGgmaBCaNytWtv/9hdU2EYx9CI9ssVimRUlqn4jZrkzP/
w3rhiXj3yMQyU258CP/YtcB9VdchHc7OkeowYFbyvGNXT0CfVoMYS+lxyVzkv2XMz0MylMl6JHeq
7meQ9LxBiULsBhWR+mzyTalAKEFlMixmuIgtBisn/SAvAMo6IHMJGjpLQtj3blF8PRD4h4AdoBzr
v8nwSOvH70H0sGCryQuC6frZ25XIWaxgcbEO1KbGzK/yyzloM3K7tkOGh7LICo5apnpneBHMfBbn
OBkrDLCgX0MrIAMS4A6ZagUF6Ku0CYj8HfMMZKpvaNYjJVa1Rzwpz3Qq5y/GifE6G++ECgJryabQ
O49FLCVIgRz8EkIh+abmTbZs6iyMLfytobLPoxWXSxAZWSEf/Vc6jWDz3LfibQ7AE5RgMhVen8Ca
k3bGG1G3OVL1ZKdUSa7It+wQH2zCw8oRpJLCFlJEOun0fcWy6tHzsrgi/2kZ4Bp9JyWz77ObduTE
NPrwQ0sYqzd4rbvc1Ui31LR53UH+Rv7hY0lEanHEdwiGdN5VVs/Musa9yV9DQY5JQumqt0ccQw1r
PPQjy/cOWcRVN0RN4zWX5+jxuSUmk8krElEdduN9vtKEKACe+S0FETRRry3XDSZDxbAB0a3tQWNR
JNtZGCaOhud+ERqiO+t9C3OwOeFIaoXi6NMVOV3Ph8sb3h5zWzMnfjAzpGGZ9IeHqfPMDN28zqmi
sdDbcJiM21UH/PjroBUcVUPfTbP9CrNd/3YhfQyVQ5oh85ISy2Lnn0DfF/hu3Amve+WONkHqhQn2
XWmHEEVdYW6ya9yWGnDBbyoyVeq8AH2rvNXcBCRp6QL9oDCIw5YqK4rL+NPnHzfCTckXjLIWmOY2
2TS9ZOqG5vcsx5RWK3A35E9n0mQxcy7jv8Q28Y2C6guKuWio2okVR5H60a/z3vKyr23xQkmj7MPI
dT0763X69TBzPQQPCGFeKuUmhcYxdxxrqvpd50NMsYvQ7Yq3Fgmhp7ii2FL+ky1WZk3zRa7A4tHn
qwTpy++OCaceId5qpQvLb456nZzkE4IP4tor3OB3aGfrIAl4Xme4ouNr7z3Y+LVsQSyiLjBSc5x+
rV6z8Cci8OzbX7HJeUg/KIyPpKCSA/avu9YJfF26ZQw0IRo2a2n27tWRfBqfSnYKnCQny2p1WdU7
ump1Ekd3qprHdimm0WX+bMxmw0U/3gjC0jdO4z4Pjn+UhIgJ3nWV4BvoNLKGmxh2xINUwLzuQ89f
tNJwEb+JYB4adUd/Cg3kxM8/qcwQ/x2cgCESw85fVTDZMRwFZq0I4x0tEzaLA/OzWWFYuFP3/8K+
/B5mTWsGB7/aUxT/vD9OH9cr9mRYJdUCZSKcIf/B1Q7TSuvcadpKkcHzLPwJCOkUHYkKjUldIi7Q
ekA3sKVzWQv6758pYVj/cUHnDaSk/Ca9+G/izoW8DJuD8OulPTzzhQ1bpeYaL18fgAMvRAPTst11
zVQoXIz+lDCcOgEmAg2Zx7LJ1ojBxTMsRLxWkP14RR9wq8puP+sVIWIJtoXH/36e55ZvJwJx43Ms
2c1aSUuVlB8w6sQkXxLfBAh0p3yf3mdZHqtZG5C//BcYE44XRNiX6uohSS89iSF8TIzrbSa8qYT/
JCyxzCvMvDwL+hhzJ2qP+O8c9PlbmMOLjlmC09a+ev0ZBsnn0IsIKNes4npZd4NCqH4tPOlISv+y
zMsuRLA5yfROSO4CLJx3W1hCfGqXhdNs8Eh7MdNxddXYAkIOre9Pie695pub82zT4HAOg3X2yUr6
lwImXa7Yu9SqVnsT8ItRxQ+o3L8KseZUPrYGlZ6DWSbQnJn+arYfvz21zDXQ8j+lo0FqtQ3J7hdN
J3DPsixa2MY7cJblqGDpDw3/REp8W4kCFNiEQj+a7ChCDuRil+Ib/0M0NWbBLqjxea9QDeBi5fw3
jBaw2rcOkxA/iC8q2KfujrvFGXXvkklDqkRXoe26Utg1FCXAfK6tBTDVo8q5Ukf3MVJ9zoMqLB5K
8o11uEGxOqNhHMgL73eMnvKxvcp8032zYzdbZvoo7q2fxCdcRbzDaTEHXehDp3bFkDp8MzxNCSxj
g14Sz3rpObefQ++a4p0uUrBKVf6F2PM4MMNjTbkspl2ixwqSxt9wYZ39R59PAtMixXpEn8cwcyYe
sTURluExRkV+fFi2hJ7Ch2gcXWFjnxzS6vNpBVmbK4WbHC6vOh7OOEGXks0kjEM9go8zOufVjtzv
mdladNHU8B177Ye3BdxBBzce0I2/wiatr/D2ob/6PF+uqJDjfcYY8GogIC1XVcBYUL7X7LtvbAJS
M9zlqMxuGmujtP5JGNmMa1MhSsCeD9FINiTjvF1ZMGA+sAh1SZSXTRYjRDBSzFLPemT6IhP0ETwU
Vd/2mXroEqaENFAmveVRPVcZ8aomVGLKeKNND6FwQ0uSinj6lT2UqvFhvKzkxAXIsGhDcuPe7mgG
MipKxi7gpC6ReougnpnSV7OpRgZQ/naZxdfE2uKuIhus3HMcoRjRj3qe2OpHWPU1vIvjnD1fQ1SR
vPgWVfbJ9USfDzE7LxS4dKGow3Su71tp7IB4+X2NRQm84ATerI2iBOye6KYa+B/Yxmc6cir4fPy9
QavNyXxoBwEeqmd+SpxzWVQN6n1yQzmFvpRkEbPp92591RAwWacbV+ZaI2wvKrGJKRrl5STSN9Kp
Xd07R+9YD+lnz9A2AUd/JFPs1k5Eqes9tnld7uYiyxfhxlh2ZkRB7rBu/xyBg9cVdmRVyZfj29MM
yT/xRnEucJl9+yQTcU4RJNIM7ix4i+XCAg5Hf3H6w6eOcaqlfIbJwI2z+encuTS46MgqXWlz4WKC
az5WeKtymiP/h0qCnFKEsz2CQXK0WiyRvBkdibcG/nuogT3TLacXVpFzGTmM9Jp8sodsR6EeJx4h
UW61VDVbA+ENVgOpDLEJ+2jwRaHhh8hc7fCCygCHtZOBDjczYc/ufRPYS1VTex7wkEXbsbFCRK0r
xe3cPCKxsZjFYMLV1vxfULlfsNO27eLdNJl2Kd17jxPeZjfeNW1H2mqs2E4p1LlEwJ7OeY7vROAr
g1eEUYt/TPRigsz8uSNyPEY/pcMDbLLsLM9V27eePIhUXC0JpFG38LwuTZU/yCQbwheSJrGpAowq
w8JuEX6ipmY10e7HFZf+Iwp9umPvQvWEfvjZaN4PlTmr5z3X0FQNk2lrfHsuYSxhNdUxnZIGGBpo
6Bg70hKl9dIuYhOotMJB7DkdvJu4LmnL22y5I5oumKTFqHBl2hG/LhOvc/BaKYhKuPrq1VkdN6Tx
W6pBqJdQVveCrzWElmEdxXQtoAeoqIlzsXJn0ChXNBBMy7Kqr+jB9pvW2b/jZ+vJ1mliWONyyCVc
+yY8BxFS8R600QIKtEr1yF/L1r1uqJM+/OXjnlBlJmkWRwqaGQXJIo4U1n96YJkfgWN8a+VeD63g
d3bG/sqKRaqH3T70kHaGlJucbS2BZrVWSD2JHrwSlIkxqKmY03fYpKXuNdul2TMD/VLYiq84n8mR
KXR8R5wxbFVm24taRyXFnR6fzmBqFxn1pvYu6MW0c23DI1bZeGLNB+badQJyWtNcBTVboX6KAGdF
2ClBdr10PNUR95g2yO6w2wGMWUmcMIWejBBt4jSNclJ/uQPhNKcrTXgZOX6TvvPyyoU2qD6ZQQEG
JMPqiD/bug==
`protect end_protected
