library verilog;
use verilog.vl_types.all;
entity Video_Image_Processor_TB is
end Video_Image_Processor_TB;
