`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Y4RWAvYjBGnG41B17t7itgqxIOJXGz4Xs44tc60vm9o6ziMbpO6vASrmn7fk/dQJta9xgzAYHoZv
VOBZw1E9ow==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qreEh1uz8fo1M7xuhJDuVWOnziZCxCJIJ+v/fW6AFrMOrPi4NhmlCaPFvlBUYJv68V+gD500j7zP
EYOO4tgNGWFba/kJsQbbZ0DAWKfUxBJC8HaZJgcrydU62++02DHUV+xRRJnifSdnQ8a1j5AxaWrz
Pat4ihE6dODmCrp10Y8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fKJ37zNFLK0TruQrvW3TtIQsSngl0S4DBB3O9RkrdDc+NCAsCxPg/2CpTnXIeg1OvnreqtyneSaX
A1Ti1C9TyeWIGqJtDFM7zRGaRlpYVPNOSpzN0RQg2/h/6GTglolb1TCgaJoYmGgtednDRawxd+YI
I0vtjukb0OhjrNB6AecZ/4oZCRnoBIn2UQuygbsl4aKyFJgCUkLB+vAKN3E4Ivz12LJCd3DjFJqJ
3OaHdPVoku6IBEoaeymD4P1c3TECpI/w5AwuPlyylE43CgZrCB1VLiYrn4rQUyd6nWp9G+7DTBb3
fMISxI+YKFTsoDb+5+uKpm071lkq3NiovjKg9Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RXkStlwcTkgO3NvOIj8FTU6oGT7F35iz6DDvF6S/qLQxsfaiND5r31FcJ0PTWAe66dT9nhYL5sX6
tFUFr2gTf5Gr+wo/ggls1zCdlGeHqybKRD/qbLLWYCic80TqeMXgtfOAKMjDzEc8/fMDq2cBIKtK
4wCu7kbvIT4xi+TgoWA1B4Po8GgPucZcOy7LkqfZMu4r98CPHSkoHKXgfSj9burC8dx8bsShdYYm
lAu0FBscwmRx6KhLzQsHxdtdaH0bF2QfwY0m2L7oPc+OPw/KF0mMXhsTvYORetK3d9/WFyrsn2ji
jpGEsJxGme/+dy0b6i3soFhwu0i6KKDW2nBWnA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qDL/Bg4amn7mlR1VKzTtu68WQx/BftRW9t2lFUujHVMDrn17KtYxSIXhRO31FxvFMseB82lzIiQn
vC2tbUchFUHQNm7x48Ac6Mr4sh2Z6iRfxubzLyk54E9TcNLZVW6TNjpzG1NZYxNb4qS3cBvszQjP
1XvCPSku9lNyRC6VqULGS4MSRqcZp5BN1u3nxEb1obT2a34DYZpp60+UDkM8U1iQPrM+jWB+qsGg
M8ZPdostWr+3WXP8FqTByio3kHHYc7Ao/PjKZQHfCKiIj2SKJyS/s3up+ynE8SLKkhMAHV3azS2i
xRqURZwpC8rIokUiegLOfOhIYLRc6t7F+RHK3Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PmG3GCErn2/zmzwtvFG44CEeJVF3aOZHti5qevMwg3XI4TYdJ94u7zwF6sbVSufFmHB0Gb6TW+90
m9ZUukyXtXMdxOnPq0o4/YLyCXNH4UTB9Z5tiqWj+lyqL8nUNIVvnsmt/pdiqTo03mB8GS0s6DUh
ODgI4iiGm13+EQUCKOU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aRWGZWJw4MnlKyg+1f5Yutz/SvHSEor+l1bqzjwYG5MW5W/+KqqIh1XcHWxfbz/B8vUVzsBCT0yu
SmElplhqMwytIRvZ9jVLPqy9+jQ2zvUGI0Zv8+3+HvZi48MD1l21ZDorTquMcfHmMHwsDd7boIqf
4zCW30Fau+H1Z7IOPvrsxZqEi//2E0rf2KeanBMEia2ecOR1ttDeyfCbg4e5UJj0DbW/XDLfEmfR
S80LXenYJ8RP/DrkJEIN+f/To4yIqN02lh6k+a74RZIyF6SWD9bEjMe3U36Hf3ew7AuW4ITCIiGA
+LeuunRSYJCoSY9ikU6OIo+YYKwqwlmjKJYIHA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
MjBWKTXfcE2eJwjypSJszf8ehUl3CvLOHEAfywiB6IrR7i0tV9oUQU5Amg3ZALW4GiiO6TkmLLss
68hwnHsWI7HMVtmYlBiBwnBII3Zedlq2MxzvLgkwDUNdRtEwi0MjWMMNO3GNs5l84lg8DR8eMk7D
pcMYebUD5mGqgDo6DVb3qZ8HXw/0KErRfTY6XUEom1gUPhqRInibhR/r3YAyt6R3n601SZqKHyu9
xxyh09EtljXDQCs3YyZILr/koFqUPZXONEpCTLH5iZUsOSZRRtR0KhC/64AB9lYd7u88mO/tfZ2S
sGSFXFaU//Pw+zVgKpy2KUcHT2FU/i4mwVjNeabsi/D2g48FIzqqyVUQCvTtT3zB+eIuzj/jtpUk
4OeUEJEcYYLMca1bmYduu9ttbdPXRXUUQD1dwjyJIfDsIQQuJLsbUGZO24uUDS1nxfIpkAQzG+Q/
J0jHvolTRpZH+t70CkSXdwMAEmWYbRWwv0SqaLU1R7GOSZKkMHg2SlREuHO24Iv+HK9VuGVTsf3z
E3ah4S1/f1Ea6ieH18ZERyEDlBBuRXWUgdW0tH1oGH1mdZsjwkGXVVCkTrg/ZhkDaQSfq5KanFJU
WX6Z5MkYpFZaQVzEgMbn0ODNz6UcDptE3a/ubZV8MbENfEbeKEV5f0ewM4pjap9KLS+GapxnbKsp
K75M0OlqWWExCaudrjRsRt9m0yDTP2Msk3OLbx+u5QtisPj53bUxyfwvDzl4J83ZCW7ooM6gli5s
7J6DcALqsaDNqIS62BQXK6VXCGEXKj7YkjOo7FOmfUd60SJzALPcx1B8Qo1g7//yE+FwXMamo9WB
jx8z2BItJoGNZGwoBN8xfoNTtAHC2RAcS4C0Tlju50JoW98eGUupglhoD63n8DaCRskrP+4x34cP
yTAz8LxzPPsIgoiLwcBsi7fuI0dl7haDVgMIMbwGF4UbxWbl26VLaxW0/n9XbvI5FUj3+b4HcvuD
V8oRgqcDoaSH1506mfg2rdROt677EpqWKqpafccOPP7PUI+pH8fFbsEaPfJ03Cszfs1h95gUAI27
hb/88Id9HsmA34LbWKxYcZbXBT/S/g2wi6dYQedv5bgwQqNeN3X5RfPAUIDuulfLsO3xZZTkqOQi
VepN9e6oFOssEJrSuXSPvTGNxBqjN6JojR5lAhB7O7DiJ+1yrCR8XBUPv5jETihOfGOgVRlMtvtE
S0CPrrd2MdBZ1W8nmXkZLooKQkyRb4wauoSVcVj/gbVJH826oNjruoYaYGE0OYZ6P8DGs+lE4kkr
IhhIcyjazKcx1/RjoH1lu10zvEsJ58ofr+5VXckI4ql6+br9SzTGCZZTyY/ir7oeGc4YkfbGvYZ+
84hKl2R/kbj3riTSsyqtBVHJRx58a99b5QAIY/ZZbClfDJjQtzpBwJOEujq1Jdx8pzJR2YbqiEAs
enPVghEup0UCUmlgqtLOyKpXUU4DDB4LXJyWOCguZ/IDkMvJ9MxuNrcG3e9/3Pss3XpvclhdJ5Pz
LxtaMQAmUpVA9IvDzeM2ObFkF9o+gfZjZAmzhFQAd6Thj5YYi2hc6itdDQACL5Tc7RueRscrUMW5
pWHHcwktHpQ9fJe0Vck+KR4JkO7SllsmgRn8U1WLGY6DTyX0cIfGf7iGMVZs6c6yCyPGLHo/jJA+
TdZQ2sh3BPJ5ELP8KlOltqB/eYqlpoNXNf+NZB2wvq9r1p6IdrSfxYqqKY9RGjshlvB6rAmJTsSd
jn1o2k+Apt76eFQH4BlIdcXRQ/utnfQg2kagK5QSA7p/pj8fMd3R5/FWbLCf7FjXiKDx/3ypixMv
MnFdMW0IQPpcdKqpCdNCg+CVsBFdj5ughXLb7fGlNqOaFSpC+FQtDVFhH09iQe3LJyCT/g0tlMsy
1DbG6us9/blx078jHOTfGZc0J0UWsDQOmPludaWX3ZatjwM77XqrOZ6/+18PMNpi6KZmFk21Emsu
RPPTw+YMz4X7Be453UTy9/6CODdQWRgN/1TTXX1V6DAsrIutUNTsLv6c6uvdw1BntFq2o8libx1g
aeD7JL/oePDt15KyIK1EUnOFkUX8BlgiHXvK83uK91U1dCGJUbfeGVjz2odN3XDCU/C8pIn9lXeX
s6L1psYddZGtjYpLKCA424MmGsyCyTjAP5oekiIlJwFXQyKeBwVovKpE9b04ZwSexNN/tAntGb7x
wU/p2rU2NYSAB5AF7NyzFAqxVDnqJMr8m9zCx6o3GlJo+tTpwPZZDfbC1L+6Weor5bFb4cerRWLs
P39fs77hzF0Bj/CGMzNSnEJBEcCqymYkYKsO6mVddc2BA4UzVSZISsZZxUs/mC1o8RAP1fYw56WW
LiX6x/OM+wcN/aPKMQRfpMQDvuB7NVwNnPxZyj/K5sWRpuo+P/z6LwzB1yxpvXyJFcgYlzBAxseq
KjGSwvams5u+0Xq25Q7dJXV3CS8L/JxQ/Mg3BlSCHGDThi4WfolGHIAfzzHrP4truO26XrNb24j9
T4Ry6C4qmlAplJmpUeODblaWwNG3zZZ3Inmx6VrbvrkFRlepXCiRIkA7qfaVFYH723sP9qYJnvjv
mRN5b3oEaGxueI//nI3vUY9E/yiXnim+VsMVcgElFcyfyabKSCHfwk++qOcp0NgCsFPvHKexzsSj
tEJFe+1KXIZ8uoVZ74t1YzLAktxvWRp9h6qYgxJlg1czA8I+zn720QlfqTrIf88/HHBka2RK5ZvB
q5SALDdzAy3mAngZCLHKrzYTALQkvkX61X4RhZ44j04ZLfU8/KVofF2uKjdeRvEQ7qDiMqyaXpaV
hdu1ooGdroxVW5rDUgcrbH30XFbFGfCponA4tdd8JB6D1tvWbPwkNKhpTW18BqbmFxyEiawH8OqY
oE+3/AiTgepI30AJi4c25ihINnFXMh9zl6Kcp1ICA9faZbDc6RlZ59BKsfld8pAQZQUeANoNWuiu
Moddo6x0QIJHod8O7BUfFmEcB+C1cTLbw46zL5WS3DiI96+a770W4J2XZSItLcfBovw2KqhLAGkn
q25InyFEHvzb367A5TZONu7wqxJDMnY4FEpnlleu+XuWZlcc5TVCijifSR8Ywa3iCMS+LFMaYCWO
fBNIrdTVBi8HCfWRlw6xpktCSY0AF6bP0AZZ2jHpEq7oxIZEbI2N5bkH0JYKmtu1KB8fJhFQZCo9
zITfr/PMMlPFT53Zts57pBUzFXlzjXPgCMRCaelMfhwrkEfC6dkhbOXBAMnI3VAofKXaMaTBZdkH
pKqqnaV2MyicXadTbiNWyfuwv+Jc5hi46dbScrl6yEMEoesuqsumRZW2BFO/z33mDbDi5GfxB0IY
7kYekx4aYOWcPRVfWx8NzqbXQ+uxfAguYsX6ehMQgTRQfPShO96X0c9GJfqi9gEq7llu0RpatFVW
Y8caziK86rnXaKZiJq1K/Bk9Zyq+Mup7gVHcsGv1cJ3En9pM7N8n9yoNX6F5PDxzPKPCFJxbw5Py
d1LLiVCllq0p9qCNkg73/SNpEebcqY2pmenv3dqWmqXle1lGJDDjIO9cKqOlkNAdGaApa5XcHewD
Kl1Blq4gSvZx1n9a8pokSxZtODz4uDwDpAa0ADDnjC1P46TscQmzHqBUQyPEhVXY0IZ4TV5ZD2cM
OY2gqMvLZR6YNcfjfLPfkkJ5XVITounHVu2tRlxYCuD+4IYlbi/IPkMgzNQVqAzxbS77npG2RAYm
QWTiCIGU9CHFM0PRyy52kG4CNyqNg4/SHjtpXrJ8voML3Oi+NAUKjIwwhtlLysdUWpokEGhx+rkt
B36k2dOsXXB68hFrhAo0SAnoodW/YTqLP40/4/GxiuGTWYEtbigb9VYPdQLx1s8g/fUgRNFgtNB0
NiXyO17pG5Y8J2x/zkV6xmGQoB4rAWj4YRMNKSj7Tb9OA2xEgnPrYI71bRKYGUmzoJ4RQvFSk5H2
S30WwF8tiY7Yok/yi0Z2iurilZ7l8O9tn8Qz8FzhnravkHmWmwDWxcljbMXpU6xPqzPHiVLGiFbc
4cLWU2n3AHhuy+mDdnCUkiNZ1spwmgoU3vgu5yG3Xjr3vAl3tPtKhhFLBQdYbIipROcGnc//FRPd
5KuS2+5YWTyz78VxtU8xP3Qf32MecmdZ4XHvk4n0AKeK0QNZCgB++a4xUbqZNzH7U9UzRk1+YLmG
fHTBhJxjvXIIqQ+BPg68y21Boh1+uSQDNhs8QxzUaS7kZJsfaArZqQBYN3aQ7axUUIChXxf47L2J
hk3QXVX6/o6xJ0vUhZaSWK1cRjsQDxChhnPgA42pMG7DzClqmkx0lNNay6h3h8XaHS3y/oRYej4H
z7PDiDaXsgxWhprylPmo7fqxuvA9tI5PA9ocC3nnf7EEbwRvILR4/WXMQIFyWGv46kWfkJfvEcea
FzJQ+yTH0Mw3cVdWK+XN83b+KxFKC5HhnOHyImeNlVGziiwXvj9Sxtqrv5uHQeW0k0vN/Qp+Zfr+
Jip0MxwPSFz9980udFBg3iy4ZRryIkXzlRs7iZ8LTJknhV2+dT2kllS6WBAtDBzJCe15GMDfdktl
dLh7V/EQAH2AedUSWkTiccvAzR/Qm2JQqpXJIGioTlPIKrg2YRIMuqR2HfPsHwwuxUB74OQaP5TP
s6TCDXJgG1iuxf4fayecrkEi+gyUgd/mb7solbBXn5zLtrpu0L16LXpeqmfBUCOcrchTvwwXY1SN
IX6jzevh1PEIf/Vew7piafWFZG/9W4WDVCSfBeE/VHTM1ROkND1+AipTgcKB7foO74WCM1b8pCL0
a/y2/kBl9qxRsxpIj3i7rsHP/O8rFP7982ICwm5xVLEoeX6YFjzU0vhDGe+4aFFOpNsrMOvXlemm
PjzScZb4W5frpoqJuPGJHNcsToI3IEvTcG84PlzDWMfdE88oa2ZGY5Yn+Km49O0DseKJAHVpFmpD
lWIDGA9/KDpBfwS9DNq6vLoF6bFVrHmzavo7PHnvXsalI7GVVkk2wMNX62RUcaehOv2bNdP3aTVf
Qct6rXGVBFLtC4DGoG18E+N8Q2wyiP8TwYedR7DisQ+EYbgTZV8uT4Wf0EdQpGiZ9JfMW9YXO/P7
kTkkYGO597QbseFfQb57Y9NB6NvTe5sJe5g+S8hZwirBuRWHy8OL0rbS6znTFqs3s73xYHXS+RTk
FJ3rKvYNNFa+IW1gZgVAhVarqE9mf7sh76QwP9KJZUju4hKr2wyRjBOOclHdGXTJdldzCzjo2zml
9fYy+sz7/wgc5Gjdc7HY4ijmi2+8wepbajMqbCHdS75SDEjfVvCdW9eNuqwsnd9e+cdTuiU49AhG
mEHG0Dp+FcZ0AZSKPdXsyYIad57G1KhnZ0TCDWY7kyVHK8/vQ7U4xfQghtURl0yG/GrCouZJMSrZ
qrzLuqe1ppwj1+uDQfWdepfmxKAFpg4pV7YWUU/WhEVyw10HdvPNpzmNuo+KSIW1impWyn82gA9P
nktRVKoVdWl/06u4YX0nxufk8nYrez/roHuZ1H9eCJesxjRPuOEiVV5xUkTk2rXy/VQntT2dm6GO
FSB588tTR27M9/Rzuw1Y68DuwK0IxoD/i0BsBCUGJxtZ/VFwnIREldeI9RKuDqa4ms56EbkNq/Ae
6xo7zvCB1m1yO+zUR6pX44RR/daC8opKHN4FHpya3CT5LVYZ6xmSNPcPWRO7+SP3cRIKulESV/Ww
JFau70nGFKcb86axCTERTQaLBeUF1SvxvXJNvXKn9rBUixVhh5OvoSYDkz2AR6dx/x8TYl3LwQwp
CcmIBTKr3IQFRBHOUcj/uGBOX/q1mfOrThWRBQgmifSczOnxifIBB4skq4WgjJmmxSbq1lKszP8V
/NVKCu5htL1zS+7+r9tbpAxpcTL0QtZHSxCl/QPDchMiC3JOrFOd6bdoPFhjv7DEkOCY06FHZZQb
filWuICdBe4UElroDCstcIn30J0ocPiyTzdVhMRirn5hkFfj7bxu/KKRRNSCHqoFVOMi3klsokTH
VPO6vuZQr2gMP3/7KzXrv+SnW6bYfBQva2PqeHIj296kpN8Ueb1o2hRSEe0JHrdyhuodKgQQ3vea
iCrLVOdO3lO8tZi4jVIZGBRN6vYGxFALVgAcIfg62K7378Cmyqn03p31kCxiUMOo5zm3Lz2y14iM
Lt+YX5LFhhhujfceH2BooyWqd+2kw01LSDJdMY/3K8+RRqHhuIIVmSMR+pMxQuzjuT+UnlTIrp+r
O8ROBQInk1SXRfyUaHXwwh8xnebFCmliduZt9JjZRU9tbgL3o5SqxxnI0/piaz8JkYc2Vny2GEmL
A55m5RV/FdEiz5UMWFGLgq0XKYBuzZgZtDsWhE7IJGUUx1xHRypZuacZpdM1cfG8YQXJP8CDkCky
XDTBjuk3qzkJaruwf7I5RnQ9MUqNmc8nH7wzKmf0qtaN9KS6SbF3RqeJUNRTeqPRSk/LAWnK4Yyj
WlMSnB1XL3aJw0SV3R69iGhLrLu2q27aKJ+CI8crR7FcQsaToCMMwLLGrsfC1G0HCf/9CKdyxBJH
J9wx+nP1D4hfyCuKAHvonttS7nIHWYSFX02Jpj8yG5cVQDG4kZy7M3K9rdbHuHEbzAg2R+N13Lo/
2SnAF0J0DQd8o/wH43bH7JQI4HeQaokRZsYgy9def5SxcYZpyoN8hMGPS7xnxcyNmRttieqwdM7V
Ue9nnDSDfgw/Q2u9GFlqlvmQ42fShfwu1yd5cr9ToPkrPqY15GBO7lPlCUrjsE4pNZyU4f2KwSXm
wHPmmJAD02Ym9bmsiJNXLY9wbclvqBWJcTEHx07Vm37bDjyTrGN1uxkczvBVjStYrIfsTdXYfIWa
Z/m6CYUS3OzodnemUs0OCvysGGmJ0m7P6vhWqKAltOi/HQzQqp59qjxg3eUs36aLOvjNCivgQYjs
Rhsh+seEp5Z7/hca+KhO9ybA8LWyj4PMjYWH2r38qxR8YdEX1YSphrKJDV1ZE3XNuETxb+y9chMh
azj8Y6CgiHr956wyrduQnPh7/AgKF3HPTa3KbTU+ASrjgYqkUGZlV08QYboDuli60FMMJaGgTFT8
Z+6cpeJYJw/H7cDySGusv6YRPx68L5HBpO+I4zKSXmqqcfvyqjREtBC/OICoTIs+2BZp5xNZVWR0
MY32/LKbaY6CD94Z8FeBOR/SE2umybvcFPhNoy1QRUl9AsoqoaEcsAZ3GjHWpR0EyiL19xoicEdW
lNXO+2ol7yA7yPKyxzqELVC3eY852Ad42Ctjk6BuaD7jeboOwlhY3rdF5xp2NgOBqDqV1wQdIUj1
nv0LURFJ5HCkLR+SRgU8JBGBSyDChesG0TJDma5AVm3bF8Pm0KsntfWB+2U8Sa+V0uPmkuMOh6UA
1PzO6hKs2ILHLFGIK7oNCGCEsws1260ZXOMU1ZJGgr6NZ1YaIrfiuf2KF5yw/vA/jwMIC4A3jThI
ZEyfdZPn0bu3a8gLu9V/5p8zxmv4NCdyHsBzCeXFtG2GL6hTQyAmtZPhrIZAx+792qlm7FTwHUGj
Uq92CavaGfn5k7CDG+0xsiwkHKjbM1tbzAjaIJVnvnMVWG25MIOAz3azA7+WVl32EV4ZTlIg38y/
HJOwODTZrRJVA5UvJNoG/6KH/c0R8AOqTviLYSgc0DpqMLE71XtC1XFap01IA0qs6xMHf4YFrSO0
J2sKskCMU0zuHWsxenOzQNC/yKaT2a1TjrnCSxfjldvn53JZVgVbZy3X775WgLppTqeO0D8Hdvwy
nW6juITQQ9PsVe4mZqhvzvp/OTef8g/hmsM3x7vOz+gwJ5CTUr9jmRbMfCwhpoNOkLFqjZdOvhWr
t4TTBoJC0250T8YXmvHuBqusp3Fm6yAolrBDFoDJoFw4qsctDnwNHKysBxSzLmI88JmhM/4BYpdw
E4ODjkVj01a5do2YiyCZNy7ZMTGTI5+5sXte6ITC+yvMdg/RrK3V2ddC9zf/R+M9o7CCbw1RqwMp
6cYWbJUBljNkPEUQgM46HutZqXXn5WLQkiio0ZWuktbMbyc4vy909BHnJIMg+646FyL8s1DK+oPm
RZU9kWYbcEdyoSZTq8uZU+flGOzTVjYcBnFkMCe3N4N2sWv2gpIh8T3GStp9t4ug0HXU9qip2rd8
RlSvcOK8sLxfmGiVpKhzpZQtYRXmAwSrLLNraD+83zXMxhz1iWcdrJG2pMI89q24N1jqfbVsqJhI
o9ZamYDIcO5ZqkTHYrwtv8Lray44wAVMuIeg1cd+oCCey84HPhcbIyDE3vcBXqoPsCtFnXPeIrvV
17gFsdTJl1+7gpj/Tcvma4shveqEb6w+PVEHETXqUvJ36Gy5tgIJH56SPU5HHYjRmsxSKHGNeOPN
BuSITHIJK3K/xl5dSaDsd2NRrNSXeE5RyH6a1ASLsaZauaOTw6i0l9DUBkiygdJMQ3PA79f717Rm
CN/kF+8xf+Zwipq0yUWN1+JTz3AUa3tfMkWDPhZnNhqyxAtTqxzQt601KvOdBZ9ZXZ3TGPaZ5hyo
ZFR+lRyKvpWh+lxrnFY6ea37vE6DZv9y2TQMnlItoca67it9LjgpWVyxPErFP5GWnXCfuH1PUliS
OGTHQOwMYN25VXljjwdkeEW20FejP4qJjKmgxOZnwahVZLhAOAcyMcNx0hty1VyJnD5Mw5MeE3bx
TJyzHLJfzgj+Is5dcysiWD++iX1NEsbP7OA5ZumpTq4YbRJCl24X030p2UTDbstm2wTqFbj1yuGm
GzpIpRwoLmW8e8EQZf3B3QvcUcPL6fgD1q4qJnlqZKsbYsm0RSwtAyGBPD6BilhUIl1haYy7rWzi
lL/tiuaqhiCXVA+77soAR7yE2PmXqnNldFapA2o1Vqi2xobkB9ysTK1v5zSwQ3GtYBZIyOmFf+Pb
ygiYIAVZ1wzxiT+KvpkRyPnpkOgFGNYF366a4Cni790+xfcqtIwtAl0fI2O33YyOT3pALy9PbADE
sBu+fONt82RiSihKL0zDc4A+wvH9GECMX/7petfAMj/H2jhJQJXmAqAYLX9pKD+6zLOaNQ/7EcJt
lzpIW8AOYYxhPqitMbUAi2yetO2bf4jnB0Y+hnSTOKxQSElGDKKrCB7UIHx62AYe+ThBnlsE6/t+
4W1xrNWywVCcoMsJ+llJRuOTfkG7Wn7P9SdlT6DYBHSoqv5b72Vjr6W4uJMNniSzBCXvNFyxKgT9
DFwiYhNSQBRNJhYCjzo3eN7zeK8eMrMb0Woglu/pCrX/zbZDfV8ZTwR3DU32eMoeqKswzR3LxtZn
5Wg2YDDC2lB+mIz++q+UeplG45d/G1TYEJ8IW1lLALcW3n2WB3W98mrOHrgsrGbekWRG5hlvpdNh
cajym0OgPdj9sJRezRhQ4eTEBzkKU7kfrWjXEj72zKhS1sPUBu79EfQBshAq/0Xsv1tgwxkc2KL5
zJahwdG7oVLIqKMgfau3ARpu/kgnTzyY0IDujnFPlfQAnb+/K9hmWVQY6OzZP5UiPm6JLfhSlVdD
GKvg8tEsXFO5zp5QxjPSyrof9AoqZGhU+dbnq+sngUlwa/NA6SAa95IrZNUZrVL7PJZ3sA5Pdhnb
lde7yf0reHyZKOAHzWbicuWKVHpeZBYLp3TySbkEwoRqNgMVDeGUBH3nyWmZKBDqhovIwPMmySIC
7ziGMY7TkFLiozRTAfUISe5BO2XZwkmBCz3sNTliIW7aTDavj3Ff+FCyr1EmNMhmioQIe0GlGNnl
LCUrqMzyiHkPz6r2SgvaGPCbvOhr/ZCoT6IYZkHDliFFXHyYIVrnfGiqmIrwPjrFCIQdD5n/DS2K
GeEH/9HsyRQWVSjzxzPEdNp/H22tT0Bx7LViORUGPMsoulfwCix9TVB14kf7PSOIbynDztxlM+L1
XCaOW2hRmmX0+lI6iw5eUpTtj/HYw8mjx/fFv/whZ9oX1EJoQZUepcXswk2VG2Us5oH51CupgCcv
BbMMkhWQx0TjAIenQG7x5B37mVvzPLJCqvZOLn6ONNtMEMwymKXCOb1V8Cz+lglVGxHzceE4R/3t
KHwKLA5pWNB+BnvPh4bjhy3pb1gQvsZfDnEp3ZN0Gr2lr2Eu3IsvKA86De9SlMwveInk7FYtJDFW
icZJRh9SMo9vt0nNYcfJDDk2/oIi/dWiDduyGJ6yZsJKKUF7THPhl9yYmeEiTKRPG9373u4y++iu
omNJAeFW7XM1IhLk0XgT/cBiAAFXs6StjBOWsUcS6L9xZlGsVjCdsj3FKR2H55BcDU5D3NP4yjWD
J+cfqOEEJO0J1B4So0hZcMhIAKdlLVw6AQQS/Gu6/kvTa6AQ99wDP3wYK1+N4XWAlRB5llrHXo7c
MlJ7UxsqQByjt++HpGJZHfsKrnkhzghLRXT8qCbW9YNSRvqngFcRKvBUg1iFGZKhdaKfNwI6o4Xy
JgZNGrV7GdpFN99VPWc93RT3zheVDvG6g6tdZYw+gJb/fZglE8qv1AoTrog1YoOAaMDvsQ+noF51
A6XoFX0ec6BkjD/Ups1A2SURBUrNF01rrSdgd0t+A54lWe/v6cw7nKENOGok0TfD/5oU4QcQ85m1
vXsxIKZHPpBeZVTS8VQhkqDBUk+bomjQdHQkwJv4G9xMvPW3i8mz0ah9cfNwMAhvTNXnrrUb4owv
S9dtmTG+OvOlwm/yyMUtulkefJs0bVjSbNk0CvceOg/KVQrgkr50gyDAN0Qrbs6dqXImD8BDtQtL
+bQCDbxDLqDa5wRgybrqOFzfrAXzr+1WLbh1vYZ4OLK/3o45a1WgKAW0Qa7igxcO1mJjXW6xOW74
4QkwDvvP6+HPWe2x/tjyFNpPCWVvNA6xWhAGnPuEKgq41mE6nJ+zjR5IeGlJKY6lFWDThhtzsGZS
9DSRKhUctQB+wGbV9jpxah9PDIdbWIMfMbMxorYO3rvlNv9PGj5RFsM/w2eIhJeidXJcR0GuX4ke
dY43VF0iCoxePTXX90fItjRD7SxWLDzdIKHeqgMYVN/BRIC4KcDWYDZrXNtm3Rqx3qJhJjfVxqxk
bjDH44nJjN6pyIRHetSF/CcBwlzksLaZJIMzeElHT38/ulA0OzrrQwrnAeoiU/r2PdOtAhle3B/W
iiAMAYEmmMZ6j7Z2Pom6ZHr77xtZZURy8uMsotJw9bxNON7pGoF59EVMSq8ZmUaP8lZvmAYbEpzh
0tXIvYjVM9pHohUQYBHVoKw4r2eWLppqOWNYsVbiKJnJ9XYSUh+ukB415CI/v3F4nFeXvFRjasxq
t9ZSPpZI+yYU00YjwwGzUZXViffJORNGwT6IcRVcX9cQonTVYeLKRfUeIKhpm/tGLUmENQrMvuqS
nXKb01B487AyOss5A6qfMSc5h5KHnVvJJIfZjEqQmszXxMF0SdN0MfQs/raO/ItpWugLcrnpElcZ
z+WShBecFXt4LZ0m66j7Zn6aJ8X7C+QJXj1hAUlDeiUPTgNPZiPC8ubezYQTEgW0m8ucul+MfK+d
/vEbKtXecMEYUkM6ggC6vScbGDG3LCF4eP56AwbhPL9/NnURihDnAtoQsvU4FvsRyyXgCQHYZ8pa
EASz8Hgc+KXyp059wvOKGrsTAB30HJqNAiWaOIkxZHbCYmqYnJRzWqIJbOV8rlRaO6cTs4xfWBmT
bwXLbNou9ofuIjqgMoTn8cJx2FoEwbHJRW62mb1xDtleI6hdmZ6pYSrxMJ1ny6Tf1yrozcEQQzjW
9KSOzO2PhmNKpfqM4qUKEJ9F5n9HXsMq+mMj9dtklhWHGuTLd/3E3X+mpxG3CtGjaGgECSnGSdDI
HHyY/51e0XU0K2irifdQ8f/8c86Ti/9yMn/dFOFrENVcPtq2Aum8Z780ZQ4Dgtbk3vWnveKFRrJp
j8QN4/o0biQWBMKRJknnHS81RDhPE3iy6clTQ3/zGVYOeyRCFB9unO/8Ik3lQ5nNppzBfH1nMjUD
0Rf/hxxcbcqKczYJ4PsBFk6NqtlocKbB759woUqcF2DDiMvDXPnSeyopXOF+YoAkrfGYIfn0r3XW
/aOL4iba7IJvOrOzKxR7lkBLmmpaECYcoUe2zP4OdgcuRWUzWpbFcOSi4jdkpeGZ9OkLJKvMNTe3
4XrEEUd7UysnrYBah0Q/oMOD22COV+s1cqgc6ZvwnUQyONC8mn5xEPGHhmKaplFv1u9126lnijaN
l30tRE1i/i6gcxhAXYKPc89cooPNUIxhwaBwOER55vmyNf4WFOBgvMLpDPUI8cUWsYm7NRcrTaPo
gFRx4EFWZ77I8tzF66+B92LYMtQwhveQDEOUFIzRIRd9XZCpo0TRWvlQOBOP6LKL4ASkW8ybKfVm
+grzWZA1uEDbuu7C4DH0TZb3uwGuY269v8SKinEG8AyZdsHM8T8JOZUYVNgkyVo4peyYweZJBRGD
DDl08UcmnwesFBx8CwKow/Fn9p9Hp5tPewVxncKSKTlwwU7L/7yjgqSLSvnyu5iQQiAEdNew8oQo
8cRSFfsB6eouEmghCYw4h2NynJKWlv8ppv9wYXOt5M0/hqavoxqd51DIZXJ4IFeaNL0WFshpcjRo
ualNntMrRce8eQ1pfh6mXb4mkr0UuiMw9GXBm3M7FmcJ0lPnmWSJppb4UY/+GifwAOZEcIMdS6Az
8f/MhFopHtNtXduuNiMDcplkW9Bt/j265NP8o7ZFEpIs54/2L8Bex1wFcDbfi3RRqvVMATUNQH0j
FwEO3gqvj5rpTLCZdXAEgDtJgFsZw2uYAW47/xu30Wqh3JQbTvJCKnsZ+zaU8SOEpZod0of89f5u
NsCSEePnnchagKzYBtEoRZqx6G455C0csD+R4YU8eF4/Aqme2zLzhLHbASfgmOiQx9Ye2Z8A74Hv
4/0RKcpwxVIy3gC3Ly3hAljSPBAPB0g+4vQw8NMRxXpjTUaNnxIpfSfPy62csdnbb6i1DU+KT8gh
qfAguX+vescKo7jtCeX3vA38Wljcq/6s5qg4JUy03l0WM50WLH+2/OnkClPCGWb8cR77X9p09owt
ttYR7HfioFP78HetFIQEZMToH1JxYmr+5fb7+/joXxcAlgeot6gP5dv4OdUQsg2UeggX5tzmOA4g
bnFojFnKg350NmBOcnQJ8f991gCFCPYRPRwroQqTqhtoK/nTGgPuOFYXTKjrDEXib/16UXk6ZlE0
XfmaHEgHeSEoCsbFY3IUZXhiQl9VWFyhDLU4ieWlfwyNSAyUIqQU46+8yenfibrFk1ip8oDu3jK7
G8z13w/OFfWWywSFfNYwT9arFN2NBQWJrZTVwHFPKodl6cIHAkqxONyBV97T0outolua52hLPGkK
3oOkMLg3mlT9R2rnWLNKk8gcY2sxTNup5AtnNmoNkKee1zH9jpeQHIMpJn4Pa3672KbQ4CkJ8ZOm
GMkTyz4NsvlYdPVYn3/of/IbMKhlFXDXxZuIzxsqBNWa0HM9eOqR1Ea4TOiI3e99XGTfgGaDVfvC
D3EDCc2jV8qK2Qrvr30giqeeDayYQCywW5znCih4vZmnjV4cXtZpA24ES0cOuaA2yVP6TYfW2yNe
t4KUVFENYveANg+k0eP1PvJiQWTAPokKvVo5hS4/brY10Ay37kVzEapYX0U7chVc1x/IHTbRRXiI
mUwx5QTc/+oXMtTUxVYKeXZWIWEfBfbegHXcrdJHLj0fIGvVAXGKGjUivB+BKyIZ7AcErSkQ1Dui
DcMJJyckUAdx97MNU/Um2eA4J8eubMyAZPrvPwdc8s9wntOpkZuN8rgir9MI8apkVM1omvcJX5Vw
8Diiw84I8R/jFtZoU9wwW0k5cgLJqcDlPUWcATYxlSI/PMXRgFV3lsU7HHXjJzRNzgVrQC60ctjG
nyyh8bO23pFZc9Lb2VHtBcCLb0qodehqr6+fV8AeWTPxUTuciMQs2txCBoensIMPlSRbwM0qr3l/
NTzwNk6sIGqB6TSIE4ieNg4q3/iO1ftm7DfMUzlXMcHkcI+U82Sg9WPiiuW18i2O8NFQrHbYWxPK
yax7m62aFfrgI2H3kncbnjUeNED48OdH6ljLsIj9RvsVQ3iG2lZa9NjizPfIefj0Ojmy3y/LXJWi
4jOf0JboqbM9y7eJq4N6jwaaXBTJcEPvPnPqm4T4AUDGT1wCdgH8/f+Xye0fqA25VDJJ3E+uIBIs
7235pineMXAYSw8aFHhD6mHfXSnyZ67J03xpUPLSCwj3SPlE2iO+b771PvkM5/r1QnOEek2ipL4B
8Ru2QP/smft7c8YLAY9/HzToS2iTOony9E57VkspOLpT4n83dClX8sbiVj6uYyCvWffe1fxxzJsp
/lAHMGsa/m4CbfFPbjuhXJobP1W8w2TmZmwj1RIat4utQKtIW3oCc09S5uR8jFayFitZb9u5JDBN
5+JQPuttVldwA7ZjBzjkcFBzstVR25xw1g4rL0sOWFAIowZ9E+VamyTu9RZ76R1RcvIxfRHsbCJK
V/AVsS/KkFNIsZH1gt//Zc9+lIlEW/8P63KnCOMLLjfiUYXlkFFHgsHOV/yqdyZPXwTf4P2vid5s
AxJjEnAy8oDvFwhQDiorhR0iKdMJqYbq0ohcE4tlyqjJaFDliQCBp94QcMq97aLyLiCT5wxMqlLD
8fwIJXe1ffrcrAbKjLiDKthWkmpHDSjjCa86Knou1W7KiddICPKb4kerdeXAYijrW2KEBZAY9Knq
cLw/yPKNT50+6DZ4daNi4kp6H/79f2U5dI+DB8qNPPwdorpj201jL6RFw80F6Llisnp29du+G8n1
bGJg/1lfD2+FY3uX9I4ifuFwuNr3Wh05sTnN/HfqRUZ2rQa5/mnfqzBGoL7OpSgS3enn+AjaIhbm
f9likQlLHVO8qwScfShTiAWlSaMXaTE+qvpj4qnaHZ6IhbEfkyM8qZrGlx6sugk20LTV8gSqr6qa
MNf20fapQ3ndLpiPvVwTkW1f65bYOezoCAFXDyDQycK/oz/9VYKnemGLYP42pbu7w+hEZiyw539a
/GmUks1cBycuRfUqTfDr/UqN36/a3Yjri5Tbqxox+gM2zgLvvPsqg6ZJRA31SWSx3na2ZyYnJLcT
5KtKCE6SeL4TraxkebbYZtiGcfKmtZwkjVVZyLQzm2/Q4BCG7BDoInkDbfmExATt3xNIp7i5oLUF
nxgSjfnFH+cBKvAubPV9wa5DloL5QEUfnA1EKsCcZZ7EdEeNOjlDqoosTkUW7HnokLROGxOZxwWL
Wvs9pQSlbGqoG//xNxY346NUQVad1sGgtTixFWdpxWsQ3I76UstB1RLMIYtuUieEDaN+gG1ocr85
QKIeBA34H3ZISOx3Ojsno5TRFWH34UT3OC+Ib4cyj3sWR8pe/biVzHCGuBnix/3Rcx1w+6I92mJD
O9k4BGjR++FCbXbxymJGd3xiEGBXeglMr10XID3FdPSs3WmCHkFP0aiGKnWpecyk9yXRVIEdLpIJ
jWUh02eYSPKs3syuW/QPLFTnCSmrdhtIqlkbrMlz5Lx4Z1vXNx29pQGl99jtbH0J1+baLdpKJXJ2
6E2euw31iUpQJEmAGLXOUlJr9R5Xn0b1zMCyLHtiTUYpKcQWonMqsgw7zn5f7Cy0eQAaOfsZRtHk
+jgl/f9pvIS9w8L1kpbsiERKM/Vpxd+s1NwFpA0qRCdYG/OE/5P3Y7amyzHNQ6nvtWFhae2Qdmax
t4eUkbExoZp46cRDecM9HfL95Fw5uhu8sPk9xaqbS/sl7U73lDQ1plfQBolJGeM9rmr5vlZKmOGh
ovW0GkxnansYBzDGq/h+Aj3yw6tsDHvJCN0b8XjZmpfVvRAvSmvw9I1RvApFf3UF/UH6W+ey17jR
vO0PW08W95/oBDbfZv6OHCwIlTu+ctVnF/9xDoRngK1ZZYfrfSDRbtWe2hTMdUmQg68OtDF7iA6R
Z/0ykgU+A/FctSFPBVq5yYuGCtSFUpJwlw6gzT6e4TlhffpBJa05uNPssGhrjYYoWxhTcDN4/9D1
pc/zSz7Eo7jflozXJ+sG9TOKx4dWief/0MJUiliwTX0CDC37I0wU+AElZaZJpo8oWVrGfIbWLrhi
K1ZOgz+GT0nO68s/07aYAMSkfvG1cHNnZTgrkNB9PZVcHg9Li9DrrBkJvD9PnhMoNS6EECZgNmvb
wS+lH87qJneQWr4R5Akq/Q0teTUaGnpWVrcuacebb4+7MVGNn8Kkpi2IbwbD80MtDJaUXTSDOahM
DJdVJRBUVw2FmuKBcxNdyNs0WocG4J4BQgf171iOYWDGcr1tkeRvnbq5psMur13R9UfD0VC5s0fo
FoAO7Rx8e2mRnQFknoM5dSvatO0akNmdnIt3zmd/iRQ8RsCFUl7sDPZvwuQelp8AMsC4UMZftUaQ
q6aL/M1aCgdlWRLuV1V8HhygPLNTBoLf0FjvVLdhzRf0rKIWe8IFgh9io701csYXlYdUyIHAv2L8
VqByy7JGLWDlYaHZ4mvnvranjzrudIE67y8XCztxcXmBeHM4HRv0/j/eacEDt+lWPbgi3cnmFAu/
QWgAWiLBzsdbDBdKqyW/xdYTepqlvPU2iUE6o5Kv5MhCr9Gda2i6roDDU/QOJqDQz8KminG2EEaQ
u5uMWyvNVRVbVCBWUma0HMcsRZRlSiQgpZrC+ghTB8PfnIfMoKCBIuH4b10M4sx5UzJVue4eVSAT
GVyWIOxFkCkHvsWsb88To7e0DFwytUjV6PsgJQwkQGKA79DCaIsYlm2Ec54GBBpjGxinr0G+c5gq
PzsE4lnQNHZcWomffGkErj3y6EOD8dFiFBcpqtOpIIGyUHrCYbZAKAKXQavVq/rOvh07+zeQoI9G
Y1/oZY4DzLmbTYMKELAcK3lQjFiMbJp02hzpLUuYXw/EDJ9fhN7m69DkTOJ2tIYsUEK/DzOIr2wz
5W3Bkncva/cXn17R9B+uFP95v413lTMuCPW+3+zs56kVxzqgScf+NYb/JR24yi0L/6qDK5EUVVsU
DhH4BJNAmk9DsnzDxHVL/gBy0bv8KTlj1H73Jq+Qlo192czI/QqkM7UTJH+jJ4bVsjXn/TB40zQ2
rz7at0nzx7WtMvyjjUiH509cLELjlomQ5UekPj2YgeuzsaS8W2nS1THMWd3qRi2G5zJMosyQlLw2
GNY4707TRpxnddqwj0CyImT32igTNj41bXBSyZxTRdTNxC3ZklCzZ+/eFAnFEijM+UKzKjByyyHi
5t2GEgE6o1zdTaUJsXviLf1Tii4DI3PaOgkNY+k3I5wW1e6nrlakW+djS2ydX3LdAEV0L57LVP5e
bwMqvSE9lWh2v1Ww4grlA+Cdjlvw4zrrjCm9bMRKotkzLTbtkM7qDDGiY1G7u14XvM3D0LUN8qja
Vmn1IQv8JSF77qzcu07Fr0hSjSJ/u91nC3D9VOFeDSxbIKVswjpd+2U+Qx2d2u5Ms1amjrdOqI1L
06dlZFhn4n4nIV/RvI66pDrymLVvhoXRFst48eNlQQ5nfeFzqD8JPWZAB7WYswGf2mkqSieViXkU
0QIHRLcoud93Vc2dehBDZ3BQ8dRL5fSoXP/pghTPuGSUWtEBp1M6Hlft7O9uUm+GxZGd8uFhfIJ0
FzCFyRPCWbSuVZii//NyI4CPhRkuE6KQbVPhzXDC5FvpECedu+bHhqo7TEaXJ2m252q712J8zMiD
WP8TB3v+6Ob/zqIJNdca84qZQ7EeNLeop1oyBECcoa00ua5ujlCdiT+n35W5GkHBI9GADFWkEN5E
2a4tuup5UCGXsmL4/pHuhwAKhsWrt8QJCmcNlUM/O2L0i/TeJ4VATS9yuqg3qE/nDRAvIVWuPNrG
BJv97HGF9Sr5QOfi9eX8aBNRjEelYk5UtWIkmq65Sc68/xF1kMzWVRztZRVwi3SPbwC1Xz6mwIUD
Bx5BYmwlpLG05HRtRFUVFAjYOj1Y/dPXmjNHhUj17p5wBP18HAEw81ae1xdaWpSuKKVtMv6RrkEG
YxfPX4uFQ5dfMT/RhQUg+gBWdzm9vfKzI6y4MofV5wKgtagR1uoszWMF7k4I9KmFHKcmFsG9ws5V
nds9F5x+fse5vEZmVzShy0r/YaZe+P9jBhu9vdAhnY3PZ+C00mhaBiNgbKOCzDJxxqX1Nbz8D74c
YPOf/x9eEh3QcDdluvvzhSiz9LJ7M1xFbixzx+0w3VzWPNVoKJV9V7oaukUPgBCgRLcAjABOf6Ez
uOz3DGe5E9albJ9S7SSaeaJOcnuYx14Zv+zXQLV8AX7crH0iEdyo/4Th5y+khIP8758OEyZpYh7R
sXjpL8qDAkbAtlVk67EIuWjjYbNk9ixmPDw5b3pQH6SVlig+Ui1NruwqCKPrdidt8hHLV3fApzN6
luX6iXTvDIh0utH1imP0uHDJf7c6DYWwMecvOds6unFRjxEV0B5SYUGfNzho1iux1MERprlklbZ2
D/3njHRF19ymhIz3kZX+x+MC5J1gbBrscbhkA6+6thSoBLHHBy685ZoAM8DVd/ejNfMUpZYcqbqp
PQoakJcX7CtAKPs/lQnTRpaWiLHeRWtjvuZj+2iR/ATLxZMRzaM1YYjjA7CYC7ZCLgvYLZvU3tYd
Y3XxK8IefS3n0hAKt5RNDvltQcRoHYQu1fpKX99f43yNmeLPDAMJpknytkjBY3q5F4jhCP2/z1jd
ViYdwVj4g2g4iuAOCHfosxp2olXqI+kdcCc1Jpoa9E5jo512sZiJcG2atKFz5R+6Ww/pMxz73aay
VeXRApyNsne/zIbx4X22ZHITZtHgYQKssXccxg+X8T/mFOlvC4OSfpDPdWflPpHvgt5tbi2uLVSP
sZDP5SDR8ciTzG4Gl/1zWBn9ZhYVfgw7zUB+ZaheF7XhWK04Cb+BswztiX7w0Dj4ioKKsAEaIiNJ
Jx+Z4K3UtEYn6AL13riq7R9kABlchGanvYxYRxN/T+kdyY6KFtMew6BIfpmqD4BkEPABlW+uH5aB
QYUHXVrg3r1yruqdaVn0ZNPuGyz+rsBiDxB4U+mPbT7o3++Cc+xH4SePn+/KkTDtgCZTi9XGvoKR
vADTm5jxj/owlTIQ4bjmMsqcnV93g0r0ZN0XpFLz8azagIJCQyB4ECdc/AHPkDMA0j+H+x9QlcDk
P3nphbCjM9VcNsSNP0JIF+9HE37dcHiuUvlWVX+SSZvyvfFXvYwZUMwlXZPNlMHQeJoM2/BjTTv8
7hcke8BonJjXjjGD/7HWLuu28kivqT/7nCMHYzn2REmro6Y6bnNCsQMF3AA86SYzT+9k/qml+zu9
Rn+5tuT83971WRE+gZth3WCX3HXe5rspKKgNYKGfphOx1Vjvdv+A4aN2x5xFzwZTOv7Mr8xyYJY6
jJNR2HZ4Tl7wxqtQU5rvKpH0Eo36r9zj2RjdAbyF5+cLE+wcGYcsobEdAsBG+o5u9V0DEPnUOGDs
0OdganUEVmNBo8Ej6i/e3NvN1tuox8LQEg+Bhqf0uMq5li5/odkl+3EM0/fYQIpQ0Zfq94nP8jKb
7V8xuFtHQan1IlMFWC+nXc9ulhxUCHELTVkX6rvxToIYmYvRLYmBc7E/qzPd+q10pc7/7/JbgEYF
j7pq0p0NJyqULiY43RwhRqk69ncdJy+dLi6n8G5JH+0l0EAaGaBNE/UGdh5CQ/Dvoi5tf4uJGIhs
8EZJ2zS4rM6Oa+3Lu1fSGE+uJIVpcEeeM+UE09qcnEkwwMod5QOBco3JntrjnPcv+ItO6I9e8i8l
0dgHVmP1Ul8ZAKuYv6Qd1p657oIbIrO45hSR2CilfUU2Y33YvaFM6uLIQoiEe+ZKSZEthQVMaT+m
fXV+MNcetlXKkefDhLe/2CLCwmyz+Wl7O6DoLhA39mpuCER3iJs7w7ArMD7PpYkwxFrAoapzw81v
vYyZmmCzLy2M3eNQg3bZEATwhbw2mkaDj/qkf59wBLc8DdiKkf/9BMkHRA/K/rfC+hY10C0OrH07
G7XUiA6ueUhkzDdwNFiv3BgOjw1X+k7K1ibG7+MLVhln4+bFO8nG0eK+YgUwn+ge1N6wsNcvlwSo
RwZ5hBAC3uHz1J0R0dVUjT7wRZf94yaH3jzw74yTD4UgoMtZNtxIPyzzMs06dGk1mbRf35xNbJaX
hiQKiZF0He7+K9nTxOHEVF3RXInE2fRPvrRoWVIXJTLgO7Iow0Yh79yU6yU58QRo2rn+XHR/huUy
wVmcqqTPRtQMaj7lrRew8sJtxqEn2CAiWbnCx92LBJy5QzXOa3y6cVquHmXfIWCwxxOCk/mDxdd5
V8QwqhDnQyW1KbNk1jn9Tb646WN1/xTfuUJDke/rCspZcs8QFF+pnQvMkTLLxyFWO8fH6CwSY8Ox
0l9RVPVQ9CwGwnBpvdPzW8a/Asq5guJXJtNwdQIEV7ISdTOEUpppZ1RAR1/MR1J6g2EOq3WlJIqh
MyiGpRUgWRJyc43Z2RVAbZjdGVtx9iBU3U6KXrtG5shKMaIQuZkTPvMHIeqOnH9OalVwIgt4nQeg
FRg9fITBz8gHG9771U1sxxGg7EBrJaHKCZQ9E0e3QHVxiif+ZryNdFRLd2ya4MoxEJGelcLzU7Ne
xVnmj8eeedZpe+BpI0qyy3ejVXM0+E3KvgaeExbDgGRAPWAWxxCCk+o7MjEa8BSQlCNIC0iZZHYy
u8R5tOl2NTMJZko59EHxM8L+HezXrsxy5NIXXPvSXUiENHqNGXHuTOV+IktHuEITQFhH46DVYS6O
qocNScP/NcnTHOWOkUJ3evI0ggeVa6Yis+4FBC6bz7nuGZZRbMg0gALKZt/KyRU3SDSbYefmbhfv
wmzLwVK4RuJJpe8dmBY8PU3pb/9y6IEHo8+zVq8fjIs5vCPnBHI5PBBuxTI0ykDYValyBit4NfFQ
ab1F9JQV05SE/EG/7Ct2Tfb7jFrakNxz2toE/VvlZnGoX4x8q1MF2/CWsXWk8Za/FfAFWS5kjge9
0ExbjTzb8a1kY1PhmA9oqm/J4DMRk5h3kEUKO8EchLpG5nafXKoiNYw/gvAqudI1KDwuTpUkk5ve
1gUuz7lb90N3mGMPXZNrYGK87gFpsjNDEKBc7sXETFf9O+eVXk2ETCFe6ZgO9y8WuOLUvBueVIhh
Fk/2JS5GPwgW/m5YkBPWr9sOH0wf9by3+rv56gyyHq1evaOM6itYexaTsGpwK1R+bTBhMroaCB/3
Ich0ys/b0HnvoO/nW07Iac2Enf3qhBHuSDuiQtYVATx8ypTSkD8EkkIoULl7Fan6e21s4/tTatzz
7hN0Ta5O1BnhCNo4tY4gwFubKKx0HH3IuIaiymnkbmnlZwUG0JJC1wSc63N6EWIWdFy3XtVZtp0b
RRHhlw/n90zA7Z83Q7idZTp4wFcDQLnRvpTrDdZJBohCRQ55fZeSRiUn+Te3Z5E2OdC/5qKT/5IT
kuLq5mpH+X7YqOrGiydram9ErE4v0mRNLLHOGNjqIttlbH84kqpKuBUA/CDHUVrYLyXUeXvaei1q
8wBqZZvFKX2ecvafp9wqEMzMsz0yx4MwahnzL7vPrnVoBEN56piYvQHjHLJbwoyialAzHFl3PbHB
vvYseSA1hBD/ZBixR3oh7ktgTVciV14YNKHcjpVZRjAd0C8pobvOcq/4C+zEOhFa52eQomOzyDnA
8suFn4x1GFFkR0qgiq7Vf2Jhq0NNrU2cWNMR+6GDZgvOu2/1qAgxz8KUUodz1v2EzzYog/rkXZVO
dR2nmAD/x+2snQru0kdW95PbTf/bkQ2IABy1njSHGCh1gSdlgTpzOffpOa7f8Jx7KLOT8ZQ9Nb8N
RFdBP9WT+OSzA3JQskdXJqhonPtgZiMtefy6Xyd9ePOan8UqiaGUezTxf1a08Iv/Yw6XmPzYECrR
wYOk/hdXr7XxOHKgY0m4mkBba0w/yy7H8h+ikMfoa9tgDw7ZmFC8HIkicyr70SPp9Wjr2wULmx/k
e/4cT/QHBL54nPyhym0dSZAOLgw2lKgWxyHOgPPlc0BgouIR1TmZ11rKRAnl80l9InPJtSQRMZrE
YbFfwnOoafGTz5jDmXDLvR+6au9GhBeOaLwHEM8yRn5FbPMttHd9pKA6t7aCaLX4r75l2KoBmkCF
9Pgf8DBYCZkWF/BpFec1K1FO1WuFP/nUKOdeQVoBSCZ2dNPe31S8NQxcayYLg/aGKtPQTGLjx6Ls
hBo3uOm17JeHLp7IuhUGO7e1kCYM0G2rW2b9+iU6YmjjgzxwgNSg3bEimi9fcFC3N4f8U4uUiCdc
X2FF2crWOPyO1VHqHdLz7HmDIoKsH1cfKJsR0xtmN51CCy4vsGlhEnK41ejBUNIqRLm3cMGGk+H7
Hiqpqi71AvJS5saBnaLT9l+XnUOVji8fstw8VJOX0rCe+lo7pVCZgCPaxHNmqIVSEvfGr6/scBoj
afkM7gZVtY7Fn9aCOCOrv/iXvWmf8gHnaMcw+0hCZj1d44MyKZoHkxa3/Uknl2StibP377GAO22L
xecETEaVPv72TiF1tcYTgMtpKzD4dDLs/EjKKx2VV0HeiET9/j9fPz70le+oQTGEWeOIbxvdSd7I
9t38O+BmR1hyo2B1S/cvg1iPWtSbhqAQSDN6KvuvJndKKc6yTuqRT3DgW4vM0jBnPCF40jhBbEEL
T+bIgKLvL+vGfjUgXfVOqIO4FZiKhoexkTzzBbS4NMBX04cpjWtO+LDTi8dZIHxh5SKgO3dDnRmN
aAIrsGzuQMGJkj6fkiuvT4q7PjsQRie85OGebQaeBoz1eBQ7coTaFSNwamxlflR+tNi8PGmJBypg
r0Aw21dalVaDOZsUIz7/11p0cwfZibikVWT1zEzLrpFbSpnrZeFhFOkgO9b9EAk/kE0CJqojCdS9
iJ/bsNehwFOpE2wKQvBcK6t+ILkFtLVLTGZ/uh9IREVMzYbD6qqVatKbwtsB1p8aIhKvmt/je1CJ
AuT5KZcEvX/3HYGsrbEYHzmDUrnZQaUDaT+jeloZrZdTfMomikuaENkwgujOUYzofe2OEh/v6b5F
iargJLBfPq+CXGoDqvklHt407/HnHQyuuvIB2BlO9hiH+9wo0UGLz+lK3AGZtdS9HCI46LTnewJL
qrPq0mUspupZaW61Qt55NU53u7LV1aep/cj0TJHLEEMyScms5mS39h6F6csiYjKlh1xCdCXgjgrP
1MHLJyLvoOLdJFqiN00ojQDstJozit3oWvxox6Oar6JD4ByxyVyGt+efSTtK6ejET5caaYv7HoiM
ID5ICzfENZeHLoOThai8NOMsPz5AztHFRlMAMYvxaDZlsR4vt7MJYLO2YDv4b87Wr+UWvBNcIjlu
d+2OCzcNz8KquU7DmRQrKsjN/DxPLQvjK5Rbs6XiCMMJF1++qwYH8iaMnfSIvzEuONjg/R+NPFK4
a/6dM5CB3mInlgKfNlclBqYVKlAORIVi3HDtp0ailyfeCs02+IvFaAmYOqftOjYYDuT3HIEItoV8
Ef+kQ/Fi+pWemYMN340P/AUfQGmeHZfHHU0/ebSor7DlOyITkLu2NzFdx987AkSMPL/GRGiJhX8F
Lz7Rc9VGn/Fm6Kyl5OanOq5uHJGJwd9B/6nXJPDhmrmQaXMGyj6+0Jfbli496xqdd5ewhVmiRiUN
9TdP3sEudVfVF4udqYu41jkKWZRTEdT6gUbDKheAxJ4wrk03phza8rMvkfK67u0lxopx3MqR0XBp
c5vRKb6XQDout7nkXMXhDB2my9drdMWv9IbM4zfosy27THnYuA1zMWS6ie6yO3qzyUnbsgzaaEHO
lbjlvnSynCsg1S10ExawHY6PWif+obo3aL2Ke5HPFwFLY6eeZjnA0q+q8Ss7XraG5rqCTa1Eyl1W
V01/6I3WG3lvPaiD0iIoBY/0ZauNJK2rXfMJhnem47acnbOYau6lMoIhjB2nDY899H2G6y+Jo8Iq
icNgdySmiLpqubrWP+zvYQVbjlIhdxY6rOFjdgwx9htR0/u24Nkw2585+6+JYlIrNWvxNRjZGBP9
9gXl6LhqSINOPZRn2iadAvm0N40knPfFksQXwAYadnwohsrPa1rsmLaTP710KAXSiiKu3k0y/Rdu
tbVlcsPfVxKk2r2LkxJb9dmPK2tKLuanGQJgFLKacTnk2OkH9eWBCJVQlKubI+IDDO9oMOvYGDv3
V/TzDogNEqSslypKOXUzcsPyy/4VC6ujIE+2MrJdSdkGGFckvBAj51pbqjikatcWxzJv3fxU6Qzs
9jYBMBM0ShVzas0uf65bebvBE1ydg5qDX6ZsaXaDTL7jSs2qxy7e6b5vFlpdIn1dCwP5MRy4YDFG
j/NdINWRgK+Ac0pd9yvvOqQhalm40QgF4itz3LwJoXsoD/btPgE1qGiak6x02eiuu+tC6cwetZZa
/5+1ElZWflTsVVsvIMuW8QZC+pOw564qLGKLD5lNFh6RUYipfZOea4OI91gcdqKFaDIu+sz3TXVP
RgPAiU/nWAWGa7z86aryXEdzPIQVsVZhLXi2zMwxVXh3JQy0z4U77mI3pZDvtTirhKj2JYnBiTYZ
amxGYhRSwy4LFCWx07SrG/92NptgHVrkCx7CUm+9Vz+4Y4rX6ROluZpNZUyiqXvE77w9zKNgjRJ6
BQeF7PRRUkVWJ+WrekhXROAd8wQSn7WTicFsejSdKljUb/vFmTrvG/ThEw7Bd2KG+K80LFjIMhE8
5yTCtWGamMWDPySPspCT9Zts3jdFFkClJ88jxEtHH1JKpUtPfBAniM5/F/bJV+zBW9BEBFuHo+/1
t1jiSdsIL3dLUcye8GoAnzR69B/y1FerxaWA38RYz07fIFwrgXuFiDlMNo7T5vmqEM9uVYoyLNJU
x1c6gA6Hguc28rJ2s+PjfLVTzP6pmR+DKSEbRZXUbtY5YaMjLeDjU+cJPqMqWiTs2U+2ZANfRxME
87yJkzv7kB1YPKyqdf0k/z3xy6d4kkq0GyhyJUT5Q6SsitxXYHFQu6KL0bF+xoVIPr/niTTG4p0W
01STq6G2JkYqtOdjgDNWQGk1HToWlOfWnsJsTwkShzXU/toQOMjaY8eeMSkQSmVOpP/TmybXG3gD
FL9uKkLi+yHoeOjVFiqxaXS1xb7IE9sou/rRyqbec/Hx8Yj1AQQC2YepObt+4546xGP+3/kHY4OH
2ozaV556eICUAqa/KsWnXDQDMte94aE5MUHc8mB2VT1n+eD05/XfWq9AhbW9QlW9zY8HDqZRRevz
JRu4U/Kpj64RwXEUili2NuvCQmFA/ZcfOaSxHJEoawBanL5ba3NYXPkJ8d36es56gmAzCwI8sPlJ
+Fo/gadiXdxfBFuZSs9jb3E4KDivdeNoNaAg8z/ZHKxByVQ0uhY3xujSk5vzJW/aGbcyZevHpv8x
VgOG2djseBVfJZ7crvPOdxRkt/hoizoIv25XLteYDa1zKdEzd1TACfgpEwTuRCQ7lm+f8HHRt0Ig
HLo6EvyVzyjC6eOZRxIDi1eHIKsbIOahokmhlbwULp8lGMp/y2sYGu9eAX2kG4sSNxmg5JgaSLJz
vanHUAW/qfbojBzPDVdECGbDgoCETVj2IvicZeh+540rqJzDvhArCAcgF+CsFKbrp0jIh0hOKL2S
pPCqR+ud9i33KSwVIP9MtczHgC1KKJ2BhMGsGPJ8ECOrIXRrs8c2Z3zEPYUyWegeSUsdQOhAhoh3
2i36jDgGnpx8wOj/d8flRF1xokZbwWkydU+8Dg/wAP8tTUSoApVtZrZeRTEs3UX2GbWHT2RdGmwn
7iUVjdIxznuQj73jyyCpbTh1Q9++wrWjkaxxNCLnRlbxaUXQMjmu1VplnMIi1IQtTk+8FJVJEpRN
FmwDZ2K9bCBVm+pfMAvZu3VCbe1uEvkA4aLcTYB6JnacKo4u/Nw8kRayv0wiLu52q+wZtAso/58C
ZAzbbkiOZIyd9IQmMFoBUacuIfpxU7pWWXSV8ECh4wSyWZovf0DpXtIKO0tL/upupq0IgtkUVRQi
wPM3FrzdQ+nj8uTlP+S1Ea2Cnjj0Rg/N/29kh7Mwmd4oY/PLtfSN9kSyq9VRDZMmhd3vLPwTDPm/
jCU1LiUojXBGDNXJchd41WayNSGSH8SEV9prO94BMWFqWpk5ZoRHCSKgySiMEStYDfb9taz0LVky
YVeiTDff6SrNZwihoBcwKxAIOckMUSkeVZodbvf6e4YPfEY2MOBjHrBI+4w+pqbg9NEWmPRCkUW6
EypIXt8YQkXvEKHBrHKkFbhpas4tIOJJsHJ+a21fN6pZmhlsLfkEZl8VceL9i3+uxzs+IRSjyKRb
xUR2zv/p1SzEB8twwJF0KijuWAqZF6LI++HDGtPqRT/p6uGv7TwOZL2E5V53R6czKEACpYxmoXE0
2yNsACUu7nRRsI1oKwxsIwGSn42wrX+stjc/tNUhYHdzZsrTOoEAETmtQ3wjSEns+ax31UVtPWyj
Pvnq9191LoDqFe7ej6Q/yragDxV/7peClvbZTgX2CSCw+AUrxF0I7LKMscHjP1C/7LCxKN15DOES
LjlKD6+1fn8iOZmEo4TYhlf7wHLkha9E6LL1B0yLzdm9XMmJsT7Aeza/McTZx899VQtG2akFxBKd
E/jvDDOxtDl809WSf2P1Mh01pgBR9/QL2JWwPcZjOCndY4+JDdbwtcBKhDOK5Xcj1MAJw9Iqa1rW
fTPPxnFJWKkG+qOwyu2tCFSDligpDxFUY8rnl7g1u00BKwkg2O9pjHozeK92MsSc/sQxi20J8NBY
kWHxelKlcEzd/2BDurq35Txx2IjUGx5vqCYaOiXAhc/G/brb6yx9W4FP2lb3uqkJIZb/Jq8iJlAv
NEfgib4gG0H58Ow6skySmyIHyP8JRMGz6zNfFQZKu+2Z+GviP455l9nj9BQ+KTLZWb9G6coAcBjX
fZ4tmi5U2nmdAdyuWryGMsNiAmCN2KKFthf3h3bbyu0lAPkZSgN7p2O8Iml78biYZC7yyOzqsMui
pGA3AT1RupYf9pjxTeoOTe5mvQQ/TqLKd7SkNRIadwN7VETmaF1QciEvmJt9M2eWRfFr+MyNUJ0l
NBcMVNb9I7Qjmf8t+BpCPVcl1keDeNN/6ZtsBYjI5FlX9hbDTBklW3VMUBOqr+o9oYHIn4A3Jvrp
XRcGSCVsxKJUC49NlhUnRx75p9rZbfSCYEcM6JiKB5htN8hc7inT6wzXFKi0REOuksNSD1cBh7hz
+KkXHzWb1ZcwFsiSbFXNkXiL2pKo6Xi0DNYEKzXB9HY91TAuF3YFhZVdtVJ1+mCJ1nYehgvU7dyq
91EkYQLuZecQBC2d4dglC6dVJH3zqj88rmmNRJqou6x4Cs4QAi5Ep1qHIyP7QhjX64k/jYchn+RD
WH4Ou1gkDO42Znu3GDoD6tBw/DyPFtN8J20fZM08LJNO3bl1BoZs/mZrTMoGPcZ1mwGV0W+FGHG9
ZZHSCWltqclvfeL3ypCs4I5YnLH3CuecNa3tQR45MDgM5iwbvQzC3lQyslaOwqQNJfYPK/+9crzT
UjoZ0ZLTTvW4Ovbe9sDkVFoJD/Nf+YCHkqHZLRcuCxPUW5n24stxmLmnn2gRqmnRCqgD872WEepP
YNRADrOZSCBAOKLO8A5JgW5YQQYyGAG/8P/Tq/VYdi7r93rGvEi1lE1XEXOlPHX5PPfqhv9aFKRY
6iGjaVfPDRN/SBwltUZ3FOtF3O3xnUAmyhFLwfAJqP63tJ8sUCVBtxGa/Mh9Qy1Y4OdoGQnJNVuV
/vvvy1cITLrfvH1JjQxqvJsd05rW6/WVVn4seRx3MYh2Z9emUtaMhkhqBilyWeQrLnjDF4wDRbSM
eyHr+9dJclJ5fExFVwvR7sgEzZ4yKHiO1+6GALFlfN/E6H7F6DhfGGrWK/0AOqSEmGNOe+ghfejh
Pi6/PzXdJQhsYYe1eyyJEalFoMqeGelLNeDmNyhbPk4LPHN6GuhipooQfvEvKhBJpdRNDR6x8F0M
6VU9l8qpNW8cQj+Ua+ZO1sJ1W2/QV7M7VWUw3rDszCycPOeUt2LKtGuI5iXGLZWypfR+rnzpw34k
r6b6iqVuXTB9FH/CES0zkwe16pLI2xBTXL/ogY4C/a2/Sx06Bm8gi0EZ/0dkUKvCFtsaskKBHLgt
hcK/YxEoVBK7U6N5C59P6E7REe+CyUFaibShQvtodCr+cjKzcLnxaFNq/mx3heGKVf1wBBoCLPPc
1YRVpZ0mfs0qIxY5xN6B+ySdw+hGqUf9ikAerYP7JtOPITDwu7NyZN/DYBgE2etLaCiYAE6ZRp4T
QRuFV+AxK3i3EJ01yHbVGtG3cih8J6x1+depsm5/+5/Hxy3YQNY/ecDPxPQTDQchvaEiDtd2VhVX
J7GRDqDnCZO08CXSMrzLm9tZ82joTvsLavdzDxUZL6GTHoFrwHNAEAtE239nmgXLVETwsjaWjiNM
xBl72BppouZzYHNJ8YEa37dFPb8pGl/J/F5Zw7lTeAyfxr5hBfnHnGbY3kf0G0sZuIlT+8A8FJ/L
R5TpQ2H44p52/gP6oL4Eo6lz4rt/bTMZQPBnxYHOxYsErTouXdvCsQnOOIG3OeVKYxhXsLFdDkCJ
PLkjzq7SerR+6oSAsRRjxtHyamahg6wf1Wd0y9bN8Qe0TxeP43HTVqKFwj6nGhXej8I30PV1Rsno
yQsb+dw6a3guYaHKp3TJeqWDBerT3yYdZglhfRUruZ3GR+poh4Fownj1MJ6Bwj+Epry25XWtsCTv
6mWCmoXTpDNEgqYwT0XNhg1Leebh2C7CGL6SKLJ8RCOy5vcZtFZnqTFOa0JVsUXbmrh5udNRfTRP
w0B0yJ/J/I441hI2HPAPDapmTcZBn3avKwrgr+Skn+8QvkMuJmDztQ5m5NZvKxDu5ibiNFmtLvIU
fzkowqpju2bm9ZXk6vlpn2d3NrOIh+GSAu3DiHWJEZAmAauNPY6sYNP2Wzq83vfyaJY5prszZg6u
MB7vIF/gh04I3FsoxunHf+EdhSLqupdipqiOBDwldFCeDtRsRj/sVmfGBeRjxSpSGRxPVnQdYaP2
uhpOrh2vLzPHZ0m3ygI3Z4mQg/SMJTyI1hawYscwKrMIEkP068h31x9hZI7X42ke8+Gupwbjboc/
Y8thhN+eDJYvkVRgWDa2dCnHyiv54yu7DImdnMuull6Tc11FuSZu3/uptpkpGqB1sqOxE7ZZmyIo
FMhOZiUSRUZ38VtZ1K1D/ZM2xiuXxRaxxhhJ60WtNqwnvguBwrGSh0eyKjNXUx4I1YDcxXzRfKeg
dAlE01hGM8EusOd7nzqRd1wMOw90k9jMLTr4Ry5Hu3M4mW7KM75K0rFj1cxgCWo/Xgy3fVxjRbdv
SQq+bQb191kEWdLS5hQvP8vX5cGB2ibpB93Zz1gPMi1zO0zu2k4SXwtCE8/8v/7X/8RFy4fEY9ep
dn10sSv6h4xiJQtpR9YzosOW1wZnmv+3ln+FrRpfCzqU4Bn4r3/MgshK/3no87m5BxvCu+tq5HYp
qz0Tg4ZAdHxFKZaJAWOqwpib+WAqIuMARxHi7OefBWxNm6RygqX0vA3frb6rPEDqyU1l871asJpR
6/5Q9w7RJZ5OcpBIDF/CZXEjPS2ut2Mvnf6+zykwgOW4OVsVKxR6acGg5WNLI8Lp/1w798+2gRYd
nBLPXzGfKRlgYFLQNyVEjj8V0Prv9mg16fGOyB5vVSTRI9/5VP9D6z3M7nUJnNyGKD/afisf+Kjy
qM35zCO1eS0vlbYzVNU4UrsBAr/tn+dZ02DeDIbHsb7o7B+zGuqK4wuOtrNIkFEtAxGbZaPapJC6
cDWEmppgzDjtWeHcz0uOnoxwL9sMNhmrV4q/uCBx1VMhKrljMgYD/UwUphIZ17EVjmjn6NKSlWyV
fvLqhW4mCZ2itJQwTCFem3Fx4gVw2prRqla0ptLSZLKrBtGir+bo3I13kaCPWUNYKopvsRUxvin9
ek8E1DKP1PMyXXunddxgbRyO4NGB54xqyN99xJjGkldfxukpAQ644NuMWDsKCiXSNsZrjqeUIMo9
f5TcXCKgj709esgGp30OmBMVibdKWC7ZbisX5n+smBD032iywSf7tGqMFiAHqbXnrq27ctuWFwtl
dUmULDd9GHDvT27VJnuqYeovDkKCQprQDqN+L/OMt7/SirGthxhzdergtwuNdqn2pLiz6sLLSjP5
mVTgMEAoxES+4NH6CxlJM3YFumqMd1du4zTs3ka54V19Tm36COZOpF1pLsCZu0qQwq65PdXHuZcI
Y3iz3ISdZ+b/pV/52uCbeWA9Oz+dpm9175E6jQmNXhxNybDj/xJiuOWlZMFlQjIxT26+PdaFnOu+
42xuPqzqYVFtBvkXxe/qtndgh09VPCW4ui3dObqHVXpY0wy2TOfB1jgoqKzGxtWNHZ7xnUPejgOJ
+S1PwCr3FjxWpuSZQlsomAqnrKrPAq4/Ap6Oh+Z+AVGaXgPDgKtbioxSMc2igFqKNqhEObt7I1WA
sYKvcf1Aq/xLHlCsAnc4SIt2zW8BeNwAIeWTvK2YE2rmx3LkuBvnlYpTmWVfaXxnp7Q/MIysMWia
4cpQKN3D5nU+KIeoHcaz6KeEkDBTTLLrTr4/qkvY56B9vTRxtcVPW2Q0Lv7jeMFJtxZiPlrOO4o7
aLfIGooNknNca+soGzxAf1riaoIjBzNTUtUMsHE5HqL7BbB8kDfy71jkoLeVF54U68JxlMo7NbMC
NeZNTEVmh+tklbd4QiNvZ6GsACITZpr9FNYwtD9J2ovyEN6Rm4XkmmF8JfNGupmUdsgd8abqFDPF
J5iw1DsM7+fcMgrrw6GGNZCWeeAi9XHxGqywxgKgZpzKmR5QV4IoVxuLWUKyPrN0kgqLLi4vEucT
rPSVxg+ThgW1YmM9H0QlAQ06ovQw0IgmLZbr7SJPTEzHDSy5dNit5zjZiCc2R4b7Tbj6vKw3cWRD
NcK7/xITp6kcVqRCkk8qgudBtDSwUIIPOaM/m4Ol8lnavlvwEHWXwqXBJS1uWPvcLMhmfKximyBt
2/I2m744YGrHb9+FJtsywPxvtr1j6VmNq6MreB9CBNCyIfqP6qO7XQQW2SdeGdZnhMYjw7G9jc+3
9VE8cZW4ksZQoSDr2ptsa9d7id7BJdJa/fiRE0q2Ktkhnj8r341zY3XLvrb+XqFPVdB6g+Uj9tH5
KgRGHrrwk+XEhKq6KLtrju3dnUJasxDRN0Gz8MA+rAU+y70CdCX2PVwEKWj2Ug64BYpWGBX6sC3s
5Ce7j2+dVWq3ft7DwUmRb3wtfSte5HJxP9TcqnX9jU9bid0Tfg11TwX3zM8mZBA+bRH6Mi6Ezt+p
exsTFKFoHjmZ4TIlSRoxugwbiKa7A3fkpxDrPTDsDLahNcQKhS8cdn+mtSSUiS76zbFUcE1Rh3+w
/l1oXQHsQ6HVKlxVeYidpSkqS6jBY42Md3CZV/eM2W5B3ILLnWc4NVx51wTB+mokqJFx3xQ7jWCa
DhRbj+zqhyd/M44xNd6OKwXTWfLwcVBSOXtyDuHUAKztRsA+E5VHfJZAMx1elXaKhHzuSQdFbcqC
Z+BESnHhisSG+S8RCKH29cyU+W8emIbYvJK9q8tQQj8wml/fSl09w2+lFshFC+cImFjr1jdxJ9b2
SSk5XYKuzd6e47jOxWNy2YyOQd0U+Qq1zpLxRS+1cOaxuuSpkpQwCFiIr30LWeOyY5IX/rdhMHaq
KOHs29tB2Gtb1ZSyagYofRiQVATE1QiAfMNZh+1m58ja+OKoGYw7XhVd0PXzRqI1rnQ8VVJ/e90I
V/A2HcQn32/6wsGOxDrzoiPhBML4roAmOqbgRUcmVqxCOuCCU1GxJfso2/xt0Zf086Os1DXjsqtR
WU6j0/fw+ngchbR1hnVJC7vUo9+VTBjImoMTRPybQjBNCZoExKRK6r9/6SYyi4ST0HojPb36/V0f
dTCLlFNBjiJK6pA/s+FdpVcfc9L7iCiPk8N122l4X9D74LICIQtdJLHVvZsXFvPlcBsG+J+Jw5hP
Zd4CeMk/1kvqe9q+4h68+FCexSnvvUGiLkY7z3spKxYZBvFuxc1xCPEMRvBLqaoz/HbmKOWfYjDe
Mq2SHajOUelMqdUbDL7GpgR6VT2sSOgsE7nKPIBg70GXovpzwidRVwLIoJf+zlS1MBtkviVvEukM
UizxeNW6+zuUSvPRF/qNwNNyJfx0jjNx0HIvaE05PTjY15RuFQmpegn11B7tJwR/2ukSvKmUcWtK
QzOLV0QekQP57JB/uHkbM/q/IYCi39XCNm8Q2F54MQaGH0M8439O1CX1NHiWkvlSDoG99E7vOlUy
0BiRs/PRAqxOQi9gnefFDTcmB5dGk4ozB9+RZUX4w7c5ceCsd/7vApNkbS5qBbz7sfH9VO7fAFHK
hCHczN5MuleHRJZWBSZrDJFCd/tDCzIfC/YW+ivhT0bKFUJ6kpL7WSPIfhTVyANi9+Z/v/uhF4sd
KZzTs7mZBl/mWm1zEjJLTmmGWIw7AP5P2ht8pFH5S5iMjDb7RajV/KrhOoIo65Lx2yjSiM8UotOb
FE1+USoybmeoJ1GX8SjqhBt4q8FQkyIRYpFsCbrvh9wV7ze6DZYw2k8NcXlCTB5TWW+hjehRaAYW
roYFsx/PBP9tgGEW89U/v9+E7dxfJX0bkXV4IdI4EbqQ66xoPf+ihjPGqRlXAIs3x0ZZKz6Yw9BB
F+7svfCwTe8LVhovV2aVLzw6wzoPMLhih0lGvXSAZeWr2B/n9t3vKrecG4KbNoCfcUlGYAyXqqWz
fyrqM7kivCQ1i3OAArCDmnYiI1sEnkYI3hRLmXStSq5yDYPzsVAerQpIjsG4oLVUf6TQEqaGtIF9
ZZ+Lg1n+jQ2nUHnu1K3Zo0aLx/RROCkaF2r56UCuhlPucSl+cbNDBtYcaoQybMfVNftZJ7ZU3Nut
8od+SglUtnMq4rYAY5pwOklvCCpKBL+iZhVzbRflyTqC9QmV7xc3Q8zbSVN1bErOi49tX42vmhk/
xEkxEj5lmXjs7OmGsHnj52sI4liAHNfCedED1F29DmpcHTiotcXYvdtIE09Naz3SkhZqivsZyem1
r1BQNGJT5NFWFmtU0fiRQsuVmsPtDS91iLX4wwvVsOVlUjBhyw1brB9ymBBIRjnGl0ZgqpIWP3Zt
BNgktxahP0d7KhhVT+aLRpqYxe79l9aPHS8MGGpi8t4JjkWeJBNeO3Asly4DxZfPjsqXEdAogxB9
5iCrJuPF2XIfBE+8F/qVobOZjaaabGm+n09KClzAvmAzznLm2NsdeE+wCcL7kq8+Q4oSpqUZ9EkI
62jvC+oRoQ3AGdW2QUtoGxarkzcjhEJjVNUNaWgiGll7oSbgDI3x7W0+hPXFgNgO93jTvPhc+0kU
DqSZKzl64b2SXN41s3AFGH6tp4owMlsJCeHQygD3rH4vgpnH6gcPqNkV9ZLX4i5SyGytA0wnUE7x
WypCCx2uJbj567eyTiQBxMytYoTx1yFHEjVn34oPH1NCVm2Lzow7fjY27aQNiGYpAz5kjt7rbSgn
2dpSTk38DSbXDt9+U/+MT1rlknGxilKRS75la3TF4gm4L5F/sV1v3mCm3xgq2K4Ced5YXbw+PBSC
qmW+5iotj4SVvsECxZ5sw/BV1LXp26fiek6NhuuaQqPx4xF0ACHRx89dSKZbQ59QooeT0trdiHIR
rLiZzynfycaJTYN2wxz/40n+b3tQ2qGhwdCLHwPiCfiuvaC7HovXkw+AXpIbI/UrWbJ7xkWSZLZ9
mUOjjZHOxUbeXXmes1bam68i9JoczYZccrOMtjNwZKLJv8pvctxy7NQUuAkg2AJqAEX1chKvVRIG
3/OKVosKl4VQ1EFpCSZUk/bQgBV+ISDQx9HxNrckjIBc9JsQehuv16NfV7C0BKpsYbho6/DDzG5E
t20q70SuZtxePV1xmFKG+Ex48lBQvQAMYNLd9tKED3dA7epniPoLJJ0AexN7JG651H67gn15vDSk
Avf7VXFTvqwbR7LUBOI0dfwGmWK8zCIvnpsKSxmLabbDR5uVzhzRPXx1KTfiynpiTTKwZsl/1AJy
DJkFVKEiZDfNIGRAxe5tSa2VXf0+6OsISEr/Wj4NS7hgdhdn5P7lBp8SR9JcUKtrVMR129tOmTGH
53SicnOBK68+cOXIIOtacQb5ad6zWTTDo6XDDTqzFBswZSaBGGnd1oYF7Xq/JzADMwOh2o/Z35fk
JDlKoSZC8sszJ3D99fyi3IDsjrx81cUfBgOtTlpZzo2ILGh4VTiHX6qca0VFsDH9sRM54pFvZ2Ht
FNAsBIC8Ff9XzoCxRoxrzZR6TRv3aSwZpdPSTOhFEj/szjo5uy3CEfn0LTAPYMrr6L1flgCiriDY
YBndwN+bQob0II3PopQMk/QA6Mf0ZAmtQHGekKNKhLBbDa3IuTmewsxgLfEgVp8RIDhjAXcFt7fQ
hGZj/SKSGjmZzhi1bGyzz3AOUw82Yyw3jHl79ljAcOTG2VMCGv68f856O61HTL58ZoQjMfb0H9JB
Y9QqVw57cnQy6eFMrn2bKn8YS0CO9Iy6brFfd3RJDri24gkX8ItiXWyvzC98hOWj2ykZ3YTiXxiQ
gIVjZJxZRxHeS0001rgocg+4F73LRSPPflbd6TOVuufEcFUZ8iBkVA+xFakyysCcSARgzRj7ZeYL
zKzkZTaNpvDzh8zqS1+PLpM8MF4jaSlgSl9CbQHZ8K3YpLWVWqqJgZzJyFX7cn6J8AGhxp5GN8EH
qeItbNBQnCoG3Uk3qZKyJeDak88ZYoHf+fHuLy9HBJfzgSZ0pdGsYDQYJ9ew7qrLZmdh4FaVdq6w
ehgXPBrF9YkkbyO1+rp5C9LaXXuVtV5CaoWtJ46R2GJUkiniAIIPnqHPaNaNIOfnlyMX+BWSUP+k
e6/6mqtfsKBwSrSmNPD4Wpsibzs8uT1If3tPJKV2+nS0TLB36gwZe1MA6llZcTzG35PBVAYW5o1u
IjPVaBp24dSJtOJNfb59UxsHoFthgoWlDiFlgGGmSFpsgql1eMvhRRTYc/BrCKrxl0WH7k/4xxwY
/eDLI5opEBBKrYMRNhOfoTTWlGqEJkxgU7A3y9wCjMpuVFVZbBcufO+qjHRQzI6/aG5T2rusjE5S
B7VXxM+1WwQ+lcWMzImhfLk81oDDf7OxNZBRqkca9NAJB5WBJzxZX+17cGKcSLSBFXSk+B0jufBw
TUn4Vv4+E/OvnBFBjfXRMuSEwe5LK/5xyMrS8jXsyyyiK2SCXhJCK8o8qEnfRsAXnK2kcA+246EF
3RGIpugxnguqZiYIfvFD3Zw5BL8bXdw349i5/Ua1B57/vyeaLq5b8fD/ZkhVv89OKP22lG6UnydX
QxKg9hi6+SARfmPIEA7tTnoyP6orK+WXkauIg2jOCbKkWazA/GW3WVCVUHhKAE6QIbb/xOt++OFe
emeYWCU9o2wJOfFYXy+XCIicDXS0PWH/5fMN8CdQBNnWgqvCx5unDFUW01c19D2vUKYtInLvCEH9
2OQLJswQuhsGsTgt89ZTwHCOq8Il5yrBRPAoqENC8hhu6ae9H+kgCh2XFrt0vOU/Sk6AKMi1XYjQ
uSI8HOcTGwcfoEbbkIvR1KqRnkbEqbQ2edydQQJAGxyc97/NbwjNZydw/DP6JUwIz2/9HsxanVuk
GcjS2YLZFGv8/rLsB1pHLE2mrQEG8vsUDQOlbc1q2aeYgzU/L8ZBPs9yfpFQh6VJUuXn6YUWRkYL
2oMwA2V6ediL7HYa3nOnY9/RRiPXc8PGVQbc+flFm088y0DCnkR7ew2uuHy78+1cbx7dcorR4xu4
SdG1LC3+ZIIt2nJvzP+nBMEKSNQk95BxBaFHzJlko7FjmhTK1FuayD0MbL5JxVEfUtOKNiEfEe7U
ENgqqc06/QsJKxKKW/PWsRjXPVeH7CgWsseEN0eUGXB7f32iWTN0tb/gQh7aZClyv6AH4vJxpZv2
ILo+rRw4aVNzK2HmhDLh63QDO7pA99KBAkafgE8PDQaTBavNr5wiLpx/01rpd4eMO3M+2GqZRDSK
cpf7YN53xyluA3S9f7N21jKtMH/CA33b/DdhE1IKkY2U1AnGXgMr06MusafWK2oZS/8zGcDazWGr
CCINQcfk1/iN7xmWguf2Vb579xEUDjmnEBFZ7HPkxgpqgPAIIe2/G9DFvlTaV81jvhAvhgEYPoGD
ivP+THU1DdXsRof4Ug+SSMHuYB3ndr2q20PUW5NIITSBlVtS8ic2RSW1XEQQ29j+N6bnwIsNPE+H
M5idd6XP6OOFNqp/sMZRwRBla7yH/z0lrq29yGEe2+lk2COUnSkI9XFJF2ILCJnFD5FifzEQqsoS
3/8zOKJs56BLiZvSZ8z8P6B3KyIWdOQn2qSELBvEu9cCTkKHoAoqF5+CcrHN+IBCqvEnELXMzvvF
g+d8NDxgcANcTmXRFe3yhpYy0vc8fFE9UriKLWQiK9URcdc1R75LaKJ4+jwoH7OUFkO7H8zTS++e
+GK/CZzEwPaQb1qtGuP8puP4KVzKP7QYhCWRcpZ/DGzfWHnJdmFtwDtfKQ4L4coJPwG74RTzmeSn
56eSujyUKVbZaASYWhG+tQnh2OtqPPaY9R+yTlhfBJn9e22eqLEyZXTEx7YhZ1Jlh0DfkngrbIsK
SZ04cVhLldn9I9/WH7JTpNWHEVW54/AmmFQFZpGBQZDTPM1HtsPW77PR5gWvvi6dUNUYjwkULPt0
wP8k5kA4jlpAZcUHcEf33sE5kJp/PVntx3o+50DrGRGm7GZikThWzv3ZaeiF2TPhn9WwCF7TnIjY
DL9i6asw4SPprCTTBcIWFbX2WCGGA0cVruRTbG6QKli4/HUwJEwYft2Oh0wxFbfH8uMG8wr5AAEa
2NT3QqIiHdTS+Y4utzRl9roYP7A0APWU91AX4EGhfkgDBLAXdv4i4YmJm4gMLkEFvVJV7qpXkvPp
KRBB0E6VtRrvzaSY/iqkYNqrtkoTSTMrZ7ff/qzWScH5MU5eiQoej7pjHA8L9cXV3LDweYm2oSQT
TUjuGkthhq9LvhvDDrNRbTkWSkv+y6Gk3z246nQEKQ0x3gFZQWxP9yRquvOnrK2hSVUMsmJrH3uh
e5biB1onhXBPuo5sOi5wymBnQooK7eZO1AngR3GsybX6BARjYc6vkkKTOFc587jVDgyKtaETtPq9
fH+uoIjTl4YKa2B6T+Xm96KtKET4W0pOmCTFVdrV4SgwR/nWqCxmAvmSdqh16SktYIeHmOwLxI5F
1pFEQ8RwD7hluXt0mt6nXEJI28xOn2trZ4uKB5e6ZTiLlqS79ie7qLEh57kBhInFPFH49DocP1RJ
hnKQtctJvQg5q/1T6Mqkm95XmU6RrtjVRaI5VgvGecLb/hTTr7p/KsZPymxoh0imbMMbCXBznn8G
e3IGYs9R7kBzJR6eVBEDctUg2LMWOk3S1r6Hy913oFW/dgkAztQsIhpKl2W8LmFa20s9+fnsypfL
hkUa6cbVm8doG8QmDLqrqeXTy93pfyxBLkgc1oGAQgt3ZR9BdogYudNZ0qZrWwWjpd2CMkpjbnA3
r4IdkcM9JscUWPwyUudfKOA3UHxf0h22mIvSldfdYH/vQyEoJo8dMWxK5Xhcd45AfEnybz/o95/1
dKItnJ2yCv1vAvVsWvoWXSI+pDJGJ6hPpxnjMFBoSDTqCdfLKZ1SgHrGE+8RJW6WFPSuav/6wFpa
5Utl49msaEa5N7WPYrTC17cnWKbxI/x/Ma+dOM4smwfx9MriujjKPYL11JE522nWEto3g57QGlkc
g/LxOVMZDR6F/ugiJO6Q9aTwRL1gE30AuxHmDLgF9sZdquxmh3709OgIcrwsZCMpa3I/LS4MPgcj
WPcHOykHdrJR4gV06hUkON7P9yRYCq44BtIPmZL1DJD3ig9zIr1d9BtuvJycQqHIcz8itezJZXdQ
Q15K7uPi+bLZ23nyNlPNCTxsPD08tOd6308jI3Lx3QgXzVy9oct5ZfzJPD9w6ScPJY01bRbAKae6
yLuCXloOUsDn/WD4KF7WhXmonTNDwP1Th9hiFQa5cs43C95hRByOWU9g3ZLBaxpPLANloZpm8dDO
5z4XqTuf0Ib3wYxku4Eg015A5obKvA5lJ1PEuE6DRbeagi3jpZov/K3LKspBjIRd8WpWdtvFKxNF
a25EuyMdCpsPSZb0ece6ZTZjSYIR8g6Te0Zak+tvTri7/XSzypAEzx2aoTkU/R9FBa8vYC7+er8f
78FoMe45u4MlKbrkUeadkgo4gGeWAWePioNdKRN/FUfrvlSt48TnrvMZDLJqPvV69I83f+eusNuT
lhjNn8SkAuCuu94vLYM8LXkcCP7vCVY8mlHbpTYCCa8mCPQD+8O1AuWfPSIvFbVBzlj7hmC08lXu
vvTZelokq5kSc4c2nsu2l+iz7jfE7lga9xlCZYStMoNkxIs3IrnPkzKFQ6gMAQmbrw8exnRGmqbl
JFUetcUZ0qnPGjQh3IF/SauqlNNL6P/jYx7chZWIbUFCaSuUGldEAZ7jO/5bx2sSZn1sdZy49pr5
eTpIfCPYIn+u7DraPnbMpv+ylrq1YaQAdf09DEyco300b7gRgXa1mh2HMMR7dy4aDeMrN8M93nQQ
UkCof94f3j6hrFNFMUEI07V0mxmp19sFNc0iUfWe6K30obQo1tspGOz7J6WRbOvE0T7tTMJq/I/y
jV8FV5dQ7WLhtXSdaWmXXIpioua/2Vd42Yb9rz5yQvHMip/RNZUqzy3Y6AhqzB4N+UMQETrnnLb+
pLefjXMaONydWGD53c3TKlGOYhplgUoxbmuyMdbx8IXwk0/nR+u6MlxExAILX6tS6SbZeV6Qo5Kn
n98eU+N0EPwPlwJztIigZ2bXhhiZUiymyYdg4/u88NdO/lBkKDCOS0ZH4dfBtAsSxroWP1QmG55R
89rLtrhLfDaLZu7i5qm4SZmTGY+7326WTwQ9Ci9dBENt1T+YFLH9nstFq6kZX825Zo7VKJzeOaB/
Ph1vR5mEDhXRl47/kuItIuWJLoRSae3jPr5MWMcdy9++nCJ/NwlcHwWmmBGTGFqDd7p2kVSdgx51
9JTH9DEg4OmGQD7OZKSiLRVLxsPBfMylCJwmsizXODuDb6hqCm2FbRQxJLraMqvUoEeOZWB28d1Q
EQNi1jm5us3aj+yNXa/OHad7XWzCuEArqA1Lqf7c0nCw3QAR+aZgv6KKb5tSIB0gYIR5ZW8l4dpg
sY+usHG6ftiriLg1D0bkl2mvXVShdESjRqpb6S0wBzMWIaQQ6QmJ1orXiyVufJdBMx2QuaUjePzJ
V5v34kDdaBZf4qsGkkBrDDeUCZpDBwJ1PT61VmcdGun8TLmnxCv0cd+M4t+zZLyzMjY8vaIApk2P
gN9ys/0ETszZEh8OkzZvoMxwEgAbzt5onbDHaMXDGq9WtmFBAlvXeCdrfuuW1UMc8G2CB16f63F3
OmDdXeEfhrc4kKilWvMM8OSs8TLZrVhENw58ssFqxFP40UD/buo+f2QCsYw/5Hq+p1ZXjJAVTnST
LMBPhr0Pq5zUuTnNgtO5xUSw8Dc5+hgNrU8UYGzFgrO/R9tJD9hE4GhKUYIEn6FbzBa3mgBjiFHP
yZolEl5IoC5MPPq4cms+e2xslFNojIhmeCtlcJvAZwmHMkqrO/P5WZ6ZKTc5fzIFzfq4WDbmUQag
0E6gccj1zTmuazyhOKnQ/7C//aZ3sylT9Uuk4/FAgbKRlBNsDirhkKSag/ptBGgmK7V++2QmMElB
qqzOBLZVtUkbaGom2kcqI3smWVREMWvZijmkmdeT1ebGQTNFSCUfgku7GtWLF2P6eIEhe81x7To3
bpDEQaGIzoQlPKSJs5Hr90BZ04EwSXbrvZy/OUQGPLF41CZzAb6Djhn2jXnatHuWGWB3g0RaZSoD
dtPPSseuTnWb8uf0YhdNP5KX/6brfHWCOkWRjw+BWJHvAsZDgvCFVOrdUyip+2YJ0yF/g+Sv6zff
58JGLPsy6NR2pPoFqRTfu+GEtsIj8430lxC3fp2zEt7NleHhzdeDc2KuiQYyhQBvm189anfzTInf
J4Ysoh24iqKFWKoNSq0W7vPm8luo/R8bEv8yy6C5oT7KeQeStmHpC0jCI47MEEJSfogT9KiOAAuZ
ypkNf6v8r01STirHL/Ug2KWKFOEDH3YKB6XNzMHBCkG2Y8sLoaJnN7xKUv8ciWQaFpNftNb0r1V3
N3p8wWGVDSm6M+pjxs/JTIMcL3zBi3w9IrE5/xqZPpv6s4oDmlmZ0CBlZyER01KfX68Xrn9B5BEj
J96qJ1UnLRRrGlT1W62/q/I5ilGH2H2h6IVeqRROFObi6+OSPN7jAp4O4LYBJq3eAUZlBzh/V1G9
cEXrt/zTFbZclTDhig/5Jy9/vGU5JDtueoDJiqFpl4DrBDJFvBrTKNv7ClEGhSGmeGLAK/8Tc+71
6HiwC2F5dmpKa8xNlkhUIAA87chtxk4Lt3FCRr+slktjcaxDzcZnjm7SuhCYwLGeAojerhaSd7ec
WD7t8NBtKfxjN6mkSvsxUZYu6pNL31W5qY++yvFkl1SDmbLv00VgU4I6Sao0wK6s5EBBOvXLWAVF
1ToVO/GnymQdlkCal7+cMJl0SDF60ztM6DSlsv0+hbRrRoK9Hv3RGI7mJBcXXl0YE61g8uolYQ4b
m3TOSHbwL4HKeB+5nSBsg6q/hKlIh7nx/BPnCGILyL7jpeMBPpi4CbSN+CUisos2UQ5nvkMkyVOH
Wz7plXcijBEgwy/8tBZZmUqSqQtuGqWiTV/DvxYwmQdF4hgc50mdy1WKREWnWurtR7yegJIJygKD
XJSsurwRumo90nJYD2Ca7oJjH06sO+miBhWNG2k1/++DvWcp5u+8Kg04LLlyHPodgOa6tk2mw2mI
Fz8SNYY/Cj3njnf9b9rd6Mu70268lQFB4Quy2wli6NoudjK6zNlxDg7P2VuLBLca2U5vkk5DCZxS
YLH3+zMlgYFduscGhow4OUjkIRHMNbL2ttJVpFPKSWpfiT/VwZFbyKJwOeZLeO3WyiN9HnmYJz2+
upIGxfjZCh7Vt2RFLyq6lTVwA2f1bUzDNE2etmx+oKJtywnrMp/ClGvFX8RVR1pSwTFJBtpYw/Bk
CxGOxoSagauCu0PxYOqR++Xhk2tJdEMyb91rLgBxw8XeLAYctHKqWwKWKCYZT79Fbo5/MFGJ05Tr
cz3I00SWq4mdIzmgJ3Jqdba7Z0ACcuDOjPPPTalh2/4IE/kY74WoQQFO3hf/G4N8uxdvUQSrqriw
zym7SWMZahEZ8LJvxsii2Y/TVX+b8zU1RunUZ9dI5kNThWTQMdIP8YRYLNwBF6vsbMO4P1Jzh+f3
cg8tSGJ7XH1uvejKeQIm92IuUWR+rfO51JgMf7nFgQLYdvJID2QVxjBl17ZVfzp5aZhkQFwhl8Hr
adRC0BbcSVJpfSC2/XvaTfiWRQnw2RgmJIDX3+l6J0DRohfVFLKn75UeZxFwaca0y+4g+W2HrKoL
ehIFFaT7N+mt85q9lIcPS7+rJIRqPFkEJm6KWFEjkkB4mny+B5eW4wHE5ZVvVuFZzUopyjQoh9hv
JnlrgTiSFXwMh7QFK3fnwNOSSUeKTwh3/nH0IqX0XGXQV76CjtbUuZwPOroHY8MRAaqwLTrg8KW8
TiLFMvEep+4YdKKYMj/6V6DlvNb3d4IZlB0+6HkVfAxhm1heNjQzPRjJHxfFuCfG6wsdeSQjQjX5
Jja4BFCNgex/ijWJRV+lYbeQIPnzkZTEJZsKpDX/HqLgUQCu0RvaydogE+JD8GPA0B9huoDY/eGT
hWdLLx6QIdnXWNUhssR6XhLSApYBNauG9JRYt1tzifWX+uW/BDds2Wmae85uEvkcS95sHHY6Nzl8
vdGDNBfgTvQKcmUO1GXGy06S0htiydEn2XhWMfLzu0AMLeGgNtQS8EEVSjuhhjcKH2ZH25+5JUDv
QAYZYhEnMjEGtUiVx59OnGlO9IqdgZk/CDdDV7rMEyy7z4hL/d8nnWpn7hsytVzvkBXel9mFeghu
4c0se7pjDfZX7G98+9V0FKl/foqhUn7sG+Xwj7XE+McfG613X9osklp5oZIttya+o3W1I+rCobdt
1bOUy9R1g9HQLCxBoNywapggMrjjEY5aMUP+FiWDghiC1shvd5GeyQvAnJWi7ez1fuRvVfbVkZbS
X8ty1fVPQqxfQEXUEbpQ2dEYbeHnI6yU6yp/hpqYRUCcGo5zJKYtwhC4B9Z+7c0hLxdCzPXnoOuD
GMC7ioXD/t4JU7cqFsZoszXCExte2kv54/wbhsPhE6a+CTznn81nSiF64zc+aX7sRBhkWmzyA8Fj
bt2RrSa6xYPsTETuGP8zUTd6J2MFlqEaDWcStYNaagszLycHMxXhuoADXktxGqYGyQfdvCzXq03Z
bki7jkxI4u9Rqy5Zt9Zkt15jH7uATBKjjgs5C0wz53oA4JBFPPR93KxMQm/yFtmuBuuLFX8N4XP+
UFjhbuk7Oxf35rmaUry5Ql26Boz+AyXoUjjmUlzoBXP89M6f0qtGYI4rxrI9d1MHN5wGvYvFdqfU
xYiAQ9e5W4cpp8VR0R/8a5O7cYvZLVSP7XQvA9lGVRtToCj4BOYrcr9reBuTbSqwOZZG/9JlQwkA
rmiRO1B+MD4ceDPJZ7qhv8DHZucReExUegrCeQgFRMVD0r3fZ5crxYN7ubTJLqrzISPAUPTb8oex
OB0COjImyCFGfe7a06dv1yug6+VGlYro4Sxj3pPjLG3ajQORRg4ZL6K7J8XP8BvM7mH+ITTWaftA
wOlsZ4QbrMTY29u9A44nvQfATeVDHkT0oAJjtAs+eaKDfkX1S5ObGL3BjDfPzZ2h55wKQEk5auMV
+gWiNXx9W7ll1g/t6weYHRWYBMgt1hJovO5U6OBu4Zz0WUy6g55aDmX5PtDQic/E1JANPh/lbp5H
MAghwcjd80pyvCSppmi3zEBDJ58FdHfr3PWTzzZEnV2SxHSwVWF3Ybsc+IIEfup5n2Ny51VNNb0H
LK6dXLQ8RKxQDluvXLxHrnM1FEYqCCGNQp/TVNE93hI+Yaf/eHx/1nrpkRlPCWSopHr9JettEwKT
YZJbL/f50cwOFFtVKH9+AJZowtrx7WdzQt8xSIF52K/bHnpneKhgl44CKU3OjxRU3n8zDLFVfhMn
XlH+IU29DCYkefoYekjxTT/+vLLKeEQeLES95saaRPkeh1jccxcTcTx49XTkAqPECixf4RSu9DJ9
ZLkbxWsppHqynUqICOof2j5EdIzUeZxt+dTPpeQY9w74C6IhPPPhs1yCi3gh7YmR8jVjiB50KwvE
Y1dk7Qw6Jdghta+7nur5bGm+umCTsBCWr0PfuzVjFc+9Dcnd4IUD28fCcoqjveVswqfCevTh5ZJ0
1utLQUllFUw36Tj6FzOt1Rsz6YUAnBi6juz2UsF9dZ1NlTIgnqXgQHlcAoYlc1M7rrLqTjG7vtsV
0/jufo9DoStp7xDsadFgv0tpT2zhm1IvicBFUR6WCUo/2hu3CLJ8iCjQgRnJfKlCDORAxDnQbF0h
/D40ITXqi+cgCSj+nPpVmcEpx8n+toODNmPMf05Guk6fzbNOc9y2WnJMjA7U0WpAWUj93buFxZbw
2QGJWRU+U7z/oF6HRsJgizpTsLV7uRwAk8uC/v+045mkeImLpM9IRMYcpCMebuGSpCt/W3eLVNTu
pJDJ7Fq3hcFRYcPTyrVu+u6/jyDpCN/HNmN96pKAb17uWjXR9p9mQ/pJA1d/yedfEX609l/kqu5W
Top0Pgxp6a1XtCwRt2T7uaI2dUkuNnZXijwTeATkVWgKmPDEXifxjYDSdKd+VzzmnFC2dBiCYnnX
crN/PHfgHQV2wmdFi5pGHJwKE3s/XdyNdn2LZ/zBlJtOzoMOvgxyaTilUuuZGBLOEGlbsMDFuJ5D
IwmXQddMUeLy0LxezHGFZKjRriJxd10ZaxSy+jve4OWJH999UBAiUIeTXvYS5K9KpfPc+9pBCwPO
2r2XlsSckYhamM7HccZ+WQKemnBtdHAqGJzsUk4lF7izoPdPDRXtICSwxdjeb9/G17HnmClZC5p8
wNFqEAbjut5QPR+cpLrkJWYd3ABRk0QESpDbci3AF61Vg2mseSqBfG4DEG2saF1Cmx6222EcD40s
siOwvfSEMTrS/b4b/tFhqUdyiolHApMOiuGyTrGs5Aw0KplrES6MmOufFzCH/e4za2wWy82Ko4GX
H5CDygvnKjVgHMTu5ljktb0efmVXIJmNOfO0CXgiMa5HKH5uf+mM4uRfPvEFBzcfIyadXWZT/sba
khR0dBI4WbzOvfcMsub9FXz9OswTaBJCNSkavKtD9xbRYxKDKDluNKvkq/N1/md0TNb7phVYpZdz
rd0RC++hKfJlI4MQcmszbz6swYQukPGzQ6EGEAUSRokmhDPkQOcSciUSYt3MiIzn4VHIQ+TD+KQl
jPkq+OoBGp+QxN7UiQ6b9/UHMkZO6m8O4el2Hz1KfRxlDcw738XNBTwX07PmWSzpgUQw76nOAWZe
FD5bC2aMHT7pU5oJuclf3y8yShJbB96DWlAz0mGvxs1ENAMmB3xZdtAscBfGsUfJ8waWLF38pu+8
Ns2EHgiXcJZ84Xe5/l0o3BHJkW/728+61pFTQExTLItHaC73zTf0hBUKW4DCFEFV1UEqb8tbKI1V
TffeaNTHlb1LNG9GJZQy5FuV9U87P0gL0XXLzo2KbndRET3jLaH19InpnZ1piyI0QK3dP3Y5b0lR
xi5xcQEYw7o0/NxWpSLRbAjMhawSfO9ckOaIJanOuk/mmtOlZ5rBGgoJTQ3PdZ81c56DnaIWWq/+
u4nUnpRCm6fS4vm/pLUC78n/Q2IW84qvQDhtg1+7xS3wKbKzIAkKeTugYjXp99wx5oSDiwT0fklg
kS0EAmgwve0s8Rzl1+NvVPRRIAFy8FXEPN2Zwhi0d+GGzXJAHR3qbDKpqSYrOYjuxf31JuU50Ncr
5BMtBKMzgyfe0JOyaAmbsX6F+F+qlmGMac7Vq3otGVTXC2dJkf19esBl7ckovzpLMcFyJ6MwxfqA
FCT3r+aLCfaNf9nkWymvDDCpShvFjEQ+uXHiureaxcuA5hErOE9XVgnM/Q4mD9f0zzq6fGBXu83E
W8579eoC7FzKqJUz9tG4tdjh4u5KfTPXgG8jFx6zU/kyyR9IoKyPjS/MRWCP1RZYRXGes2YC1qrQ
Q9aziTkAAhQYhYxVi+eLZ1lnEwhC4nUsBO0D0LzHdKhyGLNJZhfMYOx1Sx5+3uGsKufdP+dobk6b
n8LOh531njFjBgTOWro5inXd/wmQFRd7ecIInLcQ03/N8ncNyFy3TVOIdBo1Cmy1wrvJ0ncFTGTi
s0t3l9D+KNawaA4HoOzEGgaOTkd6FY7tP0crNKkeN48/bA3Bp1CimH6xEACIEL/EsKyUUdcAARPi
3fLy+1ncOA9Bw766A7XyhYEXExtgbLzQimg8+Nj2Xui/seAqZYUuV+XlM8xuS6AhWThszOZvHNPo
wHUELUMYACC58a3otfZrTzBZXIItcat0ilJiR/qc1v4ZQx72To/SpNk+0VVdibApTUrykusFQG2C
Spr3Z+rmOjJiHghBbowoeAKwadWmji9q6/eBmbD/OMpImvqlz/3syJutSYKNgnu2H9EHwxvubI1Z
tGbIlFYIUHv2pYgTuqln6R8o65eznkjNJ5tk8b1s3AgvIywCD9hb1IXSXI1q0hLv/6xsqcbXOcbJ
pm+2zSiw5j2CaScyY35rzecgxq17GxOkLPDgaXfaybRG9FXOzS9Kd85h/O42CjfeI1G8HILnIaHI
LPcb5FypV6d/C8b8BRFYSPgnqP5FDzwdpOiQdlIcERpqDjZZ03+qm+P4fMNyuy7QER/V0zSCub/E
sGBqBP9EHvN5yqcVW5ymSJ8f7xLQpAQCW89H4lWCcXQkInvGG50pN0MjRr35JhXKU2anbg6OQX6V
uYUcDPCxDuFScGq1fn1hQSH1KnRvj1Z+WGKKZWqbswQ4Ql/nid3Ou53y5qKt7hmbpf8bM5BN4FpU
6ZR5An1Q5xr5KakfEHcsROzCFr8MQJnHEF1I4A3LUIa2a5SOLLK+M+x13UtrcO/UUY0JO3Rf8Axi
pQv71D44bF3uVVczXB9SzhPZCPpMwRRdLEkQnwaQOPkhg+Wl7ABFpBuCtyK14jQTj+sIOhPqouJJ
N2AqmJTHhnAu+g84HdnaK7mu+/jha3F/XAPV9eQnZ+JWyLFuOdzSakfRc/btEg4aoTCXQ9RNU6PP
r+HUeY0C3VrF2S08ihf944NNXWY0h0+3+ezsVLsuwhdaNN9swbEeyUM9YSm59TlkDL1y2FNkEMr1
oUCZOcUkfP4sHh5ROZkcaBl16waJ9gCj1MNcFQXASFLiSTqx8CkjkQeCZkB+5tobqdkxeuSKeGEj
xIMbG+9e9OZzpvtVB1XZCwdy3dse3IvFKmF9MNhudr1IAoERE0PLiiuTcvUUoBKk6ZKA3ElYtby2
uHkTEDaMEOTtHBX0Kaghdy0jexTlvN9jpEwNW66t9tTxzkyxEaw4e5/8dcwF6y7HO3NNIEzGYa94
zC7r3dWRujXDslSP57U3glvJ24VyigjH3VJfkzYXTva2bNSuIhIUeCDhN/Oa8Bnuys+MMpFjR0cY
av/sOxOuuG5ftOBhJ/6YSX5+aOCT5F2l2yDlLyW+9sXEaXAHbzQpKDEGhlHdQgeowlA/83yxPDd+
TDKgqXY2LpKJXML/2KCP7NF6/nSBHYfh9A+LP+WS6qDf0yHWI3JPEaOD8PVKyTemdBE5WBNvtCZc
VQvpte5ynIZMxsN79Z/tcH0RlRYtAKuBcNN9B6nVY89qegkrZN6dZyEQ2FxnQ9oW+NynWDbyoJgJ
FF2Deaepbb0GZXwLW6lbiQTVn6Id80M1vPlHZYEqFrpncuzItaHEif+Hd8jpQvo033nALv6gWRbg
C82AIRo8mhvmy4mTV8TtTXcAFQYkDFgHHK0zLVH8kkt2kuegNf1U5Bkg8AAERwokUtzAAqiFUYIY
xZiHOupG3bc7WP39JImQbNLby++9m93uGZfFrirs8UUmFvOxwNt66pHyQFzTeNUnEOpr4TuXE2U4
9If1TQBYpj2n2xW1qAAfQ2lFUFWnJ5SXR/9Vn/KOHMVAub6AEEbKei1NH5GYQE2K1mzNPnYiO6Vm
pia1X84RxaeIoTB/3QeuHk3Nce2E9PKYwdkcQ3/Yjc8a7iVwIFMxCGhmmxAf4uO9fCAYHHw77ARg
FUSHMGv87xJ5hb+hX4V3DGkE+pataAME/MLP7bVHkCJzTZQQEHin14lahaPbh89qmp0abNSmgfkH
ksofnTs4fzD9BErHeVy+mMHT9DQ8dJfuFScvlUFydUZAzrdbLhApkfLURNFJCg41ea0WOXoLPQTo
1WtppnUZKGUBBflNYcAi3wb1f1YUVUiDPUpRU21sPEbVrau71t0hkdKn3Nu3VmpOhEhkQWSt9du3
CdojKhA9s5ck+GJzPVrR51nSt75Ewg0hPqhk5hHTxT/g/4rpYksX1GyWnyZZcfPYhM44rKd1pKRl
R4ZlaWfknls/JRRet93b3h7da0iETVtADdWYuSfxMABOSuU3BTDPjTN/IGQn8KvaGp1qFGxTzzqC
WSm2MIgCV+jYZQE1QeagE1J1E1dS9XYwTfyZuWBN8ZySmV0rPCAup6LdSUrtVV5ZMR8WqijPtp0f
i3cA/cLrC+FmxvrvqO2x0thUxg8jEf/HsCbTTtlnqjvmCH/XLZLu/lYN1L9roLlv5hcoFEqVBsy/
EhA42D0TLreoeMulI0EhswGupmRlRaQunA2OqgJopo3Bbid0EgvrxFefdyns0FW23sjI3Gum2Wv5
Pw4Ul03gFL+J87B+oELm+QhbC688ptxPbtnlCEecfexMbJrtQ21ZarNaYss8uXAqK9kbadU9t2VC
roIzxbnPvF1depFQUeL/BoNlkbjMY+rC+c8YflEv/hnl9KSU+7OfPzuLoG5zz04782zIi1KXBX2H
63oV6x4tLh7btck5LL7Jo18mcY60u0hLR6cFqgj1NcHMtWDymPRQ4HpDv7/Fus1N3G78TUz44iBj
kwZBagAIB1qUNfu4sHXPbZ3Clno/JQ+ZkJl1Y+mbi5CkGDDY9UOlC68V0DMQaB9LKHjxtPYNkxKu
0B8oZWC4Ix7e3hCZQykVpFmeZ8LmswsGHNUwxdJKWn+TL+CVx9oEr55cqvFBiLawpPyElAqa26hO
OsIILkc4UgP9DSTSYZjYtEJqqj9r8pDiBj1t0+YeB1nmOkdll+IFEC/lc6+SfR3ujKaRp2QqvBzC
9+GD8CyyjIQYeYLlNIHrq3bYnG7VkWTuxnW/qjKCFc36ml3PZcLLhqahsjs8MBFTGNhXnAfGTi5d
fILI1HtO2T0UBhPk+ODVbVoB/dF5CHvTbNL/jewISQdjh+GfH2Jakx2V1atw8GTKeGHQ8yFkyAYE
GTUAawpazJa04vusPLPHn598plCfcuLzWcdj7HeOAe8fRmH0mru7ieCLNjxQUIb/kQ9jxeKsXRvu
M4+oBIU316StNng/9F7JOnU/B3zxwzVtd2pJCU5hjo48at9zuNn9TgZiVkzPri98NPTtp6Z0r8jO
HhAJHjTDut/2rpFjoHYi4US80tK3/w/3v6GYatQFpB8LXXvjGEZQf3EPwi4bxj1H3fyVHVxgQdnn
zkSnodXTMzpQs9NYoiL4uE+yhgc1LWEyg3A7B/GweYrXi83iRi3lLIpTflnyUXWKNeI6tjDloPb4
y+JNTC9iHqHp+dlO3gi0rf0YTaYFrwdU2Q/axMVpQ6YhoBCS2S2zl7q2hNUdcbUs/4H/S7eV0Tz5
6uzlvzRQ/S1QpHIMw23rCwsNzyjYJRjfGHH3Dgojy7HJ6rdd6+xKzFjTtewnQ+eUZTGX+O3ihzrV
KjGF0Lcr2N0KJv0eNwCmRsSrJ1dNBQFsAqWOseWO49RozWg57dL+alQxf1+AT9PuA7Du4gCpdqYv
hCYIy0hV5pKjwCNsJfOfe2Msp5+QX81NE7MPmwgJXh/0tHnCkk7ZRjSi3yb9CbW4lsXPrJ9D7Xyj
xK9SlRgee8ihO9EajvafzV2kU4WSN86vedai+eGTfJDHE7cPaiGDBpVF1VoBA+90+0guZ8emni3H
9BkOkA1WzTW+pY+0mVnUAU7quRxufcHv40yZHDgifP5egBiPjkF3SfmUOUphSJwiAxGuEWkokTUw
MCwjLQ6w3yShhaUwAGF+TQekmK0cI3dCAQXzSsqxlVT7BeFIbyupe4LvwbNdMyMo62B3KbwlDS4M
feyHIpy8PsU5+bdefXZ2+PBj/l0jfOwPuDE3g2g/9/nttO4ZLzTFsbCUG4RRY4BhHF1tqPWs/kTg
CtqlZKYtssi4xKHEjl23yMSkDjykTCDzQfGiocxccGIm88Lt9XPxRjaXtj1EZeL0F4bDEqFpmY6G
6yKjznRpPb/g8Ka4xHM27vbFqkfrFJYHF5vUVKY7Py9ipDGtc/wasyMdJTWo6/+2gTnNRroPKMqR
JsSvCFpd1IdZeR0VsxNb3dhTfMz6MY9XO3nTkDEBu+xjvioamWoypuBojuoQNdKf4fVwhykyEcik
DG5RwWfd8zZuUd7zg7dE6QPkNcqz9r/QNOdVuWM31mbXbs+RLvX1gst/wouGCfgOUrfp/uyeP0gy
pREbzHyzaawsOnvbrNQyqkFh1Lvdn+l1XnsZyq8TWfvxiJspLUdB90JF+K501DLedestRgAnJYWd
AdC8VkuYllL7LwSy0wVUHnOSprGXBRw0rnZoZxKitaoJabM+pdTqK+AlyXC8qiMJi2AUhab3ou6+
FSB6uqvfRZPF/5yB6ktxXnr3GuxljK5L883gOolpQ+Q1csjRJ7Q7t1vIC8Ewnc+NlN2t2bSsRuAa
8Dd5BVgTKIQe0ekQiSihacwgNc6Z7IZlCbN1JWkat+St9PwBSZSv0SZy4kfu7vbGVXiKKrRO9qwm
s4S+pKIZmwULP9nn6Sj2eeJqI+khT0P83Vds4zqimKx5lTKibkm5My3xE9ngLZDG57JzBh8prvtB
3XFKNZbQWsmCZNbjrtRq0dLFM2FoHLXCf0Kv8x/BAbet5JoFCvjFS474V0ujl65u2VgXpPTJDHfb
ZHK+vFb/jFXAWyKyu1wKwYShOlJQlFUf9M/QWJY/73kSEYOOOraFd0dNHeX51rJYP/o1GeKcZuUJ
uE8J34WHoa60BnFy4M0n6Ii45Wi2Yt5oe7iUMW8DBX2hGSbPv8ZAuHTwNqGf5MfubJVxPr/QV+GU
F3w+zklPSzRmjG08QBcof1+nx49DPyXZHxaRl1fgIOQGQtkSC7tU86k2qrHyrzOxAe1BmOYl1t4s
l8QKjVaOHU1XbXQQmWLIJt2ebc+UMo2OD/toe1gRgNEhRLzDAUjaCN1MfAjVXtzRAFTdJ0C/wd3e
7CK3KeJoeRAeiDlkfZqgSJkTKDVOOv7Ap+PCpB76SIlXsxbOkUz3nshVO1txtAXPPZux63TYwjMK
0Et5VGwgSLY/CvaVs/MpZ4+R1tcZ741AwzCuQ/Ly6NUW83IGWfLHTvKW4fDByYmkvOAxh0BFY57T
QtVtLaJp9vI7NvZlQemrBsqjCd+v8V8E37KG0GbmqMevlyEceN6soRL84SGm7+xFGKOo910tXShd
/9dA1G22zZJ8vyNfSkYmFFafSqhuZErUlGH2DGyMwyQjRCPk+ScNyzYOzT5kYyBNbSYhb36/II0+
aH83mZ3XJuAURIEPy8p9ZZWoENOv7OzlRcKWhnbgJv+hcaLJJr/wUtPwR4336Ln10eom6634odGI
+mJId/eCDytp6y5bdjyAJqxOLSAiBCNh2TYAURCrcBrcfgBsTB7E2fo+ThJbFIhtNHNBeYvavcv0
PRUb1NNACNpu7KecwX1KJXAXBzZ9ISqj0MTWkpITZyFCSvLlSWySUlmCdlOC5ewekzUAnGajGv60
6OJwgR3erq14UWH4/rVVShllgtAawibJm7kvX+BCyP9XZ19H+ceNXAAy8Qd/EvbG+MyhouBcx6I6
dt3DZbbrarpgkhoMql0ltCNXedFvHWeeOMI86x/mTDDFsv0CHCH76kYdx03pEPcESIIHTIqzTzSU
4AkpKmwepAoofgEMzrtg8+4J6K9iuZ9/zsCUJwZTa1sm66BPH57Gp9C+1jswHiDbDgLrb/tEiWP6
S0WllO1KgPhuBF2+nqLfBzQxdXYkf2F+ggfZ/PHZZdq1CIJzzinrtWGhEQ4ErC4Wfu1Xcx0lE1Qx
+B1l9vkEf/4NEJTMwQWHbU/lQV3nRScMKV8icsMMzcPx67wSK8OSVzutmMAW86IF7P98hyTcZzBb
0G+2KtTQUib4Nykuhll2U8byC/QN0z6JIodbpYGUhVFD1etgAk+7nTDtMjEbFqu7/nXnUdHmPTSd
FxO/J9WpEtXefWTiOAqY28gLejfTXL8eT2b5UWi11KBBcoq45Ra11bUj4CTebrpabkHuOSJWDpvW
pWXECLL2qJkDn4MBH8oGv/Zm3ckq6QARH+9Zhbde5hrug2fLBSx93LYXDZclwoiULc58CkoXSjoV
/1LAEzRYeN5e3qKYyPeirwoa0SioKoskIedhWKf9syVTh6UgIKdzGZLoP4gN8uIoImC/jNOBLFB4
YYpS01cTTMEddbuDgDy91Hn0gUMYvRq+gP7hJoZETUGNhGOIPJ4BWH2yKBIEjmBCoGMVT0Kq7FOs
g728Tt3+m8SkBPok91Z/q0d9jd1E1P/k5TFYexduwqrZ1CQarGqwnuMa8ht+CcAOyJuBWgV0aoCZ
IuYWhX/BJqnPhLkLSdc0wSOYxk+STqykLwrltogwLxml1kAmHF31jtRcQ4P5wzedBX3L363/ZcRz
CD5lq8WKfeEdQwrZ7v4nPgI2Jif4RrEmKiG5u1a2JemIq9CmjaGVt3cqgBAUx6UPoSQ1/+oWUhvb
rB55N/TuNWSRBz0YC8msBKoj+HEKtZ9G52xFIqhOuVisx7BrGpJT/5rbgEk5yF2Y5Q3FkNnnfrYr
I7LgrF4HMjh6J8VRC61Qk969DZP2O/g+V0x+2b+YAu4C4fofJdl5HeYXxp6MaeO8CAXCOFumjEBv
UwlG5INTGo8zvbxQ9bYGFTzZmyE3hyiM52Xy/Tms8GnN/tKcuEONPhu1yT6Y+Nyko8WumhkcTc+L
rYngFM/RUgwg0/g7/dM8E+dW+VvySPKhH4+rWO6+1mWG6S4LB0cdLOD1AfJoVCLh6XH8bibXypbP
tkWbdB4orwEb8hr/cS6xurWUyjLO3o3I7bdmRoSM5lwkY8/1cUpMy1yDk4CsLSzGj5tOtielch2z
0H1omQE0HgjsEGZXQUGOHSxLNggOTOthzPrNq3i/ZE8rjEJGu1GP/hldBu/f3p7RiWx9T/TVoldh
cR9y1L1nxBJo/F6vZuFwoaNm56341OMU5eXz2UZ/QS0l+rDR/DsmC8j4fsJr7C7Lcv1iA5kx2UCQ
HChR72dXWBFNLL1h4qQfPMWKZVf/B/udv2gOU1+VwSGa0vpyzuzAHFzw4qE1eREp2oi6VxRTy0G6
b8MMH5qs/9L6DBOPdjlsc4Vs6c8fUiU9T6xYZfwL4wkh0nq91RB6PbKX3kEJ8A49D4hkK5QrkS2E
3gG5ryF7nZDJzLeSwvWlMnhBp4VkuuvzPF490oJ+AYk1GfNCM5wL6PEUEWdZgJJbD1PnGbdGdIng
oa/W2pxfDbrSL0Vp6IPyLrV72VoMUspq9LoPoEFWTR97rCE0vIVv7pVXpg/7x3PbHmILIpCpxb0C
O12cD3VlJCNELM+pqVORJXJtq5vyy2tC4lmGXBstEjp+eoA8cfx0aE8KrTn5fPYqogHD2x6pw8aC
hx2zbiKdo0hc6PJ6p5UJrxg6UbwZXwWdd2VYviKQdwWfaF7YSZC/18DCvCr9dEtj+1JVR8BogEQE
2YVr5gsKMW4LFQBHXgyFd//v8o9otk2RnQcelZilnrBfaD9PJyJw1JIzvWJzxXCg+yM0tM2PnEvI
zSaODzGKdCKAwvZWrDHQNBqbQgEnFn9P+QpuZ9ui4HydUWHjYQTZaaQa6lpTVSRcM1AnXCr5bG3f
xu4mClpJ7l3+2VvuzUBj/nTI5h9tVVGpDSZ7+CCIcZH8zWbVbSRPm83Y2EFz44Ob7Cc1DxKPQXew
t4E/shenuWwl3m6wqy75p+YASFeLSzswCy9pekKJm5mpspI6H50s/fLb6FVUfDGbDvajEOCS37De
oG2srN0FSJy6WxuE1dYnSqHLtXsUCzy73maZ2euQ9/+q2/ASRDXk3BcZTcFHmKOw8eyYdCTlgmhw
M24i6Suea6XIji8m2CW06XAiE5QUS0EnfalJrdo3f9DFFrtqRMcQy++OoAIfJCuLPPAseQLI01Bn
+81h7awiDOPssNmtRS2RR4cghAoYE6hXDAUi9fswcHaLe/bIxw9Y6HN061ZQdgH6viNYAXDTPVCk
nE5JLFxV0tJvjpuDvNYzCEe159Msn5Z6rIgP+mVhGnlVatQ3lfcQlWRLZYQ4hVxD5Z3uJd8KD2L/
fg34LuL6z5w2/81ClnSnBxh23/WaVyWkLqIkRuRUXM/l9rlrJ/XnLLrrViQ5m6GwOK0MfqCZSSX1
CdhY7LZE1DGzzYUhRX277KVBp0sR+Qu2J9pKULYvHGeFSIMzQqBvJhU0hRNvDtvhOfFUOn0Yb0+r
c+khTXuxaPhK4sfUSKikKbd5NJTlsS4/WQOT6OfnYdZ6Cu+F0gi/RRom6rs0nDqlAonnPjb4ISHl
WsSWMdecLNorDLCmV2cBHxltY7QjWoAlHxr82VkZBDTPtsejclsHy98Sv/PGkGt4NFEvwzjr8RA5
uumODi9isjjo8Gh9BMv0uPNfrkkZa5armP3pV8apuEQ2MVR0+5BrSx7p5sRRwI8frdQ7qAtSpATf
Na5uR4obR/KWEvfkuERQGD0ujswT8o84p7fxRchahiB3SoxVEYdvtNAKvPZJsj2raYJnPFpFpgc3
6wxEXDKARgHt3jEmeTjKH4ulMKX2OjBAyUfXg/zExr2s5vp1FJOglzApHZKNV8vvZcyFiG18LQDY
Jfv5SehfUFsfvHXNvtNDH8TrePhHo/zsyEYQ6uRBNy4EgdCck0x2UE+RR9O/JIwWJQy8+P/IOSvl
3JyCTHQe91vaJ35xSdkrnMeG+AMJ00mymz3ddoPsZ/NPfiQ0x5LsTdihSCojKEIG64n4udFs9fvt
iWiiy3zyoA7B7t9AnYqBSS8Hwo+vNrH0qwrZdvlJBcM41dkj1VDIUqnFOLwr0L0WscTOOU2rjkso
87FzN+JPL5L5NoGZLYGvrvrh4pOLB/er9WWyNTmTPHSyB73W7ACmshjLtO60gZz/bwrDtfrAKCe2
FzZeuE6KOdgq5r87owECyKMQWlRpbN4/0Hek/MQoAgTeUGiWIZ6qlZhwkx639/7OQEQXfbBN0AdB
uodJmF0ZHE2mJ2seWB7TY2DYdGEbOnuWg0aA7S3aqwdaN/Ni5DFq43xD5NsB1Zfnbws8NjYwOj/m
gA5j+V1X0EeHId4ZhCEzLheqERDF5d29axiURmLj/TrdRQV0kI3pTqlpXSD3DM51l9r4XikxzqsE
4N2S39ARzkv9W1ULRe8e/ssZgbOCuFwri1KlI6Hk6F94eRLkv8VaQPnGqBENNIgu6bcpQgEsj7un
Bo+kiL0ncagCsVy/y5gcf73eXyHmGELN6EhSw17CApfWDzesqxKryI30LyI+puD7Wqbz4XYlD0Ry
QTE25NzgCUHw/4we3LidF/ybcW0mJuux1EVAEdvt6r2RGxeqxc/fPKbWapWQ1uWjjY0HMlhWVZhu
/kGRkl4xFfZKPW4hQWpRZSx0P19FbXqqNBm9imaBMexeXXV0NeLHfVuRZBkD5NfGEF076EbntdXt
wsYBS2V3fpct/SSU2q5VQwr+0+duhDRBKed9KGATapNia2/s0XoSLgvsp3EOA8hAvKGhgAn/lOW8
slc44blQErbrDi18MIynmZETxkp903fpGLXnY4gDspyvO8TLeN+E2jvVOt4Q4HfMRwISheYcnLiy
Pp5UXq1YSMbr2w8zbt7lBRkOZLSmRPJsG58De4IBSDcu2M4GVSrXwzWPoOfXDhDcxeA8asaeMVNh
eLRCVGfoK6iGvdLV2ur4lYFWTY+tULUDKnvOZQ1WFQDT7NNOHfBbEdMuCj/6U20h0LHmRz2ySLz1
aVNvFKD/bWHbKPPpu1g4k7Wwyk6K99irgL+u5ehBm6MCxgJGRWIWccv+edC171776YaDC5xKToQT
b1VZmIqrrGAYSU7ztqtxi+eEjNPaoN0N/qgbgxze/Uerm9wtHKAYmlCKsC+l9I12nTQ9I2QA8QPF
o5j7A+ev/aprz7tJalWum+Ase5ASR9FJXdZTKvvkr45/VKASTUyHiaYHYyqGCHvOduEwk6WytasT
Sg4gWrSGvVlHyl9YASm1ikhVpazS2nm+XJ9EmjkJndblLNMUKCFzbSwhoAIxE515YtqG3Z3taXvM
TMIXVESkZmAGYK9wPup6hYI0CWojgewu1NB2QIUYbx36Uwvm/X9JvN3csGQuuiJbCdGivKt9CPdS
v7YqjJLYmvt4/qQlKWGJeayZT8VBUmbQrG3LcYptMvLz63CN+s0A0Ynu1mUvLK6qCc7AdreuAV3+
aOSA5zRNvgQc+0PHXd/dQ2sskVb9I/IvruukEHM81LYGAl2ITBM56SUR7cCc1lVHLSEzOFKfu7Ii
AXM6SpI9Oyqdo7CN3ewrwLCcC7E47446KQwGuntlWjZbqDzLk1fqxD2+J0m0ZXjzRItGtZ3X3GLY
FT2Sde1DjZ0tTp7M5us7RLXVecQ0YsxOU89aY1TMrnSfHgOZrjo3cQUFoZr6H1/KbRA03gmy9xS6
CRo6AKQmlwDFo3JP5aBJplkCIM2REtkmpAOAnvld7uBeY3DSJNL+QsaMLHwo4EyqY066dkT2rZsP
m6h8ZVIcCkYW0U52GwSvDaIIbJ/JAdar8C0OxzK808dPc5HVHuc+BYl9SMHPWmVkXh8ynFQm1uU2
ueXduWMd6zKU6deVaWU50vMKRzX8EZefo3kg02d9rlGWUsNIWuEmEEr43c2iHf1JH2M9uKzzsBm9
FBfzqMFB5Hxlnj0P46VowMWI1lPq4Ip4V44lMaP1jjsYFa+HTqD12cSG3GQguu1KKtUV8WMlLpaQ
qq3sEDFERetBGb8gKkZFwKv480F315HNFL5Prs4Ja5DR3JT/NdaicknowF5MxMjIiSM3QdH+U0Qa
/vbwW/ONu7Hnx411dPzfnrDJEosS/TRfzqVVo4V6jr6NBal6kUcrc/upON+XMigmYV3TiQ3vBCkD
G/uBHZQqRkqRp24PFISVW7v73yGIQDwuynL5eYYgoQVEgIKe/UW9TCrpWLd5TSsl8LqW8iKfgosH
PUfjE0H1W+aqLea/JryQ5LY53fHJzkmRpx4VXbTDLL4NDc6O3j64OseB/gcrQ05qkHJ6+ZNPn5fb
Hr+M7jBRltht8Uxki/dXVLZUIaPPY2VpR5cYN08mIXRkc5CKzvS+MhEGfOodvvLsMEiAycs4gbUz
A+QJq26+WXWf5JpQWBrHla3l7SuLBL2w8mXvGhEUeVGZ5XA+kEjJ3obzXVUJWcTXAbaBrUQb7ejK
qRFNA8f7WQNS11Oo1GXO8+WySvIEA/5YfL3YcIkBS1PbtOBjB9RM9fJ1k4ksrqnp2AWcf6mLGqPp
s0h6rtPcEoE/UWkFMgZqLhyX7ToGSOYOUrOCksAEdKU/uIII2Du9JsIQotdi7ky+W4Y75j9xAY89
LK6cu4gLhLE6RqH5LM7nIXv2dhTM2OU7iXz2KLP6YOClwYb+/3ClPp4Irg/LBa/GZ/x/QroQ/4Et
QnVd6l25s87WiOcZ9nY+xSz99FsvdFFDXW9EmW12EEE9vj6HbNM/8jClx62mA5PR6/3GrIJXUgJm
2HkI6wS3L4K6B2LD+y/7cpLgkKpGxR6uuVdPpg9UYTEpVh4yB+xBxD8UHG4pPOOYrPvMiATYJlSN
fsc3PGFEHmt0CyT/VhMnqnWbt2cRNYMZxL/lY/eLnwCAT4yO5gYqkMQzbze2QXJNe0WnhrNdFLZq
/9TPFF9AzHQSRyLUIt8lRqOTRHqEpogHssrOqlXEDYyvrNLW2IdF0TUiXM0L3YOzI+BTkoXBDr7w
730J3tLKBDYGJmsgB7lG2mZ1OgPXVLL48bFQBitbIVMKcXVJAZOeh97uZFcrSGT93dJgZ445yCHy
H5gUVBULMuugJiN9Sfj2Gdn6flwyRxKoTUJs8P2S6xAF6cfXbQJ0Y82BI4MdF7GpUgNYnvtIjjdN
2LHg0e0x0afXja5yjo35QneSkNw+yhsJ6q+jiBwVSaCX+LF0m6RO5kdf4B/SuVpkyHqd6uR4YkzT
1wX5sd5/qgFrZa0EV37CvqFWW7efHlAjVwBiutRdorBBY+UZ0E5BrD6tzK+Nc9ygpGL99r7FW7Bt
5b08UPgC8k4T1vHa73y8EDJx9oE65b3h64MqXzDj/IeEz4UEneWFAl+kfZ82bkH7DY04h5784VcE
fWONkg523DydcG1MBXo18pNXgMjBbKHem+HgtBGx93Spg2tCpjNCl8RK4D1Ze1h2jlQ530BHmacO
q5Ld21MHyRMzmi2oP3egkccba6oGXoFPZNHTKc+1ObCPIcIRppqM2dz2zSR5Jg2ldtNbx6Ui5faG
bMSbNvtpZHURxsNf/z9+y/R35mdstOJIhV3XlDxRbLj8pPJQ69lMgsUktOUHel0Wbg/NMKkhsG+k
EAAOFaLUtfa9smYTm5lybhC5cvC0VJfkHeWFEbikDj/9l5WAqGu2HmDmJ2PsJUOl184KQVX63OBZ
QefXPY30e6GslP9Z3+JDQDputcXlwypxdxhE9iadUZdcCufFT8jLqhV3TGtwPWhQrg7pNEgr+DRJ
Td7PDTTKKx6snPasRvr1Qmmjeld6j8wS/BeKgih+2kIVZmLpsarAxce6zgeosjq2OaMEwTwcUNoM
4lJk7BUp3MoM6jqD0h3Xvk9gyd1NTSQO5UHGNTr/waJysX0exLQddvo5cDdeBEanGLGzEfVONOnE
f2ntgi3gSn7GqFlMcjHY7/XYO/em3HBVzOli466rDgbFQV6dwv4ORMLL8hvcDgcSJ7dzLsx1X7DY
orQRQE3ODE8DBeY9TrYRt1gf6pYGvyG3RMx6ND2JGVSvPSMEWG+Rf6ghz7yKNXNHmL5UhYrF4UwM
WXAYau9k+gocL5q48JqERvnKlYYFZpf9XFw7ErQgZOUqRs0VOfYsQ30GJ9iVzhEYeXxQORLR069Y
6VGlkG8o2UK+L7fmBBD3rilN1t96GHE5M57n0GBRHXAlttrhFaRG74FZvWc3KU9gpw0QqGKIn98A
BN2DY9fX1XEWhSMJdDcPP8rKOyTrjeKrKNky/n9t7tuFd3epV3t+kY25v9+tVJYiu6sk3/xrVTKv
iMV5vTjdzqzwxvBgKnzLbFwP2GvJfa3DufOgV1vicrz2f2uCtvf0Fh60QX0lj6NEcpNzyjrSgBn0
c3xphdB7Hf5Vajuto+W9EUtA7rQjWUsZ95QeazoLRYfN+TAdYNWQofB6dp9ZxhV9bpF0jMTgvODH
f3APIminXmTaV18lfNSw/minjqlZJtCYX6iKkGjyrs943cyHfRvLD9xCE98tdGJJHnTUyaHEsHBa
NG5OjrfS+qyqc6tDN3Rd/E/5MnAuu7tAqnyo5IBIFPuUDB0dNTL8dx4PjRLa7UldfGrhEr/+QwWY
LFOEH0WNsyJ4J3H/+15c0C8I95ezi+/Pb/E10dZVglLo3TWULfj5SXputz+lecsfUxpcpVZMFbEx
pgpVZmDT404wWDeAfWyMLp7PrmVLaNYgVzWZo1uJIl4Yw2k6LO6sLv15ks1JHmaiYGv2CqDHl42F
0ddI5DcNvKtOYmvGcrpACwcbd8ScEIRrJA+NsvlTuu/WlLbFPcphCDWVXlEyKRESl/1CTD3XrKUv
XiuDdR2WL4Ezf+sJFtCCN9mO5SSI1Px7nihEI+2K3m8fsX98M4RZfZmYv1cGN04w+Hk/ClLgRjYR
6fAnZN/CcaYodcK8UxnpxuHG+hZkeCKa0OcnMP0ez6JG0qXxCMMR7Tlci/I22QmFEjl+VlJbbd6t
HqJMxg802NfASk7585b0zxBkR9xHPricdM1GBmhoVCBubpUCZ68uAtKVwywWdn6K1QHkWci73/Fe
miMC5ONwZDWpPJEUOSKgwKaqIRl2zC38HLhn3D7Dq50fYYCABLudfBkK38L6rVaYxDuaxdYfcm7x
A7CtfsTNHC8sRXdeZswLdsDAp7T/Rve38A9tQ093FQU+X7hCgr+2qJrG9Y+Pxg5cPw0OdA/FbzEb
c/BkJWR9UEdEH16Clsug99IkNXke2f2mhVPDFiu9y9UDxosA+uSEeY4ESiWXf+LP69ZgmkcWALlO
DSSc8PfFN6SjkNpwIXu3NumWanDsR4QZvoHQMjRNJau6q9n0NP//iAmvCiSLkjtfCQco98PcJCUR
KDxM3nbtfEiRShAL3Ew+Sn8tAhbUbR6ws8OSBVY4U4WP+1/peX15GLHb7nQ66VmYYFxKpyFLX1Ld
q9CTmn/0KBELVK7CZ/7ap8hqC7hGJbFQKkSD10osoZdCRb4G5lp0okW60OXW5QQi70kZqXkhWcpX
zR94W2rv0EZcitIVEnQIIANik759+ITxQ/AO+hrbS+MWT9lD2fatREK8wBsgMgvykA+Wn5QV1LLN
ux3JAWkuE/CbUbirldzAeuWOo7yQiQKMPZhSAcQhJdJOwq57mjWIxuTY3Y0Jya2i0KXIOfstiyFS
MaqvfXx0SSYjf4aTKv+jLvc8HqhOk2jZYwnBnCAfLcoldFIn0yho1zzJsuQBD3SpKxIeBi3ZED15
RKq4hIAtrPHd33a+BMfeHVLRD+CrkOJxEiIBDBLxiZ4WYnwtC3r3StJ11oADtvBFk+uJiOGU/jpc
Yt910kmrwaJez+3WHZTO4nvdQO9/LNgxkaTHbhpaW8tgocoO9vn+5LqVNV8CIGniwydCKgHJ/Cdb
3qM/zfDg95HE2R1cIhc9hoO7Y08oLfPCqnEicn3N2RJy/1d2Ju9MnWeXOfkbUIMR8HI/5McZ/0I/
e9AuJ/VZsiqlEqpqP3BXNggWQwwP838LN52U8RRJHMBpV7n0iq3IzWGlnkJdlDdMLQXgFDS4JONx
Ww0tv+fQK7SSAKvetLsOJ4m75SDZEuZD3YJ5KVdJcNfuxSVNvwzc8fyNUEx7nFreJNT1gOK+WpqQ
mS82V+eaPiLk+R+OER8fg7nAKUHehG1Q9JJLviAcGXYZaQggqqntTqTjoc1AXlgMqe7ptfrAWK33
nrUdc7s55MpncQ5yEDrnOaVjrdR8vkTV/ItPG9zDGVrrdd8HwWNqHZ6A9RL8i0fGlH+luCgohlvS
RkROlr9K/ZKUmimGH8Q8tti988tgi9f9gtehox4SpYfo0kOp5THPrf41UxmdQyP+zIsQUKDtYXh/
5iPl3wugk+jKmc/uOhncgU+MjWkCOe9dYcvo/USo67/DZ70TBBWdTCFsp71gxhVGXfVsYyUOV3iC
Ahw2EoSBuODKjjr7fPRPQ+RBTd7eagME7HaZ543JPlIfqQm3SUEni2qmL20HPWGfJji29RC9FDZG
Dxoloh74ed96Ey72zUKi0FwrXKr5e2AeeBEMt/GKHS4l8WRtwWp1DSkgNLuphuDAdSVReEW4keDv
nn0sQ9vfhONPynCACJi3/lFTzaadGEcskwbSpjYDc/1KSzRYsUjjpA7Kc6h4bFKk7Rz01w/yDVIl
2MIubP14/D92vEA/yyDcOhhm5TLiFF93/Czkbgi/Y8PWkdg5rasSZEDMgw8f/yVZrVK1ZYwCltd3
PiKIh7xhCCe1IKXWuhGhEHOcp2EONDe6563DO4TTXS8VSdFbtzcv57a0xsMhTgMJiFHgTGrj4Q8T
UjsRu1w0uJ/CJSW6NEpcF/2i/+u/eCyq3+gKoI3iWzzsNs2uFFulC7nEkHg/R4zkeTI+vFGG5ASs
X+NstPWEfMkmf7HR9IrYSePpiFNyU1FKHmm9wLpyzar50E8lLImh3Iqugcmj3gZCJHao/1xiB6lK
FezoztUGKUE8/+Im9EoC7943bnGMlbw8xZu4jdhuhzkuh27ydmU/bg3e3FiMcbAkmePvqd2/+6Al
U5WbPNHm/xT2tfta5/gWbcXQnzAWcMV7nKpFTfUAAyiN/DLdVBScUjTNKxL76NTJmZqgED8ot4ce
ehImeC4mf/Yb1HXIaIuxERSDD9WgRRotTdlsVfjfXax4IsPjavs4RXHDDkq5eOzNaE6b5cSSzZOB
tPDzOGzIctObkwjgB49oyV4wOGrMcf4dQkmHJ7V74hHfg5Sq4DUvOsA+WueuUt5kfCJbuhyPfdjv
6j+/o2U/iTD15AVwvr+dvN0UmK0hccffulTSi5ZvBAeMh1lqJDeX8VDuSY4FaDGtYiOQDAnlFIXf
uENuHIp1u8Tw9F2AbAM/EGhsiYT1w3+6W3XuM5kckVL7FKrtXkOboJsC9AE1t0gL5ukaSndmqRiu
F+aMI6jdKu+3LUCfHym5DOAi8kYs8hHtGSTmBvpSc/E21bJMl6dtfVsGZkBby9uGvDdfZLLYIu1d
ziyyxhzv+XcNOjYHz6gj6xRfJqywT+VOx0tdxoh3bKPkHZ22hgx/JBP+VCVXTQjkw4H1HZmB84FK
E2130/kzEcoTrjeunj7HOd4tuqJpknLMVqpzw7DgEOpVJCGdpzEa+ZOMutmAXteWjgkLRBJg3bAF
osBn6PZhwRQX3Aq+pFuFG5MXSf5+qlxVrW7HS6mjzJmaWUwFGah/p08HkkZbAq6nfiqScjS4ka7q
1JweC9byHWzAviheturPFQSKjmNyVYPVYPb7ywI7tm805GMQaIleV1VvmSJXx9KwUQUSJDqg9xu5
BXHfRYmV55Oj9DB0Je4JylgUSJBTMDBH5o7D6W58cAeGktaaNKmnZwjjEf8ORu+ZJ2adHo4Q4il2
EptWaywrZeg/uWfkChIvdrFY6+pNWw8p+llWlEVOMZ9wW742sG+5qvFAZDysFjIFdOjbzd4TL+Zj
duLpWeXf7YEiDTQPj88553SPmbYq4vzouReK7vxzAr5o4wf+83knGh8WlXn1zx+Avny/Cemh2pdc
THZ05Y0Pc677r4O+GvqH/ocE8wGMydHsxH0xT7enagx828z4vivZBaqLTy3BvwV9Z1gOzwd7PtOw
lVKjqj5Yrv+AJW5W3UzQKZ//SLRh+uZV6pPF0SOVU/NXnQeEiYrYqWkwlc0MAR9SSHwVIlX4B9F7
LAeXS9VkwbY40mI9VQPeBkJuU7l90EzZr6XlqpmIeAVLxImF8/Fp0iBAkUpffLH330MdzqsK4SK4
Yin7IcQK1j3x8B/GWQQpCNKEVpUfs4dqRgSARyq8TR0cI74QymrC8RVc+Qu58Z41sWEV+J3mGPzU
YactTgSYp9xue1lPSbE2RaxRdcXl2l0Q5yODyyPcTIQ7l37RmNLTeJ1IbqQFzSWB6MCNpWmtZZxk
/EyzSj5Os65t3q8WWAFMgqdthmV5g+98fEYljTbPkZiJQZdB6huxUT/hRSMDZeH76U9LqruXIxcM
nn7zPpU71a9fJ10JYeI+N535EvQjoVtX2lDmscnAcSVHZlTniNTy6aXxs3lA0+vvq7tZmokyNQF4
NZo5uYWdUmD0zfLHwJ3D31pg1bnTCTSUhXZmqFHj3sX88AxOWHeBJtnE5jAXBGp2/XZVxpY0QoAL
Fezg3ai8Vr39wxlRLmxh+b5mNVKPld6arB+cJWYeGxn9hK4l/v23jCaphB+F71BBdsabGqfc7hod
kYPeHQSjy67UjfzsHOkCHkAzoPVTelK7XRgn8ExMurr9UcigV6sQzVLAxGVaT5Z81fnLSZFGfSqN
sy4PNB1/338O9RCTDWi/HGU2bIrLVQfpDuIIYxq+xbejHND2xC+JXiGSc47j8SYHZs8DICpFPNOm
wrAxTuFFJQ+gDjLN3aM0EWtT40jvpl9FlP6Wb7CiRvSU1LSq4P03YT2HTcC5KuHcABPJrhZX0Ikw
44pKaFPLH8eZ5gEgnvoiGksqy0FAXWVH1QMYHTrHOLBHg+A0FrUxacm7uLJkjM0Err9QSjval0BE
9cvgDB+fc4BgRPx7M4GZ0CXe8+wLBMXwzK95jvlR3BfeotBkmRpvF4Bogri5gAOpOZqwC+OJb5HT
kZK978Nnq0UKu8gUKwlI29I+LdCvD/X0pa3N0WfOgB6mwylAyDY74JpMbe0pZKQ/oiBuT1R8gVvR
SWquksKnNJh1W0XTenHcrpIaXgqUBF0TSAd46vAd7piRV9dUGRrNuVvpxP5lkvinA1sSWs9sWgEO
Jb9J7c2DRljOebkAeSyQyb7oLfXloU32Z5UYZSo99rl6F6ka4elAkBxW/k1mnFhIhpt91DROVn4f
q6WxKZp9cNhnXyZJofV35fxXMstnYHSOusxtYOxNoxTiAi511K1r5TLraoT6y5UBM4dTvkPSS5vA
lEog0LfRZPeocx5s/yYeP1FIqubgimuf/KRrF4pN32nTcSe/11G5ZyM50PoZJQydtSHh7u32+rUa
Jx//3QEs/AjcQc23jyss+xu5zw8ZXPltIH1rVEKBPY5P5Pz+HMIxnMlgSPFujQWQi1Z/+Kqm0khV
RG+o/8JBrXKqzdyW8YE/K5wyPHCkYTeLPvsEZDwK3eBZgYEsasMRV+xmSSm188yn8dAftjf9HNFW
OqRzQNKZfHbI9XG6mxDekKrbZOw4MRUXCmMSdYEMGEUPrnOvKbbgT8+NAG6BcYrXTiBnnxhgGNPP
UPqEecsvu1kSxWmbXaDhBqazs3rTK/TzCnYTGvFi3zWFy4N24h/NAlD2H6nMya1N9Y6Xw4acrkOq
01w9sw/pEZWD8HN6S5r+/NoX2+eOWODhhPrITCTGPT1wvFbTYGVAdg1GIpl6ZWErjhircyIpgsLY
VW+Z7KZGmtgVxcbuo4dTo3OIYpQTGxoOfqoBm2uEstr7cbpsKdvNGJmWQv8ca/Klfv7EzXo6j6sH
9jHHtqn+vMN7fXzAl1KtLkytHLyOLcXwcC6PwWOHKo8xJyAWN04iGInNwisQ9e6wG2SOB6OMQUIx
qWolRVY9RExve6L+yNlxhjX/241aYm1VrD8QYEK4s+2CANMDPdFTip415Y0LiM2Glw3/XHCZejeu
a7xoNPryN9ZFduOAUvlm6eIUh3XaHlPUNvpcRjehC1POICenODLfbwrGwCboKlbrJX3JcJ68IVSR
fdVUoo95I+Jyav++bhSS8q26/LNCmFM+NQ5soDFwjci5bfD0wXavw8s5neGPIhtjy1U5rNDZAW0t
+tJ76sf/DgOVyZReE56kbehcjBtJPKQpRl5KoPHTHDHcoQ2zyd3wZl/o4myLLt8AIOBd1+6EFBWH
GvRT0vlvXTi7+EGDLy5oGVm0qq0dHy6C069JNeUpNJ+8ThorBVq2q32rSNg6+E1GIKoo+DdLJU9x
Dny/6ppz0aM62z8a/P4NjjosWUclbJI/9xZKguRO6FVKwZkbxgiCVv0l061tDh3H/HGQyCGjiRlW
hdonFNdnYxc/ybLMiy7IYO6TPlPrg9CvQmwBhrcN8xy7kTC/QANvD5wg1r1a+knhfdyMeu8coji/
TgTLFDRRsLrQ5VN/KxWfeEjCrKXpXPAI/wWy6bOHqfllCYjoZxXu9B+anc3bL64WHab0bGI89dh3
xGKhlZojRTHzGHdqJ+AVrle135W0U4xJDJi2CKOz6FGCmiJXS8nYWyM8e9F8QTJnwk1jxA8oEQfR
H7aG4YI+gUj59MjQE6LO1qKjtjWEtRtdti6XG/rEZhlYTU9PljzrwTLA3hEwquT2fxoOavBEQqFE
vJtrSgxCMxs1uhqmL0MT9CCHQKrRI3G3O11AON9JVEhuPtp/rogP7xID6Kr5+7DcYatsrcrmVkdq
DhhhoHVFHoqTof2R1fC2U/GOwQiI8tWUOAVmqrzCJmLkUiYN6IAjhxIZRdSevkXyJrAKqfmJZxmg
0522hPczbzi3FHJil1R6C0Huq+4m/uXXxjjICzNHsWkeuyBAMwlrE3+qycAMB+R3W+jl34HE94ul
R0OXFvipAmC0R3hsAn1oif1fC5aHyqu1izKojyRgMiA2EW9SWts9WqNC5xW/2uib3BlH0udLutYr
0GuwgKp41h84Xr1msp5WAhESFmktJM7XLWrW8gDQtLOXcOY4wKo90ZCBxzNgmfVgLkbHOU9V296B
kSWGaB+mj92cjZjq3wowmQncBlk5K6fLzhtZNose0OGysr+N8aAlXOJnlqiiIhxcXCZVOtPgDU45
9VCLpBAAe/dAjAfmnucrRWxVdVl4oyXRvopeH65k7XYhTDRpiPwIGNHlAZ8uunK4DqJaI/nobdh1
dPMpcQ91dnYTq8RfHtbRyzAdE/vBWHKZxpSoQG1SfZ4gqBoe2n2tsNlkowS/Ke3Q37vVecyE7LRt
f95wLsLk7jo/oO6g6DdZZfEYXGTaydxJHCZCEpdqpYxl+YbYZRg2zU/x0tQ0oLGq9IH2zL730Fct
B2q+SwnwPM7nqZ3z3XKAsBGjaJAAWFaqoFa0op9wm1YJ4sYqCohlpYpFm3M9dNXpKYgcmXjVGHkw
6i7x/ej7G8q5m3VyhNMkYZH8kq1wYfH8SPtPtWo7HVr4lygliLt9I/bHmFSUiMcX8hQTIQ/2fBof
/yv28AXKHgXimANuniZrXOOWRLrB0yIJxIuPl9puQOUpXtH729yp0roYwiVHDJoz5hy4aYuwytxr
8iCuHkzxHC09g1b+/rv89YsAK8FWocAD6w3dWZonnTe16duJ7uIUkIeUhgstwM11UdtDgjyjDYxM
SaoUHQtBO8BgyvQXtBdRJSz5/87T0H01vcu1B7jMjWsTd9wb7lUwtyhT4S2JO5cNqFkrz86nKBxx
u5xLPuRaI4UEE2fbpX7Ionenyi2D82o1Tj85q1/kNpzZb44RXk0mw8d6dawhj4vOhqsvqMGYFbKm
WXhltjtCwZ74/rdZ8HBUV3JtY2IfUgTKo7vgrDU/XDnI8w2kQh4B7fTJl/LsoT8kR9QVHe8u5086
CfCAyJi5xt9CyPS6umyoGuchLUVkKMyjGXmLQXKa/j1e7cjf/pLvLFdTzS9BWbF3gurnmFr4Y7Q+
P0/Z6OqFYnoufo38Ks9nMbqSBA4TpfRVPExDvfH50LMx3PL+IbwDdvBVjGxoAd1oMBRchN38Xgih
uJv1I/eqdyetkPrYCHzGEFG/B09NVRknYi+f238Sz33Y8/T5OPI/TAWNZ550ivkBfXtmEyGMj/zR
vYQ+TsnjZFaytVSn3vdiC/Sdyf8/2PRM+T8h9wSETaNW4/sJxzdCddtffOkMHAXLqNnSRAxReEaF
htl4gbqZXBJcGsIm1o5xfByHI0/ED6LMh5hdP08wdro9Z27uewEha5zvkXDOSgYNdfIi6e1DhEde
lwqJtwClMALTGir4rJbozZgdmiFGQYegZAfu13J23w3jKkdiKLjFGh81YTAEyRH4TAHwqULBL/HJ
LDeZFUSV5pohLwTpkMHTKSA+0bmZW1OFUvof39oqn9d/xvMF2D28otCpGva31bpAxi7/nHwsbqAA
HsMjKlfUK+b7xOGyokyxwxCqO4oDN0ae2SiKiTC//V0gaZB9wT+uglOOR0oAG8QQ2GgpimVxEBkL
G2qJfVgZYrbgQBGtHE0GDQV0rN1IV5q3CZ4ms7+yrb2uve7SGkGBgBVf0m7OOk08oi1hBjmKB2cW
TL3u22/ELZskD23QFjgKhR5+okvNX9L2N1WBTUH6yDor/7kPKBT89vpYgLOURDRgPX2O2IK2N+c7
8bwgjZhrN69KLMq7FzPXtZzZyOLpnZn/9Eq4c/x3zDaMJmFmo0OEM8UBuFpyII0Km4N2UgtDH38B
iv49PB5HeN2nNPAAV8mLmdyZ/diNec1XwmfPDi8dNhUSltI9zcVkksS6gJbKoREVlNVIQP7zMZw5
ZwyrbsgPUJw/+vE4DUsQshIAgo6u8ZJVNduI8OcNQJawSKzaR6qyamnOWo5OquqBxQVLZJFedOKH
q01FJDxOyOv6Sy37C6DnDr22wO7/MUGrEZvhaOMaUHZi7v5y57bQHuWLZMgLcrkD4fvIo6PTfJk3
1l8H4srgmuKMlTFDLRGsKC7VcM9tXRezU7PP3UbIqfv1aWPQAC4n3ISo5PLd8UUJtM8phFlEqGsj
OMFv0sR/mfJde9JAZtBV6CWIxQuOx1CfLbzi36ZLfUnBu8RF7EDligU7kpCPYNFyLqsioLHMNwbH
B2TLB3ARyxqI9nG6qyShXdGkOu+27sPhuKtz9vSzydabQxjWx7dU8Cu5QfWVZvy5zNcnTborjie+
YQ6SgbtsHlLEbxy7fnZfLX5EXoS0h2lRer2sxHZdVJaUmi9vyeLwtsWDF9+95nXp2H/KVmMuSrcX
flAXOjcilG2aYF0k0YUaY/1QBIn7OWFMM42SIN8zM4MsR7/0qjomqih7qi/vVnERWHfV3X3wVIqo
4eIJ36wTKxGf2P5QAyuoFBCjoPKuEuwZWDwGJpZTsRHY/AGs5OLjwnHzxNP7ycHxv9ucRHyjMKst
rvEC6H8eNq7+ijP8Koe6+EkoLXpG0wwf6wtFMDFMjBQSILqq39zPOj3PJCP3wq1SYV+pSQtoQMRL
0RNVLAMn3EWNdyL9Gv2jlWv4efsGHOSdXLj59CsiuyYvQ0B87x3zbgNwHJtkprKY7OIuTfA162ST
QTaX4F3RQIhT4EYzcENTZ8da3dj/EdqsAt9jLObsELtRAjdemC0zDUJTOVIZbMw2JGmOBZrmHbG1
f2f4zUXIDWZvgkUKlcr0ngu+hKrDvaoSBzkBOUoTiEiCp9p6uaDg0ZrFFyV901h1uI1QlI88orIv
TCXRuMpamGlOUKkENG7FM1UR77Y/WpDW4IzA6Vq4+cLpUsjmIYHYEqcDcxXlX5rsjnqBG3XxcteS
30vRrliM2kZKZ/BTpJfWTrUbkb6Y5hodiTRGM6diNV6mhh1rCjO0BNvfsieyiAyytz32ohuOI35f
PHRIzgWATK+GVcDzMS2zzqb2p+sVZBxHYs/4gAje43hJI0g9JV09JQaQDd4bKYn3oUIJYZ5GcuFm
CoUuYja0KpNOXnLa3FDAZaPbYFYyINEtkfXsgGLo/wn/HQvcudkV6rKbsTaRq3Z3Jc6vrbtGICgF
0DP299BO9a/lrBSDTHWc8Cjs7TjlIv8pjGiU3JIRRcD0vKxeM/+g0fkEouhBbaqTOqToYL7LSTEH
hDOfPP9MmcxcBOk+3/XW1qIfKf7f5k/ftUiJa3d05OBJ8gMhQcuH93YTwmZy7PL55COXPtEygUYg
/BLQua4tHEtqOdbQOf1XoLCBpk+pECSZ6BSXIySuncLoOs1T0RcfkM3vcDscPWRc3EDivnaNQqia
p7GRLBFNRIJLRxH6DfDqM8fP1UYzZiai0s5znczfnUWfKgSNsEbd0w0mqL+EnRSs/fkRlsnegfFS
3Tf//SEnE55hMcHsabGz8jNTfLXc2Z+Llc3Bcmw1OCbIFevvjrGkHW+M9Ixg4gU5Hoh3reIicwOc
+PNnBVbpZY3xTB6M6dl8I4IGHsT+C72e1Oitbnx1EGYi/f5kEl5V9PvxdRspVmDUPn0m46EAf6yr
OhOrxnG+V6OASsErmuTVGkeHggksOmA0DfQtJ9wl/9U24vIoV1oeJHGyLfvwR97Fo/xSfHtegAae
4I9FX9cvD6q1weOUaZS/0sH5qvPM2zO00KymTJvK9qUujMTX22pvd1GIM08WkjdGknmrD0ZYgq6W
CZ6oKG7fxSlhFdmd+UzfE7xqfmhmHmd4CQAat+XkJSOQ7R0SJP71dITEt4Min847Cwc6K7wYBg7K
OHupbdvxtV0/6VJc9QOxGjRKHk+jt8DUnDsLnXj4etzDi4frSRZCaLFXL85luxyXvy0EgMyUDLcT
1xjp2HFlp4aTsE3CtBxVnfV/ynIHA67aUB9ciWqqOVNisTdJH1CVWsXdUyhFaH0AkoHJ5Cdk8dKm
XJyHngMIJrnTqUa2wosNxCpbO0ILvN3eazvLgr//F591jCaaa0rUOqJnk0J3g98yoYUCygWPrwqQ
XTOJf1mSdNyw9q3LQsZwC78CzePJaQ0viwi/cB/cflKTos/g67ccnebvkxBfLaEIN6p77EsFDL95
OSyqBz8UR3Qg06fz0v50yJezCoOeGxvFC69T0t2u/5FzbnA5qZG+vlWjgDeBKxS/q79UST77TmUA
80jMsTNEfLlqqmtEs3dKs56BMSFX74QFnNzDyyBaKEnElPFgUY4onOkKwAaRDps/TK3lnRrbr0du
hWK2U+Yuv6MvYeELPiFgFDu8ZWTiurV+Z4WcfcsfYUxzt2VQk/ClgZ8FOXTbwTkwlkWf22rvXSeV
Ab18y/QMGfJdHxMzeEAenaLdXW3FIS4bI2OAX6rRxJK/5PwLnr5KetXxE+XWwGI8guQNpWUNzHhZ
CAs3pj5TtJDtkl1Ec7nxSIOoBZ0S/K/8BSn7ATYt6vBwgJg6Oy6yGGTPed/i8wjG2mRC0Cbu7ne3
MV1B6mXIvg2DB0iHiGQh/6XMNJzG21l+yqtwiu5p3sHmBIk4sFl/TthC+qNuz6BvPIXcp3Wvw9lM
kGWoMUoAkqWOpSxvXmPZj4296UR3gB1kp/TVySBFqcy41ZpcvcLCOs9w30R7zNCJs9+L4/MwPAgS
O9PgZhEn+dr8B5PxaC6uOn3GZg+M+akY8t57KBzmnozEz7Vr5p0oWvCKqlPd+MjQvUZmoMYISzUC
ocp879s5Y7r0WrvNPDOJ7hveSs7NyteuTfq8Jo8T46lzi3b7y489sjkJMxwkExekHGDHdY137Lzj
apa7CiClzv4ZGTTSDSZjZSjsnTky2z769rT9Eaeebg3RjCZbbdVqjYrG7LGA3LBWGXrNGsPqpjk/
dlTCxrkBtTYPLE7VgtxrmP7/wh2bTjfOc+5UnWRmLEdAsg2K401HYcpITnLHo6DBGWFG+2PgkpqG
GTfFt9uWqhsVjJEEOMSIKR6zI5k9UvC/KBjpkffeSBEQZPt8DDksr87bhoaNMSUUff4c71ANl6LX
nCsM4gXc7wsgoeUQQCGsEk3TnApc7Brxv2BC4fDBxY+ezXJvlspTecvxt16Zs6XLrVjGbo7p3T6L
ABROcgpVccQVnmFQisflijOpJJFNS962wELDc3Zu004UftJlNV24KYyR55ofIl2EK1MbL/DZWAX4
XOyA8QXjDNCT62+bvNkbHkZIbH7L59zVDe8daKoxWllPj+CnKULY0feVmet3LW4e3NtwqfvgIuuc
T2/RWXKa1nM1AsSUqqw58KDAUyNP8huRpnIMUQo/1KL3MRvGC9A6sWF8G/YLfnFoaOEMnCj425n2
D+upvN91gIuLGYp6SJv+rqNSZ6pG/nGWZmTS7Wo633LeP8RXpNkek/67391TkYB2P6fRJoBlHWM3
4oXVzwbyIsNu2vE/HyhsWRyA2OC+L7VqKD4C4fXyrQx0H4YdvH7tSKyJUCqUW2Y7wKz1KZ8P/VVO
QKfQeRN7K1/WLJ95NRwy0zzy87eoJEQuIGtWG8droaQttHnX/wtxGBaX5w6GJ/HX1NdrZ5Tf+QAf
N2c1ODumExj6idubWx3RSTA/COWD4XqMUD9/M/oFSN7VLckE8ajVvHqpwYIhMHjBVZ4nNHDoYCxE
roHxFwxDNG64RF4p7q6XtdjKstK3tPEQg9qyLOXY1Er1mqI1RrS0+nGqTFDmM0CYbnmFi8XUEG8v
L27HYgKlYS0CqFmEIk++ax37tXGvp186IHgzOeferl/HrNvKWsvtRQ/V3GXizLwFUPjGSu82PYQJ
aikLgKA16SDPNi8/3RcqmOhFRTqYbpopFab1UKaPZ9KjNHKA0w5jMHOI//ESr8v/TNcQtbdOSFTP
2VK/TjiK17qcQwyNiVKYVmjjXe6gSt2rO/ZDyM5hnnoYbtx+M+pHZB1GCadkJ5wbQOphJV4ffGsT
bcojOx3IfErfJExJSo6Hn1SOdwSaigI80TDX/IfYBKwIrlGT6weEtYmMVFMl8p4fXEOQLWFR+GLS
C6ZaES6Z06UWW5jmxHhFq0aYbAI9s4dY5kHsdlLSESP4QyMEPqvYdxF+hlpXGLvnNhPPNlmhNRNE
sNqb/N8aRBiaYkRH4+UJ7iNwWPn2Igv8JsB5HZI44HjEqzzfU/1tseVqU/Gs2GB+4udsgRBJJmML
7ofEsgLqRQiTfQ0qSpFC87sqNoj0NiJuDuJ162PI5az5iEomYd4GeVrseWZI3HS8u3M0Le4Gb/3P
j/3v6tFskfHrbBOVbCm7QAydLvhoYEBU51A8wPQWxoBRcd/aqmuriLc7XERcx3qYJCCLKi1stLEX
39w/Egm6db6tnk5qBz54yvfenSj/DR78XmjVM05d+DVk+j/tkMkpeoMKBRfKMqUHvZEifTr6TxUn
Kcry5OsjVcEOn2V8UPldHjfKq8Vbi4mTjzbnOZ7dz6wY+ylvbhT52O8S9MuJQX37QsNvECLcPp7b
fUevWPBsiDZczWfmqRTX+Ul+4qznEuYQowN2t3WQoMXilST62W6BR0TDZaPS616gytRCj3gbLotO
6IfHZFVAw/ZBztNFMeO54diBHUVlGEmjcVGVu0bRGPiun1qQ9Kfy0mV6KjnrPvQiurjnkSKCmW4N
pSpRfYtfUSyqJYI6ardK4ZGSQBQ5guaW02igy6OKWDV7EWaEz94U7TMbZpq1i5aCi7xDt8DLxgxD
pJ4glhxCM7CUMndtdN/A5uAvDe+EyLDFWHzEJ1UzRG5dIB8Cjw0XwSrIOBI6i2iLDqrpvuA/HuVc
hSZjlBxW/ElXL2e95PTGjQvdSNtUgl81ND/1eHRBNd7Qs+4FbgkKb8pkG84pZrG8rYhb5ay3Gstv
B1Ut3jqJwV3ZJRl4/f5552uZrfmrQcppv8DcUW4awyUYngM996xCUm+7fT0Ukk0bhvVEj8Edpb3C
eC3T8AuclhkcZG5k9jRnJ2tffqddAI8seZck8EBjUOkiVdYOknmnY9mMEbwkyQ+jtOqF7iKhEoDh
V5F+SrzNEtTQm9BqfrweKWugmsUMJxrIbdM04AF3QNu8WDoyAvb0Xfd7Fh3A2NbVEabRwQPht/NV
4A7hb/iJOayLz4itsZL2A9YEZV+bvgGclmZFvjSdfsGCTJOHM9dI+LvqUtCzu13HjG8TdP8pY/LS
YFwgkJgwn4SoOaEww/e4KwzcPWtlJJsWfoUEjzn+2+H1QWKxoDn+Zkhpnj5xLzuvPQ18U6/7ilUB
OS/6p8NsoAGKdAMYrRLgp69NZMxIWZpopkfLzGNB0hciL0wMz2+4qBror4ToC02drCiiIkxn0q5a
DhqErYOQwsGeUdN+k3aZJm/f7xfdCc6/NfTM1UB286IHtW2DKuYbFqwNZ6mGfFzV7KfyNt2xXKAG
RNjjxzogTDtbKiPyz10b49QtvhBiOuTV46oD5TZR0xjQ5zMbM82nhCC0A4ONLZQgttmTn5Rs/97X
o3Dy257taN+On1hJasglP7bVLzooom3pLEO53eE//RttEWiZm38hZa9QgMJvmEfNf15dXljTnbD+
BukxcOZHTZPYXuZC7XrvkocxlOH3229uDaZWnJi5HA5wYpGhReGFC70qALrL/pAeTrV993mjttMF
wXyMLg9U7FEszXYjrWY4P/qVwwzhRAWP9Fa23i+F9XlB+1UBMUFU3/1bUDxWT5A9AtF84HV0iHOo
Js//VsZwRMTqtjbuqJf0UW6YknFVrVDEhEqKu/I5S7yVUirlhhQT+mrpY2LSNwi8Z2Xxoo9dGo7f
BPqW6KCJaZMyK6qF/8qghpb7ralVfic8QtaNUnql3jkhRCnQlq6+V2uLPq3MtJlw8kqbAClQrE+L
GC1kLewdZrMfMRi0TmrNekIL8ATphTpdlO2OMIvZGFbgI9VJGCKoU6GVfEvGSx6K7Bogs6kDxBwn
EkBsbnsZ8gvYJxCsxLrnDHWcy5MT/sc8NA6KrMiqS4Scpui5XuM8NkAtg9AR+GkVG8uQnOATZrg1
ekmzkAGbubvEJxgGvv+BSqE1TPdAw5CwDcfU+lETDkbCb6V6vYcWzfIHeS9c9YEgsiWffNwg0KJA
X2jQBlSD1Sb49j+z9vMv7WqWE4nxvimdEFjzBHB/GF9eB27lriljP9B6MK4uIulzN55LLK2eOacX
rCcNAO57I58COI4/FVu6tIYcrXk1I/We6noONgZt20uUMgErvDlMeJU2geyMkeB4w4LHB3GMyLI0
H44BPC4u2YNsuHsqLzy5Lr7xjImK3+784I22z0cAR9D7Xe+h+VeEHXRbsKRQI8yNzAtauZPG3gIa
nbLWQgfB9sMwrC/OggkPIQYp91w1UW8p7KksoYcPI1nI3z71Y+x2T/DRupmbO+VI2NRMV82zgo1u
yYKxVbFE3Q45yR9SMIkSkT/mak3pmn/USk37N9lKO9bI2XcIFFlqN2NSKfL5no0ySE+K5/F01eIq
XRpCeJ3l5JZ9g1YYMNuPfEG2nk2p3D/cV+RXBTgm0H1Oc4YfkLdyCY2nzhlUMP0PWWj8sX0sJ1lp
H2M8mx3DZEJ3hSjT9HrYu7IxJKyJU6MvU6yvo0iKVAxY5wp+TEt99lXaaTQnjacDMgY15tc6yTEV
MvW8a/5lc3V/ei7A9DG4DB8nq2baYQUgf2n9qtHJ1e8/0HOK84G+Brv/5hZcKz+OHsQ294u1KsRp
JESMAH8Y1X07Zch/7BGWrBKiGWLK6bBL/hNec84UeWzhA31Rum7j71HubOXYjPH0GMTNxSJwB5ms
NmM3a+2LxmjYDxuHdj8D3Z/0hePp9sky57AzV5EidHNJim3FTy8oktRKXX3hL2nMPQo60ViwNcAr
iYzjc8NYDM0YdnZEHBhOUORWC4LPN9EcRdfKzTeVVw8WajSPLKhAodfm2stm5OT0MS9WGy4aartv
IjtD9z2KT3mNr25Cbo0dzT8VXcWHMAVgAvBndU0e1NZQEGblptulvjV4xl3pfj3tkyonwuRnl4sD
zcsc8qi6oQee6qkaXucy1Q7GlgsZSADPTIFGJk9yv4q/odvvYd30fnlc1zzPeV+8O0ZqPqhZ0B7P
BUx7gKlZ6PWeCxZvOkDVP8oPBfFaq3+BfBBbRhLavh439dUzq4JMrO7HsN/PI+xHfTPs6OteY7Th
D1nsX5cn792x5AqV1PV76FscNkHXgJ/Yxtv5YonfVGi3w6ZA61xDq/XgvXk9LWgpOF06qq2FaA1O
fQXN2bqgkzwzfPbJC0bVByUhT/aY5+mhOyWp6+y695d4P67MLxFBN69ekD1AsgJgdcpEHZSLMfSy
9MxJ8TIf/7Sx+unURiFkTNNMvEQ+NfWQgWfgtQKfHidryaCON6C7H2oq8Ve7GW9MbR+MKAY+7vh+
XnnGT6z+fb9ch8cx+KdHtzG9CkbTflj63F4E4R5JruVelyy1P7+nwvINp2HO+fDGTL+NQIXujxXx
txanC2nNf/qKhsANKYKUN+FOUsBiZ/zF4nngZ2ZRz1O2MljdAS7qol6+mGceueIXI2j2LCuP17bF
dxKNI7p7GfDVNRtES977e+dnqh15OqRlFh250j0mrVMNbitOz4vUW9NJc8tgrW8fmuSubd4J/s59
A9St7gctOpucmh2NusHu08Y3CPUhCHrFDLX3+sFPjXKaj3eCVbGIHbnDw60mGz4Z5KL9XJyGTZB9
6TGfflhbx5xWDUSxN4Mn2Jo50Ac9aK5xth9uZAjBPG8s3O/LPcdOTpb+I0+veuCGWqBissL9ffq2
eT38Zxt/UUeFJcXWadWCKK/YU+6P8IcGyCY639D+wuPgLRaEM3V9G5ss2XJ+qUWW6hm4hj3rw9QQ
DHSJcVquHO+2cyZ6QzZgwHquGsexL8ZSbl64A57QgFAqRV+xX90MQZZme9eqSukVnebPTzTDLpol
Zqgn5yBjxrkLWwtWLxAVaX60jmT1orR5WaxNKCfqhIhxH7584PBBPBvoE/fDdOms2F6Jhy/vCx4y
kGzVXO7K0+x3wz4J9MexoGZZSCnsOtZaK15MEPbyRTD+LHQ3nTPwgzY/pUk6uihNxPYFrcdnXZeb
6EDP4aqDLdAyi0pNTfFVCiDE5nAyKH5v4NLwEQizktpWXTekYOsS7+uWGu5+kyokp5mFy/+8ckuN
CLdurUj/nOy2TYAZhX4p9QyHj8+J7PC5h+nbb864qjv58A5w7Ww3+tGZtPRQSyaJU8CSY95bzYXZ
g9/+/+qOL+N/oioStR/cn6P614LpSyn46WNOn2Is5d4JbZ8a+PSMv8MuITUdXTewXjHwNR4JJOuB
ZKVj82PjrphGxQ4IuoHc6d0xSND9E8QUnjGiJC1g4Erh67qSgFTHAPVktTPLjKD9EGAuapOcNAe3
Asui3K0rnZFUAtSS7OgQBZvSjIMbE07wKf981M84IMT+8vA2aiMT1QNyQ1dnFR+HpAHMoxzZw1Ht
1K6zyvF7DXn+7cQXY8BbgR6PWdteJtUfwnI6BQi4euT4hifusMJjNg61RcFTMnn/tN/d2V5fehn9
XdrKey3FT17odqHHPwHwvVP5fGUfX2Zhf8hd0WIFI3LQK322FZ7r6FFQFKtJct7jXt5vQYqUR+rI
I0uxvPJUXesZ62NXa4SpSg39HYPwHgMTliuQhR0xAkKxcgXmtxgp4KkSRi6nAnCULIx2hUFLD5bG
8uR2A7si+RCmmcMi+3OEJWq+IDXtTbkKnRhPFMR/MOSo+1hvDdlv+JUaRGnV3JeQN3ep1rzRTc8S
AoT0vLv54DeSpLdZlXATYAQhlTh2NhD/zoICZcZmtoRvizgMuK68Udl8qp/jretSay5qLvAtGwaK
5mI8QHha+aCzkeUpA15cylECPbmt49W1hpPZ2kO84nMCUPjs0WIbeyzI5llguowrGjjX8zRsyg4A
uoVvDlmkmNcMSRrbY/GMYjtexiN6dP19tSk1TwWoGwgkSiKTpZp/jyjswzMHNuwaENyArbXe/OIT
OAlDqJ+WXXpAc/kdMv7/TVHukVnWuuL2lufWPvxwvx9ReUw6vdkBqUiMbbCAM181lohF2Q+nkZTH
JSL9siQ5oYX5MRPCNRuBZ1gU7TvaQeyTnt4GuPhNFClUmYi3Xew1IrxZgUaY1Aa1SjpSAqD6DJfq
aPg356jLlM4ZQBXk1W0bA/wPguhloGCbXWA3kD63pTEoOmS92fjkVgaMciIFGVO7kHjO/hMiO/Ln
We8/LAoNnoRliK4Bc9BoKX4tej7/otyiYk5SFRdgFWJDh6BRQc1A8Kj/O6173vgcC4/oR1xNT20M
7M8dQGalP5a48R6iHjR7gJ4UwD/kkl1qGycgr3d8JLt2vu4KdJUrFIjn/ObqdRbbCQPaN6ZXJTXQ
WLkpt+hZiKW5Z7iuYXiVJ2dYjC2TJSOxnb3sTchKds6GfKcmDEByuYVSced/RM6glx2HXK3d1Y0V
kz6ApPU3H4LoFiLSJfsKXtmid1AV9FHlBuFsvk4ZoSgaYph96hwGGcBnzbgCkHe8NHpiM4FcXzW2
wKGsPbMOH++KEH61NJUpFvk+QPMeMdLslkUmDE1/XukXLbTeKCUbjZRFF1ArO2xkiA1i/4i/6Z69
OdcsZpVSPCQd76AVM4MdLZZP6Co8j4pBkErv7Vbu9xRWJkiFRW4eO5giUusSqu1PREsqitlysgNd
8xuLzBcjH/BgNT6MRVr9Juw6xzGX2amX436rZWVLALHi5drIPw6xhMtM8BMWNPEUzHtJd6UulMZB
bNaj75TgeHzFWITdc7U46y+jqGsUvGwLte20VntBDq5hIUEPWJ+JBq0pGxUzd8dTbJx6eGrMCO4a
3ExNTeinV58mHhTryeeEKcK1iR0W4seab36ic/1cXLHw44jGXQvqrloP2iYluzvMAyX67j7FpIpN
Qqd68eaxAMs9tomS9XZn8lNtvC+62qj7aBqq2r8JiRE/L8gRgnqrk62A6jrLmkA7M67vddOvqkS5
ZLnp4ontQem0mU9qwypRzDvuxfHnUKVICkEZ5laNWv8xf6QDRR71yYo3BF5+m7FpDCEvkgIDP0V9
+h2MCVa20sZalBWfL6nr+SMntUB8fNGWNwXquQAdTt2fliBkeX4n7JKBI0TBOtxq5JqIcKjOVs+Y
znmNRBAD0TN1LD1jHA4ZdRcnonnjPO2qp9F7PjXP+pX7KQu+Bdf0CKEl/9IA0bR4ohAN+QVvCoZ/
pHsVc8ptAeNXMVYNrDdJlCE6eYhw3HBoCHHzzRIHjBWTOqyozOso2U7/kQfN0Hi9YJWu1Ne/v+Po
CPs0QUnf4q6Oh5ViLC0v8+7sAH5Mi9qgSJac4uAD0Icm2oTCAjdKIL/KAgzQmFxb2cHVBCiYC0yQ
4NGMdP6hoPoYn6tKIKEYtat7hJ7crG42hvL6JOrUYWqLv7Kkuq44NDwcBeXfDWKij+13jReSdhNC
sonXvKWkoBsgtcDpg1YAQBtk19wtE7/9AApT4xOeVVKH1ndlg1QP2gsrXsufahiYFvvPFg8sFBKk
UaGInKZetZEYrFMV+DBtZEAKPvZG0B73egSuCikJhqwxlORvYqx/yGHH90IVMMKEzSPNRTswT4Xv
CUrCafgfHdPAcsr690Q1BSCSU5PUVESgcOtv8MDLdcFLZYwDV+wftrkzm6+dlF/W3Y6MBi6N2ZFm
MiTuwrowWCqHZwhkAilehsI63syWBpgRKWYOoIpqIzN/YzW55BSdimm9Bay67tSPtRdZiOl9mX2c
9SSMfsIBiFPFQiVsWeT8bf2WN4Jlx4LzBQExgerRAmy69gDUKEn0USw82kUtHew34U7WdLvg+ZWg
zdfT45YNawqU0qruHTFMc4mRqKbDEcM3JQUZgwnLCCpJeI6w0MDeld3Qm9v4iwDmQd8s0cDFoeWW
Il6lY0TAGLzWDmtA1KPIif2/B3VMDZVzZJLDM/EMIha1+kuZribPcj07xFMGFU+5Whyq7XqDVGRc
1WPRnbP3i8GWdqFp4zSCb6Hu4aAK8eQ6ZjwaLntlWWyq/f9VRrHuG0HoEsrin9nxbsrcbIhIpiNM
XUEv4dNyZwgljptm1wnLGopFVsEaQke5u1s7Fr6kIlUqxI0jItFrayNTYXsfxsPz4yLfJ3dzoHjq
Xs7JCZCmXcWkIMjezKVr1q4c6qM8suJ0x2bZoMZtasvmj0iR1sdpD4itmZqBnmfEJij58LHud3GW
rYJV2AJqJwdFH8p9/jUj7PrdhXVkmmQkrUam6uNic5M0gC37sKZrFeYikjkCRJt9bvzhNmzp7C9A
dSrCETcpAtD85cGszV+/X8BCG6hE+Kc1SI5eO4IiH6XmcJOse7RbhDPJnuBJipWSOqq7u1rbb5bp
VrivpJ/4e6E+nHNuO4GNUnmNKriC91JEE7Qjq2rYn2WZoBYfMuSWUnGKFRYCheuo0una/BTAMa07
cLGByt80K4+S3PTlzMyAuduLKZOrodgy1yVxgyu8Lufku6GIJW+BoX0gYHYB+nSVBuCyfd2ebEiY
vBeyGtfWw07ITmcpQKm4+MFbzcHr6XKRTMUqnztNEwbR8gYzs233tuvbH16QFUtduwZC3PBawGln
xU6aclH2+pdx0DqLYd62cnVffPxXLn8OQsDDzGYwt/ryavzMh+FeqZEuOwynlQK2cfPAQgMXY0ab
kxwMhGrx8bIu+xjbN7vEeYvWQsGFQlgrnc4t18Xm+PWh5evG6uYaAokuvo6yR8T/mvO8+AzI9YKY
5xC8OOksicDigVW9p0j+INP1c1cqSOcEeBDZNXzvJeLadxWUrqs9EyugJ3iNfGrO4HurmVFwoLQz
Pv07CZQmNgF1425vobCkzyN4LfHi84p9xabpc1Oj55KlPm5ydVDxE/TGkTCQ81cfxLZhZgxbs6ZO
hNPqVckMPYAjdRdkE7uPuZtRVCuiS0Z05MhglfcdKy+v9l1yf2KPOj1jbfnB0dbyJgF8YjTP4VSw
3BAj5k4zIShvejTmSCqGNjO/YzOnYb4IoAipJl7FzVDTzrg/SrSY5fG44yfOumMzWr2jXeObqt+5
rnZc44AQrCy7ZR5gmDOue1Ynf3Ssghd4WUH3aSSMAdEj5bYROVv33v7PP4UA1ouAPMbjgB5mHthJ
wCOJ47JNGRjdT8aoM+1vAWsfMBA3dVhZ+GN9OZcJsEWlmEDHIlr2KCk/VLd7SdupVT/NLO79WU1a
2wdx6H+/WqcyfLe7/DII7CnMhqVzaRGHepORKRjAfxecr+VHt7UTIjPWo+ALqbaGFOsBiNUb9jqK
m8EMu1fs+ndWLz6UAp1iEb+VQ+LofuB2RXuJoq2kzQIEf+3cE2I3LdWkfs5qxe/XWHyi6CCe2IFA
lEqdmCEjPzKbcj8ANLJ3WoPlrTpKL9Lyd/VZ1A8IA7lYhZ0zyT1zQcqD6QKYIZwBd35Qb7iozPz1
rQh0UxRV+aK9NksKL/xaa07WT0iyBGyIeaa6Uzyg+XBe0a7fHsAaulUikNravi7U+a34buvr4t2G
dEb0LDvN8z9sKCL5m9nn0vJR+uKM7Dj/C0IZwUYWOye6uJH+qDtuvu0+luBvvkXDsw+CeKiSg31z
qalWpW6DI8qKUuwCQOiw99veFimCRKqVPuyapJrSxFiagvYxq9vyT3ogRPPbnueBfKwGQxt8oPHE
9Bi9UgMORF1KewtAHjv6Ziw2X+MHhp7JQCcQW6oKWIybn42SjMNM1duCe83W2FtuxN9uQy7jD4ja
kb3rOU274p/0PwTY/sTKbyfLXxxx3iqMFZqOGiUPTljT8TrtjJiCgf3OMZI/EbI9TyDlp6XYs8SR
jeYP684I/6fqHZCGfIJgCLUznQYTQZcuaogofIxtnK6PeMGIcwdMTdfb8h9jcw1t7xktQdFTwQMu
2a37Be8IQP1sdwGHckfYlkiKZSV1wmSxv00mHP25SEm2W5jGvJImaO237EYGLStbjkpW6dRDWNx5
IdBLgBcVmP8Lg+08pftbXne6NGK98JT0npzZZ78kv5xiajqs8c0DpRg3Ddj23o81DAMqdebzBVVh
3VSI51a9Oh6hO+NaIybkODaCSM4M3RBZwTZr6/veFl/aBpyTCYRFrBRbX5/hbAC/6EM3WMw8LtEc
BdVOOche8hM0VpvMwIM5ELb2CROJ5PNag62QEysj3hJ2Bw4pJSRB5aHUQx0s/eiiU64cZLGjid45
7AUz5GQRMDJbF59R4rmDVmqsQFiN901zTPKRBwuXKc4Ah3o407VU7AiYbc1oTHZASjq3I8F5NGh4
XYkGn8dtfR/+jzOPzEXxTGuVs4s8ZlqI14VXal3KwksMIImndegGJ8GOCE4WpnHsJ77RJ1Vvr3gU
7oEO+ZkK4yW4KUC1TcwCI8lLej6nNKnJiL56Mf/feGW5FN5UipH74RbSvGMEx3TjVgQwDzsPQMMq
mCntCbMIx/eO2jidphADnLppuFXF4nSmCoStdylFfG838biyymSyy6APm5O+v0e4FmckSWUvtfvo
y47pram7pIw5aW2nGOOAVhx2aUd6+JNsS+CGZjJewMvAxDcJ4QvyjxcIQbpkhw5Z1wKLUAq8JNyw
rYzeFBvFZgKd4Aeh/Fqtt6u0Ob0lwSAo5NSBb2qcGa18Te8hXZY877ZBeZEzMpTjShgM8ZbSrYtS
Hp9HcEsch3Fot3ihvBRdsZPyD4r7J6jwhXs/qsXid2xq+hTmUX4Q9YBkuhSYJuoGudq0L3GFtQAL
2Ret5i1AJXj0FSlXWZmIwikFoMHMfp3WmN9VmKGm7ny7Q906bFxkrhvl9J5J7qvc0CKNYD6sy258
15JWtBtAciGT/D+Qi/8e1C1xdEUomC+GvY9EguXU42TVXUXNA+8Khp4PaeZI3y3D7/nlFy0tjUBn
j2O8pZtzE5i/PrgTx+htDT4EmfvzfHBgzNUfunz/KX03PnqxtTyuqlGaAXExOivxenbI9+cvu8M2
iGj5SZs0c6d6kafMAj9VFXU7dcNp+kln0xJVXPV+YIFc8eytmLZSCkSQXr62xX8NO0wAA/0Tpgkg
LzuGSl9981KKFrDaTej61mICa32AbSDnEfzh/Yaxu+BXkGhhAIAWH/cGmbU+KMdLa2FtqT3Z4zJv
KPhAi07gBxyFEJicRIyg7xJ5AqgSenN7vtstJpCaL4Absn5cUq2eyOhQW9C7F/BkoxCEBwcJZZUa
081+8S2XYE8RnqZ9s7eu6blbO0OdhpkSBijuffAoO/jq8ZGNbkjgJHqnrY+LzQqsoYZStmcjcKC/
hloKBTCyDGpDe945AXjQba3mHcjiiG6snTiBRVXRc2B3xM1i2pQds0TiSlhHIsxVxBuYcLIWZhkH
xaFO0Yh2kuCMxwyWGxZdBfXprXbn3CdLkDtdMao+erem3fLj01xilCjFcwPj4j0uvG/u76yZwt4E
81b1ANx/3Aan9VBjAifTdHMW+XCmEe7A0tvBXwItMIhjQwzNcLHU2otjF9e115wVtJSQ5eWZnflN
fH8UgdJcxht5JFNZTeYBZvYwgNRwXFIL1JeE2+kCbEKGJKqcxIW4aCTclmnDXQX9qa40spG8jI5g
akhpLsg+UPfyz3sK6Yd7KAODmntgMpLn67j+Ml92y7ko7kKh28u89HczMJYwmq87kL77+0pDw6ag
ETvuAdhQMtS4GHjSQHb2eeLEg4OxwG6hkmpfdIXcYci+1aZIc00V6BdWDnrG/TyTZQSGi+3G+ilm
aDw24RtEscXkMruvQavWWzQqOQ8DP2yGRANtNoreFH561R5IUPC4outmUIW736STnU/lvW9kBVm4
5phRlYqaWxDVeD95SS5VMeWjPmVUUv23fAIM9ESbk4M+9n5zmQihcIaL1ev1t9GRxy6SQq8DK5Vg
rePG2vo0+sTghy+WTKqj3sw3yOGhr3z3OSqAAAd72/ebeQASR3MLyDHNS2wPiO5WSiSg0oTh9r2J
I/tp0zPxTmqOhLVNPgo8NW8JIK61cCJ4yGACwdIUxIF6SHrAxIpi4kvuc+OyL1r78KTYyVXF8H/U
UtMe5Ze9U5RAJkZS45SFRMsowLtAltM+AGcM8N4+x1UFGEeAD+NVdTOZRWE92x1RqiGSCujDpct8
vx2FVc39pH4GQGn7Ly1vp1qJexkeXWdMPsDOAaxpf4/EHADEsgQws+tUBxhfW+Zen+wZGb6dyjNa
acT2ZXCO5y5Ugv6zx4UW9lc3ytbO0I5SHXM6jUlIUQtrfgDadFa7SV3iSL4QXRMK2ZjQBPbfiLSx
o27KrpgC6um+/gcDyrrZqYTi+7d603lwMn2waEk1L4tTM9kDVRUOjblgNnEqt/ZNhguWCx+ADL6w
oCCtPx3IHBHyHXrpdXnA2oVf+B1+tZqRMyiVVlxSsJP37MbUDJBQ92nRLZQLZWiR13hQxpEzZ0ma
JQj3XMOQArIPEkBmtneY8PgTIK8pvSLlqvejgVqxOeNuxfesvN0+FxXYF5yhYoasP7HI9SXGie8L
fVepz/LIR1BDB9kHW1HG1OuqVQ83iwEMwZtMRWZNvQVloaZux1jsEriFJlhHPqYfdeIsNiyLY7J7
6wYCaps+oPz5k49L9d73gjjtxa5B/06wVA9DQVsiU+j6E/J8fg9xmIdX/z3peI6zSiXzs46eMmld
yekm/Pt61tl8o0GzlxdKWF200w49TtJLmKNrofdCP3f4PjOs4f2rqAn9XMtWQueK1EB9HXnmFvqk
wNRNuBSafoYf83rD4b5gapNPObhvUr8IX8fZcmRlNgrpn3SmoIT3yT4G6KEFeS6FsCj0SrLRUdcv
SREBxD072uQ0CTFgou16RnpAzrydsIB4p8y051qHsNWuSzJutMCsjoLCm1hPvB06kNhLHo5d5fqK
OuX/IYkf67FI9JXEue5yElfj4ekk47lFWqNSsH3bT7i4FWaM3Pw5vkTpHbUPO7tmoMpS7dCjnNda
xI0ZKbKqOHE5Hf5xMrpzggkFI11oTH+/wzOE38bK03IH01lYx3i7dJMmYc8m8NsTP2SffkOxqQqv
FU6B1J32mt0SO6ShuaGwDVx+dbU4l6ScGbLhERnjEtEC5DY6xoskNiUMIpFB0G8J4Ysoes5n61Vf
WB6hxOjzqDMVVwoh++VIe68HKnld/BfJPRB1BfPg2CEz1uMQEtorXJo6fweAI45s5lhhT6PNL5Un
D09Tsqvkdy3Rne8NNtq9XE0D7TEiw6nO0R34amJdgwB9y+2hIy4NgzGU55SbJsMAR0vJ/MkTu176
q06WyzeWpn54L2+xxriJUXipIrQrv7PXVtdkISrLGkuVV8BF8tC97+HiFh4uM8MyI/ZN1Odu41wN
V5J3330Pyd2uI+1cboTk0TYw4J5wpS76aiJ3DFcvIwuJCxiqglqPeAKNnPNBZ5eZv2LzGqUBOWak
/t3bVr1/dRYahgPSPXJxPLNuCzCj2T2rWp1el2HhXqvczMQ9YjvsRlpBnTFBBtk3aimW6JdroPKV
hcikI919muAm4iVIZ+SB/3fXXjiy9cr4vSf4v002toeBEOryKLOc3bOGIA7S6d0YRhYjqz9RyZGi
hcT+kIW6GNwmqw/yscW09FNugajj37kxoiUOJO8WBd05SxU0aDVDkDrTY1Cw78kW6SswYEXGFNP8
1f+yj3oVOv73C1JA+gylfyVPbf3aid1wcP1wwJ+ZHN4hqFOnVFAMWfYgX/VLUE8Hch+5+20g5oNY
zTabM22w8oU9Q1eaCh+7TTl56/1MoyzrhK0oekWSbf/VtDdQ2JgZJCPan7WjZI8bU36CbSJZrS4H
ew9sE5wqmUVDPsjSIZfZr3JL2exy9IxnmOcSXskkk2x6o6tYKucXQfFnCj2DYpL0ohZRulAdqPWa
DChlDTIVrojjX8s8Aow3WkYn5tHHOdrWQlJhgI6cn02aeo1jzyVx1PWWiAgcWkztzv3eBbe3T2PM
CelQXrz5/BA1AaWeSzFaPkNLSiqYjvGYVkTdjsrwL2A5GKm93Av5h+ztoxvT7DKB4Oow1/LtklPQ
mKjtRN7fGIAkXvFg03XQ6pEqtJOSjhmbaitcnQu6KeZ5bsZqoX0ZtUweuPdAymWLvEjrzWmqL148
lW1wnZfUtU57HjMeV9yvREizeA0V51lds6x3V6QXO2pWKoItir84sSfJkqYSIm4XeyFZa8cPSbZ2
TGLH+jnxs27TpafxfIlVUAc8fyrWfp1HsecYgPOSB7OuQCY85FNsfMqJM1SlSkk1PjOSpdGG2HyS
X3WFj/T9n+8hbUCXqdMXjwPgI4KpJO739ONCkoBA/WLMFIZCSdR3qFtf3Tdzft/rpLzT2STuhOcT
YDzm2Zcdcs1yFs5hzaV2tE+O3redOEHt4J9qC/7gPBlvGjcKTRzIKVduyHXa+xG5k9FmVLb9x9/C
l40Tp5YSmwaDj9pd3d37b3BF73qV7g5ZqGV+q2ShNS+2bKQv4VH+Q7vVa2p472fIYBkxkB/QzlHc
w+Bx9enqluA41lqXdj/51ISL6/TOhtxIdoVO3xe4ALYx65dwBPEfTttcGP5kL0rClQoaNM3Ygixl
6CChxakNIXjeOBaJxQL2UJZfl/NYfPH+g3BLwxcUSxlf/BYnBwquc/sxtK+qJtAvn6XO8N4YF46p
petDE+fkYrsI2FvECAgP+rWiZSL29Ih0R0tycR/0z7fnq9OKOtNy2ImtAbMrCKiDaSe67sPsbhvd
xNbOhYJWR/0IgOZywp1ZT+HEMvjVtNUB/QQZcHjv9mx/BI+XwnVVqpFvkp9YZJIQu7uMG8OMARKQ
oCZiXEGTE9EGS75xn/LqYnQLcopDHJGMSavpFOe8bGhF3VNRkpHZAF2TBgFu9zO+G8qvem7z3PvS
tKG7+7iihcXmHXPL6tpmLgkPv9IR/dmzNjv6byGxkxMncqe7QeB9c83MZpYrots5ZNM7HGn9r+7l
P6bpkGIMEifvColnKTGj3QyGpdeAGmZbhSQEbXkJGxzDsIohvv0gbE7LWOE7o4oKklaKEontb7Dg
71CmJaxpPwh1FRH4iKW9U67jDLURUSlPSzaxhZt5+csYqXodFtSfc7PvcBppJLuFc087opyyVZEA
hIptucecf5xvXkofcNQtYdvHmjyD/rn2ukoHoeOjc0RryZSB3rtb+qg2HAhysULzFolCNF3vG8LS
afnIWHEJwiRzHsu6nPBFBhApQc3rEfnJCNs1gQq6+G3CExYGTV52A6P2QGSD3y63lm/4twMjIjya
gkzaF5oexkFXYhKwhK9w+G/GTO0XCYt1Sc1CwCjs/SIWC0RTCuzlXELDwlDr3Bi/hcn1/tsNHCCX
yT45aWie/Z9YrLM03tuahBwZckWenaK39nY6/9YmGbkuyh1ylErv9LWqazXwOMFhvNmfnxpTP6lh
xIIEGKORXSNIuoBGxE+OnrP0YGh3qSKEH/pTnNjac7vki9dSkhKVTt31gQHCiLtW6B7cvhMuaJ9c
ojC7Vmq2Reslgu1zx/Rt0BkU21ay9RWe+AUOUswzGjAWnNRkTXlyWrpj58oof5suPYO0s/+pbpIv
mW/NJAG7Rbat9z/1bF5xsXO1IhEBlU+Z2WHxkQbqoKhOOyIjT3za1xgEpu5ld6EB3zcgvglgmZZc
83lCdi3UO3APPPwTWqRGrTY5yZMuk6M7Pcmfm8ROzczSvv45Ppfii1NJwhYQ0Ctgj55fEJR1zXVE
5gdEAzcaFJFwOD7UHB6dVpzcQEDjekRDodYuSbgOzyVa2VTY8mm9eIKZHdOkUEhMM4Ay+kljn4/J
hgzfU+MdLq8iBQD0qL/rK5K5D7MpMnckSUHe133/Z5xQ820qryxE+oBtPj8uUpB6JJbskq1hsZLf
e0mLW9wOtCJO3C7f4izZ99dLQwl2PJpQLuzIfKGxrv+vA8l4hamryOGzbPL5pHvaKQMCW29Q5POY
8jTmWmip0cV+oYziM+o/HqJkZfCOHXV4LpZ3Z+HAoapu0lZyOdxznIzOqkQ5emR775dloml5FUza
hQBVk66G70H+TaiGDyoEmjALmiap0KxFH8gqnOFKv00eJnmDdRrVyTlPZKtYUgIXpGj9lBaAqJQX
RNoRwYPPLHSj9li5ENfwMDkywugGJGUUlLICOkVCRQEAQ3J+fmrvXLuHEJPqv4JKAXDuBQWzJ2Pr
ZVSH7Gy20f1Xh3tMkDCY79q8REChL+JoIE3EG1BvbX3930ww780beuzPJ81KNoOdb1TqdyUjE9JE
Npyo2ZpI3m35uGy+n9adksx496PSjFU6zgI3meSqZ98L+pz3nSaJnGBPAkFaAPmmHJbsOJyci0h4
3S5Bn9ruCYqn0/g+Lf9ruBKIEPQa+7gTMtcWq0CjwSGTt9tpvxXtVPO0d7VrBDEJmX1svDfHeBht
YfNnPrvE/5KSwHh9Rravf2J+Q2IZ0202+bFWI10mCEcrdXysRCaGpsfN2ObmpDUe0JOVgMtTxIpi
UnhG4RVa5bnlXmo8mp91RwZPXdRXzYHaqwv55M943kgPfhfdAwsk2IyTxD8qvXMdhENhrx/zjVU8
bQkCSWb5PJyDzOZHOI7nNYmDb+gF8Jrnvf0UU7hURtH6ARY0jkIaLI5eoQdIEM4nPhhB+MOfOQjR
TfyJ9gqRVV+QZqT0hFxVPwQBeA3C9k30mDPRoGyjB1Ub0aaihhp+pGUEh3qzTR725Laj13O7du7Z
/XLiFzoC/svsk6gNkNDyLFOJincQy7BBpiRSqMoTNkmee6qG+Rq3BaZ4FDp0cGgGyqPYxp+xAWm+
FIq1L04+DsPl2VzgWCUWgMwXds5dpCLf/FuNl+zluv/7+rFrvD1S1/HI4eVNeiubnkvasiW71kCB
vJK3G0KQKqdww+Dkwn0j/MVE+vjBkVLmD07AiLrqrQGkK4NqABY4IUmXXLnlNoow42dZ2+vbDqdj
bo6kPWn6DpfzvfIIePbst1krfZETLB58ffEW/wfB5MSsWJbaV7knZzAOxSfxhsnF2jYQeTMJn4m+
uVvzu8lzX7gTUsE4zAv0pMnQFFVNUvdp9xMuBYQUSzcIrCxbECt465Ku9Il2vNE7+qgOswj811f6
/zlDr+VyY9SdeziV4FQpq+t8HB08oIor/WEzj+Gaku5ILWCm/GV6vTBFw2TiW60LXLgRaGZJW60W
qAq6r4NFuEtlrS+or0IrWQvFfyhqeEdKpeWCnMJxiEVqGqUw9fcs598GuCfX5g23I//arnr/aXPz
TqKo3KpEbfJtopdrSJdQ8XUrFRGYu1lvNomcj5kxvywHSMxunRPlahz58uSlsoiXH1ZxueGZK0+I
HjlpBYaRA5s8d82fagfW4nXLFWVKZIDvrQpjZidapHpqO9Grs4QCuvzaijjtY9XMMGJ4hDTc4aqe
3Su16OzxOmKnitGmEkbzfxgh33CeyGtRux+R7lazGpE6EVUInptGmy88oCh/HTyM0xXpFa/sj6QE
gzhV3AzREv86LH5yuHiy0frUe6PSMVSRNXnpgG99OPBeYvIt8cSCHu8SzsdmoxjiurYwEjoLBHUm
D7tSYqxIu3PS1vOwgDLWxQE1ytYk1mQdLbx8n+T+FzqWG7jBk3GuQ24hFQfkIYblG81ZDBw0fhZD
kI1Uka72zQqvtAI9FznSW3h7UgCVo9/KmXOUcUiz1CEYXhAMGTUKaK6zwSwoNYK74t/+oUnohW7u
nF6QmijYVA9h8cmvwoTL+Qyb+6PF79Z3XUG2pucJFr6eURJLfpH8RS0cfI9K+F954zse+CMrFBW3
GqzkYySYeW+s84lRbVz98x/SiXmkGcROgyFhcV5YANPD0Bfefk7/tvC+47YcgHRNfyO722bqny8b
Osfh9PTtdeF+l8xv0YZ5HtKY93a/N992fzUDK+5f1SDre5S8yXP3eYIvjCOnbavX6sn5WGp62c0Z
1qjrsEq/8omxvrF/HKxYLdmfbTt5tyV7bqvRmOPRqacYH5ZGOgKW9G+Q6QIPksw5MG/upByjm+Yb
dkuFth4YejKNLDNT375BWfPSG/XIJbz7YpC92eRezRwZnLsxgPpvHw+FmKbHE6V2nbnCAbVgI+1s
0BEcDZoEzr0IW64V1sROR8mOhw7sSE7W3Fps3qp/t4XRaNLesh8ILi8Y9pgLeB2zX44TKFjG7Hor
nCsZKliIlQVQqCR+pXj6Vpe+7aqBvcWHUl/CiQBtgcTg2gqVr0ijZBmodVxwGqi3D8YY6Of5Jwry
4DjEB040tTV0KMGYdJib1lNoZZx3D7dfTsGU+VO60xGbMDzUSJ+axVwtgjiJsLUXJyIksxBPYd90
gfEWIYT5H4Cmgz83QJZOAy+3GD+lLzRXsjDaoss78Ql3n5aG02vypc2ClJkgIWEJiWVFmQDl9mJx
v02wgWRVGIZSv7vG78BedDcTHNP6S26BkAad5QvSs8/0lPUUKhoWUa0x5qhV8s5Ydjx9V3yJ7ToV
teJLHNtM2FKRp8/gSFk4LuZDPER03bYkxACNC/4h7Ff3clIYjy5Kn0YMBuEN4ASa6lFTr+Do3thU
0p30c1YNXpLt44zNa8saHDDl0t/XQqMLKUgp+O8YRXfGLYNifiOhSNQctu5B6BgQTRzbLciyR+ME
BhnvO7ReEGi7vlZ5rDjQBduekTK+0d/jN5w5jldNkuLIc9+h+Sn2zHJRrVveyNzqHVN9Evnm/ol7
wG22FzMeW267lkEh1oTw212sYqDKiX/Z3WxtHYuLSL+LZ9FqOPZyQxdFuImt0nIaueKzM7mHwJiu
Lp+rXjanqLLyOLSVjoFVLPpS5XvS7hf3IUF9kGRPgk4eKwwVoaAna4U2AGoYVpsYhTIFqtvBOf5E
NkMAVpycXUTPyznLBtg0xdPPtANNzcfPsFIM9Ni8ywH39PYTT3lTvnhzSXGMS5eT4qcv32Lh+8uT
AtRWq8SBrhcfX/tk6V5/9QsQRnz0aKYj1LLo20R5hod4FUYDcILR/y5I4aU7z7CcyL/b98c60gi0
Xbvd2Ipwj40zRFrhWc9JJbEq2wSLOe23e6kJsqAfrT28jASXl/kmJZ0Zm88PYJfPRKWGJZkW5ABP
mAc+iid8WPvdRTzdMmLE89z2oypW+jRxC/Z6SybQM3AG9r4IKn9EMgGu3F2rpHKNVMzGAdm1AMbY
UqnfDG/Gb1ZSViEzWa5644rEI3zBoDB3HHGj4bdLH4U89tdLJU41A/nxwm9qGLtdQPAYVn9Kf6Vd
7YjJeqNO9p8PbXZlev14FZ9M7Qn+RNSIxufNNdoxlSsjXn7JnJxzFFt/kzXNpZ+8eQP0mKF9IDY3
/404hJb7pU3Sd+K6bQlIccefTdOskg2jVq3zIYSxONDXLxe4BpmGbQubZ34Ij9JZpThvpbR3P2z8
0PJEkuoUJF7d//2ngFvlhW5DOIm83LC5a7AN5xz3Es1RtsfTz3uJKU0F6eN9H0n+b4WIOLYbo2va
mfcf6b3kiftnB+Fdu7YC5vgjT4NaVFDxLQ5vO9L6hdIEWqmM7lHemKpSWT1HFVfg62ZFfevu1JCD
r/RC+pZx9ukf0H86pKBXn03C+z8Zgk+eynGTyRrCNRFpHmYan0CEin7fg3PTs4+yCARgesWYAUDM
nFTuuXj7Q9qi+ru3zWxRE0Nmz2acspu/Yh7N6ibJ6+EL0pu60XOEHgmM2F95s+lvaJo7zJIEkhy0
Qnv3OJkD9rSjWC7Yd+axB7qE6+QRxIXmwWdf2FCrtl98k2CnX0jl1LbzkB5wCjlvcEyZl8Su5y7A
XqPT3H7thUn6XGzQ+KGbqVhhXW0PH747cDG/lMlFHEQwfPSNQsSvmK0ZO8NqUodwDhlWvHcd7NFG
vLT+JbugAjED6+X4cmb+yHwGke4ZP7X942Wh7Bg/0MZTH4XKauHPjtP8cmrseuAPHwbDQLpxUEBY
jK8C+Vwzt5LSG2F1NjJueheXVHwCt6Pn0TxBhfML9FuaakiVQkPHVa0VGKqQxM0Ag9UzJkGYd3pV
vTvg6BdYXBt6iXsP38fKwAX/eHQr+OP+B9VM4cNjfN55BnccctcK2Fp416cHc3JimF9iL0Rl+MpI
0YcUqbl60JVmMEch9AEvfBRxAPAiuC1Q6U922GRw++EWJ4Jku3A1BqnSW/5XTaXAgJY68/ikP7gd
Hvnv8M+zEtCQ2jNQA3CnOUSjfdJFXJCaQGRRzrQKnPWrHEBJKyotTWOpBDs75VK7lJmUUkbpCxrK
qIFMGrjqetBo/COx2WeTeXoGYg+83TsnrEGfCifaLHuMk57HpKHoJzHU1VT05FWCno9YvebaTL4b
jJFKATZh99BI3ID3BYjB+tBnLFVErVRUCnxNAur++fWKuPX+AVxEi7Lojuz5PChu+ALNIeG/RdsQ
fwCUZCsxPnweNmeLrMKHiKaLt7CgK6UF53day1kraeluS8Pn6DllKbtbUFEyeg370MDV76fvVjUV
p1R84mNBHxTtvTHzhThGAm1j/LOHJgeWhwxhWaslH+z3CyUpHRT+KCQ5TYTvNYmao5iQsWpKd69T
ihmXm05y3JZ2ZCpwzrbm9wbJDYA24P0xs7T1Aj8UJqK8v3qHjmrX3FpEBmiILGEOir6Yghd+y20L
mWMnzrOcJA6klRITfxZZIb6ywQ02YUqmG3lacFXLidvQSQAQkDqmEUCBTVXzDhBqJJnPuZr1N4qB
xC4mSDZg0HHBUJ0xo7THVozdHc41cnKCqjk0ZPCWq4c1UZ5QLc5BHMRrqlFkipWsnbZM6U09au6b
6pjWEtDJUR9gv0AsyUNIOpuHGkGS7mjJf2nUHc4zzrGJxoCkfeKmLpUKcxveuF2kqznPUwvRPVlb
My/IrXew1dQEDikr9vucqInh8b8Ay0WYS2y5+aLxJti3eM7smmYbD3dsOzlb2/hnkBklQ9wE27We
Lva8DpCLr8fHxNMRh63mjP9goE4qykXg8cgYhqxioEzHaOTrMKGvs7a9EsyZ4z7FKaHNNSE9uXIc
8WJtvl1mx+rhhvnw3SexCn0w9bXxFnJlYf3HSgcFk60qBtz4jhAbc0QCnit/4Z2psxKU2k9pfJHn
MKcixoHT09KUfZSLh69MS1zLRpsDWk7qm+DcSkJhZ6Om+028udhVM5FUPRYbgn1aQsWA5VfGFcEt
f9b1Yy77fUvt0O/PKZtoH3YSgmCyxd/72cxuOnnC5enm+h2oZhVZboAhC2j/jFKhZvDR26VqbZa2
E6u5hj80NYgmvoM0lMKYXW7jQczWrQTsWnJI/w43rjav8I0dAxOxtgy6CJEg0DAuIf/D42cLLyzz
MljF1JpbqJMMwDmG1OEh/+3VCGVQKBoZVPViFG2dG78bZUZcnk9YdujT7mLS4fSMbvj9fGh9ryNK
rT4TRA0ojryn8UtH6xtvsnqqpvn0nq32F9lkMoNwSBrBJflylyoWpFVoJgAIY3kWnPuwdckHDPdX
Y9IUPfd+tbmLr+4TBpKieLy1fLMhLr7Z89RZ3jKneGT3+6WF0L4eGK4enVa+vJCKYXuV1hJvOAYR
OrJil6Pj6pbr94xGUOE1SFPs8AhuNx8BBCl1+QpM8Z0IQK68T8oY04mutXZwzwcPExxH4ydQq2tl
JiCZN+eZ20Xqr0Gua2DN6hzh1+Ga8wrXIQXCAPcMTWE4Mo5aEsg8G87592M+8PPpNb6LoGgnnwS+
Mys52urhmBWsXz3BIEgq/eazhZ0iqVHMS4vUTVsu4hBYaXimh/7wNjHghmUNoUaYYrKl6pALlUPz
np8Fvd/PSBOh8L0MLOy0bOra7tKHR/AB0HPPoSZBZHJwcJ5k04+FeJNxqoQF01MuIyAfyBYfV07U
KpKgqEBdWsHtgQyzXCnZCJHnufzqn8AOhTGvfdLV10g6kfBLXKEC9+by/bs0txcSIYXCnN//LWHd
dzAdJFz4GPUoy9Eu4jjtq0HEyau0TE2DMDHuLnYKBPCMIpU9g5L+Wf4yD/3kmU7G47kYF3hhmOvN
MC82JuVgCuXoZZccGZ3RPvAjylP06c2tYGUEMERAAYikW/UiNH+BTvPvRia4QIwCfoxBPhd1vvpb
FvJ2BCJ8pvy2gVDnza3yzuwZNGtq8DdZ9KiuKQ9e5LczxvkR6rBHSWlMxTBiAyg5LANiOgtrSB8c
oj0nuIxAi7Uw8qi4QQiDjFrvZBrfS0WpFYce6Y1XpspyevmcEbJgYQXRG5TSeWwf5OWjY0EOyitR
9Z+nHgeMXYlqRZEJ16wTxOUWvllDbFmy//2L2G27OvsTiEPv1IbegPAgl7jLIpv9I4BWj9sRWdPz
ktvVKGlByIO21n5mglPcTU48RaLPAfpNZ5wuTnew1cf5wtaha5fj1Iy6cl7qjOY6vFOmQtDMBeBm
J46DkldsJoHMYA3bPIrwu7f++8pmAJZm2irQhji5SHBv+vn6Imdnlz54ZCem4IobqD+3aM1R0OZz
YusPint9m+pFvWZgdKXUDNtP8Z0+8D9qozNhX5kYZrK+D4k7hJQM5PoQfn6TBsR2pRHp8PbkQ1LL
F+b2GOxL1jgKBbUMLz0E9WAFfeInLK5CMgXD8Khxdho4ty5lu+AlRBbqzQaEiHn91I3J+g2HVPon
NPpy6toNyAbQi9si/agJeQbJfDtfM2co+mu/5JaQRBuJ4VawiniYZoi1UTXs3UFTOowbRaQTlfkI
e0h2+eWHCQmwYEPhu8APK4jRZXPqrNsk4spTNaAGfFCA1aBBqqJoueciV90JVxtKNzwg/r2F3Ss6
EJjZGm8IgK0BFOdLc+KSe9pu5etfnhhGzkwwx2R22/3SB7/kQuuN/lmCQkxg/idHW9WauEXj0cKJ
z1o3mByh6Ru+v2+UxosINDzjKxTWNljVhdqAYibtyjPzreoLekmLFGB854RPIqIhySJIkx4GXicP
fVCr/q+1XMlUEcebp4U3L0gG+arQcIR+NbijJ6PZkwuqNPtrr7VjWBwbqmBdG6RkmnGG3Mfzks4B
OyIdxQQ85svUbtvzRJjrKoCy9pfnN/ZXdMDG5VZ2MxEHqeohGH5bJRrsf+E8fX0G8YErPsMOOMny
53F96bdsWCnyVn9HsApipkR2UpgHxtzfZoN/NVI7jyDPryhrL5ipAw1sbAgXa2kREbtbPdaEkOCg
8zzX5CMmqg9bDOFeCHxKKanqYgwm2SN3gXbACPfouvF4kWhvlGqEFyw6OWRwmafvmJ/95RrJDt1F
fMP/bEgyTK2oh9Nn0dIhtKA3JldLwxDMhpEy+wWGGtc8DUsiBw0zSoBh6ULDCEySHFAypUtsZX34
D+XEykDj+EQODn3rX5r2qyrps8UW95mejUGI+XipHTfw8GoMZaZHP2QG6AWzSdOEtLdv69FsLjPw
1giI+5RzIVSz8ouEJgwY/9VqgGuDl1MnGxfKEsAZNZOSc53dNUcQh5pr6D5qRZ+fYXiEmcQCpHSd
7R6lDlCBt+s/zSmRRZuDcS5Yx86YTLPi0px4B4Jruh6DuToKwSb4FtyHZvyyogMgPUWU3tXX9slj
/FZnQbVIdyzEaDcdI4zUUIVgd5oZ4lH/o9llAs1rxU0z/XvM5V3YD1MfxdskcGpCuahLPl0lb8xw
O7LRAp/3qm+RG7ixsDyTsu7q9FpfXp97Z5irlKH8e7adUqh/263sNCBDJMkbRDjcK5nDoi0wgKp2
ODp9mJcsPzx4vAlDuystVJPGhuJC+fP8lWmOlrIcgi6unL0DlhrcD6KEsiDlkkrUhKSi1tLGOU13
067areJRTt47cFwCb91MdCFyZU+EQtwK7ZH88xqPLWkwzIuz2om2dX8gSQ7xictxB19GRn8gVKHj
/7+JnXFf+p42sUp9cOXuHBfxyi5MvrqGC/cl9LLD5WZx+lVTpnmO34YFvoz+Gqjykc+lFA5ytdOj
xaWROnq+T5nNnNGzEKxDZrPFu1Asn96ZIYT7dmcMjNjVbcZ9FsW8jODj22O4eO7JlYaUqnC7L+rV
hoAQotup0sz4eXsZFOANEyB1UxLsoQIqKWtJyE2dvoJ6PTRv1vcwPq1K1iVDoVGGvoUVGZuUbi31
6AOrrnbvul5HzlFs2ghwxfsnfyaWb1fpueaN2lDFpjs58HI3XwdzO75ugTl2O67zQf//hSKZFnVd
JbGENymvVeFMjbsmuZK8RO7ivTzxfR10WeZyZhIq8OHGdYVm5uRNzDLEcym4gsRkafVXkvaSTtiD
b3V4AHTavTHjnXa/p7BPApt2zgoOnyfuUScfOqYkW/IBdFof7vvh+o0g27MQDtrAGBwk7EGa6HhZ
ekyk4xxrwsSkqvP/UVimXdMQ9brIgjA3BMF5Qn7V2+03g0XEa4sYJyMJYuxirzxK0m4jESab/WxA
q2wNOl3q/tArpqo//uKTGR7mWqkeZ9Kem8MJJnbTIrH0oAS4uEqufLSrwyZhBKvBFnNjt2h6Hpml
N7gnD+6Pk+RD1IFfd9Jjm9Xu73j0Sa9fiWT6vJTc6dv7f8Fu+x3EgfZfHAeqToIHoxaSpKz8Jvl+
w0tRRA3dbvsTxX8tMrCzYoUK+JdhQ/InRNjX/8UWuUC5/vYIzH7FWajPjKhpVcY4o07ohfE17Hwi
KHA36Z87rxpVWyNV6el5XHPIJL3xhCyj/KL7MKY28bHi8KyFivQF34dld7TIWF+6/+i9ek7DxrxU
I09QK3qq3ElCU2gkpNcL3N460Rm293t227sHJPo3tWjyc31CLYIB1eG1fiDjg/O5qvvBkfwGhscv
mmxrJTaGqepduRlHorRX4vgQwk0vCxP59jk0scVPMVR3JXpfV1eA/Qs7+rrSmWMYWWOnqmOpzw6M
XgSPHBjNJ0QpTbL5ieLjLEyDQ2CAxk1FjKRidyn53IJip95aoAsaGxnc5pwUdpJRyAq3uwGrZKAr
ho7+my/CEFjNzVpM4zl/y6D1E9unNjTeLPi9/rtaMnXYIqhHM4mKtOuh76BDkjG8YYWTnbV11Hsw
5+7kRjmCrRUWCl19cklclSuxWmsxbxxltAJu8SZrZ4e4pR4UvXXJJpWHkUJsrDj6ddLRlSmSzAR7
juxqBl4tOjzP+kz/JuCAe/jkH/RptE+DInnC+DqL2VRzamVS5/X608uOsa+Y6JOCuffZHRQcSD10
xbgZhKoYH2DNfKW9wNcKzN8ZVLT5I2B5aJkkwyD94QUvYAF7hWFFwJantK14N6/VNDb/a+ndoU/G
XKjQD0w1A8QaP6D+A/l0cQEyH+FcT1qgarO2CAoX4Iaey9ruucMWpDJPrZ6EvKvQM9VqLFX6kTz+
SR968p30kMPdWvI8pEKli3b0mb3nCguA5hMg08DBP5iFxtf86IE54q09YvFMCIm6nIGFPwd51Efq
o1HOBrvehB7Ze/DsF7NsQzZWQbtNXJc3uyCUYfZYiqvP3PK0vhCs6cZWe1waQ6ChY2vgYFhlHyan
IxQ33eVqfqSRkxUCXSpQHxHVj4XMB/UwRgZdu7SuxsLr5OvsI5ScHxT9/5m9DUFoHe7SKnmnzTu3
6/cL8uKxanHKl5C4vjr7LyrFtnzebFER3bhAhw1eKpvOPPaa+shyVqPC95y61kE+IocDbSQzOWln
01fSO8aecrICSMcqijifvLNuRafIeW2JRH8LQqxfRmarBaOmgEky+mA/mKm2ajs0UhxdBrN3axpt
SBAY/PV+cBW+RLEqlBdGGhGLRzYSEZYF22izRFizKxEeKEcqYGvRjPRcTKodmsKyQuQtX33w1TR9
1tj38Dw6TR1vmrPVMnLD7OgZbXmiFB4k6H49a2TUmQf+uXGhLZvgSkVfoCx8gpzM/910EZxRtKGF
225Cn8aXL9wXGsj3vZDqSQ2bdbWopEauMs/Mk5oDcEerpSbRDsfcyoTTJ/0AOjSpiDpuy5aP0GDf
VD+oNo3GUNSUlOHKEgUozBLsOBrwxfSOxyWuAUkm9xpk02WG2abEmgunuaTqaeff6jtLSoEZhnFz
A8XoccIlUMfZnFNtrF4OqPEFuGB1dshsPFpoOrOyBvDXeCj0Hk5CGwX6t1Ea10XQzAJis1tBI6ji
59DllCzIZgZ29AkubcbvYTgLSlTbY9zLH3v7b6nazk2w4wEkrdohVlayEbD/nbHeUtZVP3K2FBjb
ct8ihs63/Cdjblecg5AZi5fLsotK8ldG7r/gFsIFbKmnstDLM0a8AwmFWGqFHjeYXsSP1LA5LdrW
M0fNdHTGU+YHl7FIFvovmbKk1wwNKz6IcOpT1cHGoJ9ZwatJpRjtZAB6hcfAia7JXkybxFHO7TKS
nbCq6/RK1Ed1qkGQ9kjvfEo2aYx/7T0i7dMmk8cA6av2/5wNa6VW+9YPG4ylG0GzCeRWF4tJ5Yar
XRaoYYK8M9wbOsJ/sWNSKXxjOx+v8ierpgh52/OOWR+5JRBLGWRRPsDd0QwM9rdgZV9uVtPdPkgE
eqmQXxon0Az7BFGSfS7l76+IeFTde31R+dkJ3+tCUl1/4aXaz+9m2l6M8aKDQQf5A41EJT/LwxgA
5gCr1KOcnRnbhQKqhJ8BCnilLTNCZ4kHMxO3LaIjEBl0gdBFVEk34CaTF60JIW7odVbqYT+kkuID
/jYcduEq07J2s0VtIsPqI0Hml/MHV4t+ZA+wtBfmwY9xsXBVPAfVBQCHN8PfYlSysDMnmsZkRZD1
5FRM14u3luJZckfPnCV87YohSGOPxOyNx2zfU76Eljs/QsiT3Ex59g8Y76B6vXwf3Skt7QDnoHaw
9coWqfehSLsqjzf/VxGe8eK2CS6cvB3fCIADS6prSRU+wj+H3SOEWJDijzz6dghv1RBhJgttAL/W
Vu0PWJ9K/NMhthFfz6QpWQKkarJcr3wlWXapoGGclJQPOI7t5DFPlZFGLWC/Lk+6pgEjDnYPJWZ9
LyHXzAcHBtSO4VeO5IIH2sCUvCghW8pGPJiCWSzPzATjTr/mXH4mMZznBgE+wfKLuV1Av+w0bXO9
X0473KzeRPKT8AuB/E6Ih5k9Te4P7hCcaY/GhAP8kZyr6ZZyJXGrenoGNd+ADH/DoCI4U+nHANKE
z04JXNLt46ZCcVOxeIhdjKbWHOJh9yy4CmbnYE4YeRbxgHDcmVsoZLPAifELAZ3VOY/uAuwRIiGQ
8U3t4oOMQf0bmIEYf3/oXeG8W1rOBmevsuaWy721dPGfnWMV10z9iNGBtehierI9BoZe1cPQQzEq
Xsqih0fFtHBqgLB1zCJSimSzMkCkfW0BFy/3u/IbHaAhhyY27zrttHl5MGXsoP9/GDvyYqShkbIA
S2B/8j1AFAX4UGYhV9/8vpIVhEyN+NByx8ysaevDC0Bfd2LYTvEsW/JpFkhTAjVaxaIRcCN6MXiM
y0XUHGdAJu8bMYtH7OH0UvGKMrh75sK3FeFXZkdX2HPzZzI4CWh0HZeTdGAM3IXzcsTiG3ldW5T0
7G3WgLSH6nFNeUo4iZLc4xQ9jpIeR4+puIHnbmPC9m55aYJnWFef5FW8LWRU9sBK1GK9qRGxs+ov
5NaNuJ4jtAEqMHPWkZzteyWmC0ipu4Qrud5MV1heAMXCHroDSlzPfu3yAx+cr181Qi2CGT69pneE
M4hwrgP00BcJvK2gAKFc7hl/PSQGMUWZnSLMJLCybHclHIa0lL9MIsrFZ4TGhcLTF56qkrhzUmnI
tdde5wT3MsTmtSnhI2QJNt9CgBm9p/tDWTxU7ODn30RnttdrEcNaSeCZNJ42aeH+foxBIgEnMe60
VvSPWzvq5ANLw/2IdhYHULUozUfla/jDmCDsROucjzItl9fiYHVAJIgUq88rEA/lnsClIpdQuvzD
17L1zIR3amGHHexX4uiT5rfwEfiLTOOOdQbjICrYbaZj5gyYdlY3v2ygKNllTwPwxmGnnKNtaorj
8e/4PK6TRNprNXncYpK10UIxgrLYLFGqluK3hxYNakr97ZXrQ9Ar8icSuruAg7hur5ZZZNZ1Eb1Q
Ogaj7iFKYdwrYL2qLLzE+H1rxJwyqD/Vp0Kjfrl4FU2iil0ln1Wz5o4rMxPy/YjUwhzEGywlPqqR
w8MQd5jTvoVJrFvl3jMO4OIXd4fNqO5rM46zX3zPi4DTJZl/WuLvppWUJcvFVyxywneNqlns+4t1
pynNxiuJ1qSdOo1u1tqNaCmz16gCWUsaleYr0kOzbmKaoiVgJPC1PW0cwtchfBEKur2FFEqZX5if
9DB3emJiSELAYIAGs1QhStnkSCFZpGGpx9Fo1GtbPCyKEGUN8i5qCFtwUlf58/xbgtm4a6rZtwg2
qDxdenePjmYeXu7j82Z4FkaV4xM1KgGRwcD85c//LoYlO8dTiH7IDckOVDstrssynGRm7cpHSgi4
ghesd6Je0at0RYt1Tzpfjv9XQtlJoSHLbjPTe6i1lv1il2/5ZSziA1TLUDDf8btG4mlS1CJ5y2ok
tD562e7O+Q7IODHXYhOaANCSmpkR5t9zpNod/uNYrKI9qoAlAMIDCuhLhkXZt9C866TrtxQloYKX
hNy2RAl0xN4Fpljk9h5Sh1iZJ9XV4uE5KpUEZ4KIwgl8fPF4r+KzNQ3uHsa5RT8HVgQaGSr4XLZ4
kMXMM2rIz51z2CLy59v3sqDgQfr1YkOwz0QQRdYRJrGvWoZlBoTrkHoqX2kSXWKiXYVoANGJGS50
3uDgOZtcQrZ+hU+fRSd8TwxlQm2xJm5mxm5t4Ve1mmdnjpFXQD2PFND6zuaY8Sea9ru4wFQyQkMD
V+oKqM2JRhQ+12mqfHwh8mTOcKWZT6cnKRJFE1E/51dWWFehokXRPwPgqQZ7Keyprm8OnIUEptqd
zqPRiY6rSlxKE0vbhupaKCFzN/DeUNThI9KRgF26MPoxRjs0eec4pnbq74jM3GAa1RIyqa0l+vf5
9mpibuYBQ96t0xQicpUih89V/P0pmMJgWbw2QDAemRQPpERt4A3Eyil0Wx3hW/ERMMbnCfm3A7Oc
h277yxzkiBDE77OCfOBoRXszBK+Nf/d05HFL78hAQAyzizYPi5vnARr69QEMQf+TIyTvAPp7IFpU
PR/wkthQ+H2Y2lMYb6QPuC6xY8vX7s7dCDgxTpDSFQ8nnj3pWVOL1rJnSwhsXcjJCkAZ8mO87f+q
OK3aafXqzcQAHrN47CuZAfOIjSxxNMDoq/5YadNaftOjKtMFCAG1lOxNfe9+4KM9xY2nn9WrGHEI
KaZPmW61u4Lsr6APzCu666xMRnLRzEUdptXaO6trblNSy3XwNLNq+1/EaqKMo2t8GByjPD/QbEJA
a5to0xJDzxfeo/zEUsytsOK/TnPBA/qjpeSJSfyTvdjHmFxdc3is/zoQOvISumCgYGPQHl+Jpf3X
d4Qxncr+ByoA57voOlzF9nESSpTtY3Cul9SZLegy8Ts/KzF8t6RiO9N7SbH5ZyX5zY9pNiXt2sca
S9eiMzKR+S7zCaIeSbBzXgLGkKzN1hqGzXTAu+W5SC1QexYObkwF1vO4alNakH0LChW+jxOCXETS
RBJVExKWxmcZrvae8LFigueB25MYYAuak/b2/kaeeGBPB5GtWzHoYKKSc+p9KQ8NWEzmBI1kFpaD
hQ4ILnZfD/y6Woph2PmhEeTch9znLh/NQ4GZR/N17Ie0gUbO0siU2KKGDRdkR18ljw4W0XIRwMM3
+k+if+1DYjFFvx6y9STzarWHGUAfpia8Jx15hT7mlg8PPXLDxCXHHPet0zb5Z6+G8kAfMLzEFFFC
mghCMJx2Sc9elFtQNXDTonirXFNzTk983GV7DrSjitKAw6Z/5XhurWeka4h4DCBQvRIrifr3l5xL
QEpFgCZbg3CjAe8DlVcyQtRrSRmNa8T5/Dk/aWa1AoBsnS5I2N0GniIpSA7iYjs31F1s5RtoUD57
jIjv8p8s/F5CNHZia5tLtxqbdJqmHqFdu/RLE4Mm7HzZ1pB3/N0mbiuO+X2UXu43kva9djuqnqQ6
O3OmC0GFU0uHq/MDBzKlx6bYqkhF+ehrC0YMIFz6+LSUVFsumyq3N8iJiy6NlJlYXhSf5V7NXSc7
Wd+vlJpOZBICX9vz5Exn/3g3jL9Z9LUOnYPvoEHCIx0fY7EJkO1FcyTE3LLnT//QoCuIHzhZFDbf
GE9gVaNbgN+z8oIFbWOLcA3SRndZ9r4CTnc+B1FOYN7Cn+AXLwRjwc6lbPjh8xfunNN4STdy+2jZ
sagy5Gxa1BtWZE/heUONlYl5dqGWoZ8xgOdXGhMGW1tKZz14P7OvSFeSWhFae3kWQ6eOA1wmYSWP
LDKElt0y+og4FWeRjr0ZCmmqqRlGRTeMOPHjwUO+cMmMsFXV9mpttcIHkYI2/O39CrJcrdQf8iIe
lFuwkwdeOZPC11p1Xs6rqXrwN3H7TGnzBzSgtXNrB0bUr9h/f4/EagzTtgI0DQvXE8ueTtBdZ2jg
pN1gVkxtlLJyPRCjdTZ4768oo9E4PjWcljYJxQBc6mQ7r0VPII66Qc8AQheIelxoGWQwZ/i4K0eu
Gk+W9u9U0zEgmQDPs8d20Dd5mx0+J8Q8iYbGCw9ry4d/RpJDkw2HR2eWlU4xTTXMn7XVWCX+yUkc
77nhIpS5lygx3+rwA8gHO5ej/t+uzSSGwPwalE4vG76+qSjkxfoM8FJOGTtny2+ALg3PBBY/NyO/
miu4E8u+kaIFlExIYT0+5h5axa233OMH3U5+/z7gDrff1nyWvCt0v613w5r1OASAZWoVcXWYtkQq
I5aOxYym7YyZRkwjR/Je+YOa4CQmXNaq5j5zHUkvfxKx5BEsxpCcc9m5DiPNA767edhL4fRknkfC
Q5OAujVrjkfJNzdxQAnpNoXfFr6CuojpAxwUl5+S7+5+5SDczf7Yf95ES620gpkAx5Nyc8VdNWhn
1tWJ8nezi7e9fkYbu2IRWYEw24FB1MkhidNRUFj4Z1aXmg+l/2CGoIps+NSHNWsRUvAnkdIibzzP
aOf3eh/OmvEr0pnuKB4jtAin1VoxP98LeVm3Fc8nJto/DLMDaE4G4e88m9Tpwys99wR7tB+i6tvX
p+3uVH3pY+6Jv0njAyY2OmauAoEP1eRiPkaea9gVKPP9Qx7qecG+r/iN4Owv+eBTJtSIaNoVNT2Q
vSUpnvvvNthnOZSBEaHM3nweWzj3dErstzDT2q2uNQCIKGvfEskJqif6x5bEJk79EFyUOHhzzbd0
g8x00uKtq9KHr+pl/MlEzd+xGlh3kLcujjC6fhijck172hD1zs2Sdt1XQ4yD2O06LuCzi+CBaWN+
TZwhsf78Jki6tOIoG8Red2EqnOe0QCgnnk8Zyhw7CH2oME9gZMa6B5oyFdJIBTHqfsw/Vt9/WeK4
J1tMgw2KSyDmCwCSKDu9EPK41PET6vRNVNYWPysIgU0GGV18MnAmoFqlWlI8kEcGpQiubuxurrHL
vKzCxkEm2+MaF4DXb4PqmxfkUuaC/UJTeeIkzFENEtRwHnZrb52G2/CXe7CZTtpcTGUmBM1lvg/K
ghou1gAdu7HiGG3HQlT1eMiH2G+Ftw0LEnPi2zqIL8jp9yEFgRH2Elk1ll/1Ik+njO8o/aqKMc/k
X2LlIghhvtr3SvEVvEYbEretGXho2XAR+ATqA7gp1HaqO0PVxfXErrmJTcmrlMKrtYZQpJZT9kUy
kgtX3NJthL1l3PyhAr3uO2RP6olZBhgWAgoSZ5/V6zqzGzsvoom3N55WHs0pVgpTFI6MMnx+rZez
jRIkU++GihLDLsGsmpSUVPpnBfHFZmSzdHz0DE96vz+TAJDO6nZK+b3FIcw1eoin5oq5aZ5q137L
VOsPnYcdkzsnHHlCDXs/SDDbDtDlmIGuBDr2lbar40+c8k1zSMYrnOff6SVTNJRE18rYquIDn1hu
q/+fwFb/VqkCWwXK3OZ5Bv6NGJ80mC57PSdd848Q2/hIxQ1fXEuJLJxYB03iM4onToqxGslcADn4
2AqGdQUFmFg5uqg+sYSGxgq1ipi2bAg/tVdP5DZRq7/YHC52t9wNMS+uzsWIWDsh2eMUr5sKacXr
rI6dLpglNKH5NX+fhafBfhsTmh0tR9/F+/8s4bnHF9buBOa2AqcwgjFkVJLJnB5UD0njxUeQzPqL
bW3L6mOoKSCCsjEe4jjpF57YI8R2sM93BhhVXK6VxgJyZreXm0JDRvn86cgukk7TK8y51XzmLAcS
s9XRx1D6x9EcihJBOj5dZYPpzzMxHQOiYtG9hOhZO468vJPkPSyoIOIuVlsbd7632WVAO4ck2GqX
BvfFeFzPq6btXKZN0zbdWpfvn3R4ZzJi9zSIEhqoHNAMGtUXHevFKi7rZOAjxvoZaq373/XSH/rm
NC1JvfONWQQfGNNzkUp1KqBtgsO9UYQGq5lMLQLA8p3vQUefgW6GUJUMK1uu1t/vwM5FPAiN7Wxe
UzOh6rCaDi/yBsrf0J5OPjf3jra43cVMAkpD8Az3nnAHNLUIy2lhRWoEhV5hbwV+jBRrQSDADC6T
oJ5jccaqNJ67Rnb9WpfKmy520fv68ZhrAiXQcoWF7Wi1oLhknnINDquRutdBGbfHu4dlA5AVVSJs
AMGNmXEeUn9mo5M7QveNZKyX6zM/pLNy+oSO+fHB+ETvJADOGnHk7Q2b51qaaiQxXf9wq7pF0FM5
xzKyVV9i6aFUP7083o+VKwYFm/nvoWn4WNN03jyaTrywkkkGZ9JlqnGrSTovl1LzrkCtTx0IOEoG
PdUPiq66ZzbvCZ+Ilfb4K4/4Frx8Qdy1BiJ/KtOIWkZu9iR/+9IH0vDflJ8HeJefX3oNqfQg0+MC
8u875oBxNA6X6zrwv5UkGV58Ac7l/LafNK/d6BlkcC4b+7nf/GTiYCnT6GoTsScXyU1ux9ReVQUg
o3C23ogVjF6lFmniR0ulQGYe1GZr97RSlzXfsmOBtWG4g0418T7u8HGfRQgR+fvElE0Jqc3yhL/z
ataO0CZqp1aNcOblQvvwqMJofSSqEmaIcSRbsob0cnq5mR7AOJj/ams7hxjAwrg9K3YqWIETwzuB
9YjKSb/yJq58j1ljvULHVBiKgLEh/6MWotU7sMJFXxFyNiLTBAOCCNfrbwrLqQZvMLP3U9exvw+J
aUxBo3DgG1afQ4EY0Knivez8LyDSOxAHWAZOCihoXsQILgxKaqr2fXOdFu3OjqRsjzHHl1UQJ5ZS
mB+8biTOi0whg5MAn+eXemXvpXF4vFlwynsI8dwB5+1x4XQzp2heOjTCYsyXrkUCPFGuCxHvXO7c
fLkV6q+v5RuYSOnCW296mgOJkfOTPEqIY6noaX3zNBneo+Z96zP8GHi+6G6ydQmY40z9+EE15Myc
alLLfJAcTXP+s1M2jtvRtSii18iWzSVLWnprI4/fA6Dtu6iOYfgNUBI0mEZQiJsh/h5c/d9fszDe
ymA3NYtfxTWUkjV9HHpm46LNKgyazwZ7GvXp8Yz1l9uvZ4UYBz8Eg9AUfHBzMSSJxgjKAJ5ADMam
9CHhkQy0QmGqCeFntofPg53s3tjtgPR6WVH5bwd+p5+43MGiJk3YzEBo6LJ2rvMdRcaIlYIQu+rA
wOFl67Z/POB35Ga5bT2aIiB3b1Xb8t2WNI/ocnHqZcEaC9nCrx9d/yLs0qK2KKOjfBzGi/G43bTx
Cg9D8IyeBQvJUjGq6UclQFBcREh8atNYZKewAMPkZoWT9cs7GBTju1zUgXahpF2DYRwWsn3x83/f
EPdgI4UyDhpi7X1NxwAY4v1edGfhaObnbxO/EdwE2JqRCxNqYiNgfY2JNgpaTPoVODyOQS8lspdf
gtS7RONlMt/iIBMrJhjJH717Ds9yHYdaNfCOAfVSRe9c6B+E1Yt6jbGM2MH0QcCov1SYk0+Hl8iY
i0GCj7m2qfFDB0zkQzHfwPsi3jj1ISCPuXmZrLhqnHs2DQkkhlNg/i+3CvSlwYHlaS0fLuBfau0h
ETy3ybdVVLhDPuP4uUP0UWOGe/x7tzSXDkW21PX5ukj4wpIo75K7gffEH+ToPtxp49UMz5bkS+jY
uqJqwN7+38C02Lv1Mccb0VZ6gv8px6h4htH15HLgnPIsXDvGCcbyYoSCm34tqJSbGz/yYksbLtOF
9CgkpKHsx3H9qELXU3F1QvxSquFB4PWAHpb8e+iLR5887aFEMF/mUth/QkjiP+wYbkYoD+jYYKgo
Fy4W2uWm2CbDlI77/Wp207E6eFskaA/H9i1Smtt7RJXOjPAdIOxv7aayJLUZCCPuQUNYHKirMYmn
jHXPT0vWEnbJrSu99ZuH1VkAdoxCxov3/O1Ezmc46LC6mWvzPHxVGz4nX93i4hpnS6l61M4dNSVB
i6K8ishMaKmP+uj6Xl6QapmER3ewE7MpN9Zsb3H9bhtcZ9DArQCaEvHDQpjO/W/gJ7EQSyfGSsRZ
TJvYIZoFpB+PqDQD19XL+T5KEbjmvExOuOyMcD+gRqSn1Hngk8ZOSQfDmLag5xXwFp7OHazMsQgK
2bEtyikALZFEd9HNCxx6FYPUdbb9LvR2zKlS+QtuX8jgVPOmuj9+In7QUGdIOaVZfTplLtLyDRUQ
I6xMcKMB8dMDOZfdkCOh8TusTM2pS4vRghyWsibWd0xWzrwbmDIjM/ZPW0xFF+BLdvAGLtgPnOyf
uvkdZl9KMXhdPeS3RosGfXyGuN+AUXXKXBzE0boYGGmEIvRG3yKG5jEuBxr4UZh5a8Z3PIYkpnQX
G1CGkAltsVXnO3GZJYYW+h6nsVpDAAS+wkDnZNKfVjAQ5drVQjLStFbgtDGjMtXuddb6wIMWzBsx
5GxpDq2+3qHdsIKWR1nhTBOmR2IYw52Wt0FWmV20w4IFqKPrIuU8GQFxxeONLlXbsn/QHf7Nj4D6
6LmeMvhQ2Tjz7tnQvCuRvQgnKMcbl9rlFWEKRek6ZksBi7y+UxBe+0/b02ro7pWtXEFDQx1KfmUl
dhh0N5X6/GI3LVQ+qoRX//dF1dWcs5aYXI+4Fh1IjQTxoJAoL/QT6thlRzIU9ZDOmm4d0s6FmjY0
08UX8p/NfgmILgKqBy2RSXbO11TjByjDq/EYBaxG72CywqPmbAHYvmQlTohz8g+7H1mr4cYlBku4
muh1cfmxtplttdaoeIzny0LowbqLyl7j09X9OqvTeCmiMTrX/lsS28tNstV5RDPxIsL/VqgVb+Z8
J6BBsIqvyDIvXQMRKqPnwzzVncBLhU+vg1NcnokJs0uJzRIaW4npx9l4VkykNfLUJ1EdV/op2LaP
S2VG0rqQeFSWhLAJBNdZcTh8LE4atBtXEKxY/L+p+v3iZHFGrmJSSGjy2Tgdg6NMLOzhATz9xd5d
ZmGZd70RWIf3dHjPM1qlKoFLU0oS82ob2uqaTMv784VVki9Jg9ON4TCOJ5hNPQud04pOO4QkIw3K
XL/XdSQeXbijwrcWQnx7RGWZ01J6CI387QQ2TgGitogBb88pKIHN1XJt+OXRl3bAT28+R0Tm8Bio
yqJDwfMAWCx/buKsF1f+VaZKEIJJ0h6pZ9Y5/x3W23pPGJ//Uj5pjY85HRTTrpjoC/sfv8A/eYxc
J4JWqPHG9JfNcwDNIirOZVXWgW0Ch08gWCRsxuYL2pYg6cBAObN/wwi1YwBXp/2rtknLCWCHwLlO
KVkM1haFea/9+Ex6yeC1YimDpyfIL+bFTLl9faAIrR5LyETKwiNQsGxZkcGYGFjLLpV+Rpby4Erc
0w2jHl4V/2hO6jYmQDPv9lc8JMGA+LXOUgYc6QIHfzu7D9jz7JjuxSRYwY1aU6OIODoXToOYjkf4
t+5WQqus6gigm8uLC9UonJMSRrp83hOX7MDjjFEH5Fg5gPmO5ovopJeurufz+DWB37ngMYDepMgT
WIL74NEAW6QP47yygmG3Kd1/Wh0BT+y6NhEo3dp9tmSqLHj/U+M2qLb89rZzQIic7UtmxgRl3acO
wOwhlfiNoK8qAndDS2X6r2mj3JaKWumFNogEaibVtxLyS7cS0UfcVPAi/iSTEmeuv/VlEFKakGjD
U5u4n078TEUCrkQI3/2Py/z85fmghYT1mi0lVISxfhH7019SluEj7crlYV8sCzCAwLZBXe3kaPmT
av8w9Vq8xDFVlT9lmt9LjU7js0h2gpenHE69Ax+8Q1+ccZEiGNTPhf8nTiTq5CQSnFVzfCMgHjTq
tMSHquWoywApOxPWnwNqn5zgxecdJv/tLUjNRYip2yNrmiI44C4a4VncrNyMWzkygqxpTK/oCf1I
HqBMsO4SDdCkb9OUIW8ynfDondKsg4pISmuvSJqXhRpbLPSDZdD2aJA203/vFieU6c++2PG7Isza
MU6h95L48KIywWIhphWj7b8WcnxD7a12KZapa/+DI8GljyzFMZQAVA57mf6jAuRCN/qAyWPy372W
XKvZHb+BBpZwaA2vXqmi8oaO40emf1D4nuD3aRax3RNLbDBcEqEwr+tyoGI9gdUu+C2Btpx4U/M6
r5bcsCRIOvR5B9Kjal+1wCWRlasppZ04NUkK027eOjA2bgJr5Th1/5AktnSujw3RszmH8okeqjcd
qNih2KdXrW3IvinK1r67DO04wH9pDPLemJGyHU3CxLSJ0Ulb0wTVJezZeQyEsuk/tU9I0CLOo3jF
T29CXYAxXI/ktYs3PkIo0c1TF0uk1oLvOkZZSFGXA88JBENZ9vQ8h0iRn+QjXKGEiBaTHzNCulQx
8Sknc/YYzReDwb+lbTJKL6if8ZaxPZK2p61I1A7jOMKGhz+aSt5+nWGGItFCrkAine7upvtg8A3w
DhIYOb38LczzOUufEMJ7fi7DbnDyUa5hdQKB/QQfkXIGMWkOITu90d71AUlBuWQ3pW5Kip86sv85
UpPVON3f3Tg510Tk48ZVsEwpTcjSsRyJKKoz1snDXVM15Y7Sy7dWMgoMYnjyddxwOTSF7+4Hf4+Q
GE9QvOma8EhegMsuOrofi8xP2Wu+cECXUQd5HE2tCdQc7fq8JlLPlBVQECvHnZgtAzRG0jJXIzQV
6n+5WVKhEo+3kTvKxadH+2THTYB5oB4seFwgzKqIQ/xxZuV+CqP7FS0ru5RLvFHsio8sW1YfBbaT
J9vJc97Q5WXT6M7ROU1cGj4aPG4gIkWE/W3avsT3q/cqDwA70P4/ApIvTANJlFgF4PfhPjoMMIvk
9uA2Mdb21kVNsLn2HeqTEpdbr2INcXU1tThSFV6bh83QaWbttn0xOiou6TWzK9c8vF/UC//XAVP5
4/VhBhnBKluAiTjJAXqEt8FvBuoj2Iexihyc7114+BpSt3iW79GUIqNl2nAHSITzV26JLVGNVyHK
BD85XwgOs6U95lyiKFB8rRUlOBff6w/IhksZ9OM9OnpeiaJuC69KIyZRi2Ohw+prGJCmF+XTS6Fk
AtBxAkqJO/P36FM3wtp/KZRMspLqXnrQ85Aelg5H3WYKKvtPlZWdui16zPqK1dLwnCFEEeVm77gn
QOWd9VwVaXI7W0ERIg/H4HGaYv7+fT17eQ7/wRk3hnWomxUQJwWYx20VDakVp3vRWtYb68nlgirU
xBL8sJyclKINUCq529Lywcgbp46PZfhVc9BUBN5A/l4BP6DobHLakeM7CU7DpqTThPcJu3xhyo/q
/DcjGZegNv4wJhYnGd9nucLRO6IUHzbb+mBzyoEZ7VFMT2QT6IOy3VNHqqc8g9oLCpf21R3202Ep
452vUvRo0irf7C174XwrHk/vLm2GC8xvr/z9DkvID75omIvwCDF5wYIJUwfwZYSp4TsRnKwpOTqQ
p1rWJICdCsBlLe+UWs8Dy/9wOmF9XfvhIYjR0SJO9cbyiD5XQbM+4EEsv5jZ4ObCBE9t4NJB6HVY
2MnHohnhhHeMawDGGkOWUEEidb9/+VW02d7zmU6MT8EOSCPnL5VFs+MdBXb/SA82ptfZ+Mp/qPLQ
dkALje5bFBKKK/i6spb/0fi4j0Hf2DYM24gVFY40CJ8FCZ9HeDX70S0wfKRYZ5eiIuyck124ISUg
kVwuHyyOidrVZSN8z7+H3CAKks/aFR+Qfz2OvwDGBc/22Q8q+SnbXv8hyonK5CJy8wg7z3GJs/5S
krDXfOgUeGBSyrnKCk8CKhAVA/Lu4nOLJoPZHS+3VrhwmnBKY4Quw4vMdi5LPj4X2CHRbJo2qOr+
DA6jDRgnqMeeGnSrdCag+jcXEnZ07OtqSYXA6RnTUbjuSwBUTIkXBIRP0M5gL1gSGmbSMvLPC4Wh
w3FVy+kc2+KeMITFDaFJYLJKCuyONoocxqopxC/hewvPGxEA7PGFhZwTV2An5LBABTnDfRLASBRd
PeEkyl9kLwnBA+fPYR6RbtZ96X/xhcAoplZ2LBibeM9D5T3BEZosAMQExi/GY3gsieuZmTak3Dbp
VwG/AvUFVWYQpY0DX0JuP7TRdpQGm9weo19A6s0ozN5IYQMRr5yAd+2hua30bG08A+EkcQG87erX
tDigkllbBFKs7Yfqz7vQKZ2uOtlcOsohRZLqbbZvjTwwoSHSPTRr4h/OW8CNH0GfOC65fLePT5/9
UFKSthWkH+d6ybfh1g12aL9D3+IVaGlFtNPqlKDrl9Zb0JlHA+lhhPMPmwnRiqjWiZyewgzosjgQ
kUuJxRkGrlUTR9Y4pYlCQaN790CdOFhT71coOrmRlMC1MAUzRqLK7QIrFBgWi88AtPRdt9aqBRN3
DYqe5V7PAbxkcAsTT8GzXMDi1r8PpPywGejXcmIVTI/Bo2qERvmvE8G1PzbH1lKZv5EQC3kalgjB
lH+sRQ1swgfFmuPablvXi/K82BcpKNJSd0hFtGCoICjI8TBNGoQhuPDhOXS7KtFD9rZxAp90rnFY
Hn+/5wIZBL1eIXJDWhhW12yUqDNanpfvjUzdg/+ce3e5yZ8Qy5+j9qY8jNi5sSRHZfudHjdh0Pjb
SSL9yBf0n3eeQSAHIfL0UhLQnhwG8pRkkhQlbOyCWDbVRzT5aqx/ufyGNisry5AsC5QuAC6zjAOL
Lxz6Mzpj11GEaBaI4Niy6MHSZzljdxUBDu78AnTgSRODoEFF2VWlQjIR1te5//pD2TcXGtys0ux5
9vCr51+X7VSjIoo295sziGT18bOhiALkj5x4kO490PZhtj83RoSpgN0TkYAB0Mqr4jHzYzCdyz4b
5B2VG+3XlPBR/YJFlYPWW2nPKCcC0MKCq2suDYpntHa6sP7aTG2GjvvlRiKWZsQUfi2O+cNWfCHY
WV/a6wk+T+XE366W9EYQhxnG/6bQT5nR0fL8d5czXuyD7IPdUE9PDTC+493DyXuE5Qxd/P36yHzL
6ZxXGXfkp5gPxl6O4qAPxPOSpShqsRbWraTVP6VqJ4oVlEbvdCaHHHojuiqhz/XP/bDDiFW4NxXM
w5Rw4XOfjZAnPo1PuQ4x/W9u/oybyuMeXi1HRpQGwALfg7YIGpDbssd2EM7jF4Ei3mciDnU6iQQ3
im5dqQVW3tE36D13R3hpz93XzCqq9x9pmaHBaKN5eGxV72pkSVBIxr/412wXvdFzJvh/QzIiJ9oV
tWxSJMX+Jmr3vbbtFOdNgMXga4V0QUrpboIDh72nOWM+LgziNiURUkjn104K4mICfDQa245oGIsT
ASMAGZuk+kCQpRf1WXoMYtGDr8v8vxurUnNlji3IvgzvjYcr8isMOC2kCL1pD8OLbuvKqUR6V0SA
f+jKxAra/AcHMzkEv1XzhQwph+3HFsW+tSXVRPJ+8JfkpIew76Wo/pEt1wPR+Vrn69aDfmpmS1Iz
SZYldmE8Gw5dslCWu7EMJ2YruQM6grhRf39snstcnYGjJ5HyH1CIbDaxCCPBQVsm0ILOk1wT0yrU
etUKX8Tv9fwV82jBfmNkDuiSmsudzEPFh2zFLCXP6l14/+DdWKctQq7hIEI69fFUKH4/xcfezPRw
aphRG5HVBjn2jqT6ffjxD0Mw3ILEv0Puz8iUrqfx1YHkxXmHXMYmnRsOhDWIbm2b8RZrn26b95WS
SLGSQv8oWLFzmKGSnQwmfzyfC+FI2L7GOBC7sBGPW/SgpoJMw+VefTmYePsIDorA5KsxxN2uzgS6
zOQkrFYgvmIeCodiiweuP8a5uf1z0mtuTaRDNY/+RecFm3HLT4nGrTBWrvmAvpXRrtpgLFPouc9e
MrkKKfElZlWpcGSh3qrgv944cUmz5aoeExnJVPc3mtoKuCqSdfa+VnG5eem5aRtHFg2yDiOLBTNz
ACE1inEobQw1c7tibAjtwLHPX3o4qT6E5aDwVfNXXajhXthowhW3CNVNxAfhS2BI9dnVX0Blh+KU
+pikZW4a+FXgMlM+DkIcQtwqAqcEjA1IAmRWLwdPCQHAq77ipOiFKced69FqGP7bcZuzDDrK3dg+
NAsVtYKVUm3BQl09NuA/Q+nOk3DhxkdGkQkXec49cTCLJg+VX5+6sEOSb1H36LK0nyBw5bJEEb9N
MfeMUjmS3MU4anOSjIZkNjhfcpMvB8rMU0DvHkLziYpC+MazrJF9vjdykJyYYEBWd2i9mO3Zk8od
zlfK2GjX7kyRVn7bmAI+wx+S1ziVmtpoW5ztvX+cw4Lg020qS81m46bELSn5xOb6a6kC27qJ+JYA
x6NjluOWJSAkjHcTy4K1dZ7ZLKRnSbhJBVpzHl0w0A/dPr5RXWahVpQW018N1K17BnD/s6WICQwR
SY7il4GposMMYUWmsk9xSijXC4T35u5a+pkAvwSJ/INagJktm57iRZcceH8hA/xEQBQHSZaXjsPl
I9rNVHqNxqK5FIdf8vXVfxn9u6T44SOC2zv9CuIvN1qhYaL/N/f1ehJZI+FTf317fde3NhfFMyM4
Eq0ReKOQL2E0t04/IJI1ieuzke/75Dp4st2w0KO2QN0B3KNo0J77KNFQoPkLiz9jzDRZN6ov1fg3
hw6Dx+NhNRhdhzwUeOC1J/28lk1MedXkPqwW+owktV5g74aUvMTCXcuMKbaG76Co7v57o5eNTK4a
xQ0gk7rEElYADwr2yP4i5vBfzmPtneAvXLZdW0S2tB8GcaeWChvYcV29fJQWjmo7GRM74wZvtOF0
QGfJlobGYmhfCwi5YfJph4iIw6UfdjaqSJBnvj/AcnGIr9kcmPMZ+wobLVmkWidQy0FZ/dlD6I4u
nNoXNw7NdW+a7To0bQhBhpjXegLpQozLHadvZ41GlQ5WY5ltnPDeYlVvj51uMXcyE6lLU36nwoDZ
sMzedP0hJX+QwCRr3NN0vZP9b32DEiBji629p1wtHOcbgZxoflzqw7bDZAUAsmhZRkmMC69r5ztz
N/YiGCkiWn50KVRBwnufY8acXdh5UlDkGf/f7GWk1M+Inidrl47mx4lIRtq5zK5IHlCONXLChiPG
qiYEXL3YTIjZE7hVHiNlDFLRBJZ11W5+gP1vuHFMxPI/uFAu0jSeeHfFA1wL1OpVAlWDbhAfiQxI
aLOcjJpa2DZgHc2CI58/lnKHHdTADQ0kqCdaQDScp8iJrL9+/emIVkoojrASmGjdoLGhNyBx9Mr0
l4ARgfoTbF8zbALenNb44h9M8+4WqIxFT7xKtQ3c5rxUrPKduM1cua5XxbneyI/GCN5KQhmdHCZC
Vnc3IHLzEzq9/iuHvh2hsklFNVS9S8HccqhtQ+KyxYI9Ed2SwA85Cv9rQtuypkhc4FzK+TPTOpBv
S5RevLaRrzKvTiQ2rLFHFFuctMaZ9n3O/bKfR9N1ygGieNM5VW8Cz7E/sc6qp2jc4w+RHb/tynQW
g43faCuuwYoI/Gvds4JD4JfQhpC1KkFcFb80lTqVN3du4MndVFz5aZGNmNhX/gl4KeZN4syz+RC7
NxBU+jcvHjHMc50g6NUYuGnYpnQgvAKRt0FVYMsyD+03UX9VjchiZrhTzTrBjPs2m8YyCVLa+fed
iW/zwWF8Jf77bBOPVJ11j4qTyBBkT9pOfiXkCVUOaE63KfL+zCZJadw1V6y+RxY9y4y5hdu5mSvR
sAnHI4unfKuSyxS0cL2racEPaOsfYnI4QUtvh9wY3oFcG3aibdto947Lk7iNteXlgo/p6tDu2ckG
YVxmt1sHU92G395iIM1XUx5aYi5edwqsBQuoy/3QEGNdH+gmxu2Av6a+t52+OyYHTJVPAZsS8afC
6uJp/B1YMqj79og/mxVdPBcsVGuSltBJgngBDd2K6hKyfYNEZ50X7oE1gM5TWJus9XIR4q0cCFtP
Ftq/gTtmPxpv7ajXSiwnqBpvUSpCSqRCJgypqiNO2wruPB7RYHNijaXTwds7mSGaUSNoCyTLR7n5
6Mp9aiMO0llupxUVwa3BYcvja4ECK+7FhzeXtPJu+wJqfwBud2OGk3E4xkHtd1Gg+zpC6zJXnUcZ
hgbMZnu+4Z5o3Di8gFc0Mnrx60Ok/onAMSOWMtSAuTAoNLEkNRVnhAqX+wjs/tFsh3iUAtLY5vSx
1fwgj825fGcX4B3kUTALI0BKqD3OktOMU+yPkoeegr75x8uU5LNitYHPWG/pwHbLMR2aG3LEWCWu
8q0hByVjknGN9s7bCBn+jZmwFlrrvH8r16vUgxt5UY1JDop7iQE3sIj9xHbPw3s9zOevo85FysiT
RUaMa41gOtOW3Cbj7sDTcQorBBhizKXcmRyT8EEQR2tKYzRM7liXS4tSnVZAckDQ7omv4BZwbErS
rnIU8w4P9/f+3yC+UDm1JkRe4Y61i6K6x72591M7GrGYGG2484o48ORW8kSem3MSqYe0BeQw3ixA
LIfCHBCJsSxG7TgH2BU0SmIPl7TwkD5e1HyZaLCF+QqFpmdCx+DFqv1EjnAR5q0x/qXo40xzcC5q
95cZX0+nxEihf5YBTsjr91Deu3+xBkS/JNUfBD8Rvi1wkgnRdAg1Dfy35d3G9RfcDo7/w/5pm0Zf
vM6aaoEBZxbl3dFiUOEwQsgUMcloojrWCNLq6h0NhyNKpPOFuH+YRBBJRyZw3VLpYirhi9UEdMaM
Uols/Fnl4HgjFy/q95bg5cl66+SAyE74Jk/HYnVvYNnuqo4KJB+MAACZ/8moc3Qmt7QT4NR2bH5a
+y7rOJua067djQNPiJL/GbfLjFx9RK/nHrHgwhtk++6wTkPEUx4AhFTexYGbRPqw5DzSBzhEBVjM
GaU9yQrr129bciC3l3OgsprIOLFAh58z9/pflxSiw5KFANjiXTEY8YqNcY+lbsK56CRIPp5Fr4wm
cUuL4/YgG/gvf7Ly+H6Uay3yVJSW9QU17mNKrPuLOaoP2GWgTIxtWPIvw5v8IxNntgv9L+dIwatr
lf2DqjWuD6GpM7Uwp6DAXQd8LDC2e2siehWLoRq2zShC1RbrrhxvE9LYoybah/eYm6iWz2zKDWqr
lMUvubqMbsdrWuhs5U9AIPSnPXLMy9zMZm5rqZvltydov8HFhVwT5sBB0Vic518Sz0L05kyfINVj
rUK+vWnXF6f05Ebwk5g3q3ApWxBzu4FMvMCmngu7uGMqbPQZGAqt+2sbqGNs8tS2iZj9ojziHCRN
xPODhMIbplkPSjindhnbcbDf99A4LxZl7q6EJ/HQ7J0hPpH+1TqDL8k2+uuXxxYW9HHN4srg/Yd7
mlKxesbiWcuLLDf4Cw2DvAetgOkl9QOkO0C8YT2oYIIf3DesvbZuD3RuAd/agSi78snLsb5lUZHL
FweRJoP9mmlpACnczGLyfsKs1jJetzmC+QSGnuuL+bXGQ6Mrx1ekmUuhauSxqRFB31MxTWf6uuUS
CJybAOHUXUMzQxPsiqXh1FL0odjHLWdXuKZmOKKJbyGQF/HsyfyKpHDYGab4l6Pwc/FmbY0GvbBs
lnbMgBUnSYP5jnfAHhYS9Nf+ICzAVv3mmE0LN6tubXxdTBmedZCz4g7zW+fS8ycDBznFPygfXdTj
dtgZuM4KclsRvK0mHZNQ3X/hjrS39cX/zta/rja1BtDrR45SKBOC+tsG8VFRoaW9nrL3Po/zOaj4
fBxQwvUGhXVGTtRnMrz7nQE9b2C4x0mmmaXKnamqFPF6wj/ecgmq2WdUTkqMvVt3/aI9MRTK6RZy
1kdbV5euhb+pl7/Zfs/8PPDqkkEt41DdGqPjFbZRPIMsYitvPwiuQ/ItrDaZ5yfJq9geaHzLSrkL
aYYE5GU9CCRcKoTPpsLKKHyznzi9HYP14KqqdbzqEltHdbKJbRg7GZEYpYxKAaVpUofYpjgHKqDW
mCsl7f8qC+VSgz1su/9Xh6QUn9IV5q82ilkPANc4j4EpaItHXNwR1cmYxtdjgzVQxfNlQ/SKkR6z
sOqeoUSm1JockaSOwLuy/cbjhnkwdM6nq9nqeF1T5DhoWHVeCJCJWgud3bOs3LQtpw53BxsppXFL
BZfbmYllqo82qze8lzdRD3c81TNA9au8TJMT4MlR2t6YmepEgD7Xag5uqlEe5tZSllG3MQBS8pWG
1DUiiDLfAIy8V2iBGaTDr8seb1QBrpE1ClNEcifjo1e5gMthjRDnhb4s5zBoQuwjl0aFMQKukl/z
MXzI4uUWYtV0qN7HauOjOV8xunkLhiuESdfq/njsm8NYVR/56hIKgQ3OkeNyZW5Ads0w1tnWHQY2
HMKKQ8IyNiy+JSTfy5aIHIJO45UGQiNx2bUNF7okAaGqIZ1krexAr0pu9Sse42eDNaSAsluscYLR
YED3sZUQtcahTL/BxttAHPzLFghncreIZvfvmsDtNnzDBTcWP3yeZ4fQPoIIR8j0Y3gH8PI5P9Xg
fploFHuBoM6z3d5i9BHJQt09570pydFm6m/OECtpkBaWMhxNxPfiNNEzXmF05av5jw25JFSIzG1R
dSjgV7GAqP7gxshc0Q4LiMlFdT6OK77DvVr+iCXJHmWTJsCcKH9S3eqzNgbmUhG7tICWnnI294wN
98DNACcESfU72XkLe+2321EmBQWIt9v8kO8FqmormaSsWzYYDEiM91ayyqR3OpLfiO9kv9BXkQuj
8W5vxwsPRsyKtlqg+p0diWtA8LHmnCRFfk36XonPp+BXkEGHWT5xsNKVKNF+BO6FnAyTRUCeivuh
1onWBcyor+pZx50JGSyoWtx6uLd5S54foDLMS6s6doeEPezSdVClG/ThiTRxAbAtD7eUYbDnogvc
jronNB1el6jpWDu5OEuKeJnKAl1mWD+LdOGyQ+z+qL3L6bxEBB/2WJN3fFe3C18phn3iEYo97QYy
Xai/kzeMzGz7HWvCPsJoX4BXp6bh1Rzc/Yg0K2ezVC+2rho+sBGECb7IA/ElLKYB7VJBOtESuugm
esOG6+eopEmRY5FHgvDtWMwPaEadDHeSPSqdQLzeCs4KNbm5Jd5ewXaOZXqtoGY3yu1RJGghsEQR
1AWQMFhAElFMcqx9qmPaUdx0nZhWowWIZiHTVJip0QnS2XldqDedqSGXaN+i1djYOhLtk/1FhBPI
ftmTbw7nfhdDJUoHbxRrvSkjVgJtMaPpjNFr/7E8sTyIDZdDPUrh5G8SCT6dQ/VqKDltA4N59pR4
MgypoFaF9Z2loNJQw/rpbMveAokp6rAuKp2auc/aIeaGhtHh0PA5Wddr8OJ/m4sArzTdgYYfpPPC
WQ5j3A0bI8rPBcledUaP2+V0vUBJH971fzFLpxK7tXQjEhPRmwbxvwmdwD8zPDUANioCTLcox9IJ
b+6iBNOOrL4VhjQoDqa8A1PAiJYQaHIqrdgXgW5YLMFjhMwehiGzEAMjroP7qVOyedw/OwNEwjIH
wJlr+dfgikFloBfKyPO/frT7gtD9KdEBpyrJVFjU7cC2IEOaKV9h1euJ1WjBco7Upjvdkv+XWpjF
8L+3JyJIMsurTaz+zzx1It69BFX5skUlzvKDwF0bI47Ik4PAuEGp5KcI5BixmmX0/dFPxOmAZZJr
f4h9sm3F0x2nW5cWAscQiS9GIp3q2FCVN8Eo3ztQF8FuHBhxZpneZ3KzT8f5mUJP8F3RD37ezfWy
crvS/nXPTlcVEzUkj+8PL4Otf9LDu67a7B5akKFTsNRoTWE7GooNhB2ePGUS3bjx4yVPqFxfisHi
WvxfV2M6TrBQKDHQaEELIRUjpdttgE0oda+mgxE7q/+bTZtRfp7ZXesFa03EVSZIwHI8+Ar6ID9m
0oXyCs1qC+XYnwGYLGTD2I2I+Q6GLMyyovHK4JkX15USfdJ0vTm/k6/cS46HBXURzPNnBZBsk9HG
UcJxhU2JmiIHK3VU+IzXjdwUFQeM9x5erVD6N8bVoHJr8iQ7l4cyx1G+pVnH8yE9VhmJNwaQj1VJ
5z/4alDes6cVTu0FPtSisx53TVWBdl3FfZ4s7gG7qtMbCwjJnqit3n4JMYSlI+okYnbpizbGneL6
iyY7uSMoiRRK79lVj6MDRxcxrsjc3q6EppsZKhEMyMplqsVMbF26Dp5sagIZdT6zzr3cg4GZ0rTk
TjzL9tQ0FDbsVCcoWpRl0AGTCN18uw8zud1OSQK9xx3ol80Y+c2ZYjcihTmSAPo1tlG/0ZBsjVja
jFklX+z0zRqrHK4EDXmyUm4en9sWDvjQJKav6KwKkdDl32nWPRj/dt04XGuWj89gygUN+tec59+T
i6nHETxEMfCS8jw4WIW6L/c9c+mP2aEBqsWc3afvDjPKqLp1/MyI9qiyfkbGs9LKjYXQnDtvUUps
HggfrU9uY1pBzWDGH8VRDV2CZo+52KfHPZThyKSobenozpkcLqa5CDFwa8S/p002NX2O2mzEIF5F
FQ8ATVYjO/ExEhI7tZss4Q5jvSRHiUQhVSrExxMcOoU8zmIva9wUAuibBCAm3u3Fkxxw0zECfwC4
iZNelVct3963b4JInUWbbOdCV0r9USnefeqelxPkFJi4MhjsYQDaI2Y1uU37RC+key165ehmIkZX
26GnpR0YrA2jJGvtScYylKMGKAJvtK9Qe0bV5NTqxVsKPSMaPDM3MFNgUEMlea8kg1ZLzkPW8OWO
50lQlUSVA0w7553SBdU7gevdxSj1ofPOy/j8Xpx8exhJQncYHAxw4ixmLvcOZNkrlXFepPveQzsg
goD2LgIz+0PX6GqVHKAKOglPVM2Q9ht7gqwN/f+3x/SRJMGf0+ZfHF979FAHg+zoJWqmvCajINwl
xbXQChtojhSkisNcUTjRKv1wYZlc4hnHLA9NHrnGS2BU+DXNByyxHJGuNobb7kOm9u2lUupU4duD
72y9HFSqGbncyG4ToYp0j2f0zEQ3M2PWHqNACZfuzFM2xwawml6IegWWJpy2hAHF8anPckidcx1i
pMabWNnBzPOWkA69kpBYzx+1fTboEqPF3tmL0RsXivJ3aot3RhNCpYnXrQL2u891aXmcsXmaIiHG
1tNRcvqCiTHxpxXaP0oA/Pwm7KPMS7D2S4jNABRfbqRlrnTZ7cqXpKZ3PvAzWPdt/kq9C499CZfr
mi51UerFIa3VX4rJQwX2KzY0mmiHehxxo5XTXZ2uyCKl9MOIuSc8twEXxJBtLIv5yEzMfU2l/tCK
iwGuKxU9oo+kIkrqwBaD6haaZobJmHN30lwm98kFuCfExQLO8X2WbMBRGHywTv55o8bABxkIXDip
qeP42Dij2XY/AQC0XYG3es+MyQ0GHPmELQoqv/Zl6bZYemRmckkIxWhG9STtmdicWJk5rE5W2I4z
JWz2TxV1k+NaDwLA4H1Z48rg+46iPRDXMkg+GFCoX4z36KGyoY9PDEITeoY5Mj0jzLHHzA0i9aC7
3uDxmNDF/JwjDhajcJfTgt/XVtfhw+T2DeZHNxviapxCcSA2bJbUrZDaMRGac62+AfXkrMVKqjzH
JEqWfbavBwssWOPjPy1dKQ+yV+xkVMe/RkxP+iOdQA+5nGRVinKtyzp2PJj/0uOAwHS5qXMo/+Pm
5/YzprCeXerK6Pgteri+W+/p/DNP6uFmKoDi/rVy3UQ5XRGI+V7l4FtHhGBJRl4xdcpdx9Vb9IX7
jnJira6MKSZ2ro3REnh5VKfkU1TBZq56cZ/nu/4AEZX1PnxK/dzge/Am8q/Na1z1fbOrhBE4WVoR
ZddVOJHInhecaoIzFnI7/OEmNITpA57foCDv8Qi6FZIaMFehqACTf8UP8dq+Zze3BKfUJaVg7dS9
rTr6/8RvxCD5Sao2n/Yv9C8g3IeGtQHw0L2s73m81qjsVniDP6A9hgOCAtfFnwDAJjGMUSv3XdGR
ZpNmfi4iPG+OtvzwWR9T6OlIy8YE2/pBfw4DovHUHqEx73SoXoFZSBTtS6j7ehaNid4othApP2xZ
Z+v13Eko5t2r7MCDHFgmgHMRnMB/Ii1tmGmXxEBZGYCC7sVakFMd5tUfDh9xibHlc+be3EiehpC2
7ce+F/4bUYDnravIKEbxO7fkCbUSOjEaBXxzfl0/nKHFCWSykyV9AXOpVMwivn+lDgDJX6IFqoJJ
jkPkHku6zBqOCcvAc8+Zo83xpa7CqXlKa4LsY+2v5eZxOdJmYHuvvc1Wgi7BvJ92DFocnvAeFaX9
ERhzYHYk0y31i9kpRnFjsvB9/cJ6z93WZN2Dm34YJXds0VpUNNwfEd/0xVDjh7DT6JGZDYRGhLjJ
VNHNXg+x1rQPY/5/VVb81zB1+Apwq94QFhSbB8hqIQCV2xeH++eK6h9Ny/yH+a7TdP4D8rli/f1b
RPQY/QPACV7TcU9GzH6i2AAarCoqRYNA2rUR8gMW94rI6PnWsX2eHGi53B/auqU1tjdR/6ntmo53
spir1UhrgACuraAO4tCSLGiQDEOCRcMH9pmD84hHOMhtrRH4nDBNglxpktgKNdlidW8vS+BwfdbX
7G48v7b7ZqmQegXEvfaDPuSyXYeyfyJvcD9o/hOzWqvMyOErIAPOT+d6Dyt+oczvuhLSEQsYkVip
ChYb6c3mJ1jmntkvptzKdA2f1qtLLAA/qVoj0tFfZn0CZdWzUnZ7JEkUt6kvM9L3G3W7Rpeitgio
QZshRWay2zsNMoJPEx8jNqCRxDb3b2oOQMw+XIN+hbVfbPxLctP2Gz4czjc7rcAhN9mW4S0X+DHM
9OPQFX6lOqmZFYDk5td5oXcXDUKYXqfOtSoHdQ/znt0GWtVu3Pe2xcugDTLThUj/QO63aupN1c5t
765dpmI/QEJzg29QTAy7Ae2umBLBKWteHMnxBtl/aSpwN6KNVvLb86SoV+Adg+jW57ZD7hLCVi4H
rtc7e3cgHWsYvQu7/4agv5hAszqnesEJgIrubQN1jBVxYF3pPlJznEioW9I46VSEHugogLIC8EyL
nTLBfNBZ3fqVjna2ejuDSjgyUAbtyp2LDlGk34CvfCewgh6zcu2uuI6/LXL/hnrz993H65UgoqBr
l5UU9ScJmWlughjPuAyxCPkwAVqp5TdKn2OzlfFjRvyk2V/F5MIebO2blokQxzU2/DOokLuqmJTR
9n5PXkbWQ7tGoDJaMT8DkpAGfmW5BESodQxVodhgqRXFnH/m2U4p8y1Q7NHNobF2QtgmhysbEL+v
Y+qppL35o3iTrelcPdWg7Me690i5Wier/ph5BDXxOHYFQQ7M1Lz8aHeL/yqKgzRZcWJxD297oF/j
t0zNMI0wubYJiNMRcIYWn/deLFRcVuMjsFs/VxVm+bxlmEXzdn6/cgXINlyBAjsWiF8uzs6HLEU5
ERPLU6xCsoNuM0PTysjYidxdfTxjHbwFht90SN8OS9r+ylwwi9XgG50girNfaRsZfCSCemsC8THw
8yyocjvZxMAtWOv56EoQmqQflkY5jjaA5HT6MgEDYEw+lPuSLEqJB/1A1K4KdYNL01Soa2V4I/X0
F0Mzr70AnQq/oYpr0Q6ayFXAx6Q5/Z5WrGDJrftEIGZUaZFRJIvvfvsNnucmOSzWKMaoPxyGfNOJ
K58C0mJjpE5gP/VY2L2iDJFZcR87NXSS3YriGdBI5Ll0/Az8T8IXQi30GQt7IWsQGYhZueowmUAF
WIGG0zYwZCGNz3uhXcRG36U2B35dR9EpLu3JBUKfLyQaCz6zx8t7gVehZaPzVdpRZAVV3it/+fUB
w+pDYgwOMmsPfKOUFiUAcv0poOBDaswWUVhlY0a8pl7gxbKn6WQ7OiSmnJgeS0Ypgo9GbPhB87Gq
tea46lxn7y3E/Dbg2QebiUSbIdFRNAkxJRNr/EaHE45TOk2a01Ql9evdsxVRA+V+6pQPUrx9Ce33
iG4C6C/UCef8sC83QbWKT2yfvJHdJ7/IUvEQ3Xu1Ij55ulqPE4MdysD2jrLvp4cCks7/2ZrQdkc3
td3JaBz3cO503KgIMPgDNXes9/WaPutZPclCG9oNLUHoNEKvR3o3W9qVS4EbBopAVXBSsDZCzito
Fap8liDbUsnDJX5sM317+KgUoS3d37ihlr4ecogGUyMFFiUDto+bRmSIi2+CF5rAmAwwG+CH6AsS
mLENdAwbiugCmDtfuo47L9ZDY5eactOCtUoZ1Ix2rxmBSSNMNMfYuOAdZhW3Lww4om+07+5x7MEl
EMthRVnG0talVi1YNeob7dVLgpnvUstSm0ndDMvn69oP6eArmD5M6eaC25JvEMCxAdL3t3UiKwpR
rDe8A+n3vRxoAb2Xe0ZXZG/fWL8tZa0XUAxr1t0oVR7vRbST6A6SfkeAKY86UktuW1Po2i2Mmk76
/EyEmibPQhwo0yY/gmgkxtC94ZgMs7TKZKw6E4V1X0cwywVCZ9M1j/R/Fw1gZ2XaX3uwSlPZ2XIq
NpNLdLCODbcIvk9YZK3r4xmhfEcK01bxVxI2Cm+sQZtwwZGXP2u+qH8naGIjURrGP7ua2YTzHsMv
cfPBkPYYRim3rFe137Ek0pMcR3dpRHCA+/Dn+mKudb4QektcwDDUGkVFb+TxfyOFPZZdXofWboNB
DzfF00PrFnylJWmiLVFn98vYZiOS2HF5H8ZnECV44iM4DrF/3wk3q2e3HTjYlTqXUWMe/3CK0ZvG
PWp8XU0WHv5YLargj4U4MFhKEkIT4ANxYpMeDlKz7ohJLb7ULRj/YUECL+fozrg3R9xvMUGTvbe3
pt05ZYs8NlFp+gob/90UhCaUFvCQsYn5r2p1rvjyrjQUVAufFKyEjuYn/CGUJ6EYuej0TPhIM0D8
yr4hK10oHv+toXaWGfyKB2QuitWlGcxiTnFB34ZmG7kDhRzq2UujgAVFN/gpwE5j/oM7AXF288Nt
HMVeB7Rl5uVqAGl8GkBAb5W9U2x4ebekPkpd29RwZsxgaxWhu70VjTpDyt4VYOq1omyxQfgu7Guz
oJlD++kW/3n5OKSb6sr9K+oL9cFDQq7FWp9lgmtRo9cImHcAY6CgjR4eXiGhdeIVwjBWvPLN9aVF
qS4GQjstH6Y3Z1XnIyqRcaY+yvDlVAvK5xwu7fRm3A5QyfwxSTqSQWriKxqNpwwIW3HozTduqU0G
uzv4GxGNiviL5YZiljFZcvwZTxg2Ry3OXqVCku4qgje9xce5XdC2Bj4glChBmZyPn1RS2eOzzfs+
bHQVlqCvV7zIhRThaHtEwaL7t+ZUMH6gmvksjEE7qDJ2X+q1Mx7xLsnlKJhP7fcvSYdHLpltZqPf
JPqRZmZ6IMCNyhbz2YBUrOwGPCcLVkRmRTWXXZdtr5qdn2Y9pQs/BHrOOjWSIZXkbH0T8YaA15mw
LEO9JiFD05Xw1ByvsvLlC6Jntfz+LsfB/fVyajYCBv5oL1KoxKl2p/Do1uIQLXtwL48KhrDVAn3A
LVA5ZXdxsHjIIXi2sRDySaxtFYXe5Tzgui/MHKLvPzyrpn6QxH6JpTsnkx7sZ6gGgQicTOWTQ9wz
oh4yPYfxR6itzDzZM7yzQM36X9fp2Mx6cFghwy9c6MZaZ6v7lufDP3dmxemRAbfovpQOLdAOSd7O
1vggFjS5h8nr21+oeejA/Y1R+/ebbSY8W4P++0Zf1MVfsg3Sk1CdDg9mGI0OsF8LlIQOdCM0Ou7S
P0aTd5uq3Ce80BdyR87blf7mkIs8zsaZuDAlZTVnSq41dpDwUAU4M6+/5uABGfBkqXBdmAkuH73I
tg/TZ3FfFMv6mBrL/zWkdI/cxBXDUR3iIf8BU6E0tqVPprUH2xdybHFaDJV5uBAXiUfNfO20p0be
AWy5cUYHZyRlV7MvKC+8yeCeLPh/HsjzOaLjqD5OX90amr89D9IrGsLSJkg/lD6HHHv3Cdf897Xh
lQ+Ithamnyvjl9oAyjDXYBqf045i8trfr5KSyOdYKVUz4Jn5HUu3pk9vkiirnleBRbOtsVlj4p7T
arwF7qNXgGeD41RHLYO+OG9eRu4JI7NZoJLGcJo3ypBcVPZ8ZLV6hZ+a1EqpJbzq/LcO8IXpEdZg
Kzjgcj513fy5mUZwQcg+qRIQhWCqdSfgyQLSlqCpJpJgFCtxFfExYQHE7BcroYsqYNA9bQhntPdK
cgogf82Ar/vbw4EmmH80+nm03Cm7zQJN6PItWtAm14wdQNhTaXoGb6Mqtx5vAIRs1Ddt2G6lT6TH
gjFsiaDT/xlyqGWafqrMLxiyRcL1NyH3Ppb+jFMy6Qqb+xu1Aln8plTzolKUlACJqGA5ANEItQ8E
kxVFeuro/pWj/bBbYUrIgP195YlTHs1KtIOA02+SrZUqYwKJr9Cw7r1itjEg+mS1X0RDGAGyG3Rl
vlpXmziFvMdINVheedZZgJfQpJXwJD14ZWhB3xznyzW7hCx76S+PtHxn2okyOns9KsQSuVf1E0H1
7v7vxA0Atyn2LfuSu9RBCbzkzxcYrQz3rbDYu/B4qMA6POs32zqORC6mhZKixDvH33+gyznfQUvx
ryV2NDjSl3SusnA/0OUerDIfKNSY3TDB1Io8Lx6Is6hoC1u31wcuANQv1ZDqiYxXEnnrb4d3abMA
D/5UcrNQzS7iHIClLxzeII7FqqtZCQDZT++nuwWB5uEfW2jNFjq8g9Zayy0yCGM9v5hWzpeaRadi
0mluVxJ9LRInOH3J7FFMuz8ZUOmcsHJEd3mN9hTm8fQYX8iwqWxwX8ShHcsbact+aqpP7ZDNFRv0
gHGMXbbIMIksSmS8ggy1P9zHRohObbrE1IKOLmucIlNbtJrSArjmX0eZhQoZx2ZJDsatHYF1Ym63
KvpangAFjj8IZhe+5fMnnZQ5nVaxoa1gCRzGQI82T/1lZHdC9Ps51ZTiislD9+MAaPN/RkJkmlT3
SVYaKAQ7FG2b5jVxfexUhdEbAK5zEVnkbp+vYwuE352NG7gjTKzBOPl5SHayz0tpK1QTg+VIZiMi
uWpO3zlHhcyQ45JOsE5ULpdGssIHIVCH1ftaCKgSGpnqb9qFzh6F7mMxWqzPB+toX+Ys03bzyQ9s
zwL0wQyplT7Eg1E+dxKLovXI80wo4Aby+IwmNicVVbHSXrAR+Qbd+9TJJjjelfIPlhF9t3jtQxQZ
p944mAb9PDBstuTvfGtIgrh/KjzUkkP1C33izeOxZ/n/AKy4bQ8nEPTKU47tCzm1MBTidrPkLr4e
IQmedRNdhj5Q98IQsay765ENbp1/KdD9Vf/w1e2Wx8LUH7R4/3J6E3ZjESdvqZLMntZ4xDm229NN
CCsevYBI2Q+ZADATKLJldWLQMhRnKPGPj9gp5VL/09JWLWdZ8HfmUH8m56e2sQlIZFdnVWDS3B4S
CQe5ANXjaJNNPU63X8aUmsbRjNtPP3p+uu9nSQR+VpzJv4MV2i6odFyRDtZ27/m7gvouqCHe1kMn
GMmQ5rAEzqBOVzhEdnqbZiK76I6p0CEwVJ02wJltYW/fcgxU0Y7XfkrkWKA4dqGIDm0h05FJa9md
gf0Te5Xoy0EtemFJjJ1r/w/P4AS20Uawn8ORtii21FEf6C72lflpBHIVm4Bf/mH3iWxYkqYv4CVl
r8Vu3Tt/zp6OntOMWo0/CU4bxDh8EhAeZoLJ3ub3OaW92gmDXjGmJO5yzSdGeE1r5ONXBFW/6HBP
O4qaNOvE2IgtDUDr2SjqGzyhzkWfyIKN5gh42b7rHrXOUWlCWqsTk4gkOV7267FEYR9L3r2TRgx1
fJSk/Q6IZHoWz2WSufzWPK+FFQv46hhIDGxUlh55RHlZ8U3ZLP0IvkNxu87ON6VOLpmhUprbOHsR
Cp8Sj/JlhTLJGMOtm7gvcbZCFaZ8zi56uk8YtBQbVSUMO7JPcd4jUJwO08yMKD0Ps0KN3zQew8M+
Gv5doVcj3quApFCzF1VXiRt2WmS/9wgzi2F8Uf6YyaTcBbSCDQh6XXp2uDgoiXo/5HSRoldRrIZt
a8utGJn6VmNT4aq5q8B3UPV/JJfSdwY8b+ato7i+qM4EexM5jbY7RAXV0afj2X4A5hiiilySEdKc
1gVfzW4CP9ALwQ0n/GQu4j+SfXT4rvW5Q+0eBt2cVcBPJAv3Pmps8fwFt/J5wVF+HH0tVSE3p7+Y
wnLD79aXHshutFBEBqNAem9PcHbSljCvh0fXgfMseVBQBK7Uw0p7GbjxJD6LkQYZlZqJbE8Pby9j
qj9e6+YfEXoxJAZxmY0yLlQ+0ZstxLTtq9oX/fwomUvy2oTad7GbI2DRlZrvhASd4s8PYaSJz9F6
UsczkQRS/C8I/Hths4EfiDBZuUpaKIK+C05lWPHGw1D2b+9TRoNJh5/nfzAdq7sU0eEcbHHWzq77
jjed8TavpfbRrkpD/zPadI4RmpJZj1/YvygEL0+8YpLfDzL12975J/XOp8p0dPtm3vhtFo0nlQoU
CscSWhiqeYX04+pR76BD5pohgAGTMjO/apUGdfmuOpJ/9aYfjDyypxAfd2i5Q/WXhGn+YJWYDrUU
v0jtpIamW1o77MCRY8k1Wjyp1QyjuQjVMm1bRvaPBgSAmagbyNjIRg3azKM8/u6ucaqm6MQNbsda
2nNmweVkQWrGJX7njwl9LqXlOqdpoEmhwtHn0MSjY8GO/Zzwo4mTncEb60JKZAoDMaJs9TP+TehA
i1BhjXAgPdWX3+gNWafyx0QbImlnaX0jtFDIipxCL2Sma793clg40VVRe66zXl3ebDN/EmNYSy6K
K2S24xOT2nfMdUlFRMcl5ZqiAY3a7pYx5bEDxJeFwmSnCsxfXuTftTticAhkr9kRXcIHScD+0J9L
8DLutxr9P/PVe6MU14fxCa1WnHCVCZjMbgiQbTaCyqSgsdArmjhg8x2j+7JTIuwM79aP/i7B7DX9
k8fBHGdinkO7KbjjseYHJF3MoNRhbzgughzIGQrmxU9XV7GeRuw9O/pcYapE4bDJUjImiqWO9aae
uyPdp3Tw3lDJ1nkxV+rIOSj+CmVT5mAnxJ6e38TOsUCUyJD7zcx1x3ZoBtNZ9058pgmDAB6Nza6q
Lz+/ET/OmHlFRN8d4OVCUKbaNkKnZMYV6u4ob+8S+JmNTVkOLBbxIvTlMUa7tuK2e1qhFOK6vAe5
Uliv/PKmjeKiE7rco6vY0VVFNWO0eWu72x6U33rby+oscshg4klSiFN3Mh5VR1qOAT2qpqVCcz/8
xgJzvtKcvRtwvJdRHFupKp/dl5bKC/WAD5bzHogewU4DEarbTdWPR04Mg4AHKP+PcvSOxTQ0DNKy
IsdIjRzleet06bIoem/kAUV3ri8kn8oc4Vl7n76tbucqWnJ6PSNzggx8mp7Zj+Hz6qi40V/4P4nD
g6GlyXIt0a0t3NFq7PWuQ94XuIIpcrCXQmsSlz2kcDeq1XOa8gb9pC+ma1TRgoUpoZW4YCiGNj8k
HlRM8qIgSNx0xTLE9WCAdLraJ94S92+nHKosaDqWLzqs68DGQ45zNYXfXY80mKNcn3IyGqqZem62
A+0EAV3Jl0SqS2s8VBDIOX/Bky8Hcq8sVkCk8SO0b7c6W3k9frFNNv1ViD5FHgFrpgEAkWccqL8p
nXwidkzTEDq3hB8dwdhVZXZ/F9X4kCDVPYqGLcapomxiJDQ3ZioCmoXuGUPQSew08eE1J86a3UbE
3sWeiid+qe2cGG7wPvpZ4SVhjB1Dy1e8U4iEP2vEAo42HEbEH0G3MuzuQYvR+keN3/vbGXiHExOh
C3DsaFFb6xyO69g3CHItEV/Z9RXcF7+Kkox++YlFp5i7J6NGl948CIPGaVvAcmFV/N37CFmSfLPC
bxIIxLVChgpoX8eoEFPSCz84Mrof5VY6Jp0OV3fORKwDMifIgOQyJTz1cz53NNjZjaZQl7sN6uak
VHKDPQFF5bcQhUnPfskhLbGiUnygeym8M3MwnmFyMYCf9uJzrSb1Rd21GSaYT9k+fqHf5J+cJdor
7396kRpxXiCmESo1GodlHHrF3jQrwXPCuLAb8jjJMQbllT8NF/OVfHM3a+5EvhvGmiHo/0+ENR4e
OdgQJFjeMJbYk/VNa6avi/BPPSMW8wlWuuv69h4iytEdNLEXySe20NEHLwfbw3zmhfSLLRH4GoxM
QSZT9DQ7IUnhZYfxlCdUVeDsllMlZJIiRHsc715/N/YWB5kUzNj2tPIk0QQWsWsOmQ0JkDMJT3YP
QpOI8vBlIv8Un97uzHNlmAMLbRXOmtA3X0hbTKBr3NejHywXY6+/qGgkV4FDvPxisJ6KI3lodycK
Mu0E0sgiSevBXF7c4qWvKjKAaYvufeNd3+xlJKzxZl8/bZwSYkvGHKFVzT5boYnyw1FVSVI/HnPc
mTUmkhoIEi8nMIeDKQjPnnGC8Dzyk2faAbu+kVXBhhqwyIXU8XsMimo4wqTijVgWDu6c0OulvNyb
uXkof1kP4sYcxzNWyP85AyXHjKKYMDUa/eACu2zgw/ChOdratcNyJXsfFgY9OrkGeFNqtmIC7Sf7
x55aT55fQsUdS5ymgupakXF7fY/MR5kFf66WirNltMQskE88WZXRtPmwRuIczszqbg4OaFRYoPkx
UJYFIFRfKQshOh7249/UI5/LqJIt+y37ZPTdfUVaRdhjniPHb1VSww5yzC8j1cwKRQnuRerEnZW+
/W0XnDdhLbuYJiMiJiBxeanymlh/VI51txr1QTg/KhfipItQhK3Lt7HKzV+Z+zZwtzCNKXrDPcpA
vDI/I5bpAHpdl9tz9KN3ayHuOlp7qgyCnwNrNZriI2rfU/n8Arxu2+JhvVidPRX/80ZIaAPLY7Io
U3OsDm0iR3cxGN4vh0BcJ9a7xfiinhmNzb6awhNNvEZ75y2qQSgtsaCmrAYcfU/ZIR103zRI2d02
OsUSBNrD2mTKSyNzH/zfhNQXxja87u2YKkgLSgzmif0nD0iRxi+iT1/grxzr8BFruxvV0QEpbF8O
512BsFZ8Hw1B46eajZQPjs7PAWwhNzds7FU/elAnYUYQFMdqqY+n3ogzMu93awc3S0L7Ji6qlQrP
vxYuPNWsXGFL7zT1qugPxLd3cyutNgM7XORlXDsFWd411A+vgpAtwYXw9EqDxQKUYxVtXFcH6ZtU
N9/17fZY8idhTkkXVMwHRvSPQHDgFN7ZhXeCwCHhU1Tf6BQySA83EnLJGOpSUXwo8fv9QD3EUkB/
BRh2OPTkGJ0AOwcXyGJCdZT+iaPqWlXCOzR+36mmPar5CHEjudbyAzKD5wJVRRFeUk0eGWH5uBil
mMo0Hss2gmcGeZPjypWjB3WX99g5WjKZpmb/jo2n2MWLX7GiXY7o/BEl5E66LaOD+SDTyu60QPXg
sx8Bjh1x6fJFPBkhStZMnxCEbxyjSyUTVfvGME6UVVkadlfoDttqh4EEsVYN+WgWmESeqx+xiTrI
lcd4BN5zU3Quq5KBnlWQgF8soBRu44ZDuQjsNTgiqf+6giBUmm9Misn3+wrHc/4Wo0Y8mYWJj3W5
FnTOW2sdcxrwN1UnONVKHghMYDlbv66bn61vWVDqUTXiBIKfN7Wy8jY4ht9n+axUD8Iou3ryq5RU
DO5fjA0BZ1V4YQvYYiQEoXVBStkz4z/xS4OLdmNV5v7ioiv0ZPtIcDUDi6czBelENWwy76QUqpIS
Vtz9Ml1pZfya7DL86hmO7bulb2AEsvJz6DM/q9ZmYJFRUJMCPhz5s1KHbhTIz4tpWI0UgFdr4NoX
HmiDSybdJ7vFA/rI6SyVjwpGNyyx+hHmm7pwVsygO8AOBJfpgXEMi6ZZ0PcpjSTP4C2bc2j+Uh5o
zjqAoY4HvPy0P279Y61Tfb4I/oVKUUKFIpVi0cBI6vjOS0pac2RL5pRzl7FbDIt5blbH2j/66VYG
VxqFId5H1o2TPPY6lS1AsEgLR5PgS3dULlkT/BKxEGhFWlBzzTMiJMB0/j2m5GfAT7MLlUw9Bs9c
EBl7BCE3un2yRX06C3ObgLZAdbzxWUDSAkGhbqfSW27QxvOST5+JQJRL1LP6t9qJrXCzASjM++c+
BXuZeMN9AykK3+VOsN8zboPiYZ/lNAi7/Phucyp5Xe9NoUjZzrAd/oUHQNohgBLnRfzuA5N74eWh
ijeaqSvA3yJmUk11tWaNBosZpLrjNvaBv/hQiA2msrfspVSIbjfVLalSvWqRbCWjqdK7fJ87d2W6
j6tE2ufj8Vp7E6Bn2KHa9/Rhxew+RpMD4CfW4nrM8l/VlS10C94kHHlNaPHS047gt6lIV9FMGVSy
xME2uGdJFX6dgPGF35xWk0jVXzAOvnSPOp4qJvLDUVaGtluj0bJNX16JxDJJ3FOILiWbcK9FXdrt
o1/AWTHnIKSLc2Kj4vXk9YectXACNsS6rnJT/qM/8jSAy4cT4r1dFznh343lOTAj5FqvmBDxv7pB
2jD7chLHKjVreYQzm//bBVuFSUo4Zlf5CD1Eo5I3sru87GWKNVzCX2muq4I3HW/PFpXp4zKsIAxF
XQiiCWfk/WrqfvwgQjw+5A953J1eccplrX6EoPNJToywP+DDKpbkI8jPpHMZtJAaesh9a4sdcvB0
9OFBZXlUPcR4SVPqR4iKZuT9nKSdBNhPSF5SmY1EveWF+7fBmSJg7Eq0Fwxkoqp2N6zDprbLFaCZ
WPk10bK/QlPSsOLA0z56MPbe2NxQUWBhJEEFsMHG0DCDtlKEA02tN2qfDGGCwUMhepNhIrIXa0/C
sL5RKcfZwWZpu62rLDEsk8dg6OdIyHmZlLWkrDc9p8SZQOgiitAbwT84dHBn/X++fawm+gstfAXk
nKaZQzdHkD4/anraGM89dJhQ+SwhjctwvjKiTo4nLvo0GcwQizNhfKWbL/Vxnz9RN9vs5LkAgXRS
MFpsVHiM+zUwFU6U37H5GSP6tSORJoD5IjDdwQq3an6wxy6JA9YgIFU7+/3zim6mvlCbCI/IKHS0
J/sk21SlnXjAOovPPz2pWNOvhOMje/bTRuW0JBBqN+nE3FdItoVVGPl6gXJWLDKhypptRnStGeuo
s1Ycf3nWXbdET1POmYNM7Oyl3QAY3G8N5rVhwlA6+z5600BhrvJpIeKwH1FRBTSzOa1QLNghMcJA
FnkLb6a1DgdTa+y/29ueEajyjsRt8ey5PCjpoHwqIMDIu2iNTl3YNEHJDZO2YSqZiRrwGk3ux52T
pAA7lUbfqkviVAVaKKAtDJjRtnp0xjJlo7+QqWxM4vdV5FymqDpuMxJ1XBGnmlAdVoBvG6g2rpd/
WkkkeclJKUAXz70QdHD3nuicJ9EyIxRpVaEpas2Eg3+g9wjAlKU4Qk1Kwl+VG2Ka4MnCTTKJ20td
ZAuKaPdKhj5HrJa45LdRbSWNZvAAGYqD0djgwqBgofGQ/kQY2ZxYbbfixmJrig1gvhYVCPT7akAR
a8zFMoCGAvTq4DBrYH9Nlzi3nPsgkJqlihpqTRhEtop8bmrxfgjO+pm7IvTKKNjtRDzYm0cocTJo
RClfKPtuoklP9O4Qr3cgCH8qeaCkC/++ecjJXcdvn5Kf2SOQUKaTbOTegYylaz+S9jrzcPf46qmD
ee3DlsVFII5CpKVr46kb6ISqqPrGlyv73NuW7bw+ohlyCPLdBymf4tauQXRAUwefDw+s3P7ECqaA
AzcfGtHoFgnIRzdKeKs0NVrMY+QX7vPxIyXVom7jO7VylQ8Iuh97JtZycPwEWB6x8CAh7vAJsE/6
c8G2Q/mYFTza3VlRt8eLghYzadhB+RtiCr1DHgMFV1Lxip1vP42ufT04RTsGKiWkccVFMo7juNdq
EAIWV2ZcRK1nFM5+oWWcHIzwLu7BFi4Gw5znfKG4Pbo+BX/9eDeWEYdBtwmvCbYMj7jaOMNwEU0p
vkDmQTVWkw2R/hQqhaUF62VDYzkBv1fp7xZgaeSGRvRqNfJX9BxCHALJ4WIWvVwOZLEWZUM1kKyT
ED8qGewKBxKPuAQNXqfFOoewAsC+o3Conp0wlUYBak3/RI5lqj1wqqWWtKFc5yetVzCXJiOigAWW
XTDkbI6YY93RBQrtP/jqVftSWjvsQuzmdxZfveus+FpE8HL8BCZUpoX4FA82CP59R5j/kOuzbygu
3OSXYTKiOYRWOKTvS6bejtNUBhUIDNLKUMtho+VCFjS49hCI4FRgMIb8sGDsqpxYSg+TozuTeBSa
PrDRgibi/0wdGnoGrVVWThZtNTawXNVeMxEHqXN1z+CDf6liP3xBd0k7dJmEn362S1hvmkXwpDrO
8uvZ+GWE/ckBIjR6XvmSujQ/0hmsCRQH7KPSm2lgOUV+CpeJIP+GYoOZVcItgALkt+V+aKSPj6hN
d39l4No8io/kWy7QN9ynz7Yn06I+90aXsDv/9bHn4aIHzvqDdvDgjkcgcpDKCOGKl6IHm0nUNlzS
2qkBYQh+abICI1FV7qXomqXTosLRSN372erm6LEeZ45/LwKwGT4Yh7m7lCW/zOuElgcmBP9Ump0L
R2F0J6pLv4p6bh9W98oqtMazKlXgHTgELw9hzpXThYKV6WEoDAjdrO3u4CPT31k9KF5FlvXYXl+p
yZX3jd2lWITjiRw3YuyKVEru+V/6CTdAaxRojbASmGXhV0bM8MDn+vD69d4R8u0PDPIiy5DLO7p8
7qoAbfeTSJPnd9raflcz8i0k6FyUbs6AlStr6fO0FLF31w3bVEUWhVIKXXigqN/aT/tLAzLOLaa4
ivCszWbwKqA985L8vWeiFuAXH76HnKFRpwLCIryRmI1Gr2QNTFDNHVUZ27JpCa/QgAXdu5mQECWU
de3gTN4SHNgYlytSEmmTQ89ccqnmbBekJnxdes1m4HMU/Bd0FNAUTqUbamoZ25GucSPzKehjFr1f
Iw05YQ71tKVMnCR1HnJpwwaEY0+w9Ywt3nH3ovS0DTp1AF1bitTI40T8MjBqa7GLEAu3RvWI0YOZ
aZEByqF0UzV6RTFY4cOBjKfswGWFSqYPx7VZZuDuLhhfZ8p0KpNmxHh2pHLtuwSXpeWjxK9daoNR
Pm9DkLvjL+ux2pJMBJDgoUPQMQZsOf1LWDQAgmp8au8UszgZ2Cc8JE35FwqDLbvODCSvdXY09g5l
3mByYVLBZfcTXFbg/KIX3Rx5K8a8Z9GTfKxDKlJghKY2Cv1/QEOZ6Wp3ohG1FwriW5uedpjEBJH6
LlWgZH7TR1zdo0tOCL+t6F5Dg4qL6g8aA81ZxvwuQlZ2NtoowQRogDNrBAGFn3ebRn2CP4tHJ8H0
VkU0GqzLMOFGl2dUCWOJw/PGJEb+LL3nnnbTbGMPIZCcb6Kjb1KsHtebqP6rmsPQY1//CXa+WY8O
aE/2m8rhuo2On3f6lWofX6QulWjNLpH5bBD9D6UClrU5/WNQZuyRjyZPP4U/gWvKiWx3Kz1UytgL
v32x1C7FWudAOJx2gZHcMqkDWs9l+5pMqAdf/YTG8AxWxRIRniRJfxL3YiWXTE63z4GBXmLhBHZV
Zmn4R1iQDsoCdNp6/lcJPmroDqpXA3uJQzPzWFER0w/cuLMPqA+BOn0H7sucduVJocB4sEsrGoCy
l4iZPwC/ZxNiAMKv408OEOEu27JUw23clrQ4WLuaOZsqO3mQgw/Y1q5bFbNuCu/BnhEyJPP7zIAX
lxd4ARQpfOUgUFww/Nv19ftVUJFF1X8fHAFSrm5CMA2njfkLipL39OBChY7CWiZgj57YLv2r/4LK
tbKoN8/OBdI7jm2fZq8a75ms0Cw8GrwcGXA03w2a2CVTRNm2qR3M6y7ScLuZVUxvxSAQJjxUYBPD
YbdRx36sph0GDhCrkOHMr53theDAbxMtiL7ezWmGOlqqcIYbGJpoDXJ+ctmWpdAez1q9D2mIvNEx
Ate55M4nm5RbjwXvW03KHiPc64VpA9YD5boqQ79Nu/fSVRGBmosCyruRGG/4ABrRUwhFY5Q/04/v
ZQZdSnQUtoEGWDqJzGy9ELf50upYzPv+pQOGbW+iHkvaPIw9y82s7qVRYVCu1gl8WHgCJ3jVBcdR
aiceFwzTdA9RUwSbV3w1AwOL19nqCXD3YjLWBr/O/Zskhc487oa8sq/cvj2GYTnaIMKJmCjM+FjU
cNBVkeuwfzy1l/SxYhNjVE6I1gQ4qTLglDe4mGL1VySQBDXGMB05LlwdU8GKbOoxdEtr8d92hMcg
IJzJqXkR1kEMoJ51vphZrPLhsXUAM5879gtv5KkA3LmGVB++fMTAyG5PXho+fH7rLpk5XvaiPUW/
fkrswNwZbfNhK18bMnsvxohNW++PpxgOUadiRykMaMpfgg+oM4joE1rzu0vLx6FlC2RrH8PpNrFj
uzsm0uoJq8hhc3ZYceMeDGyE/BLsI89qub4u5kMNzKU4/gRB3uTbVV2rm/H2FsJZDO6s62w3uBu0
/Y5cOYeeAoXiTmE9nU5apJR6wWSyrIskXRDovqEyt1UdQf+HOD6kksh360uIxsxNDgRAHT9SA8/9
7kKyHOPJPgR5Y6rbq2gmWbDgmiRyVB5JOXA6CAfRdjLwgtNxLYzaKUQe9WPL1KCKSn+QaT0+2syl
Xb94Nm0E/4OrBGjZZem5I3VChAYlSF8adIHJ44MqqzKIHEVRe/7josIwvTS3x/k2AVJPe1OEQ3XS
Jfo97ZU6/Yc/kBE9QGqWDx834AtZ41n87S4yfrKYw8rsl94CNZGq4td38r24sqLS6oqR82UiCCLQ
ANVvQLfcBn/kwu8tPNKfWQ81E07jV7IujtnEnXS/unE4FyJoRsYkJOZBaakyP0NYJckvxfbV8l8A
ACw7sIi7iFmoS2BxoOPiiJnAgfrA0VwlIuYnNGwO6LAic/jyqNA3YAg0xtHPVuGCgM3YVsaKgP6/
D7Q6VUhaMESf3+F0qF+uojl1Tz8K4WXKoEnuzSDbNoHnvDtLSZMOzuIzMoDwDfdu86hA/tOIp7su
7S7ne8J1eLGUELIhDf7fto4AcSakl5qmrSXTEeYe5EE3iC9lGns5RIOKctra5PhnVsqL2GQSnHnv
Zy7GKA+ErvLTLC57JvMbaMdVYv2uX2U6AivmG5kpQA3m3fWJUcvtvm/a4rUr/uckfs+Wc546a/6m
Wcv71xozcP/BGLeUCF1blO7l6v/9MsmFqz46C6iwg+vtV4Ks6NwQDUiJR2njk0DhGDtbAkkzCsuE
HMP0dvPfEf715436LbeTjtSV4IOeX9D6Q+qhqbebNp/PVpXBxhBOf1DlIRpx2OzASomlWHAGpSiV
6R5Ni4gUQcgbe3LutyAgyG7kEzFsahBeS2tUl8R6dlwxuPXmYywvPvToZY4fm7hckZQBiy1RgjC3
Po8htcR1EHWjoG/IW5uRpiEdIwzSys+l6K+H7KYnFjDkxQ+zA76MFqiejSGo5BufGh4gpaPR3nve
G1qXgjqFJOGXv58xG0UCJyUYNtk21wmTLff+Bv3mWkmDJrXE7SLl4ZLkou6zLfNYnHbd8akbLufm
kIscMjAjvcCjfgRJtfuBOvM+lcDvR8T+Mmag2DkMNBayjXZ0LYLlNPgA81E5VTUsgKkSRAMoXbc8
g8IQYCr4ISlg4rr75Hdcq2b+FqduSGfhpQcwY4IH+q4rsRiLoSTYuSy0+Ri0HFnWessd9t5BvEVQ
jAFfIY8zxfsz15Adfv5h9p4PCSuufPOMEJ3MqDPnr7r3IuCnLNr1pjewlUPNv8hzG6hnx6NqzxyH
OI01gV6NN5zX3CFIwzX3Y9RRVA2qapAN28Ejoa9BQVTQQh2Z1NOrCs8Ng0+/zJlwDRXlb2FyjLkI
2KrbtuEDK0bBwtRCqkGnoedmwkNmKi3KA8+DHx21PcDuBEspqx4LRoyimhbusGs9sxx/rAf1N9kC
CGm2wsvh7lK8EBFpDz/oMV9INl/8YBmHdK8nM9tfNp6d+9dcPfvx5TKWKGYKvLaciaPZF1LM0FzR
ZSOJfIJeK2P6fQ+Zr9uJTpuUwmmcZA/yZZNn03qozaa70sN0OafvWQNZXTPSfg7THpoN4MajYu/D
fpXCyyQbEEINLVWyvAqZUO/xRB49/5/Nnjkl4xFprPZc/slGsEJRFnsN1DoyqzlrZc5tehZEBSdy
q+rbt/GHVJl8mk46R2n8vf+Q9mWnKVBM5S4cAyjLHwSP4wOAtx/muyX35OjLiCRBgy83LLvEk/LQ
RnpF6AX6Q1aDoeygJXRD1sTqinTS+Dz7FtGBsve/KBKyvfyd9RMcaYGgjXoy8e5JqU728iCH9Mdg
51Nk6yzQ1bdPfa3F3ODmHmiXow41Pdsn/hof531ohIDyMzagupRMR/ahC/tjvGuP4YBr7N+E4xsK
REAmwbdQOnZo/cBoIM+Z/HhqLTsozFBwVwoSfQT5PuFlztKHQmvy1Ml5NroRr5B5xtcxzkrtDbQv
VUoLJNKj6GdRd3S676EaGJh2CRgLJudi0CUYip90BHlgOLouD9PSprL7oaq+0pFPDq4QgBgJWoYb
r8BCni/3mlRb3essrD5t2DP40nBdbJdvflfQR2RR6Byw5FdieMgvEaErxd8jsgZu9TfNVMt5J3qp
HXLS9sLyELL7BIwyZdM3opIYxVjjGugs2e5gnMq/qu4wUMADBIXpbfnWQTI6aJfswlD7urVVae/F
24hvGlw7WVPIx8ge69goqq+BOYgp80+9csZfF+bvsyXNMzxBYoOkA781J5dRkwNFb7MTW53KeCv3
IvD/lb6QF2fUKtdhah6IeqNbeCuPXidzneFq/V26O9tZ26f6tJnNtiid/K5r/BkaQ1JO3WjBzhD/
RzwzSzw4SEeKHPQqw8XX1tU6rzay7VUvVou/EXNnbe3tnvp4bWbwNoC+QoilB3XMnGbyYqcojK+Y
Joczag7nP0JOxLyOX6pFSOLzN2NJKxN/pHYbo0cEI0w61azdM7OatxaK7RhQvdOng7zF/Lv/tWAw
FuzL8t6bTSsSEuwWICreUdvIIfILI7/7p7DtapJH3uBr0ysZNgvPJUcFWZdxZxnk88d6MIl8MCwp
RlWbZ6npDWIC9TfFmJQ3ZTEivf0A5Ve1Pb/Tk6+T/Z7084+jzjJOPO6409tqbzusSkdFwXy9Gj3v
aKQMA5QXmw7UvEy2j6hNre1POoSy3LmzeuEz7FhHSc8KX35BjMwvy85rUf+Oa+JrpyEYr8PdAHRx
+8yC9NKccE/ptYMjHs7ncdcMgQOLEuMuMYqHeVX/UAu+WSIBIJE+Bk6SVFIdsbeRNCZKINCVSZh+
SW3OIbHh98i7ekeZdYjEEim5+xqwoT5LKSZQXGRbF+E+XemdLoPpkKENilgdn5P5B5y3nXqHBE3W
BFpDqUrfKfKsuZuP73ekoEerfPdE/nybTEWIALV3JmT2BqEIgPXRt1niwPhnPE2SUxgQua2WmUfs
+q1p10INPuyDnrgWP/6IPPa0sssobg7XWZVoDT7yayBv+K7aEIykAOrdvd3OEDoGXafLkW/poN3S
H3qSc7JFIwFiXxzlUJoMPGEs5Ktw1iChYNWzmmoReIp2Rx/AL7wFT8vW0Tp+6LLtdFxJM1JSjfIO
PwTegeFiNdZaRag6sbh7UlF01YLYYXGM328+nOYfJhyE0FLI0Etas7c0KaqaaDeMslUxJjuJMDO8
mPJK0Hh+mZcbsa8hSWPV9uhSn8ynzu11n+FGBfvYqWqZ0h77dIvRlKsjUMk3zpyslmKMhC98h6WF
uafaPSto3xZPuR+EN3i1vMoksjYAwszg8cgRYDuMLPgMORw/t/7+pLC0lc2R5boxcluNQA0Fncy7
X4Rruc1eCKkuiLYnneIMgzEBlBiNccpT6kP73weSoJdjwAiSXPwR3MTeiwhz7fIy3OnEbdKZLhai
V9bWAmrK8QlGlmCkcv7jVbWs+WNOWpZso3+SqwZCMeJDZ4/1QnOqB87PcblOjFZ7nKIHmxD9HH3C
NkHRwZMMJ4V/cQoYZpMkLEeuI6F1cfx7Q9VZA94ucaAQMfYn6mur+mUyk1O6QVRmdIjoaG5ZueD5
MhGKz3KhQfPY3kV58zXK5OjKVrdeqZOQTBXKwCL7EWQNrzz1QTOioaKYgjFfUlM0Dpe26t/Vjfdq
9y5V/Ivv70yknMgplY1o+weLW2LlkNjZRB5NZ+QWwWwZ3/5i0I3hXePisdzyfixDjsquehl8GvE1
MC9E0mxqnncPQlPTiTxB2ieXOim2ZgmVZK5OeYNt1/4lqMZ/KcEjFafY2IaDrOXdboMVMA36KPZ8
KhRRhewZn0lS9PGjRFGXsBlmEv632utRXo7qj8xs1oCQ/626itDK+lOPVoMUZTO0wB5JaFZQreg/
QbFQI6c4h4dtuzu2/tFJr5a902bV+jpQXatbvKzt0z2r/6j+LQkgScg3+09bhGS8omJbYfovrt2s
PYlMHlliA77EzIFweYB0qes01gsjKJVtNeeNIQOgC4Vrli/EzqGJ+AJIvYmAL0X2GYqP9ySAi5+q
iE8rIDVUw3aNrSVPNfyZD84z4tEuiPkuYgCw3l/DSR6E6ZTpThDVyw8j/osdHYNijf3p9//IGlVz
oNwXpFCwVQdO0Sj8LA/GJHIGrvLE2VxedOUY0E5M57500RSRWWqt1GBeeeGTZ9UI2+2yj+sZVfoC
5LIR/gG0/INTfqfrzHxQ4IoaeThyw9wnaANKVta5qVpKXK5lqs0AGu8IfV+bkltxE9+sOl4zrqGT
R6akZkrZY5q3ikk1qGkSZtQAcxYT5+4nqh0WyXFG82l2Rac0Gd8+sR38LaV0pMixR2O34VEB6rPk
4Uv/NJTDvRde3shV4fG5fD7ZsaWj/vYG53g9MnmwY5UIZbCgZoOnZSOqsm1bc5CwhRlRahDw98dn
zlQD7k5KXT+yLiOw2DOF4/RFmWoybp9b93/O5jnzzJgylBKn6kt+pkBemL7f2lOqqq0eXV4xXWWM
nJvdHGEuYcHfLajgLihlHMcPalatYlyGqr4AMvskViOnbf67sYAdp2XQD47ESe9YXYjK/qdq4zXn
JoaXhhqgyhBtAIDqsg7vqzGC3SvBJuz/m9uFEVp61zIi9iXiaozr56XS2dAc6saAsFSeMFjO4ED9
jIuYwm+tbRGy+rr0j/JUzyijOpsmhtG30CI1199k7A93BCGcLpt074Od5cA8slQGaGniQBHLfKt3
jsxb1VfAGi5MfBPR7Ecgh49+SMlFmPuYEsegJ+lYqK3e7KGcMQPcoCBvJfviHpI/Vli5YXpSKeJ7
JwgJ1vyAqJDzQBE3PN5V5bhRJBVWqxbJaCN1IprLBbt2yD92wI/1aI0Hm9YlMgwk7sTAp3odVcEL
vt19xncn8fClqkx8Mm8SLI43qLb9h6vaG/zsZffR5vRk6/vDzghdqjxQSOtXadqaNlx+pD0T6QmW
YSeUeM5u5SkuLMD1a7wUNyrzk+UQ3nQhS/paROA+8GdpbhnDieQjh4hNpMh8HV7I6lcvL7c6hjqa
GPKzqtqrDrio1Y7yhVFg8jQXSIInG1LDFblIhf9qhTO5FEBB3ZKRKovWgz6LbVM2MQcAWrP1rA+l
DA4HYVRlADmig/RTBbZdwQ/t62Lmahv29Tge1lFBg6DP7ifl9SISxnzdXfWOI7AhyVqz0+uDQVKZ
SnjPvRggI4Yrm4vsyemf0EQMaoEcmuKjG3LnV48xMmwrmCCCAqfwBDjxe407EauF5d0rwDIqHlRG
bXkTaIqdnzhhyjzdF5Km4aUR2fsrJDlToi2xQvfClegl3+TLrhUFfegqkNQFQgfplJVL45Yxa8UR
LGrXk0A6CXtY5sDWpGqpY2Pdo5xDDF+gCMXUdMZQWcOsjZQzAxbA1M9M1IxITL7unZu+QAXz9ved
QBdetPDAbxnj1Q+r99VRIrgbCFoYzu/ti30Sjz4RUFZJqRfK4yF40cOD8aOb8cSU1IS5s8eNq8x3
nJSkXJtvBwod8Cmel37VoYvW4lOrhiqJHhVBqwn1pRkViY3EUgojdVEQzOvQODkoE1tS/jGS0GEi
3kgYfltMcoOmoiXsZtLwx5Gqk+GeaR1mzg/sh9Qed7eFL6Ty5Ibc+drAJoTpMnDo3Gp82T34agFG
Xbii++qseoGCFl44ZfeOSCcmVpBA6z93DfLGd73xQkovsJH/BKlnOfTqESGZxlyAvEKAf0jItZZZ
3QjzDaA943Xb9gur4Syo6lMVav+H5Z8sTL+57SPtJR3tbm4v7UGCQVYfDDdnyipb8d5RIzd1fbdQ
3QhPbavZKVM9y6egQnU6RO2d3YU1aln9HKlsAD42Qpb/0qHzLeVte9dyhgc6QGyX24GD+YuJZdPQ
5Va9BBYf6HhbEEqnIhK7WdKtQ0Z6vEkWHIH2JNI2E8y8GDLlJlKMOIkx1xvSXoT2XnrZi728yyCt
JqiYrA3SfGXPMx9Qz2XiIjLR0g5BWNH5IW3Flh2NTpT9vcOekX3pc35TkvKvRag9XbTwQ33mb/XI
W2szNnuxXMAANZeCTQne7sFq6mWH5vblBMAsaG+QkR4JQblVAtEx2mY+EN7p0nFopHwD66fCTTZ0
0VzOEti+Fj/6oLACdFvTF72csaj3FummrWCvhobKFclJanJCEZ7vrKqyO12h8rss4wrVQy+JWwul
sJ0/KY6PrYrMS8EBJaOR9bshLAWnYu+1rTI2UCbK9YSNo1fWI9B54kPK2FAiub3FiUhMP/f23xbg
ZMAy/EaqbotVxjwRGUAVXNU3dHsvMdNF6LF4KO85n/YZ21EVblvc4oVcvUJ1IFeeL5niVrf14YMu
fDyMx7oWbHyEh6bSPOHD1KXXqn0DftQNnz/5qkOpNdqtl39MwRYamaV2buVG+CU5ef/5992ZsnOF
co5XBGviReRP3nJZWOJfyxjLb9Wl5ua3pX1lhHEtqL5PIgJbNUjxIjPoQaDUNdUAWs0Yr1KyaQ0W
ixUT1uFZeiwwPWCmmrqEMHeTIygZN0JkxEIUglJgwibKnQRF3r2AEaecK313PiZu+0Aogy/IOaHj
XB0aeITDozzUT6ScLqVw8yyxE6cTUShCWAdcLQrUXlqTImtrMm9HbokPFuBUq9008KYoxJNU5FUR
NtKlNzihWKszraSFScGSu3iYr7h2ycW9VQblPvVkLw88bk3Js2eMEeOa2a4AFpr9+shIlp8kFdfY
YojHbPsKD/tq0R2gVC5jKVRs/CFeV/USNCORa/GJ1zi/llm4KyEVbGXGmiPw4uplel2z1fnMZLK2
q+5v2ztjApk/GaENvwphJnUkFlnVDD4x4RyiVO7upyN+bTjWKxiDTYlZbW/yDgwY/1X/NcxjsEP8
oJqf7wOyZxkjQpezdXAG3ebObC9VBG5XbjfBUgszKJQ/gff3Me6oFPgBaO7f25lxNKpBCxgDZmyE
Ry0Zxa2lDaDVSY/BCNqgdf7l78K73wve0+OA46h3tKSbuQbH8DM7JaDDymTWqRNAxNH500thxnKB
jRu76+wDzbp9s2BKGZCNbClGQx9zSMQe83lzDTaggxG7NjNlGKHfN4IHYGMY0cw8N8v36/n/Hqvw
MvwoJP7xTDQ+dbtlteB5kHxJcSLYoObaxMrEbvb+TtYEaF1cjdUXB/DgVRsLBAwpcbOTwQCu1yYF
gp0s26i+5ajW3qQh8PdTZ2BUj/e8qcQmzZp/IDGOR3TgGr5f2cAXAnFiNnxYy0QiLNdcb1tyCj+/
0lSuXJvy8Ck3Z1MGzF7ADO7DzwbophggW7diY/rFBz3Qvgp4SjQ0CGO6Jeplx9xBCsgye8WHtSpz
/G/VZieeyq1v+U7ZuAa/fQqjU8jYsnzGQgtgFDqM8elWJnkoRGwCanI4U8h+JzoLgL3mhZfKAFCV
w8y7HRmXIZy4dTSzyVZ6GBw6RQvtiLhEGjOOkLczj4rIWVjIp9BpzvwvMz8gIiULZBq1bm4IPD3v
2AzYB1SoEj4/ySgkI4Tde7grEXuEwL590ABZQeYJas8tOchQ2z/AcVXC70qPMWlz0uucYZutfGVi
5dCa90ebRLdw1N+DnvenOymTVAigt7EnHa9Wrc4A2UXC2DjZoupXhyqFUAhI+FsdbMubbRmL9vKl
fAH/+YXWCB0Q4cJ4IuMK10+c1VWmtQJRUBEtvq/KSr0mbKAxUeb5/MtKZS/QOVsfiNjGl2PIljT6
hJT7vpcQJsCNXewcJYK7rM3KNpJLEjOSLIHzEa+JYch49hU6m9hMeSg5oeXD6j2bBO5m9dZtpBzm
hG9mIDmmI0c323/hcj0FLQtG9iiHN/EY9pW5xqGuzyCf4h2df9Nlp9yybafeHKllmP+v1HSEbTC1
0mNEnL2Gl7xHGSDo+0u0cenOIbj0dXXbX9KkyRl2DcXImtYRLHef/kTz4jhubEKxSED+7j/X5HaV
PNIgIp80KaSRJJ4rL4vjuXZq+3MYtNLH4+LQ3maYzFNPMGISTiyljNjSh9jb45E1nO9o3azh509B
cTA7bLltM2YgrmjMlHlFii3GeYu0immO4VC3oga6Nrqephuua1wLKu51ruv7P25EaSfVqXUV3HHA
aLKgFjRb9BfcKkIOlyBrKfdSJPL+CdeL/X2/6Vgmf79715J4Glnf0NRK6af0YQKorLlzpaRGRcjg
J7jeKtlGuMYuwKablK2LbDw0cOOgKI1JOGQ9g85kEu1CYohC2C+bzhwM3SWS2ReHeBS6MBnFRjIg
PGLu7Hg6oh5ZAR8QO3mpfY4yr3uvihMBWcXp3G6UQO5zE6BQfFOeQd6fdohe6+23qB7ALD5YOLo1
W0GuPELFQSRrOgFSEjBG4ep6ItrXhklmHQ8PjNJDXBBitJGnop89JWawFSBrikJ60c6JgalsWE9I
27DiqWm01EKLliOs90m0oOdhFxEzT5vtXxNGOG0yoyLk/2tidvyxJo1jjPnPmWz7Iw5WDV9tM0r8
27cmsc787y9QhgFCqMbxU8uwfVDoSLEHyVBRr/C8X+Z5xa0WsVZlP9l+M2PfuqPYNSPkOWXuWuVf
pPay6lyNf1rVSrX7f8kMSHSX1DrZgX+da+NueV5kSHBzHbBPoz1DZnxYcxbUWYlb5X8PDrn5WC9G
+paGa5hmp117r0GpEnvwaSTnw2zutfXoim3uys7vIfhjJXBosGSL80oEcAI50kBOqCSl/0By18R5
S0P2uasM6UbqP8cOBEUfLpdO+8ZKvwO/nOMuPoR66/hLx9MK8ZdF4LiEznLGSEHpne8I8nZuldhD
UwZgM0hHhVJ5BMKDWJpx9pdti1o/PQ0myVLbpYbahVqkZ0NHKJeg1HxbJw4DC6vxt/5fx7hsn4n9
uMtXGbknuQ32yRKLpNTZJLqRAwDxp5BJTr4fEL7uaca17JYMKaWOwHed/+vc80iQnk8/STfo+GCf
Ij3Bxj1Z0qf9gJSeLINWrAb2pvB9WsyIrsbCqLmetTM90KFzYJtmdg0IMdKtYvjc0m3vEYwLAaJM
YDnR4zV4xq+fkjeJ4rYFfI8FiBDSrCqy47J2VQmBUlzSBUibcdgRk/69mAeeKYZM6e2pUscnSeLt
HK+ELKq+oou3/rOw9t/0Zj2h9mXKWpBLyFo29e5fPTrdgvS1P+hSetOnEEeqOf+2uiAkje4Nzcfy
TRT5yiNOfy8HQplm+BPVGuVW71KWcrOr1TgI0489U98k5KOdpy+D11ne4vwntTy9K18b3zrwN5S5
8P71tdKPdImhsmYk4M81/lQtYIHYXV1PUoQ/eNv24PphE9wIxVr1lGwurDa7y7FzKVoe29/0qWL7
o+A6bPZcJ0ViTGUqt7lA4fG/cI+5nfgkFg1kkTPqbfVHnWh1qfBY7ETzZnxreQpeiGZU/7B8IW3+
PSIer+lXoc/HN8d9jz51uDlBOReucgaG6aNF+JX0yZuqC9AaiguDjkfhbxZyi/unqaHvXIq9u/7N
dCLAqu9KLtz/D8zh+1ueMTc+4aXEJOFJPVc+8qUHD84twj+GnTfwNuVm9gH2Ug89RD2EpqPAUWOM
6BAK0QXPYyN0yB3l2kVBa4rHeewx+tcfLmmU4gNiKc+Qz5cjiPzWIApv9heTU8ErEV0Ew2fyVoLY
0IrMh0rqe6T5kg1+jUNe61vL8gwae+CZLbq54n3cXSA9g347YtVXfD7hsN4dKkzqlQGg0LdSBuSE
w5eoEGbKIyktSkoK1Tz88Al5OntGuA11apnQvKgNrnxPVZhFWJ9FjOrcWdntESdww681C+D6iJB3
49VEcee5kdPNjhnP5Y4i23Ng1YaBXUE1z3cbtBY2fnUr+LsO/gwvoAhlMhNkiVa2Vo8drwlA3anD
QcAWy5Gp9qKqnVLzWmtLiHCkmJHPxsK7g0p6P2DZl37KlHAfSue7oSJ3VUvJH//hCWxfBRRQK34K
VhFpByNDbEoqP8FsQ90Y04yneu9JEMEZiWrY/bcwrn6nLWqAR+ERWxjJB7R/PDGW69JzpCNQemPb
sx5Booq2+eyOi5QA6NWASCjUd1hxlfHwfiAJlvFpeWrALIuvygA2MVPEHcfREq709cOBPuCUk1jO
wclqp66k6JA0Cg9omVo7E4pG4JD20RNL0PolRAksp1U1Xrs5DZqmmFW002Fp/m8t5k3KmTu4UiEE
WW3Uejn3PJKG/njv9lG2RdNAH0Q6e1y45M4r9EGE4YZVDMZGwanbpbJQ8aCKKWIPzhherNENln5c
w1VP0qujfO9RUijeeONEEHLhFUPT/G3VWNYiRer5nyMezIb/BVODycZtNcENXoP8GKWbv0qN2Ryn
lzGRyKzV12vyKwjV6Z6G3IKh6Qg50nhVH04u2fujQTaxqvfiY/gB2PyXg7BjLEgtUNqFbzXmJ+2I
9BMzsJ0smdvstBWUKs7YrTWzALMOQlLMinW8wmuFe1nFIjWDyB2wPa1TggH+OZzV9KRQm99628Y/
nTXQy344o4jOCB1c/uulVfLLBmU2qZFSEK+oSW59AywiFBDMqSh4q6UjDDCuzY6OMyhIl0O5LpgK
Gu0cfc9inHBf85zWqm2J1dHC+KQBF/ZBEEGXrK4mt2MFU0cuE7J6AxQE7ZiDweVlBruu0o2aSi13
N6m8M7V+jlOd+KNuVaEka2u2F9yT23n/TtXAac0bBJE8TPnXL/kgS6FITHSjxzpJT1hZAJL0ePgk
DCTPzTUbh+zbwGD/xvCHArrrlFfW5jrOWmPhNrReRTYJKV+ra1F2casLsxkKvUubVyIKzHAnJsT0
GHpfpR8Czc3lruiL220ihzu5OzI8TFflJEgagPCJR1BswyYL6J5e4BWm9ReVltfXlvy3ZDIqoepP
90+n+fTLlqOqHx/Q0P53owoTgKS0esEJPO9nPjCrGkAu9rtb0S9s15I4eprAhEEVoQaFJWLu5gFu
0qYlIleyfuZwtBlRoPfe6OGNN21cq4CMoqj48fS8IshYkrEgAPFsZw2QhJ9JUHhWhglvOpBl4SR/
b6BOGzRRQSTgN6+1sokR8hMVsxfbAv9EPB3aoqfUS0il426THve43QG9wYQLz/Ao/5YT0QqLKWnb
oG8a1mMUDBslfcVPTtgNnBP2YlZ9qCT1XcVZ6qi/TmgQwoj15X4R1UfhrknQYdrA2W8dW1CCPvig
bhYg7CGUHFM0Pv91waEFgdiql74h7hBB7lDvpVQ5n0X0HmxhzgnvHGsWV5Ds1ECIn8zIzXAB2lB6
8rnMOoe7iigCyY3dYbrpZenl+5gI2vN5DGgqFmUMElMvsGvho7C9JYlfmgHZO/2PTwW+MErGE/xi
EfAfIRHS0s8R3nJcR5MKsMnnpQKelSnJfCdTMLwI0jV566xj3DWUxC4TqFja/0KOHFek6MJ4pnUZ
hvRrfSRUY0nQFMbOR8hNDuqsCTRFI2dZS0xme014OxCydly/uqtlrb7AZxn9Kr5kEess0TtYGZme
dLtkhy+7PEXosAuTnBAsMAkgS6+VsZy9RqNfaLBAO2zm6Hmy98ca5lio4SP649bp3WikP31ZxdvV
fXe7Ow+/rOcRU9qjDvhCsycf189hd9KRlMokVclg6pj8LHvSBK6SIN2te7tm20uc6aTxDzrWsDJ5
Ev9WSRpQn0AitiujhdyIfwACZ/CsBe4iDNXLgTqMdtF4rzr1LyPfgFr34xWEuly0bG9z3UURdfkw
DTHCuhSwHF1pTa3whTPUgaxzCeU707xGxLY65QSbZTNxJMyoJ7KJJDFiL0GV2tvbgP8UYIy4BMi/
yLGLRTuRkluTz080MLvS6h+7j3SqsIktLhJpICLLOAiCrgS5EPB715S18NqasvvBsymCrLaczd4O
cz2OMtQmq0nlpnqJAYd72EaU3Xm7sxkjWKbRf+gnyB2yBESLnCMsLkJJ3pLSKyDD18PO+/i13RGk
XWe5p4WYa5cq3L53khcuPGzhQn709ESg+yN4l43wg0yl+wXLcR2yY/FeZdOXz5xaIHZDrAEkyity
Fw2S+sdYr1rR9rfg4rHX8SHm1pQYxb887TY55j9y6mSgUItimQ7ibs4/E67WwZgV2196YJ274qJ7
MiX8MKb4JWHdjstdyfHYijzsqIBE/IGWsWkSayWDWe3l7BjjP49A46p2+9vi+B4ImXDWIZ1kbDiu
4UayLpCalaqeTCg7r8SPmNddTH4HnWd+9sHRl9ykGLYTXUQSMvkq41FbF5bEx3KqIL2JE+Btrtee
QJ5vlVAbkTRPnNO6dR2SKr52jMFnfW8uKGtt7VFhcUyONbCrYi7V7zMlBoAodymOsvSzu208CJL/
49MsevAuqL53DKYN9sHOfO4ZvBMwSf9pC2ZOxFiL8EhMTS0nUj2gV0WkJHDSznlcP7GhDdgIkKsn
weEZbf1oIrZC8K+2EjE6bHzQWdySbRWcAWBGvZOl+g0T5fsymo5gFm1lkvUIw5ZINFLlGy/lVWN5
+pla1jB/4SYnk4c48Tcd8e35HVYMiNhdvDxCUeOQkR2UAxnSDnYd8iiDso+ITWqam5ViV2E8bHu7
FyZjrNCAjdCnReKWAghnqNMQRb7/impG4yU45zwbh4hvaqNMqLxtYcMn1oaiZPv6Ih+58pntUS/z
QLEN5C020KdpkSTsh4vM8dPkEO1zxUZM1QNCkkRmLY6LfnTq86JMXfHBrVDjKc0UOogPnTTVL2Z0
w+01znCcxZGsc9ZQ2QPVDVStKTb1zXbslTH165MT2Twf4d6v8QbIG4jADH4Fyeh+po3BBlWJc5ow
NSPq2kahWKAOAtzuPyChKYyGTCgk66qnTXtaYNadeVTwufNCPQr84F35nz6rcQZu7tSMV4cW8fQY
o85YYpHdNXEBWBeD1HcV/sopiEytKY8eXzTYiiaE140MkA49boBu9fwFldbxXLwahSgbrWiO6rUA
gWp18hQ/SzZJLbMLk6uqDJd8LLAIYwAwz2t76P9x4pJR6OZf1WVkEAMx8P4JPGk55mvjxOfIxmLG
KW0UBelMG2R9zOkWZLRrysZAMwOufqXZm/0QbosKbiGaW4pDCpXy0WGp7YDYkjvYDf1+/C1goFzG
tHKOBjZcppG1Q4gzXlyc13y4gIqOrasrdZCeprxNTFCuWf6HeYxuLyazwEqanpVPPYmAtzMLaGlo
mNtszr3DST+qp86uW2d71k2FbO6vsq5oSZJMWsGEb9OFFWQWwcmxyR3yWcOWuoKhCh7yOPA3YByy
5sWwS+ZK++GS+MKjQ9o9j8vrD3PNJbHPjgAq8rugN1WSNVWMypEIFthHwA/eKMR/kpAMusHxxT4s
sbmWacdQs4kvDasQz/PEwnRwHfiDECchKtIyVP2vOXuUS5YqS89ins6x4JySYnNyOXIzuopU68wh
zgsgopgLf/nwl3lhjj3YB+QFodGI0r9gGZdFHTfINwUcUqJizsfefZ+ct+LIm0cLtn7qHrB9jHsI
Igokq/GG24t1tCLIlYXxitfAWehXMYhG3bYKHOx06mT/L5JQqLtMpVo2D1xWU5FTf+gv7YfOTf6z
GQO6ERSzhtiL7ewX3KE0ETydzc3O/mnvCJy/kzfLq2u23RyUXppC/KhfMjBL9JU11j6JtxIrIWWo
LPMnJkjqwbqHoVImQuzVbLYdhaCkNtn2AtK8UoDeMvAguw/sR9afWJbTziFTF7f3yQoOEEsUQIOP
v+qzsq98gK7uXjgT1/3FGd8gppToeLBCuUHPbzgXo9YQPy2bfxEZW2E9SksaEcyZefHOydoUfZ7e
BOTWPfFuVWCBZN3XFebc7ISZ98HTjrv5B4r44IcRlvW5PJV493xheK6WPdBgo8ju1KVCyBPMZwx3
MMToYt9d4WMTe/bEWoYeHvJnVCVGKpkMC5txIHaubZk1FJaKwSZADQ9XkC17EuQ+jYc86XWUStv7
1XXM054Y1pL3+cXzlkFAgNhAgmoXRQ6tW27D+m72wi2HZYP/wuWYFkxv3l2adgCu+8R57JAhoBFY
DyMEi63pJfbXujaz0iSFeJCds9VicBaNm/DWqaW/k9NLa5uqIsXPhQxCi4M2++h9Xs4bN4R1avU9
vOhyj/vOUvD7gWmPMl33rPuqSSYqlGezjw+i2ULAgp6RmiEiZsRQMWKEvkdYY/tScyNwGknYmdRp
OUT5+uYbFv4nxHIbnJI12xamJeLlxabuRvbQrsaN2opro3Ud8Ya82zJpSgAAosfqY9oRT+Yx4Ql/
nwWHPq919OznoAWn7c3oFe8SGWMgAiFqQ0aOLMXR54Jy1hVPJhHy1iJND4QEwoTyGHeMvzHaEcMZ
FmYuRKwE2zW5WJzfgAgFBmx98Kzz8DYgTg/rL/7VuSqSDqNGsOcIZ5BHSvsf2FbQASX7pC/L+b3R
51LwymES6Yn+UM2NUQKJ94Uk134CpDYgkf8LsZejdTlz6Du0KzHZZGa6TmJPYmvSWuUmetB4vgMi
5133LON86qliFo9pisYB3IakvXe6mJpXd7lmrB35SoPgE5dd1j/H9eQmPmRySgdxH65EXZ8PYEh/
o/JpgqNFzxeJtrkM+ZG3IU2HNMXJM8282LrJRwZtZi9OkjfmrnqLoWVoSaGTWJHJ9acP+ZDBAANs
v8Xi9rGqTpHr6kqmorDyG9hVHcpE8vmtSPir9zJf07xiiNcw6Ui2NfCoeeADejWi+NjRWVKHtx3L
HvACUJnRMh3aINAIprcNKggIfVui4aVl5OLk6eCdTOzKgLzjpk/oxBlz9nhGG1LMzczUgBxeMVnT
1wVd9gumcEjOLpUN6Mjg45U82+cjEeea88PSRiFboZ7nlOzpheMvfVBY4c8TlVAj92xpQHI1J9ql
X/fA7NSmFUF/6yJpELHCGIGbaintJd60s0WkvqRZ7LoSWKf3vbclcAkKUbxWkQIS/gPGlrCzuZyh
eDoCLGR2f5Ki0lysXxUBO46/diIvqUI6MfebO2igBm2MRs66ZIr+rjCelmL87E6HT8Qxmkg9LPRK
vVyCtZ91WTDTkZyuYU+bGC1NP8/0NvTGyIr8VZGn/mdUX3Pq9YA35DHmK/riFC2BvZwBpIgGt072
DEqAh/WNopyM6XYYeeAnRQmdvcLgsKN2dbGDdrLkzyGknogj3z3/004kJACCdyAw/q7FyXNHY9RR
940e8K2LrqeJn8n/Yupev1eEWhWjGZ8cBH0k+7RViYnCPQKPtL2y6xoRpm2HCtZi+frQ5PHLMN8c
YqQvBRmhRvFN0CS4eQRpaCfRm5oqBg6d/N6j83SkmrA25cL35YuenTor6e8BNd5q/2vxgHP4/ZzQ
c4B/j/HkChHK7T80ysn3EraZUg1Aq7OVf3AOrWUBjnGieK1AckyfwvzRqZ1+KEfq5LWd366xG4GR
J+FZX3Z9BG14vP5Iw08HKq1zYCshosjhUZ7oLckPferYzfCUWCpZOaBxg/dt0/GloGvTVcYQYLlZ
+E1vTEfy8VgZzC8RiqSB4gKv6Y4DzxGtAxrk6BEeoW7emewZDpukjuy0fun1n7xr5WH8Enrbu0rR
ESYqn2XpR0YoB8rcCyasfEQFu/L4Lnf+Yic9KPQ+rg7uyu9LThsIYBs5J4DcrobARctR5gNWwAIb
MKrCK6Gru/eFgIKWRljJQhwiDWO1X96R71OyXlxUqf29WVNJVkSoiNiMbHLBuRB/Rv9EuE7Xt5Mj
BvqQC95MICWJHFul3e836c2zIU7nTYu4JIVy6NF4rm3/Rp4bwrF5uD1YwdUR5wjufQ+q05m8XSGH
FoRr4gNzlsPVxELaTEnS0PiII0UPsbZVlbHG/TU9EfElImfIr7TbE3Wjcf80XKsTEGsoY5048AE7
rXCfRVU9Of1xuutKbJxAaYiE7jswCRYQ/+17ktQYVmaeGIZy55mG6HUbBynqmI0BwdwAqw6Ht5jq
8CpeNApIqAruo3MxAjsoOmXgIBepmcl4ye1SJvKkCaetbo9Pbs5w1Dda3ZO9grySQFIVyat84ihy
X1uppzEvlnb21rBS8fRG3LZc5dg0kvkOYMypHpgaPcxEaIKMXx7Ohg0mjGcBNp2Wpicu+TOCzjh+
KwdTmFB95L26u2eHVwABaiibjdPVo2XUQkB2xw8h/sbpild/B0gGphjiyFUvS3yzEsjusJ8ZiwPT
Sb01kzRTTem/549rtR8wKNT4O7dkQy4DMAIJ0BzJqlxceRoezCmfm4EdrIu8mzRg72JJJcrHx3GH
NN52Ic5R8Da4o2wK4p/Mk9V0RL+hw0tFpioSFI5ae6GnTfID44KiipQ/Kvtlamv62lkyqtZ3jWZO
xKQM7eB5ppiZ4uLhuAA9ZCKKqK/lUfR/S0znPCyS+jz2zz3TffP1S8V8Pars/pqjLDLJiN3lbm9Z
SgrWJwi+gu7DoZ/Pv28UgsCwh8eZS5GKMc7pJa/KXCIsinwMYkrsE3VdLJ3r6YqDCoaNuAAHs2/G
y/Kw6F+K+Tcnl3HlCwCdH/aDySG40dVcOG4rnYXG39w4uOzilzHNS5O43HFCI/fo5P9IvXdcLzBt
ttgBGMXfl8njiF8UmVz4HGh4SybmLQpsAm6TAe3srw3sYxVhOnalSNAbaFMCgKKBnhBJ03RXtVbi
bUizz9p1cOTRu9XxDlfLAyv6tgO09LMCg2TVjkvyejJnRm2wFUGlfIOEPqVekpw8ZMz8KxeaxIQT
YLn51WkYEGIqYLbGOqHmA8I5l5XWjnNH3pYWoWj+RFqLrKubbxsSwkjcDQ8bPip1xzyb8j/r0qn4
h2zLG0l1PZ3n2fRJ/0qXRf/CYrqLcZddIX4EBjFI+Ti35w3sSZta6bBt7YEIrgTQUda0G8Ls/LBN
MmitFIHt03HS4mRno6J7tVQTCaaojPH69uh2hwW2W+sua+HAh0O07ZKjEmnPLgJ3D//Ki8E+82bG
8vwUJWhKwQ422B6yWF65TReJDGch79fp0QqbfiON+tvGZ9ZJfVmN9u2l+rEvX/Awt5U4xd2rxTpv
NWqMTKJeXN17Nt4pWpZuAi+6Wtb743iUi4SxMqqnpq+5Sxaye7D63h3QKt0v0GbsDpXM0K0eXzJq
vfz/LA14VdYd7gqPo1PPudu6Eo0awyXBXktEYO+TySONvQ7vL2KGngIXs0wqzrSqeLDSMHslP1RT
K/bU60N+ypt7gu1ASOBCeKxHXAKBzyeLVTnWNJKim3zcijeIl/Dj2rCLEdRlBzt9H3HIghIilPLv
eUEawuCQ9IIgjX10a9o8g8NwddzZCVc8aPXnjkxdjfYmplX3l8s+AR4Mkzk88ScMTG/J16DXZx3B
Nf1b4MLVU0aEbIAU6ZStxwI+9ka4A7d0avMsREYlKUIo4gJe4jJ4Fz/URGCeizCA2TrutO124aef
9hkroYvBw0MTga/mv2AxB+sT6GHduPM6DTzfDm/9/Rg6cYjs1p4ubFIYSIHfkwqbESQVeV/cR6xl
v8qw8YqMrd6bpp5/7/bNSvRWWx2UgBimVsHcEnPc7KSW6HX1fsnUgYzIXzQITCZP9BxsciY5eKaz
oIEPQgKk4T/1Q87NH2jgURrmWFxrpRMJuKpoMS8PkBqaGHcYW2T1fDmXkvAXIslZCsBz2ktfLaYF
7oubkoXinrzsLA2QVgWSuMu9UktDDF3QlLX5+ZP7p+FxvOSBFsY7YSKvgFawBLtofE1vamqesnyz
h6vs/2qd3B5POnW4qc34ON6Z7cwFKXzmH1EBWCrj5FHQPAEyKyras4i5ngQ+NxJ+6MrQUnY2K1/Y
gFnC4OKPwqui6fpuO9ZiiI6BkeyW4XlPqrvI38N54w3xT38dEJoIWRNKc1OvccGd8OfQWj+fZbjj
PNtYugbOY+rJzI2/9MdICvSpWTbg0/9fAAa1GxZgxtlW6x8z3chQPcxVuI2KInD8XBgGgQSJWASx
u/nM3CeL3JqlSVo0RMhsZYOVsCVLS3Ckv/ii3/p2kBxfBrHq6LfaBk1rp//Zk8GOosdIjqgm1env
5iMf+/AqCpnqoP4pFaux6TmbR7ZbR6yIzjzTVEN1iB+BRURUs4RbSvvcIXHcjxwnDml7hkgEAtCt
t9xaCCTRg6ypK1S768r18i//p+uvdPAzYIu26cEumMPeBPNd7q+DCjVnIUS9ZIDf9xWEwhUW9Pa6
NTXBiF0hHM/EqHhDPPVW5ySPV2MkiAChjAVbNfe48HLjOTC65cNkly8z/4Im7akPG90gF7aEykAr
7QF4fNW6xvfGV9EBPOKwwEMC49CFeCEQKEU4WXdgl3bVbDeO4YJRKS5ws4or6KKUWWumZE2uBCHJ
jyycm1Ef8qgLNDCUU5YynxRuDRbX9UrOHlgw4EzDWWM0hGsEf3leKtnckUSYrCuIlBY9BPWldqq+
Q60z8CBQWgvpdTwbalHpHDoByqYVMsyCXbrV6OaZdZCuB1GiAcNxfqjI8/HzmENkilxvU5R4GcN9
bmHimS8GWVJKdrcyAZSjgw+uO3e/SHAtuTLyU96DccJeR8M7ELnGKOoiIoXPTh0Pt0SS8OnQLyH7
TjcmjrIz7JN94eCOHP7fpJEcUNmU5saiWsdQWhwXBqtwJu0VllEObISW9rUWwigQvpg8cZq/jx40
ERisvrWEukGEtnsBlk6ie0bzSa10bUTA6DqgL0WRJAYFCFcdQlCGHVk8JKUQ2TunSrt+eP40DTCY
AeU0+A0tU8RURndUZeLKC/GOH8XeKByydzQo1xl+FNtrI+wkZ8P2eelLlbeVXwsQdaWl6Fa8kK0i
Ccsbk67QNf3vqWMt1VAfcZTTneLMbCmGB1zRKOos2tFcl2zI/H3lUDf0mGKQ4j2OJx0k8z+xr0rD
2Ktp8ueLcDMT0xBA85O4zn+UBP3YpWASG58orOG7Bhu54nSyw0g01KMGTK6UtZC4C9AeKeujn0IT
0XAnsM/w0jF56ZXoEn9HenFdM6XiqaGxyRmpNInMZVmtO2OldbxYwo83fzI5y8q5YuytsgBcQBEs
zlIr5SHsdCfYOqWNl5FDCJ5dCzoGIrDsHAY6dP5P+TiVWnTFWXCP+3fN6AutIErrcord02gxNPbf
BiIkqD5RM+moSrSGOQGrNb2jT2z5HFmKEX04SPaZeV+xZiDxlQgAT0ej45XrTfqpkb1eVHTKxtHT
L3pAfMoJEHwA9Mb7AyUsiC9peOEPBp/F2MSAm/9Tra2Tpm6rQmK26E5Nxoo7Apz2hE12Jw+gATBj
k+q1C0UPDVk7rQvX0Mcd7unhKbWAPoFGgRe/XPcsZqXY++R8K80vy+ynFfLhP0itPJPZc67WSK9Q
wjNoI8T2yOdNply9rD8hpBBPgQFd9hz9YR/gLPpYxff8RTOGadctjolofK9nBdCovsYuzeyknLUm
Y7l2EqiGb1z7pqxOmUCbwxD4Mf4wWOB/Co759sw07CqDEcGZ3uu4oVKsr5v4OQy4nNvPLxUEval+
uwYJU3XxAtEiwMAwZtr3C7XtYWrTFLjES8juA4IGMX1irKs9X1TuyO4ympqdp2QTIR4yD4H7t3Xf
5PCO76uSbbdRSn4eZg4kGwqFFO+ySVWhM1rBCO++UxEQdh2nDJQFDGA8Zm2KeQZjpF72wpNHEAET
BsQky1zN+lq36YRGXrrB5Z0YVI23XDK8gLHM8TZXL6E35c6JKz6TIFLlnQpfy3wO8W2Xj6QvXgk7
JP4am4QJFCSZDLIHKLPIGu9IP8nR79aPsMcl4sPX0PWSSyVA+hk5aFGU9SndrmmednzTg/RH/yQS
uUdXMUPwPAmZkQXmGcOQiXmWuZOtndVshUgtlH4+uq2pAFAqgdnLh6o3y1MM6oht9V79AInEjICM
SyzBJpXjUb/bMNksnUkJux1d6uiFWgvnj2ONY9gHIR9JddS1IoclUkkSkYNm5zL29CMzfv/5fZAH
EqnJPauCcA103lKt99je+4Cvkpn1jJxRjvAnwLSDyfRZkXiXbIvlaw/o9jyZgsdfYJAl95epMF5j
B+WaopFNp/ZBabhi8hpTaer6OPPJkKZJWZMC4l48N2vYojiXUYzUz/o/b/IedSlp8Kc4Id2W+v8u
2FAHdI7OUrjMlWaMF8Za40Bq5MFawLQulBcorqJReblb8TWtPm2dAyG0593nldQY6gy477SLzk4Y
oqcU2TeX3CfW0vPbHtyyvYJswIqioL50Vbsv9BeClUptIQZ/KDK2rLDwpV8fkivTvd/Fit93n/qG
Gk7v13PDME3ViL3AxiWKGGlbzsUaAm/2mLl6akoezOkneWglTy5tu152P3vV3cUFeFKU5JBsySKT
PVcw3Y2AJGldKMPkAJE9hLDwXzrAKvCAk0DaynQc1STfJLx+mbHUgTAjeckYaTzs683MqBGA8Hg/
sJaphnAMIUsT9MuznnKGzY/Ve8z+UEck1CVhxlWLOWSX/z2LiC5jYzuQM/TfOKwUQlvcxOBSSg9i
9Af/UZ3stheWPSoDm/foQJNEwPj68kYbfgoJDyHDbMmr3QxGKSkMcvIwShgigXi60WdWdpRq952i
ZrQP4tB0pnWb/kH7jOzLN8+HKRth5ygoECrlVF/HgxvsaMRhSP1wOVXiGr2pD4+0q/it8RUxI234
7OxLuqxXrzGOg29OXyVgQCORWdKewgJkT0G/VCnJixc7ugTbYXkE1/nvQXavM/JWle/MWkWcQk9S
Xkxquz6XVQb/oEsjyVmqL8aPAlD+x+CWBiv0OXqvXLm8IBq2zeeCp5ATC5lNRLPBUstP2wXw1uWY
YhhYRGAaTeF2PPTwmsUAgvX+FpKMyhTYM7XUcvSptjjoDWsRO4JWICaDZ074hvkJsSYZ8Rc2e4Sv
Txxi09hTS0Pw+4PE6/VwT6jWrt+cFsQcbhavVREUvmgFqlEvI0pYjleFgHM0Z+kjx1akXaY11hId
7tV9z/O79xLwEk3YGz4lLfkhi7FeArYUrird8ivz0pas49HHr79XBQsDxd4/TvWmBEL+cX5PL65D
6XKD1gQ7AzmKUdzFzgDMoPbcGo/bJTOSWW7GGyyaHYTqYZ8WZtDjpr9Rr/titKxNVJb6WXwxAA7Y
KTQVXRwDYB7PiErXDTy/8eRwDSTq+knrymKsznqIkdwr2elqW5GQYW0m2hZjoTXBT6L0TxRDgjPL
f9nX4g4nOZsuXqZ0ttem3/RkxpLf1s0RMjTZxhvOW0VFBjAV2AhgWnJZ3D9Yzt6XhOdzgCO6iVRQ
vtLty/MYpQ8f1AF/cfe936kuH7U2XvNVdakitDYWy6bq7SFxT/myAijG1sOeBsZltcgDMUGM8yl0
5qK9rybr8skQotUD7iFzUs7Jvgk/f7r3+EcKNn7fZ7JNivcjH3TdtVIwlY/iG3hlBCMZ8BKBqtNP
acdx9Kl1yKybkmFSslVVdzh+sFpcncWIvcLnaAJjBsKAYGFjeHWLjo7THKxSohKLr13UVZAXUA2U
GEzBSyyaVE10FDPIBvEY2w9sQFSG/vDLNaZBkOtwxcMBfbIh6vJ29AabQRN0a+rquA3FureSM8Sv
PxSuf+kxEPU7892xyEjjWnN2YqbbGxSx1AKC8UJtgiuxM5Lk0fe/WcJuIedbu3d+a4W2FLQQe9cC
kd+P+zfp19kUSF58xC1eLq/u5dH/n2ezJxgYVJ5SWNgOzUCfrCB7XRcj1Zo/JeO8YEn82YiRdlJR
gNbgfCPmvxnyj9wSh/wzVlXXDxq1fLcT7ANtJKqj4VXG+HlUkUECYAc80NEvKl3CAO0V5zcw7Yzz
YZuryzICp6LmpcGv+Q0TtbFXvjgi/Ml1v/glObQYxhtW/Wt0sgMQU5aKsXcsb6F40K/Hrw3X4qYR
5XJ8DA18U64mVjCVBwtwO4NFeh4otg37U++bc5gFYg4cjR/y00v7xbDhomB3JDnthUpby/8v6ETR
x7KhGCvhF/kO5lUgZoTw0JZwuGf9ZLfjmEhKOT44sA1mgUYy+p7RccumFFP0/MxPeZrPWzehVRY8
CUO3yfzP3zOy1wrtsuVxtMmDYHas1bwc+W0eQiBRZJyTlWcSJ/iWo1wkQRRA5ZHB6kT1TjUIsJUS
UnUx19s/uKoM6NS1PkkFuBBqkU4PdPSHsRYDYOyOrf9BqyWYWpoCNXpu0mUah225F8p1vYgt+rsf
82DMzLDZnDgzjEIeeo5Hl2TAOLlSzScxbQ++K01Z1kU0CXJ5TpYmf0qPF6wrI+/0T7U9ZrZjkba8
kHG8U49fC1Hl6L5Yx87Oul5Z3yYtRygafsbSg+xIQB3LpP4rnRBSlwU+Mqw7YCycg8i/orPCbsGJ
vqkQ0/aDLrjvfi+QOrrkbAIXf84T3kfwW76UiDsmrSTDdL5nIxx6Ac/4qusY9cK/Sc0Up3WJOToD
dmDzGi0zbV9IoLufESpr8hz4jzVmS1EN1noahAnyY+IVS41l5ATdODgoZ58XfDKEYZfWuBHBjKND
tnXBUPZCp1nbTPG5JlCPgcmSJ9M4U/R7dy4O/SWkuRNqwMbe348tyGN2qsJU8LLd953aH5N/h7U4
o6BcDu6lhG2wwABLCpy6iYcGQcGDHUTShfybneZ3HQuRTZd/u2IUCwybn7TnX5p2pH340ZZV1C0C
ie9nnxa9QTLVIbTR/zAySTh2z8dYwDtKFx9siXGnosOFeMShQlX8SKANx5dtBj5w3avh9Y++Oar3
shM+HCDp7/ZarzT/5CtP+XHf9ShePThSTWvxz+SKKZ/jVtzK/8c0VmfC8sv3GsgTa7U41esdcaMI
toS9IgXnKlQlJqEwDEki+A5DzvZ99Lc0QnidE59onzpGpM8n0aUALSUuODejn1O7Y+qWGJSU3aJR
ysWSNwHGCS7dd2fUbaL031XSF5HYg0Cvk9TKInriqut1kGp/4Q4+5AX0h7S1M5oVYQ9332UCdFJr
uvXS/PkvCfvtMtdGSvWamHeSycBBZ+yLYgwgPbT7tjW1gxrjgaxAv+m/CV7ViMTnyUW8vTITWaQp
+8GbkLStkuQlkhB2S+Z5GJhnwOsRtO/czP5nT4yOP8FRwsnZxgQAAqIWj7RSurFyPm8PN3upoJ5F
TTzC0YGn7Kbdtpc1bHoLc4ycWRidpCln6pWdjQ4ll30n70AJjRGjGO+WqIxA+nsaorFdy1DrnCtB
NjjGUhEWPC2pNInBtLCbVTUUjgXqffjY2pY4vm6eJ8Ib5QCZor3WzVAHdfzlNtecGIYDA49Mp29J
ojxbPBai6ncVQXpwORoOKIL2TVw9sRWrcm8bvk48L8QtubT0F82Tp1e6VOXsuQoWGY/7Ys+fHoLn
O6hbg4MrxgL2de6WuMGGLmY8NgJ1AUGqLZ+pLmO+GHBILxIWF/I/FMet+aMeHT78lwf5NIr1mbu1
51FZOvG6ZoVeDgZAZH3kXuxE2Li34No1Hi3mhdv3NJGq17313TtMlzQNdtN/ZBjRFDBmMJIZbSXW
Dsb/lnv1Aq2tCJ9lF2EnnOkgo01s3Y+tdAPISb1JST5T2wEpW+Q4Ozg4mPnZAuNnw5kQOP1LH5+N
Joc9ce+kyJaIQ1WaPTtbLPPzWhLW2H1tFQR7nxIK3m3YcuqkshX3CX7XtxZVQTz5HTeOUsjNAWGh
StHhmgW2a+wWgZl2y7tMS8RBpKi2yjITkm8py8qkAya0e6R26doCXhV2P0590JtsnrmZsMQoG0FE
6ibAC8qR+TOtSwxKoI476uVtivPxxM4a4c3yBQfG5eHc63xkFeoyv6Isto6m/FnAQPCD22MOiI2l
CdJjPnrabdaGbOVEZsGT0bU2gYDauK+UUaIAtG8eJ7xVbrRQjbI8kSZ1Ypw8SWuY2dLi+sBdUZ8t
eXI7O+iBfHRdDI/SL7EsgEXXnq8hWK0Kv0lUsNRDK5hJ9j2IUaoK4GhDptcppyZ/Xz8F0R15s0Pq
rNv9DosWBhCp8+KDtlJeMQgBYLbgN6hNdexo4nq3udowoQTHueQoKuC4LljIKU3oGqHiI/RLoa6F
4XZKhQWRgssvcxSc9D/JRujJBwfE0LaG8qAMLs/jhHKKuHh31Lfr1ZkeDzCUloAx9r2aGlLGal+l
b2bbp1wIFrB/LlLtmpr8C4m6PXalu2g2YKBSwXhDXjX2end5JNpH5VLjIVQ8/6a6g3wHL48jU7cM
bsB0YX7DYMz9VElV0SKPGdP0r0FoRfvh1H8sHn9ISDx/ZUx3PvYQ73L4ezc1rngzKZipOhwU6Tj6
Uh9JJnF6IOhg/xD0wf6g3FKTwYUl9C5N5ZcOHjwrZcBEhrdvcmYLAyGNnhUDBa5+2AOevQFEj6Pg
myy7AjSSpkarCgjqlH+Y6h0IdcNwasPTBKsVDaakcBcjHoMZxe6qRNypnFe/O3SQpN1PnmozIcZg
KC28fpW3bxq7VBpniOfdZshxTwOPkHcLUIFZ4zHaaLLIBWxApbJP7D3a1f0nW2YnlymAcU8noc94
E5QXJ+9lsGwhlZSIjjLRhcb1GLJlbg1IZkabwX2xwNBydHmqJHoGzoSttmCFMmFTRQ337YOGNwfA
taaXoE24KG6YTnrOjCe4XZOSFRduakNDYmocuJiumqtqkXhvpPSr5qKzUzT2FPPeZ6OKtR0cq0fF
WINtsvdTUysOkHJNgr/Cm8ajgdgGGyIYTkLDxReCkqFPgF61SKCLplwSqqOj8HF5BWYgcwzh9RZi
1rgb7xahxEh49B5lNch0eLVS1Lw5BVI98xSoSqLTqstXd8uGYShDc7AQVSZnXsMpHTotTcZZjktL
icQAyRP8uI6DUWy5u3k7hwpIqWUKNzswaN78liK6Y8mfCOhcwnAJbwEx0bnKtzrqWyQLhBMHquo4
jWhfN4c3qbeW6bnYEo9+bwxwL/xaVjEywgRtwQzeFIB18IH8BuyizBevawTFvPP5xBp25xgDIuA9
69bJ4EkP/f9nhrLD0KTO97Lfy2fVRyMiXDnygSO7kjM9ArYzxFOGFsZd/jojm/S1I5CTZNoQG8QW
3CwfS0v9oFx6HHRcKQ5dEKDh7sWkGNznn+4xcU3Nz3Lyd63/0/bgDksEJ2AZ/qKs+/aSgM+CjUTU
Ks1HhN3xVT+KWBbrpaYEYa3ngREmlsF19gxt58b8SzK7DeQH8SASolcaILTP4iHCc4KhZQDVuiit
YPi7ffgqibrKBMWrYm7ZKfXf8uZ4tnxirR5JkPQLfzNIrlw58L8ObZmx+bx3xs0OCVPAuGek3PyP
MuBoa3Mry8BgC4iSByD8wlEU9r5d9f/K4T/6O5Psd60GWOZlxlwnBEahaeMULB6aS8jIaLWTYTTf
QFx7a/Y/dtum03J4ayZogJpmPLwx2D0KcNs7930uwvfQRPo12Oak+p5C7UiAhYdqMHPfBsQCPzyW
VfMda4XNJTMIHd9r/ZIcTWv3AWl9Z/APMj7sBY/jskE33dV7BeYSGPBY5JEi3Q398dQE9jHN82T0
h//KbSKmxU48KoQdH3PddBsYcd73uYtHarWYg195RYD9KBrdrPfPbFiNzGiQXvV3HEsBvgBw13Gx
mOXmcDSLUipx+sthgzfxpJEHnDb/stybeUW5GzMq5A6naL0IP40gUtldPRMD3Wwwy+vN9/5MtDmG
t5qSORdhGDr+iDaY6XYIAnZH3ITadzHeOgktVcS95afMGyU1wf4ay17rBYBbR0iV5V8OAA/shUSF
mEy5Cs9PnO8GjS6XC53F3v2dh/6S4t8VpWpW3TuubbDTZGcYw3jIShkPI5XYS2DGfrPTFMIsTVL8
sD403J3IN34/fI7KB66uQY926GKaCchlm9gkZzCZIaCF4QQmAjQofCOGxugffi4bOcN6LeuoItH5
LXmdDDKCkMz3QW8JQ42DDb+2pPBfb4eaBmZm+sf5gQzBCKOjevdpTaEbL/X6qIZ8GAioEHBkr0Fl
C62Xjz8f/pwdM2xNnwAhZYRwgRrhNkvUjBVNSLxdi8lV5D4i4HN+c+LjEOh+dD9t9oIDRYABwste
sJgw27lP1pyS9yrdpKAHMfYuhRSf7PPPLiF7h+f0ZeMOAp2UzUFgvxpjWqZa7hjKTe9RSutjGzZs
+U0MzPxxLgQc4yMwL/YkpiwKhMGytkI73PTxyisQzXfgye0rxjUZmIvca3VfdqkS7rjqZMcTTKyM
w5k5IzQVAp0yzeHmXsu/fD5fD9E/KUIDvRAcfR3glyNGX8HOioXy+S998oYiBxVLbKnl3Pc4+1xa
fFKBLvGxrx4/hSuOJqQ2cM2f/fSvGZSEVbcXKsZuzGV9d49g0nynUnHoi2qQw2/1FrV4SKzp4WNF
oV1P1esMira3FNCJfvjmIQJhDiXoGqPP1eanSJdinKveZcScFey/jzPBrJx2P3QcbfLG6nT5WERZ
haD8Q4JBGSMtmE8V+7AjsXTk2rjNn7SNqklPk7PexMUPdDsUHqXvOC2oomonLXq+JrrRVx4X60Om
autHJ1sTqKvDvcu0MAsJXMjEuVwqVKYHpN3RAPApAxFZYGq4XvXkui1nQdcIZU1HqyyfHJkEnlwP
T1/sRSkc2jWHdYOt1+yLYl466WOjNwHlClZsmTUscA/x0vRAVyTkTiQJxnkhfO6UBmTFz2LdGu11
hc5WyCSG7nJYa1z39mfIc19wOn5cY5OblaDYOBHGhHApea9IHREJGAWQnZ74cRxwPqm2hCGNWXZ8
VJt5pOxXu8BiYHEKUR8PWLPx5j5uD/9S7u7qnGAnNOruKt6bDWuQuN1ZYLEtwTsZR07cWaigj0gH
RD3Tqspe9WJ4YR8QNN7Q8nNCJx9orSSbJhk2tvcC6OOUVzgtJ8X9gIbQda7ETB6D5zp2+qCrHm4O
cN8kgVLPKQwhuTEViTkfc9Lf0ZxJgGD7eEubNj/FMUHcTgpnu5FZ3cLC+NUoBDRCRQtzYVKcy5wz
xCFOUqyRV52G8yHKA3YA5bHtVeo4+BvNWPkWtwkXX/wsAfESB1XVZeG9VgezTdRYGb/0ThJo8g9E
CAFDcNVoR5ybD9WFoNiam1T6dE3aSKl54aXrMUmKa2VZBw+BsWsqCZTHk4kjUw3gMsKWfB7C4hhH
edBDy+rMIM4+neHq2oJKu8LfNq4WLqO9UV8O+geTBOjVH/dfWK3r2ri1AlC8b1QbpyWs2X6Ll64d
BggWoOcXIwOsrCD3pRMTFfyPbMglBko/055uaMKIsdIS3Uh90hu1dJ94DtBBEGTXTUUMQfpGiPkk
oYQM5mcDc83/jykpKgmglRdl7GVxDPIKDyS9KOKgmfIkdzFxoM7x9fXK4tIVFnH3I0t+KFngyz93
UKVmU5P/vDqJV+n7JreyOW3FJvWIw93E2+Dg0lS/PsK3QDDWVT0qsnQxyrz43sQfO/E8o7q3HDgn
7V3zz+rqAvfvIczJJWbq2JcE4yQlp0MtoD0GOZyV+BS85OUyaS1AN0HLRTrJGCxltkIwawuMc+t6
N4j448jHf2QownrVieRGK2OQ8XjglFAwQX+2I3Mt2zPz84936I0Q6ntVoO0NFp9qFqUw8vC4M4gQ
6D7WNhC1pDxwpy9E2KvfZbfJcmDcBJjJhZP49ApPy5T/FoPxo5wLj0O0tOT7BSynnDFN4EpmTu4v
QUOe9KrTNEemaytCRARD67Zsa79+/+1snK/KTHkubVK+MXT+v6LnZjIJ8lGsZWl8yYZdJof3Bx7M
nlxcWST9nkSEIhae5XJTyl3T9BGiAT7WoBsg7E3mv0p27MXeE6d0/m9RR3uaI/BY+smoJ24vfAz5
5FmflvfzgIit0vqAGQo+DwpWeFtsHHnyYJHMh+Xx/KtDQICfNi36rJebKkpo10t/ti0htD4Jw6kJ
bWeK9WS330HmsVwqZumgmCX4MDW1Uh1jo/sFoNYpThqYkDNMDKtD4Hn4/5jjCEKu8Etx7qbpNj9b
73IdJzeryfHfUu4r+c0RCSP14sbw2j0hVhch21Mi7Ov3qq+8UUtm2qE/N0uCdElvK4kzXY7XZ2KM
Jtj64YZsZSIsUCDWcPkynQVWg6tjlzt+nC7g1y++M6chIpFbsi0Xg/sMHN0utMkkkunPYcOObfCn
/HxZjKjrR3dTEHFJzvVnDh7OEvwznnObW4orfpLmpv6EIXArLbaOF8eUklkrBOAyFZ2XrDy+JaSI
bz+C5NmThGWe6M0UkjPDIzsXWoxZ4sIzvD2aCxCFi/zTRh37W9ZpJJ3OOhg2UUE9gw3VFucS6VgF
RqP+nMQuIignUyYC5k3YxjfgcI3euw506+WQyC5B4hG0eEqwyqaTLQqMvkle5oN2TlInxi82CIQ5
RFaFophRgHom+drVvjh19Nzd8s+y3hvTyDAe8JnJMV59G+vSqviCH7aMOzsivqqDDtcosnEuP5L5
59h3iocpHl+Ozie5ja3INmsfd0yiA/B778tXJo0TL5sZhdzsi5KcWKKKKkQTNqZcOKNDKAwrREYh
EoqR8co3bNmcCjs9Ecw+sno3Z71PzF3D2GTDsxHaifPyHWcOnOsn0YtFwvsggm+KyQ8h3A65UFrU
HGyzlzNm3T0AKXAPhhlgkLqHWtdTen7yEkCzWq1h1r8KhEBW10psEsIXmUOXni/7c4LTsv79PHXZ
AsJt9XFFSlSyW3ScacyuEJYtNxkX21tPabEhYL0e9XLF3qkGBzjJKk1OyFGz9VMnK1EBFL293VfI
6uvipGS8zdZhpl1ZNSb3CD4LPTr2J2X0Np7fTHkS/Gg14Pk9QJE8hUM4W67HdT/NcWRJKvDX6rF0
A41l7GPFwYJ3yh8QmYDIvuIaP8SI/E0/HShmx2liq4qBlY66VRXf0IaVyZ8bgM3FbP1KGdvfckP7
r2eB4sGADRpKV8c70hyj4sjIxFkEdap3SVTS/wEvlKyFDN9q38S+Xl1YMRZiUqHMF9xEvDcDNy9I
AtMDLeUhWqhfKsLyyw8B+jcT1Qmd12y6s8odtrM+p6yaiQSolL6YkYuV63wb7wU2vVxmH6oqdJDa
hzA4SSc1xtfbUqCgFQpaW6FG4bdaZa6n1RGkBuOclkMT12LW235yM6TpM2PkBgC9pNA+DAQDGdL4
VNHkzRGIkXEu+h+GftqcPifUDMp8F2vnlsk6tCJtmH6JHtF5T1jeB7PQG+1LFQs0FvfywlfgXjI0
wNP8aVHdVGgslylH3jMLqu6s+51sXF2eSzqYr9hXv3Xinbgw923MGPrHjb7603Wbh1o+y0UKloIM
I2afT4ZJjUY7bFdS8MmoUrpbeoVSHSgZ22+/TuE7je3T235nLcPPfxEgZi8XtEQpz4yVRn/03jGh
gWqptyalb/iHHG0L4IEa9L7Yek4AcCd1EcysfJDhfOtweY/djOQ0sUFkp1AO3Jqi65NX6GxwGQiB
7nkf8J8HasPqhtGRKqCUuQe3PbSsH0a6MszkG+0VGTAzUBTmnTraofz/XCof+4WxikX3cqpWhyp1
4cu1udDRJSxY4SyiZVAWQC3ZRBIEwbQM4xjnxPxLNBFkAy7jJezXaINLKByXvqEhmf9gUMVECBIa
Nic/SwxJ0b3rZIgEZK9AFjHoHGBwc2trgGNsRsIAy6/2KOLx3Ys+CvJjpd+syeZd0N4nU5mGCfbP
TZTGYbfV5/RyNZ4Rh7DdS4xby/hhxacIRXwk97ZNv3aeyWDfwsdl9hGLPFt8CBrLuzp7HBqJB8Zv
wvWJpGuVR/wJE6exAZqn20bgIGfJLoGOOGam1cYarHIpnhI69M6gK2wjS9wRh41iCj00MjYboFt1
tlMXMMHKTKQHkY84CQW2KM9eWSjRVzSP7ntLXox5djoJ+Td+GqQkyyH2Yys1w68o7ma95zkGqNEe
yhCnJ9Qa4YR+89EBH3dDOSeHnkL8ccwWJh8h0GEH8BaSeR3BKzeQ7Ow+ZThU78FqngSx169shobk
oAp5dftwko23iKa5qD6bR++HI6qTmtdVDqf6X/xLuivwWHuMFd0E2NhHAhznnkcR5lh8Qr5bjiKP
1YnBlG9gttyUWJIuVmhZ8r7dbMTCV3y2A4rSNZGqdajJKHBw0DGnEBkk0xkn8b4Is/ofcDxD0P5n
5XnFA+Dg0edMhwF2HW674vDINouPytlEMgY+Vb7OFcFEcIGpOEx0RTPF+7y7Di5U/0FN5gkQhcJ+
eZTz4bQd8wy50JSVl+mRHAt6E7xAfHndR3jjfa5lesffkkH+WDtxClHMefPuSL0hTgIK6oJ1nfqZ
//RPFl57EZE+gsvIL7U6o9ZtUsdmV3GIzo/sVaecvjTD2a7QSmgXpxaX0cxHJEDb6FBrpX36U9RP
hQ0nH2IWMYaK97YV/Zq+nOGFb2dvIfsaYLaMi/FoTm9fC6GCDZNb9PbnMy8lUZeldt2lau6zK5TR
hPQl0/dDIlSA16hL453J1bDTpcS0J+RuovU2ocFb2CErarVFDNvqQbMnxBp1WSlqmtdVFF/uiz2s
yb76en4yYqyyJ2JlUNNb6ktZnhkMtIMAYgnsm6Q7LYF3XQmFhKzu6ZhmhEPjynNkoqyEqFSWwr4a
UV2bFFAG2SXV5S/ab896NrF+oVr0T+CrE0iK3wwIIbHT0wQlEi5k1nCuScXARzcFnVqYl8kyqytz
o7lbxeLSmNRV4oP2yvjaqiXZW3wbc0Dh8BSC8rmr/dj8/ozAJn6y5EAec0QeIOnLwet2DamSe2H2
4V4ExcTFVFJ2K6145LEA7PcB8KbDuvhZSJYAlIGLpH8ocKgbLvRxDGthnhFqyjyKB1oUW3M9F67+
RXysiZNNWNEFLWrUxff9CsR2DwtzBSyep7Qn2BUtbSkL2JE1BQ45Wn6idPLG8qHlsOcuLPO2LbO2
C/o7b4wmr8+T86FGuODhVPJL9V12ddqFOBcdXNKIp1zV4MePbMhm/veeUOsH+OuA/hzppHF+4uuG
BRBZK5o/xhh4+NaQXRkpEtgGAGSeaZ7KWIyvgtbkuDE1Oi9iBlPwzHv6CMtFO90Wrs/kD7Ghcogt
+aLRbJSbq4VmAEOnuirAg6T8uNRMNpeO91t110IfzJXz8BAjTBx/krMmmLjBnUN+A3F4P56TeiSP
tKNjjOdaGtVeCKQ1GiZ+W/l0fPg53iwymMsBR6Msm2IPUOsbxveml6KrjuMgvzyOIaXTHxfIhVWO
TBajNXsHwpajSxitTt0YVtboAPkYk4r4+F6wTCKjnMmTZNdNN2ahrN+RvYb3tB1/6Yyc7NWBGAeW
rIv8vVUzZX0exuFwwQjqZJA/aDpTct22e9u4TLopyf8Wi4CR3IJO2yBPMojXfabwst+rSG31UE6P
3WAEGxzZkwCBmWNbGvuFSJKzfE5Fy16b8R9Yhl1XAqk+hinnb48j7j9rHF0pWbxCNNJ+TsC3i/bn
cRcc7akM0/Ll964bYbUrs14HUM/oGGyfGWNRd1DAcGxHGTOFU6EaquU4ChAqReV3wyZrRQH2iVrR
Q/YBg8llgGKaylVz5kjitOhS1ofg60xc/boPEc0mPrPNCKtyA249jOPkVXAuNN2qAgzHISBurtRz
wTbWt3CpwRl06nNSmWL0u4cwe5lqOI/GxL7nfgSU5ZgEQzGnK1UKSpcS32JdnvpJypP/p+4ew0yb
2EZU9auBT0Db8IBQTEew41rH1QvUpaK8+A2ugze6KIUqcXv/h2TCv2iKbwDtgmU++FVwNZ/olg5j
Dk6NbO9eecCPWNwN7IpYZjNLpikDdlionh7Z7T4TD27YBIzXHlbMdRErqowR2vA6EE3MAjR+fEjG
RVw41gJSKc7n0Cl9xXGLj+L+fuFTaTLWOXQGIXXl378leuF9YIFvcJIOHhOpcaUEJQZNLVeW4wNw
z2y2Rxw6M+TlYjipXHhvrI4dXLIsdYNCiJHB3vmKXNLSJ2ugvhIUw9K0NGRpgYIx/ytG4NV2lDzy
Mi+EDo/zb9NQqJIWFVdrV2shfWJlyh8z5/ruUES2AdtfXE7zlxc26loJ3kiz5RaNJTVehjcyUOgq
+uyXLV5BvrtY91XCdJpqfE29jGtTIIjmkzSRrzZlHN72C9Rpwg/lfL6DWNPklVN9PfsCzEcvXTd9
Mn3lZNA89S6TgbcJrz+CEjVaMU+IymF4u9wvB75JjxKNMPq8sfYOkCOeu6xgf3RLTJAOFO/jCVrD
MiuKU3MyTojZb60lrBvPimrUxeumyOdE1sz2oV/FpdwPfcf43uILMgfj9mOSnC2EBz5Tt3kg5bZ2
1Vx79cI3rMYwtsIpk+XXXgFlDkS2IIf+kKwUKMOCBYuCW9fJeke+G/vkN6l26qy496uMS1rrn/0a
O81AozyggKyI2832Uab1l75tGPaAw17AA1f422/38m85GnBRKMoG5s4otNseLJJNeyu06fVh7m0X
seaBekKyj4eBrk2McBPVkBckJwRjOzLaqHirYGbP5A4c5/MWTBd8xTGvxm38jR9SxWtCs5oF4+yZ
UvxWFbWr1iUGN4RphiM6zUxfO7FVe+4zP+9PBYXfsnTeXSErXXsjDPf4ifr9A/gvktcpZVRXvxAw
+ub7SHM0JSskbnkuopBE4xGCJ2zEkpapHYj7XYpMyHB6KjBCulXCzwUgwODpQ6WtLirjlGYpRgrV
E9wFjG0CBqxtgx11wFfB49pTOvXGI+N5y/sNWi4aAZWvSXiDEwDgo7880kwl971UzN0ZVfdwAxuw
ouGwdcjB4pqL8uJFhFs0K1AnckQgSA1epefBAEHXwT9TOzVg9aAc+DIJH7flodNua6W8UoZAj2ku
Lq1JUGeWxxd9gOF0FnhWYKniLltoiq1fIrlVmDaep3iEXaDrxIjorbfTQY5poeQRSj1lWBe+Lt8V
g/KztmEwmT4lYR3FS+aiJ7Ur5VOQpiXLkCRMcdoNA8estFG9JDpleGbJY2xj9GrX1pcDBvgFMD8M
36LJomiMn+lWq2Mkd5evT2q/TuuL3UYwc9O/DZWtLyPGbvX/0hW0BUAovUz7Jr47xSg+T8/9xu69
FypIxE0Va/zLdbCyp3NGCzSy7cNx75Sxx7mwx3YcmRq0FLFKYixJ9HB+73KI9YnDgJRbcAFiUZ2w
r4f5EqkcJqfapsViHogkRFLwmipIHO+4ky0rJ0TWOnVyQOa1UvsVdoxUsMlOUbUeRV06rMVsMUXQ
VL4jVwIgIxEcDZbG4mnQrGDvNtxU2IK0YotbXGugDFl5W4o3eUH50HJwdHxOmbQ1x6TT6Tf/gPib
9l3UAHHNelSXDeEdZkUmYuO07IwwfhBef9QOgXEg8wIe+5wdxWtad1La7WB31DDME7LW9eWPaCom
ph3fEuhd0GpOP2s+mr8alFs/oGcf2GvachA9T8NdxVLkFNxflSz6sHmZitfIkuDBeLAexlqdLebd
TdCubsGcgqpAipTWfZ7xi/mVXj2mY994OFv//0IVs5FgDwcs/cyJfXeq0MUh3n6qw9K19AV39hPZ
KP+c2jNyvKuaXaBHl0ZVu2rmZLNuloU9QZJlOO3AdhDzJaL3G57M3cB5w7mW8wpYNLyZwoYYu4Me
RfCljoqeyre1bNzIGl5vVFLaBEP4QTAvq8h8ZJDKKIw6lbTFDUTsuexHGWUAm9H0XwzgoslecqL2
6diu7idjSFrQ3ap1JmSd006eh1fzALKiG130Cg8aL1a+XUfomMPhXPq8GiGOfTY/4hi+AwOolyNj
uTCJAwCBtZlsUXtqlY4XLBAFNuUnX/vInD0IBp0VyNZ6/1epeOgu+Hy37dkXXnyfSC69e8YteF2L
hir3Zi2csz1nT506nrLlU5ZMslskeqqhfpXX94KZPaeyqoNBHeFKranbl/2UN/TMWslP/fVffF89
GJv70IUH5SgXsqeeG3XApMzOtMT/t0KFlt7P5nj/CO6sRJAqvWQOoH0oz1joq/8JSDWD9cmuAyjX
H90QtHzfmyhErMZmZDp16jUSpMXs/P4YVKnPxJBcbn7sTkUfo26ub4leUQeKJVpXs680lAzddCbg
qi+/tz/78oATbElCGr6RZmEXF3lB2JMV9Gm8q5mVxC8EEpYXE1WbGE+xuL1uUpOnknHLParCdJ6g
fee681ecTzgf7l13Ju/HE/PJ3uC3TUjIDmjd5rmdniVR7MSkxp/Uvw45WOPgWv8ppTqzAchOfT0G
YWXgVsWTcaIf3QVQi+N/mxWLENmKl5BkhuO3jOnBYePbIRlxS7bKylDmuSioFh0frAq6HEvlRGyi
1mUpfEqYKmat9IWFZ5m1zk8uKrA6WhAW1IH6q/vTMp6u9qrdVlkUnPlZRucnqrJhXMyS8s5KeAWc
9ZQoy08+bX3vI/GDPoSZ2/bvnPgoWR7JMH68FILEVl3Zq3vYnMDs8l1HAkq2ImxYSySiQOuWK2B/
YKRaX45GMuQ0RFdBVz7bAm6QF+FBhaBj0tQlttJm1vIsoN2lT6z0WuGTT1JHjcZ3vmctr3cMbRrO
KzHTSsNuoH7YUoRD5pllgT/xRfz6tTsYvBlXMC5G5X7ITXRS8PjXeqRHvrONWSv2GGGn8N6kkGYH
m22L6xD6yxNJ/0PY6MYoaEF1+F4mVHBnePUGksjmrOhNwPvpxlc3VlYH/IU58Th1+tJH3fRJ9SSW
NJ0ioXvGGq/GzlDP167BTKmcpZ9CiPqSwCA/GnC8gmmLVOX+NUMdJxDeMDneaFaEYuA25P/XCha3
qKv/U3aF+PFkX/GuOIgmE9dUkMKiS3Nth/CepRQcqjS1iTnr49714f0gbi17YZ1I0gt+hX5zzDNr
lZgrROCyGZJyofzw0R6Af+0RZPcIrTJO4IkQ48im7hJ/eDITi2N4pnX7d3nYnHW+G/hfyjUwqLeS
pOxE1Ri4rsNufNLyNOYg+d0FquRODl4hBNLNm81Gy1zbWepLVDO54MG3ycZkpF8YGQEhz/3tItEk
ly/JVotHNKqfpKopH+KfOheHwYY4YrBL9k7rBu4CoEEwiI2Q1Kb3ww17vdJJ2Eg5rWSufpQGKqmE
mf15b/4EDKhgWkNfyvqaTzXSaPcHlfQTd2xyWU3d4tQNn7RU19wLV5AnLybsfdO0f6JgE0pGfoYr
qfBAaVe6g5EA2s/kWAN2IAwfG8S/q8ood0yZ/TwvzJILtLEVAls1YLo22QNZlr+4e8fl7t9nvI5H
PPjj1WZmd74g1u4hmgy3H8XtxEQk/3TcLruopmfskgJeUklQT8sEkgnYpSvE4vA3y+x9MbcEn2/+
2LQDpoTRrxWLDUCq+gzopbM2OtBqi1Palm5jkF0IWAezOFUoeNbAWtjCMlVPZaooMPrPplD79bOK
gyuaVZ/+cwqgM8CmCdTOr23cvaGNQKSiYNA4ieTF+ZeNE/E6iCcGvfMSFrYUNwhYXd5baAiY2e3J
uAKgljuPq+q3DjT6Gbk6u1y7DJB6l/Tpq0rxCRS1eLeox4XYjVW/Ra56BAf9Py4g1g3h5roRUi36
mQvr2FcgjVmH8IvRrh+2GCc8bU3GMa0+3oMbr0X4dVoZdEvWDge/K/oCZvuQcnvY0ydCK3T1MIYm
QPSHhSiIT6rudIMBo3B9lYgNR1BgHsWrB+TliR2iy//jdLgaTSAuk4MsoS2Uqsls7o6eTjLijSMA
5P4yXqmozrZAqiR9xqh/dRPi7/juaO4eCTpMqdX38iNuZ6b52KAL2a29YRL/ISWR1/rNnSnuJshJ
XCILI5IFfkgINwvHlaAtjzdCim2S5w04+lmLZRoas9M8+ygE8+jnDaf//d/vhYKIktOWGu9/JZkJ
0dKjPLziv0bys0v7xim3+No+nsAupjYyKw==
`protect end_protected
