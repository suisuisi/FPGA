`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CvmaYyJzAT4gGJRlCkE1yXt5Lv9gJbr2gC0wBzixkhI3TupXRLTg9s4Z9WVWp43QDkUuM3VRZjAj
RVnqESt3JA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHyS2uxRkJ6sHR79RwG8dxYfMwySDoNzo0ZpVSoiAp/93R212I5J1LxM+7EujDw/cO/x9djlyxbz
erzC6/tIqQ2nS2hUZANmmER9YkiA1RlXlIqDOWo8pOFHNj1c4jf7Zdq7OJMDPvKF+fLgmk5Lu9Y0
15oIyfQw7L+gXpW1qEU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cfhh7YIOGyVJiZpd5j8xa2ugbHZdDDpkNcw6vvVCCgnGCfzlen3wlGk0omzzJqyVapnfg0aPFCVf
eH/noQVGu1bQkowx0JKcNE5x1v5DKH//UNI+lq09SNF0WKlMcTAGlNSUzO8kgVv9uNbKUHDXodcD
5iGh6bHMhVPSu1QKpTfJlIMd2CMz0JfDQiVbfTaAGKvrQhaqVte7pYpnqiXM7povPwt/ntWHBH4s
XSF4J4eDVLMuQmQNy3vrqFdEUqmQFtLWgNRpG2fwo19Y2lRzT3ux5SiA0Iv55uR6x7AG21x8BZlD
JC102ufirdrREfWUzlClY8zmr+TUHpTF/SgPMw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWceDgHVHZAg17Yudaw03bncVn75AJ6y0RYlYeqdZU3kMG9E1W6q5REaQAI7sMZSrC2g0zavsx4w
utskoq80P2avoebtdvBfjr/nBCQqUN3AvM3GSk85froboZgk4fCQ8UtEj2Qk7ob+ox/md7d9P9dw
2YULi+eG04dUc1g45wwF0ZoZdARk7Ml+fXMnm7zxmvqVieAEsVq6ETZN/P0pwvIpAakLTayKriGC
qcrb1S28bOuV+Na/FX9rxN6hM5aK7vSdFqja5GGs32r9UVRIkX6i7uqS9pWQDR0Qa31W3z6wrRrT
+2wzEwNMDKYuWVIM1FQo/Tp0NKa1Y+kyjahSGA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tLsJPLnIUk5FSxPTGLkNhAFldHrP7oFH8h39nfqyEmnC/AmGzR3fePfCEcee3I4TYySABpWhyXIf
m1jGiCuHfIpFkF2EJqjWmBev0bD33cbw1av2xtJRFa5gaQjxChO9URfjedFvCQWWwjlxejc9nD0N
O0V2XUDQxd573YmSBuByzshlxt3bujEd6Xeeb8N8NI8c2ZsfY4693LGdb3k6gtY9ZEoo4XuYVt6n
S2tNFVJTfQjyBEXbuCPqpwGf6bPdy2SKvTE/s4rSIVTO08J6bXDaEOBUGg13XVoJJqrayiJRVuQL
LhoiPzgOqS6ude1uUaMHE/SN9X/vt/6uOsOl2w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jgk19ieS+ZYiySHKvgAHMus0OAx0HPJ59p64LMaYK8CyW0wSM8LIn++sFz9tsOBdLj2gb8IKpSVr
SOX9XXXM2pQFSME7x8q0m+EPg9m1+ghIpW4bU/w4zVq4NBjYydZCI0Hpy+X3op0a3+eENVEw5SoK
4R/zOL7aV/2nZ//wkaw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L/BPRr/PHH5da1O06dKRr5ST8eskM6lzR1UPuTvZQ6RCsFEjTD1HgyqjW7/ypnIq7V5TYDC553+Y
rJnEENzDc6RSpzenrYxw7NrURpUedIWlCc/PEf5Zq9gu1ESkpND7t98rc+uiAz7zsn/pHD/K50NR
q9l/gcWkOCgArmADo1Lw9usrfZ8ECIPKY2kLxeTYbh4fsrCpPQsQUk4NxX3N1Q0h3RRUCdHSFc0O
lvGip/vd24OK8zXDMaQv4fPmgToFQMUvLrJXErEUeRlkpxkcX6g6Zu4RMWwwmkNIfZHpc5K8Q3RL
MMc5rARUSXbNbpf28H3iyAMZ0y+EgI0CrKwooA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
/7f/xDmW9E4evduK+G5uD+6SMjICiIY2xy0XVBgq0x0pL49qw/QwsQrqhjqtcQIbX4q8bzXbPOm7
zchoRNRJ9FLEEfBG+xvC9ANZnHAuFA55mqMpYhUWnRZIzumv0/2KLiQYDQgiLtnqmOQVJj35xlio
zO/zsaQ0NAsJJs3HMmPWuJf2cCj7U0pQNPNNrrvTQ6NbnXInYoojpbWTL5gksG7muLWzhkqfokNl
ZhZZtKsyiMgT2l4ZdNznlhwR28bo/ZyomXLNNl9pVX+ED9OspyL2RQJSIzp4WPoslixFQsDEkyMg
B1nMj+fhu0qyBttL7UTkTdWu2L93YH2HnF7LYtvOq9CBQ3uHZf0ui9srJ8R8Ldu2oH3uhxtXeFLW
gkAT9RUrL4K80xTJR405gg2CL9AjoRUSCtsxE54oeWdP2eexRXrvx1jNpgCvdEApP8fES1eFrWl5
fC9WSIquqRBCm0PPM6n1ul8Z82Bv1jFXaxHsARcM40l8ijGrxSFZxpuFmDi3yatYMAk5yE4ED8Pc
Yr8hOKof3qdd7fsj0sgmc5TloyemHmbjCJrvRUW3YIJRjwfAelWf36afjDwICezjOs1PkozRq1h9
G35nCa/s16gOMy3vqSrLFnKr7AmuYfNr6AWJ4b3XeocM08MsojwgjpqdK8emeLjfy39+0EwXbQ7O
4Ppw7ILz1YkfGeaXpRUEAvNOPDNIBof+mEruZMiLjV4wfDzLyPXbONgGYevh12G52AMjGpowGpXX
d80Dc1VHZLACeQ3qgBCaITyV4B0YWrCLu6X/2XA3h195JzNdJKnYMO7SiwWuJB1VYQOfzf0XMXqc
u+GHOmMj0dSaO0vhGIlTJ5ToNypcMoPeVuffjFEycghuH03m1tE2L4GJiJ+MoVhv7Y/zJEdz3Nvj
0upfltGo6tl62LbqNS3PJW+VbKvMWp7/zPXf0P+eh65EwE0T241wreeEpH3B3Ey7pIbUq7JbH0S9
yUHRvTGAWa0xiDLQIQzODHXb2eeYz2ChrkxpQMag+zl6BktJ6rilsDEEbMSJshs8moe0EULok1gy
iZJHlB5UN/1FHhiA4TFXumS4WDSAsBxIKSZJveagx7qmlBRe38DOln1to9tmZg845T8CehNvHkOC
7w+n8VnQBgWY0ryEMzUrbQcGjLKU9fzUkPijc1n8HJfJzCkPkh9IZ9ZRUSyhW5pih/EwL8zROC4q
qie8Jx8BFbmaR0sgJtlxw9YuTNwIqT9ZgFsAwOTO5v/91b4sXFaoyPe/yvJ/E3o56EcN0JlMDG7o
lwIIG/hf64Qc+ipTVjY93uQBounxezz2uQWyWJIWwJ2guaLt3TADEjSZWAjBfWcr4yhGAfi3SFOC
4amTS6KXlSuDhYKujlNajUVHxHlmphzWVuc3IyA1HXEBLO0FuMUs49AAly01uNppXzmQMIKWeDVv
XNL3/y4OB4F0tCAeq9aIjd9K3zc82VJ/+BFXGinwZCEpwVLCbLqACERnUAZhi7yPZ+GUCRo1cbOL
nT3+f4QCB05fvedzgfOLw6JkHns5kRyZKnWQR4WaSyJwn8+2OY/uZ7vgni4lIDid1M8thPTFQxwa
kgxETJjzE74gIUB2IDtsJeYKfDpPqPCf3CB+siWCc2DYhXhkYevebA0fIpK65Gdf9W7oPHipKjH4
xkTowq77zVJBk/b7kVqISAYSDN3HOktI1QTJYKe4rmNRKpcLt7r81ry8xPNfFjB+5+uYODKJn2yL
8EHO3UeiTiuVUlHWD8+8Exq+eEbRXIQz2zar67fuXvS91um3dE2bh6Pz+mwW6o2j6vFO4lQnE2UW
n2p68VcqxIGzA8BOOUcASinQYAnwlM5rh8QVBWGR2PDZftGWSCVinzJGcHH001Jiq57nwsizJh2H
0DbBYGZDDfWBufslU5eCJLUX8LgMa4S9e+39gbPMG0Zk4fzbO3XOhkLKa7OPLD4fo+W9KyNLgNJq
ikIwWtclUeU209GpoOevHyYSSmyf1g31bhpZO9ASGc1JCCqjkOcTTCeXrWKUUlEzuwu1WAcERp9y
1r3FAVLfULFbXdn6XMtwa52yQWd8lPzphiQHheR4tVncJMAbF+lAns1n7KMpxQvawnLrSlQG3ve/
dylCtLxGPf+bVWTFCU9nIMI743gwUVhdnAqdlNc2wLPxiqVfhTOzZUevyK68HSS1idcQVHMtawsQ
s3HdY7dgT8pUH/BClb0Ll97wBh062LFNkQNP3yM+Z3XmqXxtcVC4/jO06X4QvNANfmShWIF+8gAY
D5aVS2H/nhXRvQnmIz+fjTFg3+XnqaBI9pBVlA2sw5SUmA7HJLQf5dWCQpmm/lnOqho8OlEWKoIz
g/1gRLyA2b4HoH08mRk9vxNUepv4T267h+hlsCPp/VWkNiPsxVQeG/vCdWfLVLxsOOUpyRGT2h9g
hKrjT0PTwotqf5tLFI0+2il1jKT6tL1dVVbko1PZP8r51VcMBbKma2BV2Bv1CLCP1nuElKL7bUCC
+/HwyOfk11X39UT7fwlRuuYKM7hNaCbpM3F8gpVqcPc/8HxxzYyvGyUrgyu2U19gtTD3CErOffei
LzcIADW8d8WJT+HRGMWh9SNCCJBW7/7bW5aUdYapDox9udW/xCJ7AUI+QldZos9sn+yNhdWzqUf3
Ag4Z4Iva9Zk+ms2AXCIScSLS53XVaBn01880e/YolXC4b4xiTGb3+7AeK01Hh8vNGVUur/jCUoU4
Y9WPRYqyHN1aBfoDOIjSgdwrGFQHj2haQ7S1CFSryNyvWO06ZbFcV+rIGHcsDbZJ6E+ezjSYydKN
kQzIef1XTwLhp6VrXI1fhgqzo3YhxWH9ipJiJ6Bg5BKzn0V1c0wEkva98EZYZ0itdPVja/1c0FOM
C+GuFgTugHXk7rRcim4GHuzgoFfKLOZOmWGS7lXPfOQeeEzCvGOtnEtUSb8pVopmQv+M4EyIhPyX
Wq5pdzB12Mbe94ctAbistv5/UNa02UIey0XZfou6TNT5XCcmwR5aYB646jEHe3MOWz3pMrq2Fs1z
QAv6S+em8PjzbtHK2bdQfsWqsJ88htpPGvoqlMnZAJBD+sJM8nHWRHUd80TU3DMtO5OlKfTTuME8
wwctIE4U1lijCDaKdS3JrwdNG9fERWH7xnd5VkAqSAECrAvNsEs1ms/2x7MQuOF3FxLFVeF+afVo
r8+PAH0twLxcDFUsgiE9Le2iW8jz3WFMqFsp1uvMALdq+/oCfiaWOaAu+uOFfQFJaoPpnaCYdgrW
M9/l5Z32jqY+HtRt1qnVw0K44Lulu9aCLSgK35D5HHHzcEf7DFBqPPSFb7oNuuypNODie4AJOaog
ZEUK0+FhnCpSi46KnFiSdM+W6pcefnaAjUHpbEAFJYQm0PQgh+g6YhYzWJ3mlyGSbaAMFPWkZgCz
CqDC/kwmrTKB4URaTbVGhm1DRs2ccXD38wAAdRUkeH7GHtxGUZNeFdkHbUsTEnKjRP6A4YReVK2p
IiDv8P8F6ZPnb7g1v+NLLRMAA0pI7m5kTUtqtQO6vZLua6Xz5EL8FdArsV+UgonzvQ0p29ULAbjm
Pcg76TR5N5Tyl4O4qXyOPpIVNjK8W3NcSVCQyM8mvB4Kus9oZPdgOWio4+WBs0jjMMqMog1rhRfh
lu/oU4Ks17bh7YCSa4B0Iln/kRcs6nl8jNAP/GsrhOZegiHDXVlmxlwypGbqDbSyg3F/RjS2yovM
K2i31wtM4jU+OAXY8AdzjQoPUtT8ZQoB3JVqsydDIeDSHLV/zFEtRZucb3u7Pbt8JmJbriK4aNJy
1NcX26mQU+6NoiyVxTZVSdkywUTX74+u0WHahGNDEybkSSwyHEgl6XhDm0kdwfTUboYqVvK+oiIQ
vH+85Q/HREytZr5IksSPGHTAuKl8hlPfvOw8f1sjk2UHbbVfznBXFEYuyC8e5tTY60YXfuviRXZJ
enxTVj+RC5va2NE+Kls55NV/ICGlwYSxOqH2dOclt13i/w9y/7OFA+GB/8haDQAe0pBDRRqOICNk
3tCkgtAmrbGDC8JbztcdegbiSR99wftNOzpjLEOU6vA2sv8xysnVsaja2i6abl9Txqfp57+g2cpg
smqYNteRAy3ZF7KwCBudgzhwDtsxl1BpjcE+CW7DMwdJ0VynXvo9ku8ePeHdzmJYhlfxuhEw94vF
An8sEJyOF2x9wsr/jbm0XwNnFYu68IEygTuEHrARlk6sANd6hNv+frkTEACfJjnyDwlne6Sl8D48
A51UU5RwdKlnohnD9nlrUsiyGhLM1DwheBhj7e9B7jtr4pmyQIWxTrt+CwuLirxRAE2CUhttHoYE
8qwHh+XnOnm7anX5Ioo6hbOahEKcCAqpby8fioCn7L1uEIkjJZiT9Ykbi7QNAsinwf3g+qb7GSs6
DOfQ+BaTaTWFzPdR5MW1ezUD+6vZpsOD3uQQUAYLd179AV5y9h87QByIqjc02sT2kssJ8ETvRQt1
lUj2dmj/UjMDf002Zmzfm/KQA00INx+sXKCHj6R4YXbqcTJLPS84EqJld4Coa3K1T2CSwnYXnQ45
JtS8CiSEmrJnTqrWfJfqKpMnze84nfYzTisC3kW+9/TH3cZsIDK+O9ld1CnwaZBnWvmqzLg7hyFt
J3o7YqOCjSlw9TpRwsbYQ2hE/mtMgp3wstUHY73/thnJ7AEa9KTnvV1QFboODyDn6L6RsJo/+ORi
f9V3CCmh3r2XmaQel/y3GY11zwm4o3aZ6hhdJFkF0N2DL8Zd48HxjoWSSJuk6xs+WOQ0iFgNjMvH
heEeKTL8pGL4+FT5G4CVIWSzkqRhxRTh6BSFzpgKBIJcleAjHX/rExYXD7VGwcUeVnnvEPYyxxrZ
2qctf2/uWC3yXGOgZiCMt1s45qubpMLAUR2eZEA2DQOhzR+LNrB6tKRwk6IW7pBfeF/te3UxPp1E
tzzzKfDKmhglKc+fxDYTIZXl8NYBSjRWqOvNQMGGrR/tVzb/1ITkxu7OwhsSwHY+fCpVFTBPKDq2
faw3alywGjjo1R3WzaHHSSVaqeejpGNj+q9eoR9ablxJW21R0YwmhE5WfbGFGlDmFg356vb8q/Q6
fY2dPJ9U3kW42RstH6dv3L7SOXkRGITU99A7MD0uFASizxtVexQOd9JTrkVjFq8FEm5LsbKZKZai
uZ827rLuD8TZUpFCu0HXcDQ/AnrrypJtTZ5RH4xXvVCYjkmf9qPq1wH8CQTCCO43vHoE6K6QytDw
bb4mogqx9XcNKjmeubXupnuw/TLtqvc75+bwPnI/RvxR1Az9y86O1fUih5ZpkMHm4DHyvGQkDFM7
ZhcR3dl1fgji6t8t77bU+/BjEAsQ5neTuYveP4jaQFW3U5wZhW9nYjLa0UDeSV8equXBLyLFFof8
VgbDx/D9e/QNY0Se7G4aWCbEoVrp2Ai6rtq1KkZ5bMSdWZ5jdAkD733Fix8Y7jnmhZa0Ej2XkHZx
JBWNCqX+QW71jNuvHB2hVwWIT6siS9VVh8RdobM1R/JuC8hjTVWrBQ8/pwrcQ9SnvHAOoTrGqaGM
WsZddHusqamHpkg+6eN5A4LYlIK+oqHFupnO6PLIlTtjtcKk46wchb831KMZ6R7I5cj/fLpgsCld
OjJYaEyDxT1OaLo7q/+VD2IHqBbwZmeqDbg8OGJdh/6ytffvoqyAKVxD3aJPg/yxzFITyc0spD1y
JMid4wzMjlZl/2VYVgEpQCArZNxHOceIgNLCd23QlukyQIub/PdBSHmnHLk5bQClBMImVa1RunhQ
QazplbHWd/2aFZvE9rYByhQfz4nxdwj7uOpp4gsbat3U8t+Z9XVTLfLuHNNKvMG9yDhU9Y8qB9rw
f0KQXAJvjTlqNw9v1nYWYho93i/+tE0aMDsWu2G4ollIMgUrTGMQXvQvdDFJZR+/8O8OLG1QZbOo
mtvDHGLNAcMXrOcdp9ODn9XD/A+1CBhdVixlFf28pZg5qe9mEedww4yIcIL82UkdQ2b4k9aHX+X1
PtVoInBv3Yp4xZlqZEVQDBmAVZiv+PNDQVE+Wq9tUaYpPAXYZ7nDz+E98moLf6dkThvu7ixgj2iv
D9Pqb4SpzbXLAhcuSATBw61GJy+JBbh7H2L0/rlzxQZCanIHVOE5/S4OjtD+Fd5TpdgDCNVvsovE
kAKhrtw9R2vxTdcUtpLMxn+YgF15vEO0Vds+8pm+kTTPyUi5wd/z9WcRBoSQPmeBDutSinVZJFlJ
ubVXUdI8xfhuV68ouCr1cQSN8LKLSIF7uTKqZcYj0rhawFAsLwJArcGU1x/I+4DflRYm9hlDYU95
MMDMtwLWHxIQ5aOaVePsKfFXpuEACJZk6f4cNllXfsuGfdi6zAJinpYiZBYq/RDcj7OH6jzm+5J2
tvmZa3zvysz4whtuxKk4LgmlQHFGFNd+oNm5a/EDsue6yz/kjAxZw7JxLHD7Qptt3igRozjNxmKg
SiR0VIhHBGKnItnhCVYfjHDikL917sbeg/sSJGbNRTD9oWdzNHOgsP2DzKzsEMF6HigsHEs5n1XB
z5HPED0MUnbuwENl1gPQCbKxBDIG8UQvguIqiVqDwcPG3omyupC/Snbn4CDUKPjz2wPK/s+yKxYr
ZDgctKAp8aYO5j/zG5aDErfm6k4GAJymN0yHOuvARh8WnEOPbyfOCG0TINxgb14GazJAWbRUq5Be
KoWJKy5QWfqLnHEb/oaNPUjkgSiuSoG4zHXdORnDI3e1wdFNR55i7sj+76KLZe5FTrurxkUfUj3a
Ppo8H/GCXCPvZcaJ4y2/ofMZwgAKp6QEhjVV/SNXNFmSUmxwfEpsWuI5vdKoFGEcxtNNZ0TzbddR
D8Bj2akmri1Ij2kBzmhhQJgjb+DZfcDSyGEW0VSaDnnWhYbnEcfLJ4zKFk7fekV8ZaA4CTACBfZZ
9DX4NMZaocEnkqL53URAPC1LdhdQFNFoJ8FXO0N5TZeFMiFOyVRIQmfz3/SMdNoz3J3oPNgeUB4O
YlYKqwP1B1q88ETxHApQqBuELU7V1FgcOnjavvV8EXK209KzWfcUzHOZltmwrM/OZ6xgAqiSFO8I
mf61CodMNeI9Za8ArhTVbHe58UEXrPCsbG1O2tSkiDb33FX+dTfk2DR5tiQ27CkJwZ7cABuOSs83
r2sbC2WWnrTpZtlk5oaCAkgU6WDTP+Fh4PywLdSnJJl0qXmQ0ZeCVV3L4irYXbXS7sK18QbKkOfq
4kfA+cA6ezjZw26M+rw7M+H2HDV0K836/zSvSqtj4Z/kt3Wom6RjTSQEwG2AO33V8qWFF6EZaRkI
lJwFwPP/S5Z/c1OgjRWrqWWMfRMHHgzNASY3mJGHEfdvd4dIgxjSQ5WeiIJd7PuE3M+rvY4AYNwm
Pth+pcofPK5mwS0LKj/lTVIE68xfHphqUV/ijgTYXwnbApgKN16AjmxKoYZe3R/XyQ3VDXh4rZo+
/gbXYRboQ5PGfxfWwzg9Z2yT3/puI5LXHOWM0V71ee/JUoFSmQAzu/P85SJdX6dzY4YwFKEfeRrG
FfuIHTih16WEBvK8/mJEYRU8fnC7AgQ6lE1dDWBHiC6THw7cISGcopMHYjDuhIGHQ6XQTMA8dSG8
lrTfzLxHCKDP9xKDjI3KOEhEw7FF9Q9AXbJEeNbCBSBwv2SQDfarASSiXhqXwsAviJU9FVSA/AT5
mmAEoJmxh4x/M9L9HSvlnk+L0bXV9SW5g7DbV7MO81gJouAdU2mWMxOb/8ihUWlaBp8T4RdCOsnB
D9UfeCsQ9HAo45xojiAePt/0AhklzgeQgj2Wkx0AIAPkhMTQF6QX8tlzwyDh2xKq02DsPbOaqyOe
kyrrVFhOgplJNuH3mtJ6islqLzQ7kQyDPlOs/lSHqPltsjAKv+sVmlXLCEwqRr2NG35ZQnXDOjcc
uN2NgnKE6LMEhkSFBJxH2hKvzNrfNy0JRllOhe7MS6GcoYMcO7fMLMCqKNNB5g6Lsau6os1Ufvkz
x6UKe/jIonZvxwhhdODjqdfDt4hZ+axNbQLDbxDEHEPBNc2C9F0qQqhTqbpMZdqzrTrKqH59MPqE
zTpsgqazU3KjANlJoSBrBJ5ZGyWUXh0/3d8ZwT4MFaSFaelX02wcS4kIL7+n+om+fOpbMYeP+h0T
lcD4YrTCNjmdw9AJ11E0lQujp499oRdjSQ0iSqSE65w0Go3JPnzYZb7pEMErtovbPJuLRFne/vcU
lXggWhT5QLvVmxMOz631SeEeS4dZEN+81yWX7cLeyusn6t4dP8XC0P+eFZeYvQdVtxyYOV4s1uPz
0SuZBwREYUGWGWOvBnV/A6vc6amq9+GXNcWiBtDu5bVYWvnI5h0sELO0nPxuWqaIsWBIoawS/jMb
0b7OkukPB9O0UpU17zjPVUfU/uzrVyzxDCv2p0p8juislk5L0dsAsAAVci74AM9rDe8XoJ1TcgLM
ApxamECJLJY+1ol49zhju+CNzRtawJ45U7OGdD7LdhHpuOAkQB3YZyv+uR6isPPirsGTE4mXNnrP
WtsB+mSmGhu/RUgamCfkqM+FgMhU7wdyIjwTpc5omkP+hhfG4Oax0YDQxzx2C4s2ssRv1KrPyrjJ
UsVwErJmIsywjW0mS+/+kmDYeoOKo22Z/peCVDc5+uXJtvRMzidemJUGrNXL//PvrqJFuk1iLyNu
2/ZQQXq9iGGWShCFlwzXIPQRRdkcY/TYZ2H6bmZODKPyjgDOFLzMkYFIJFChu//upjckVp25FR5q
8QylyjKafOUlymanFHszMVYuWOGtj5JeiBuFW/J31y4b8fnrJdhHW9QFJYQCiY4ZST7ILkuYw7hM
ZcHqdwBV1ld3nFAb3FwANipHQTqFewL9IanMGs7Kl1AubqrvM3bopO9wgIo5VkXPn1BerBj6C6/h
ZIZ8P/yXYwh1tHYXwXEDMUwen4lojYd9s4iJ3xzNIWvjeyHBwSKwKZDQUQhaNgUDsU/IhJk7sfq5
ReUJ2y/ovaBuix7t2lEJLjfAmkIMLxRBpn3YzWT5ujT00rzozIiZhmOBORgAvJB0msE9h5X0rZEg
jvG3UUphT7ZnycasTn9UQSXHCb6K1h98xVEc1T0G98J05KLjdpln9LDty6QDbj0VO/IbGpGa7hTb
46uRF6ZhF2srPjXYBDbKu0lgi8A8BxpTCK6thWinbyvczcvV70mMeBP2dVxsqszqdRjgpvQ/u9w9
eZSo1cvUSgIuc70+Gnywg/S8Y5CEidZoleefmGZlhf2ajJxf+JUwbAYq0nbJlaP+U+67PgrYY35C
gGl3it9EOJ0tQpXNu7CXf4R98GbyrwV4Wf4aOtbPupHsmbFg1iPNWNSr1Acph9bjuUDl2n1/tE+H
aD2D/s6lmifAQ8abuUtry2flLTT617o8Q77mB77svhtK3phHYCBKK8PkJxXGj4Ximook8lXusWhS
/eWqq4D2LmuYFZ9gUQJpjEzJSF6axLaUwfwKOr7bpxLUrE9dKVnTEkPDFKOWSysDpoY6I538puYn
8dmTOrKU4POIEUwTP97ANaMsvLyyc80otmctN9N2NXvSQyuXHBCN2e3gumjrLCr5RUZ7FffRBQVU
gNqrxH7Q1NFhzxns+DZxsjsjwPU31MLLQ7QEB1SpOgYzIIcyVL+8l0cbRy3E+3KCh8sHPhE8LfAg
CrYr+zoXZpGu+f0QEBeRbL7GR3WojhvKn3fd1MSt6uuOedq5GMmddzcWBnKkqlhfeWXKTQGebn2y
hgKr3Nrp0ewJqjiynJwduQimpMRhEN0bgxv6XMZMzuE2h1Uhg069N4M5g9yjcE4MJ65RgSVJJ2TD
CBkBbKMFJph+i0TlN4T/I1iJCickb5mIAFw2UHc6ZZHT/wM0a0rU83vBMeLdvLhPtFT+EUSVdRSf
aLbEC+NWk3bJcPvxcu0D1UO0AQsrldifzssjtKn7GG81tRpB1GH7xlI5asQ3zLN32chlkjpxVgq3
wokDp7boZA81GO2Ov613l7Mm6riWu5PDvAtTP3HOPGKBz+djpw/gMWMYiKcgdpMkTYRFBcqwpQL5
Ss79HGe9VtcnGIDORBVzKeNGzACx90cUZLxlJSzaqkoaPHLe5C6W40ziN/M4RzjkcVIpBq6SCwh1
kONm49HrYVhxPat13rZ6uVYLRQBpWF5HhxHrFLL+GncAXCF4uJp0cqaUZCNQ2rmFBspMs9UHzLWT
T1kMSPoDOpXj1NM2Nu6Yq9UEiETFVK54kZ8h1cimjIjwheuMrfiH2Ax34tuWMAG+cbuHBMuGTmKN
SRpZxuhGUJhCfwQQZHx1xWCluX+gs+d12m32TLgXwn+fvbSDwEZAaDCvGYsHGbqyRp+duW9dh86i
NKkckOvEP3kQ/YLV8vgfUggIV4Hpo/0HKTMaoe4c2mljJnrS6znAD0hd5cs0kGyi7diSqpixG0AU
lVt0u+DV4VTDT60m9V3DIDdhVABWPx/colI6pun1Tk+ncfrjNhoWwim1rgucu2n94tAn/Jsf2Q7R
NHnb4BqR2tH0QiA9psaf0yXpffgIHRCFKMJuJkanmPLtAAGjUjS2bDceocgrMtftt8KyCdibauWZ
SSgHAX0OsBsIGv2Y93Ttt9CMravirtQoqgT//l/AyvBc8RmJ5bCW3TpAtKmkiA5GJ+IfEEa70OyQ
UNxR7z2fWDshlRdF3o0Jb6BRqzGCh2dLEY/KY/IexwxX7FTjvDTiRuSjIlCO6LP+Ks4saI3AivmI
l+AJsQMCqCzifGjJVvz6A6wtZl4xBGvEMNBYcAloWHaSXfwnCcecLn52NHLm2H5t0L7G9u2FkH4k
3cFUdqDFQe3iRmzSS/VoForBmwQ71m+MtxtXqsXX7EqsQkcSO+ywbL0PdZCF45GKvf8ntws9kePj
S95WyW2M9MWGLk52vD11ZR8mu2pi1dQwoI8vYqqgj1Ts1FXa8TVGRxb5uomSVgsCGnmudcqmYERS
JJD7FXAkZBDvOMd0tDg2OfnetkLNoQO435KAx4wVNvJF9RuVpaq+5MhMpJudPZe9BrKWWCaKlDLm
bxWj0pwUs5LkcreAtRw2/BP9MISj4XDYtywSqKC1/808Qb0diAuyX7j/576zzee8PeWqyBrJYu9b
uCQb8YLLCZUx1r1XaR+cuBso0FzIII1I5I4ELWZeuvd+3OJp67jGlWiqES/ref0NmSTYp9B2Mh51
x5A7pxfP/U6kgbz9DjIMgRc+NkWTZBK8CLNqnOF1SPuUKxovKDKoDRID2Gp7AEuXX5hSzDzwERMR
f4HPcyPM3CMlUsvT6o/EzpXQPY/+fMLKNIm9IFyL85+JE4E/Kgu7ikRVnAZot4kfkTPUg3o1naS8
rtibT9ee7llVtMTw5qJRcC/Jre2Y+iZMWIw+U/7ubMf+u/DMzhNrMqoDrs7jfArUjYF1vo8oQ+5c
70Fk1JfEUvxmGjD6h12qBR6btNr/piIz2uncsA7zyZyOjr0irwJ2c8GIG83wkd0aCEY6F+QkUfG3
tyohns8p/QYamvEi92j+1OsokGtDFa+HrzeS7K55go6mO8rLRe1cvYraSp/bnrW/IlTxbCZq7ETb
VVMzCQX+m62K6OrMbQq+fzKPIyZilLjbGT8L2jzhuAISvRZ6HyiFYJgfiI6m4/I+0gx+NH/Rkqv5
vOvxSU2x5z0U8uwqe3jJ+ziDUYYjGySoZUdYtDk3DdIYrQ3EtDGdizYS4COp6CdTFoNULmsWYYzL
cUEzwI2p7eNQqGFLqvHpodvUOjdV6dDg5q9RXa/J1K9ouW7T7WIXeup00p1/YMfvYIuzEzAxq7pj
YGvuy0/euz3FiivOh6XSrerysTLqeYjH6+wjZt0rSt2NbfHf4gJ14QDABqt2M16s5XMz67ARstjS
kB57OPOsFPZZGj0+xo/Tw8ZOZP9IsrflRl5LjZEpIL3BcpzVK6c1gbsnlYq+HzgK9lSPp2oewfza
Y/Rkr+mAZ5Yj81+nJoLNFxuqfmIFzu113cYridOGfV6ZWnbUkFi7H0soWRSUBkkj+0eDsKXVaUjF
6om7UV4f8/Dkc7WRKdhRivqziAfzKrAGp9e9nXLDY9Ztze4fthpfFGy05AmIul36FZfIro9DMUa+
365oZEDEJKjbGs0gUSCO/0Hk4CFfYpJFYRE4JZzhVUK7DbUCmSx4LbuntkvEe87KsUKOegNVMrY6
wMJMKOjsg/XUxjUSuYKSEVkz/78x/LD6RBztrgFDm8yPPFEpFw9oEV2cDNlJ0wswUq0COgmxuDJP
3YDzjfFMNICzK+l6Wr/5JN3LHXPHdwHQruh27dPD8jMOcuyVRDNG/uoFXbI465OiPueFwioYl1Z6
WorKFgs1RfNW/9mRNka3MJzAHNZ17x2YVQ/0mPuKtzQ4bKt4pi8HMcifMmkjne2Gy49s+W/vC9oe
dqLyAf/XprZVbtdeCF0PxnXt3S8ig0F+B49h6/vHKxzinC17lQ5wmlr/+kNMSq+IQaCZ+NOrdGIO
POv4Ma/6bEa+J6tNauXEXu74m1zh6sHis7YIlAx9VoGRUqoNwtbpZyolskt8VLttIGqrfNDnq4DW
u4A67zEJmYnDno8oGRjhy5rV5FYt588mXwVqrc+1oGW3fyReiig4PqY/gxNEzEEF6TpFDelI2rWB
HQph+/tpoTfNpa300MtYZ17gNUA5S2Q2DhnFr2bquHzaX3T9cbXBpHpfrb/5phgdqHvHoztx/l5S
WUqRt8KvRCX+JvTekW+li2thLvu6o1k1S1mtPF+HFGLf5hJ/u9iWk1HVgKIiSKsQb+FNyJNmQ9LU
zTrp8vMbO6Yp7zGuEoY7MdfkcKMVbAp5oBe3XyI1mVzQrn8m/QN41MW4H2yaaC200gLkXKubT5tt
CzZ5K8cdJJSuLejjKDv+vvuVR50rGijcUKe075gKHyg21DAAYSRFjhGOlPGC+Z4JpP1pA3nGizRW
AHX2r92/T+Eafz4RYPnPwtoKzlkjgZUtDOUJvfyyfZZLd7sKyi8cmNjAiu2nNnmBnZNFBnd5/5yG
0yiY0NQXE0u37iXINDjWFV60CEnajNrxwIr4M+2Wv5C5mCbsgX/L6fp4+YZjnjEo8ZuUlhxxySnu
cRUtVfgXTJjuXSOn3XyM/SsM03aj5qyL9e4VM8VS3xdZ47JxyGE42jnYX80EsnQaChV+43U7wli5
IOZi3pJ8ykX9OdPUNuzJedw/AX0ngbXWWo2ji8TBj32r5fomPyV6woZeNa0nSUy9SDIjCLICE3h5
0cuKGYOPy54E4aXAIxWx10ZKiLzLZWLFFF2faMI2QHlPvidp6Dyk6AuJVNJH6hB6ZFSJ8L8+sPpa
YAMEd1y5i9V2qnX1va7PW0EIco7B8LURmRs8QAwnWfOSZCvvGH78ipalzQZwH/Ino26nZW7EI9x2
dTlK8HYbJbI7NrSSWBCLeNb8CFxtaPQCKIZ/2R2Swfgl73td7YrpdCc5YTI+LSFg5Yiv90vm3RuZ
Bbt25PXTLgm49M7oeyzZXgPFI0iAIsKCfan+q/qBFjtmUvMgaXOAdHpls0KUmKRtq1ZQnCnCSnqo
YI7FLOZQy+Er0HfyhWCYpKggJIZofQ5/uvvK9OlK9f0sfpWyqfdzl2S5zD9qhq5obyDINvgKyIys
PU3dgktmGeVgBm+hhpcNN43xKdlZ5eXlRIQSoE3NX7CejkpvPszewWJcDiB5BBVJwLk3Ift1YGH0
72ZbOzNhY8F8Up5NGK9huijcUlfVmPxllXmEEH8lgHFD+MuufjCKrgI0UxunPeKPnP4b9b6GvSKY
fwEigVKshwcHDcvNP2gZ8LMLCdfKzyhRNtFONZtwuxdZUG61rZbBo8G16akHjKCjyVLWKFQ5re36
lUCUbEA9xWItHxekdpSpWRIZZnpAgnAL80Rd7lN543quc97EQFdwpLlkCrZOTG6y6Xg1N78gevSq
r4Tojd0DNJgT0qS9KWtH3n4lrzRMeBuwKWQZrDHk7RjLAIFHbLVD0m/bM5KxFymlPPyl7hLvRIcL
ZBOB70P8CMgorfYShE5oZiejHIKrGo8DKuzQgH4ShoL8/kOpcY+4V+Ozk3wTjxkNVnd2F4kfhBMX
elD6BsyodEqMZXJSLoMmi8BDF8a7RESSHWJtQEHBvcs2SSX+5C2E9SLoVI+ycVS1RRc7iiJUhcB1
Gig9Y9hrjhUGPcqa5Lv92u9/HrHcojH6NyWpbQ7CLuwlGRM3TrxI6CI2nD/pNQWv7q8GLYFzuEh0
tEmfdxt18GOQrf1vdR3YmGAu/tMYsUCuvlwEdCwAZOtSp/96ddQlU5PdVxNc3Exo72x4h1zUvkei
Qe/yW2jrlxu5Lq1VReJgBde+LJ+MtqROk9uw4PdaqpLUR/DFDnfkn9Lwz4e+HEixK2HKnLlUnpp+
4yW0Tg/p8odaNwlscp25F3mPFryL5iMTGiDq5r1MmQSFboIW1DudRHYUJvsIJepypsT7evcBYDFk
CMLnvVhGLUnIXMo4l79SNh/tXiZt+U8BdrmpueHPNUcruCtyNKM4msFacLl2Gaxpt0W78VKomVWY
1UKt7VShsXNDPKjybNWa0o6mOssn4dZp1OUZdQPa+RINOthQ7fEIHXX8fJuwVBIiYfkVl/mODkeH
ISq7FPVgfldbNqlRvTtBulWNkRLaBOWk1Dzu9bYcPSURLTX9rYeGdIg6Uk8VjKP29oOyvpInOhAr
wtXfwvwmjDkR5rMfdmcYnBPyXlL/HLw5HEHSZNZHnA4RWh5R4hBo0YhYRDIptrV9RjqwzcAiQHzA
x0gZKqXpqMhdCbWliTZ7DF4fYJiZH6yDS+kIkRdH3NXhT8ko0dooiQ8QyBVoZeomKK4wDqAC2OEK
6w3QanZHaeJZPZl1ZLnazAfy6xURn6qg2G9cXNynJg9wclieZMg/53179OHWaBnzBy68cJuNhVEU
rCS3EQbvE54T1hy5I3oGdAoNlxcMPkqDyDR70p/MhPm+bHHkZl17J/P2IGjPQDUY2xhtE1MP393E
sIwsOIw4nf0YwpsWtUlJtiKau+sT2QOs73tVvo+pRjGRxvQiXPc0/MA/EB+0hOjdnKaaNuK8H688
vCTjXRLByQxbbtwAKiXqPykinl7NnwBUHQ1iHv8mok2YmJUgpjKzgQ1nHo8zVa0WC6wo3AXtXBi2
jDz4/+/tEg8Du3aNbuvkwUouARjz/Q8LVEFwFSVe5f/d4DSmSnOw0xcvIY6lCAHZieYEAr8PJZ4a
NusJwBclKjIfPr5y9qwrR/aFP9uRRui58dV1tk/575CG4nWT4A1g3bhh1pG16l6vZAng09cXTY9J
mQ8Qooezvx05vlQvN8r/MW8kEVb2f+G0aQFJsfkoORlENGtT82uYs363Mo7jyixYFgZzKDAR2wF5
8aweXSm8jfBevmo6RPaQ0gu74xKKTbEjJF/akK4onVjR/kcFfLN9ez6TnUv33bHbeabzHaF/KV2B
lhQl9sE0883lkR17eG2kIH6vzJhXPedpfRPpBUH6mr0VYI53cT9i3+taTmwuqgliyyWaLOFinX17
bjcHUMRY07/Ksi4x3MVv5jg4qEmjHrMMgB0VttVcqFoKh7U8kASoq3AGwlwuI7pZ5WYQyyrYrIsT
CY1U9BtxjsLhqAA+JyCLJ82Uf2lRRjgXrKdN0R1k05fDQtVcj+LaLHtsLXeIHZ8f2AhhBKuAuO9D
5MqNMVX+nyhZJ5ZoyQa5sWk2LtONEEkjs4wM8JSlkOmamhluqzwGZvX2rOFEHUXK5WRygaNdHpAc
UvKc+U4ei1QU6uLFBbo6Lq1rhFriCGPJtZE2y7Qqcouxx1A4duRX82Jyg7UTLEOrUfyVe6ZUbKa9
TFt6ZsOMGq4weWRv0udI2l5InSZxczKXIARQ2r0/dIjMsY8+Yimfba3CHs2Dcg1JAnASLUbFDutM
pkHpS7HbNpatyZNRzbiRHUBdBpynAS2k6qaZSgiOFkv7dJrv+HS4ZSElD491dZ05B4Akh3XU6FWl
dQIUdqJYFhYavahc4sN3DebZKYL9hgQ4xzlRsioicBayqUE+XqUwb7+yfjzrRyMU6TzaiuqI/LOz
dfagCkdOrEse//eH1T/ypZY6BUrCtKYc7X0wrCCekddB4EE6KXfJBOTmQ1hM50zd95h14vEeRLyN
H0PlCadoe8z+6+3F0AmaxB3aoBl4OIYauqVDGBupc+jd0LU7fFPO9Eih6NoBMVhDzJ4URLqY/+Ar
HE3m5XFSGX0lEGGstqaUPcyGxwnO6MTezEuDSB4uKO9TA254UqZiEtqEznKCts1LPDgFhENHqSfj
jPbwV62PWAClaTVziOD8koqxiuqs366aMehsZxMxelAVHR1Wym3il6hSr5g7rbXijt//GrnvsOX3
zT0U1M1oK4KjBPKnlnKxaI/egA1FlxHHv/+RFCNbFuzyh9Ql6vnyAjMku+RSCNmJG8jRjP8POmqE
BLtWiSLdfgSjyS/18+9NHzETmfPkZjSodGIYyYQ1zhLIQeIAXS+RtUtejUrO1P/iL5JEdbMKnLOO
Qy1AeObwk3gcjqjQwK7RnGKQqAphkGRGbHxpwVuKauT9VHEBNnzzOZErqBvXu71c4UApvTS7QC1X
0xMuACy0QZQ1Tiaugoxgg2+W9c/6HddoxNe43aMxXatDtXvTB4Sln23egP0lyWAI1B9LbZuej1zS
SEFfS8eyZLNOrCsbXsZGZglrk5WTDtT0YPR4pSVTUjbFtB5IWUJjCfoEihowY5wlFA79S4hFdHPD
bd+iRXTHYCIsG9U824T8CiPNZFX1KqAUoypEmFteYhYPXrwtDWkDMnRu2rOkXtIWezBSvtMicQDa
YXWbdZEZtewP18koNEB9t+uAcRy6Pl8arAbMG7gJl21wk2aHHJ/iBZEJeYOnMdo/H6SDP1d1T8NG
BuX9dnz4NsJmtaoOzv1qpHZ43AuaAuSXLSbO1GTNvB0JfX1CLVUf3W/OArdo57dqRsvcv7jbxiWR
3pTrMSi/raI0bYQ2iiGMxpUxSoUDEchRZWUyzmgAzxQUR9fd3AsIRN9UKKb8xPUmcGwo4JHqIZ5E
2+kfJInwOyqlRmwX7I2qFZGVmRErFNA6y9/f/yXcxEIeGf3JkkJfhfDhcgszhXk4JvaJ9lJFyPmE
fvdV5/uhS9q8hNfLPKb9fD+CEjwJfgNJRnB85dbfSoKOEiSGqI6CvSlIgj5z1nEWZLkUOUN3In42
mNn4gnbPt/x7cdRoPR4b7v+z2VMwITVMhC7C6g9oT27SSO1iDqDDOEnlQduZp9NIJq6irJ9coCI2
FhJigJyHJzClJW/OQGwR5RLuQJuElcWgVUhyMwSRPxYh6nQe5cIjRVC4cD4zvqe3mrHYqREd5znu
3OeK3kpeQvMkl6iV8HextMTt318dtgOqFtUR3+6oOju8FQV8S6/rZw5DG1BHtPxdDirbHjC+PiDj
7oKF8XKtIZjR1xeLGo1lmOZPlA9T6ZM75Ol5MSU5ODR2LiMxFa0KnrG3wrnaJA3vdcRJMcjPlEqq
8mzudtJlyk/LSItPx8tDvvF7NERfqRUQm8GKBlnMPBuslkjVtmPg3dBgLLrNIAFzPLveHKNinF+o
F1YZvzRMUppv/DzM27S1QhAEAz8YcVPQENKEBc2VnGgjQThyqUT9nZskhztNwKKIQ+SP71+WRERa
I0JXmNy23qyUSGFQ/ktX7x/+FZbCPDMc1jp1GZPxzxK2vleUyWF2oAfqwpltQgmuwHK4veRaHkAs
Qefda0QvYebe1Z/K7ExjtO+PP/OpVPU/FXbuXzMc9y7rmvMfq7w+hx/gBBKtDzliZ99sAh8ckTKf
nIyfLe2sk3Dq3BvepNuJaFuuheJtoEha90RgumJz9T/BYcxw1+u/BdlKZtBYkBF0qutdInhBSIda
CnhKn8DXwBTKJurDfKZcPd8W71esfrsgybPNlUJvo8dPwOav0pgJEDedz/geuzNMLK8pXVKmM0Xv
vPLzptoQaC7O91EE10iZK6KOijXQ00ek3ZexE72B/0ZlXEhhLIyWJ9pfs4VVoyajzbv8RD4Dy50V
S7NH6MRUwU4VwnpK0+vRwcgpURTxCUvPLGaxHPD4J4vmKd6tgzyBdRhnbWtmuwHNdmJFm9pJoF06
Ztr8bW9YaipGVG3HuZRGb6lzx4Gj0zTqPidRgzpJl4IJqXPR5sA/W1YXzHoUEkDOFJdcETEfsjzQ
M+GfK+CfFE06taHebIJz112yoQCo0GJK0LTz2ZVC1asx9LbqyunlDzBuy5vB8d6iyEaCjHYyfQ1p
a3hh0IOuRH8qHaGQ2Icwe9B7i0Uqtur5Ugfza6mdGNwHGqlsH67pwc4SoFEvkLh8B9TyUz8chTf9
LyBFEDa/PIJ950eOYIFDGEOPmhHyfb06p910UBCtk3BOMR7Xrsqbz6hlZtgEXBk9cOhs0sHnmoJf
cgNO0IN2eR20kug17BfLPVvjX89ZcsjUH1BSpwH1Zz6l+FFJm/Qn1b1GhDEZH4u+0g7LjHWtu53/
HdBYEDFsDq5a0wsGu2TJ0JJefNq5/WfbFr/KtZJM0oXN7g54A6lIzTdt+jQO491ma0PGh4UEFYXe
wcLCC1CAU+zasPltHmguscGOVw+CTGOb56z53WMZp9sdSMLyKbFIwjmG12x7Y6zR/2WArsCHAJTI
Wx3WSKfvN+xGvLcNk0Sxbuc2p2T3lBU+9EAux/26UTCRGMLgELNAueNBE1/wB1JGdfI4N/ZVDxX8
pH/0k/OfJ17KvUivt05yBxLxg4aZAzGGyk3OgKxss9UJXlY6jcAr9trZVeuDYvbIJSvgbr0UUgap
s1aBXbmrvPR1rUQpMuendomWgRBV9H87604y9/ZkRshtztCbWoZAWSu/KLVtZgG4fVBaID7JqGo/
uhnrL8S8c8AJtzay0fbSw3rmY9sx2pdmfeVC/EYtB+TAyVdLzu1WAsqmJsuNzej8QMP14Tbneyfw
0YRq8paQx9+SLZdo1Vgl6ZuAjEIivtKqyZ+t2w2waPWPVML/QFpxTld9iYqm/rQgPlQGpv423y5R
px8exE3VdSKZVKocYe+ZX4DhocVCfM1JoAC7o3IFFk9JEp7rPgZebH7CAkUGbt3s8Uw2TSZIkbVF
FyXRIF0WW2b3i5AG1Um4YC1KbJW93kl/ia65HyNy3RcjSmJ1C/shTNu3FpSHJLWeY2g3vDYliSoc
X499fA+D3NSS95a0RdlsiudguJ9/7+3ruQ00fhejTH9ay/1gAp1rTzU0GIJ27cq700dHzjuOBNiM
bZHRg8Q+UuXv+B+VZfaQx+M5XNXwn9tWDSsYWdAomH0RPhL7SVm1FsfQqZn7Ev2fIzsbDct6Swi8
WJ7/JdzaqTwiw4xn942RjYSwNtKLfLvaNett4t3K718FwiAjh7Zc//jLg4bRmbkIk/flMg5+Lm1Z
qQ0OGmLUxqSIiNa+cIAng2iN55pr2D+QZ9on8ypT/iMQpshlUYQOXcqV4AZdSJ85SwtSKqyZZE6q
hF27yvuLqgX2KcXv/WFHuvkbrTV1pgJLBfHCyla1rLJYwcbHxWvB46kf2gxIxPe3U79S6Lcp6Lm7
CcgtD0KATpySyBmFKw7zAeQqbwDI1MLXgtkXRlQtxNN/6ZFRhER7o0pPzvQXX5Nls8kGmnKpvGXG
gVj075/PJwl/2Pj09mndnCA/vYfKsHCvx6uaJNo8gZ/iM9bR98YD1KRMdkH7l+taJMW+IYwqw3GY
4gwtJzxfVAs0KsTFXYHhZUNDzBqvpNWZJAD6kv9o0A3LTDAYBfKTNL1ydO0wZCefIePrApB22iJG
+xvAu9F4aaivImhgj2Um4LxVshr7/pmGsL42oZFWaARtfI2ihBgFbqT5+6utHTOkMXDNIhfp4MLP
NI/nTYu0pIr6h2gED/YsCujJHIi8HYzMkYafUxNvpZjNW2hqna8AlH4uYyirgNcRhg0yalGhoNjh
X79a9F02Pm9kWf0c++qZtPTRftqd3rt6ZG9E90GUXwcJNTiuKafBL+yyG5NmDWVyGXSDKOeevx1H
38Eyz/i54eDHLdDPm3cJfA7XC7FpHmRl9uj2+RRVtjiYXiXqjGbp1qg3zy+va8o586af+c5lPd98
DWQeZLcNv4tsuz0PYIfIDweegCAzfsR0ZIRiiVuIs0/Vyf4kW2DHiLp6Nz5E+u1uZ3JjRIX7QV35
O8bLeKwCvROH4PuIBW7miYSLCSU2E1RTlHCMuP+SLHodkx/flhRCb+M12MdQxra2uFlyyda2qjCu
JjISJWJP/PDsPMK5sZVouB/LoNANf4jZVeCF9bFGKynGI6EUEYURxH7x1jHSidBXa09bnhMjWZ6v
5khRyqyeK6sFHAbY6Cvct8pSRrPZ86vvXEKjLyMQjtW6RlszBLsF1VaKSK010BXSSBfR4rSOAkiv
4zFbxVqZjzXyVyi7Vh1yhQurO/0D8/WZ0akvIExrCzVRfno3lsSwOGy9o5a/qzrRO4hqzWU24ngr
AizESFkPMRJv083bgl37r1SpRvJtkEJJFCmsdgRZnewi8s+e2jiUZXajMA/jYUn+EsNsDywqi3OD
dxGWacTBVlzW0w0XS3h+Xwv/8DgkKhpynIen3dzmDJCb2XFM+ldHidTXJFq36nlpyYaEPJgY82sD
lOv/XKMjVyJvHhabBin/f9hN8R7DF3DtJIOCWKEvC3JTwScSZNyNpwuew9eZHKufEEyhshoLgcaw
NGsMFRVCejzxvJgbsQQhtOxFpb2mRlJA0Dr67GBigvA7PffEYIwisjGVyXFLq5uJw/X3Yk3fNCfC
9XrFrtPeSFzsSGmbqQXI5AHKAsH/arunUsoKi8fjp6PVrQ11omdkBk1/ne6Rg1EF2QgIBEHSGtyR
tiHjZIBEuRv3K3xml3ib3pdSIhxWjVLpypOzZ6Lcdk75zpe26qzOvLxB+B6HdwF0nmmSaJlS1r57
1Vkq1XhWJp/3BUXMbsRmGmHOZBP5pSAfPoDnsgFhHkfaKMKIPQmMzHEBpDaHGJtgwXVNABsWhGdn
XF+JxTxjdy1JVr2l7lBi7bmRIC6ndYfLq9xNVJfTDAwmU7Ht+oAH/oHF8h8gI5DI/Xvk/HxqnErC
NyFunWZY8nTTl5rvf3QNNuBW9R6Y7v44Rz1PJ9/B/sTXnSQn5sqlNe2cIqVzZdCkdm+MJFm1g9Td
idHWSOcIv1m6dyjDWPt0Uu6s3HhEZfR08k2aLCCwEh4IzIyqlboOqQdxoBoqZ/XaL+VTnZQP94Az
hcbCF9ddNIOqxp5UnxgMLL9uiWOSY3SRr90vidXkmn0YGCU59UzsxPjJ3k91jjzib2ljhd/M0zA5
5YVU9CEllUqTncn1hHEsghQ0osERDLWLkCWZlV3R3NP6oDrJysBCHZAjf0b9RYoK+H/Q0Ds9TFmJ
pB7LE9jh6LTdY/QyEFL90azl2cSDn4v3hBeLFLjaqxnADAUt8mAjE/pfpoOQemReYs8htQSKKq6E
MRFYBdZNbrFQ6A6rGywEfbj8WukTuEYbFW+x8VwlZYbWEEbvl0RKoBipTr41rx6dkPgAUp3P4s0A
vk7d3nN56b2OsfRi3O+GgUd8wYuRNu4YhuVbLA0rtZ30omvUkS51YtQHNJBFWSP2EFvQ1wgqawkF
0TEaYqvKNjkZbhauNM5zo4L7lVERs8nYKDVf3HVTBWW5BeR4unhz2yKnsIVIr6+gN8w6098vSYfp
I1AYzLG+J+PL9IUbdzObE0t1Hy96V2CqxCf5tKYtw1E7iAxSZe5fxagSkYu3JU01w+X+ShWqQhNm
lz7hM03hE+tdIOa5991mRkYtxTXPyvsGmK9SMN/JNXTawF98UxAzxtm1c1RVFih7VeeDHDTEcLZr
bVrht2jGZjbvOLCwIIs113ClF4Y7BLGfPH6dVpxzrH/32JzTqSWpNzJLSHbsa7h5+J+qzPlpDoja
985GuE7W7MuFl0qLLGHNf2tekPiSsFvdzvBoGYWOmlCBL1+iWeJOgZ5Ry720G2O3JcBE+a2SZ2Oj
jGpDK4WIAWqp1AwUZ1GZJ8J4aYWohFV9fFuh95fiZ87ZumqbLPmm2sts56rD2eCwDa0H3zzOXA7M
KCxALZ0jmUs7uNVfMO5OIc5dVePK0PWks2scsJ5EZ4P363h6uAkFdHJJeq0s/Jl3CKZRNeifuc8X
mtJ7d8J/BavakJBmFMEOUFqkM4TW2DDTXuSa6yHZ9Mtp2UmvjCXC7TOVN2E8nGYoVr90Ku2KqaAQ
c4FV66ZXqi8T/yYp4itennfCV9jcj7DzW1rvhSqaY1gVhnV9x7wQPBNa7QxQQyFb4cmY9yyXDCGh
ybEvk0Yud5rYKuiu1n73VUI5q1+EKaFUoUkcxwReh9t5kZmqrt1PSL1f8TmTXmSuT9DTaL3eVIUH
6c+qRFUPEx1YOuxCAzMiguDp5PBsrnrvXYj31R4JLuYSdHgdFXFpV8SNXXXH44KSDFgwHSyA8gR7
TADdGE29Gh4tRjiesK2Fykc2DugvrhyttT61aSmSqOvVp8wpP8zw+E+VfCWlsGKOW1u4DwfKL6mg
nhvNXOlgoVeHxBjGxOCCICXDgrtr3zkT8ghtJlRi/6eDlefp6G4IFoV+xkTmtsyKv/C8GCbwvF5I
imrrsx02/kMqtZrb721KjydQhpkjPiT+ns2zxznsRPp2ACLc5/Z+sublU0vP+Zp3bvZaB2tMNf3b
SQK3L0EIDw0Tv/H2txZ3luyETybQSgZoUpG9lSh/P7/1KaqsGaxC+v+gL9jqyx5VI9HbXsCL38Yk
33PAmC4/3KSmSbXJhL0Va7PBurpTYk9aSoN8flZy6QOX3799rvH4de9slIuF+lMXwe07ke8EQ4kX
mJI1bFI7pbBI8dG23zrLMSWUUvnO9To2qVCUgqzo79yKOzRs3IY+cAPDfRDsgA2kkIKyauIIf/rY
8cqNPQetGDbghy62fA+da2F0K6b7YqVP57BI099bVr2M2RPAVUrfcdS5HYJEURX46PV+XDrlxpEl
D9mq/fz9inYduDCXTAfMzueGxRt2lDKxmZQa4QfERM6hzHP4HABfFncDSPDpI5+Y0RmTRXvfUnHC
Akn+YEeaiYebDV5sdRvQY14pdbKwvEwgkMAauFr17xDBtrgnhYp0kILO16wCzvr4T5XwOY9eUtxr
PIStQegfCQNVXmbh7xyHek7maL05Omn/Tn2eZWJVplxYQsHA3bOMCHAbyRVQd6st5eHfEoT5/fzr
M5AqLjOHoh07/DxVbGkkaKKuC7r15eP/c52fW+WNLFsnx3TSS+Tu5A6Zllk4RVoHtKi2uXc2sJZT
LpKn3uxTeMR/abhD+0CRaWh2ffCHlyqVA1mSouvaW3d/JRXEF+Yi26p1u1ES8KhUZy0afkC07kqb
XeAj2UT4faNphKLIx63BvOVa37G6MaBHR5VMY8MxAWFRLzQlwXtWFkqNr//lyn7Pq4g1axqmlHAD
Nk41BzNINloLG408nqL8b3bDGNV3QHy1Sng8VFJvHNAWTXTHIwewokln3GjMpFuQ4j7zGsbrcFIr
Qzh/TIsUpeZKq9Kdu5aphXnZ2g81ly8wzrY7MjrYdd1gYVPu/bxI7WaBDWb+W0ho7Q4HHUs9R1AF
1lm8je330TLd3GhhWfiZojUKdiCuHKLEI5h8jMOUitOI+uLjyiLHzMcEu5M2uNqD6Ha4ZdRi5iI4
76WL7gZ9YxlttrYDCZUNMBfwWY9Su4kouuG+W9ppJSiwisJtc+BSHr8c7fqFqpY7nGgN6/kjIIpj
bWbzkUv4IvZdM73IfvwC5D92hWMHxdJTnGk7pb5+idgNJAOAkuTZbZ/h3GjjcAFlwKoAIQKvkSIg
L42eczJ2qPWnYPwE4ya3HJhvW+RMHgwBSxWTDVSTeCuQNItCqhA/sGkKB38/n3Qk/+hQJcl2bjAZ
YpkLkVfAZWsfkKGYQcHxuvw39iVExwC/uBca7mt8oySEK18GVrLQiKkBg/kljcoY4sbvtZUdBb9V
daWIEbdNA/LheD7Hx86yci/PzaqU6HrF9LK2w8rqzxnmJCgt01WYqYG4qfi10Yof5pvZJrgFeIjj
JK98WeB2EndxQ/+rvkJn9qFAABkMgAC+uTET8lsM7PaR9xXnmAHU5QjtdDLjCPHzqyC34B4DgmV4
FIOvyrXLawLPfNtjhcnuzydvhH+Mme0iTKtH5vPjlBtarUp4rZ8crHals5+vGqPrRbxPQr15cLRp
ON3E9Ot8sJNCSjsdLv5nVbQSVon1K+rD0i5fLQXh/7Yt2vmFnPGrIXUZz+SMbL4ckXH/4wqKSS97
0IoC0YEDlQsJzeV2W3ZUzMxyf7SSUDYj5D6kEqByJd4XT/njlV1TbxEI5GM6xQucgIcF7omeg77k
Ie4XMsnKJ34LmgrCaKtpU5Yc1wfDS+igHJxP5Q+KMArFwqmOwnoSa+tehfP9IG5yBg+I9FpRVPHN
lTMyjFQZZPc8NacLepw0xT1e9rCHphmOLwiLy1eukdWRH/YWsB8bsQQDZq4uFkn+lEuAW+IpDEdU
J1xtNQzs9jtqQYEGZSu+f+svMiOtQ97I/GmGiABw8TZYbS1Gl7f+VQMmruyoPqy36ovNfROIp6IJ
PFR+jlwERD1PqgSrTvNjR2WN58NPUvSmy7UksnDjKL3WAsFlat/HoJSDiTZ/IXywdTjoDUTD2gdG
Oht6Ekb+rK4UtNR25dNOiZPP0BFfh482GFjRwFVqc5AfXQex9/JnnerpO/xpc6kjI7Tsc791OvnD
DTJ/JmwthnkbUcs3+NSH+LP7DP1BtunB0Fulgsya4I4AA2dzRS5Ii7pXatyqfd3IATogDAMy/lhW
QTesJKlZ9tRs7csakZxIDCW9qfFrr6NlQLTXsYWsAc1z5dhFVbz82yPdKM2jMBFstV1/mrycOa54
JmQf8t0ifTCduSxBFrAJaZqHsby1M3W6wMTNGPcmefnDwt2vQr/oielSa1SPJj+oKnuzCiTow478
UmGVBU32L5M3ArZ21/cE+XPYeQxRZ6QzIGVX/efSQ/wT1GxCjq7FTbURiBTxKtllKQij1bpBDSXP
hx9W9afZvPR+KJVQPNC+zlIgFwOvLr6fL34apzjUxoa4/Tubj6kXzL90My/MC+jwZ1tR+Kcor7D2
TKYrEK7v3tugHeJgEqvjJxUxfFdNOUt9hGgvTY+88mA2yWlgOUITcKOnGo/PN1dKbViK6bS+SKkD
eXI14S3AsdokS6v+TBR3H7irtcmFbarwlwbhRe30U5kXQvCNnxpcKT/+cITLYuO7IyYn0szsUb0s
yl113Qjx42+rmKSNEv/zvvhBgVOn/XDzgKhilvDxi8sw9XLahCWf6FuSA6hilOWI9+Z5FIvjxtRl
z7TXC0/4YCKzpg12YIFADUMSGlgSAu+vy+39IY3NgQtpZtZQnRlXoBA7VRlKyYRL5PCUbCA3E0Hf
8tx0oxRA8um5IBz4H4QUdUmAH2kQGW3wjcFhzwN0L7HnErDfO3rxwjcm58HR8+Ge55CFdBDup/xU
BqBglwYF99/MetDf07hQ2gmrfZj5ec0M2KqA8f35ggZH3WNJmR2TpqveaS8FJd5oOmo1UuPaRNq7
FmLXxJYXBZcyv8Fheh9IQfs7gRuSRsxa8CbwR6iWQUF4WbdsrFDPPLXKCe8EcCMz2KQWXB8reOAg
ZqGlO0JwaNtBh1CE7OEjf1839TzXNjDqEnWi1JD6LLFZMV1oTbNw0VTZEhxYk+mzg6dmaiV6YMFH
6Vzi47jGtJkIweBpzvyAaZ4b4ABVLd5yI/CGYAMcM+vt7TyLCGS4YhJQsSaWUDNg1uZ5EWnjly5c
fb7RkDGOYuGT3qj5rR//exLhSrWh9mNYzMXxPQFskKQ5nHcrwz2tdaLVnoQpzXSXvg/AFdjG3Kkp
tG7EKh3vxzDoxmzg8ZYtZGP64de8hoaCndJduKFgpQ/PRcglI3L0PdSCRztCzMymsBXRKq8Hgx/H
TJKq7qDwpeqrdTtN2/2H/DiWFnkqH0arSrt4E7brR5dOfoiul+EfkJ5HJnF8MSeGeaMYqTVS0Fpf
m80oaZ3GLulCZsE0/g0xifjhR3bbS5RnlsOc+bSKOrArHG5Yx5Tlbw8PbEp/OTfToiltBJdLzL4J
3rouh3Np5To2MgyksEreLXvhC83MTjrz5qVc/qEWUVLYkm2udSKrCxy683mh23LKDZFQfYNkzslO
ZASnmUzk+uKWhTuX3iAHKuZxr8US+l27Chime7cjduf7IU4BC7lH2bZdKBqxt086I23b4dt8/hTo
vWfl6D40go43tG+HKdRXvyntp7RX0sJ4Y0wN1fQF2X7BdZECRklbamUge52ILB15UpnUWFIBgZRo
qf0668KruefCSyJJ5d70W5HbncFneztGhb/Hh3Y0UQ3pX4CJ3PJ+sdq1Uajd/aY6m2XH6dBGb0dj
jhGQtMO2Ha2vbglg37diHzivCROId6+9ESTbdam/d29JmFZBwWWycfg2Hl4SI6qRg9wSGCS2JCr6
lGMGrxS7wR36kRVSw3Xha1oWyEnvJV/EK9yBXtHo/QNg/TcWCIx+CjHC+ZbzYewu8KosKyQN60p8
5+Gx59TlNkn8FctM0xOHoJYUUQN3KQBd9sV3VccUFK5Apt2Uei6UGsGX/NQovRWQZPITuWfn+CCC
1XiHp8qY3YuR5LbOL109lAuZyIPuwET6G6vKUSlQIgM7z+r8Sa4skYYPtMAJj6UNUFHbPYWNWJ7n
Gryg9CrQlnHzfZARCl+aHGmsrmwh8rKVVdwbbmv4lJI311pAc7tXLVGIvjO++IWz3gO6oVZqzS+6
10Bd7jarJLxM2NPzkEKF0vafcLX+0/ruP1ASWZmrJe2SKDBYKMc8lsEqvFZo8REdPpHibcG0BwkV
7CyWsHq+m/787PDSSFaGaqoCE9WYpi0i6Xk+zhh8dEcnbv9kqsU6vE8SbQgbU/hAHDiSmQCQaAWA
tjj24yF5smdwngCDuLRbGQFEna/gvuf5PFlT93HoACK7WoWnqcyMMY0YD6YeIfRSvmTU6vWokGKk
E86vTpXAaj4Qom7ZdT0i+R0BYHPMgnBM5/6cxXHFGTZEjTMrc/swc+QsrtwbzVTBCVdKYRNlMG2d
X9MnXDkAx6eTfRG+Ku4w0BJtVKbwmlzbCP6VaAnbt+Hayt2+P+bNRKGfg8yGQTD6dhKI8FmTCfpB
5tAErAy8TQbg2Yo48N5Pc6Y2QhvLt6RiyY7sPRN+IBOb4CdC/C0bhlE5ZG/3Lwbo5iZZUZ2pDW0d
ZoklwxxiJgeVqZv0Y+zvlryfv89980cDwJd7sY8wNga/NXZ39I3wP4YOOx15bXXB4hUI4xbQIV3L
Eky2qDly795b6Ccl6S3TIVgAxJGmAhQIBoCmGpVajdTO8jFNCD76xPEeChvL1RcQeKmK5PT1Kxq+
lhcoZwP4POAgUQXxi0rlHPa4d0pLQi8T7PjaznUKC5iqL6Yo/CMVMr2PY3UGth/HiSsWSFN5GT90
C+sPWU9JN1ifCS3CXIBB++p1lueuBfy2AxTZklpvciI80dhyvBfxnCiMS5u0DjUEhRC6TcxLgd+2
qEyqiDeB7oeVTBZ1vhHxpz6a4CkLuqQvb2OiCNnEpll4UuSPqjgajs+9hLdSOYSXRV4N2A8zEjKt
Ll36/iL6dhWWLIEpqUzxOtrb3uof4q+2scUI+wNrINH9B2b404zmz2li8VB2V3G50XGUC38b4NLg
yAACx5e6eCE4Zt5Rcbv8NhS1n4eGflTLHb3kNOfOYPKAf3RL3kF/8PDe2dsfRkOgu11KQe8rJfcu
5Xbiw23sffU7KJR0U6Ipj2n9boElCkVVBoZT9A6QX8nyAAnG5oZNOaGGk9zCSWvyNvPAGzsngxeI
sWAMpSVc+m1XtjGrQ9+CR5rx+ujL+5CY4m0nuXQnEwiLVeMJ+qA6JysUVEjDMQnD9X4aSL3ipKaC
vcArg7KhVQ8jscVtXJX652wcPnhwNfOq+JjipYOD3ZjIOZWtkZ/kx/TksvlWkZbsP49ZejdgrAry
60vo70XWTCZztLXO/QHprgMPQt1GmojmippLQd80DEh6Q7VPGbh78qS3noqSUXh/DGJ/PF+myDrT
PwnmU9oSJD1sWrFttVuHjrDHHCU+tPyM2TYBrAqzpBCTacsHwJfON/trFRNHWMEAVyw0e7BUXpqE
zzBQKbeUKPSB+iUUAev/SaalG9XuFQCg4msaTVCkdr/iZvlgMfCwaeb0oBFbwoUrJXZ2niHmcq3o
i+vxcFEiuMv9GZdCgcNQqlOnXf2AHcpbMm2uzuYddMuHGA+DLhbJ8EIfPAdjwgEgZRXxjKmyMuPT
dzYcjGkl+wD3NBvE6D4FW58eVCUAKFoVlBDSTWPDaTQqHyAH97JDILZTYgoIz258pNEQoVlDKoxr
gD9x+89zXMVaGyhkdwwY9u61J5VS8kKfIUbXRdE1e0+RwyonDaoDdQJI2d0zBBOHu6lm7JWvMSJ+
HpqbuGpkk9yoALQ+SCbI4MGZm62Dgp0pem6BMcI5v3H7X2jtUb9RnxZaE0pxlRRWmgfHAeFPxoSE
OHnkmoGA3Um+3gwaevKBO70lshDqr5ROzOqBX7aRqjpibKmCXUxi0yhclNKXkUZrCJp93mQDYPKt
CeoaPMLHXlOKvu8AezNhUtosCoe4s/WRf/kKDrINlAXv8r3aCU1lXcc+XuJIPBjo/PvOfVMs+Elw
7EDof1h3MgYVMmsMmq9PHcap8wHjxThU7IuALXe1Q7u0TO0RE8x3NHeaBHwPpQ6X6Nu31yQfe8Xz
aO7KJ+3CwqaPLRjY8A0jFmqtsCQCfNYFmi/ZzDMt1Z+E+tkKgOGoxu1zOWzi6hDf3xJHcOLS9CvG
5qG/aD7DBgRBW0R8YtSh/G86mAUZZYBH8IFeuVyF1W+1bNFPi0JKw6O16F3fJbcfVTPmPuPc1+BO
1cdwUHkSr/RBCvOxsn1L01FwJkTUVr7z5Cj6jmu3rLfYzPOz8do+BZrmvfLEEXR0C2ttozQnLrKn
1GkzOpDztaDfOYHpgMOzG/P8cOhilQxyt1yc1KuGr/7qfphyrLiFIYPX9GkICePSWHH5pt71kEDL
x1EUP0CU6KZLeGtCSQ7AnXABU9ddvV05i7jI63QqdxSglPhPbzc1hoLlRcZhRfjrzc6Swmv/ZkL6
FCDpHB3kT58OAs/e/VGkvporqlU0jaOmo2bX1csC0B+Z2uAzMGJkIdQtWNLMECJ4cUlsoLPmoV5i
rZEVY56wwcP3VGkWvcLQvIDsiRguFOyBMlXErfdu+wlbtMrVzWPJCUsrwJnRonzcX3nmb7vuxOw+
iJxrIDyS/oL/mmQ3T1vaN2Xru6GJrOyIyDJIMNNR+sQdt+Urx7zsQa7u0KicHk+PdGP61KV2OGPk
WLY5U+p00zn0wtORLiSwmIBlKEbOAYuTG3a+jswvi1u5N2CwgJG5S3DNGt6MYYAuPDbu1XZ1AxBm
+Ud8wWQ6xWPWAFVLlWYM8Dj4Zqc/VPr5QCYWo4pxabiefwzWGGyCgVTL3edRLAQu3EcflpzIh822
efj0i2ERpawXCbGj1qWHu33QeR55WBqP6wqB03Wx8ftPUevSWKIgIORaIlwPqZpCFoek+QdI8kh3
kVA7mv5WVLploJaIzODHsMpUc96T8MAPBYoYo9SHXR0NYsbgrGlVd6w9C5GCLoXTg74H4nHic2C0
h/c9ZMUyd1VBdUt1nF06HXi772NBWplp46QtVpFJblTd9mxaAfvOgo/t7dAyphjo5wM2PtSvNBl5
YcQXeUg2dat1wzg8DOEEh0mEpeCWewbgVzjJqdCbQElmcFB3p+TaF4jN15CI+Vifm998IBQmbqBr
viE/quRSdpTsbk5h5Z/ReryRlZqxMpaVVuOx7qIQ8TGQ0aJfhqPsy0gDTN3fXHe7IFUTeysd1VDj
QbqmsHZUrOvJDvRNQdLaz563tfiGg4P8YKPTAJF2WNiqEA2ZI0JGufs1Qhzrx8ArkiWy/YfF+ATx
lHhud6BlstcfggxEgFhu9C/dGxPdO+cWzvPQasouT15v0xx13YlltkxIrCgbRN0Shhmo+26CHvkj
YVw8Dj1YUUXrMn0MJetmtUtemTYj221baP9NTp0pmhxaYmmEVpmQjfmhIR9wn1oLZKtp+YOa4H6i
GWPc5FbHOl82zAN5e0oy5nCInc7noIX4ztYSOB+cl54EpBA8xpJSYLVfwkUh0SQqjLgXw2jMLAD+
I/1agvjP6T9CVh7HQWCMyKz48ZzpYj5Pg4WavS9Vx48fjb1uhahWY5FdVqnGIAaI0yIWEKlzsR4L
cAbqYsA/KrJy5mKMHjWzXTPXFWDlUHjReDN46mK4wFi7LH00Dp2GqMNhfoFcZp8h4o2afZy6XGD+
B6ift7VMX/7bVMR/wzAmtn3xqapZ1iHXX+kAg+lxZ12xCT0W1xeYxrHpofmNjDIWk9UmSOl7hajr
YBxQFk9p8EVR6BLeSWyrqKv/DT9dd6/GXfUtxM1ht1IrkziFx2gFwn5IyufblEnVdmUFBCM47Gd1
fI/gj3cc2WLtCvglO+T2ie5VzHUfca86824M4BD7r/DmwqJJ0EeZJZn0K70qqBF9wD4kepzk6lCN
VVYjv3TNXJ+5qJZ5l6S0Oj0ksiYAoEo8x5ufFUnsakZsaak1MesQKMxqrugMbgMPSKmjE9umnUi9
d4lp5ta8970jUpZ8M4x63MUIhCd7Wo57cBm3HUkmdyMnH4XDxxkScoNVW4uASLn1OlsDZRYffSvh
Q6mU4uX2gJGs531NqOuu3gXd3f0wBF6E0k9+I3UY29CdVLG5lGRhDUFV+Bt3MYQ/h+babi4oc7hc
gxTRABgiRubf/5X22YFhTyg/+iu49lttKPB2aD8DCNmNZUkqSbk2FQ81mI/CSBdnReM96X9QqD+Z
xYOSdTVZfcoMVRaKb63SmjxTcRCQlQmAK2vr87GhUjiLZs6+vBNxd5QYye0QmgSbCzWr90eINU5Z
HtdJdBQ0PS3z/t8THOecx2I1cIOu1r/F4Kkb+GDlzftWl7wRA8qCzb1rnGnTxAgDyAlL1YVgoUsb
LZBwZiiiCeaKnoAGXZjhJEhNtxTQmacejZUXVtAeuZbWJFSrYaMmYgXoqD1rH1LOL596iPYeVVCH
roTMEbiWYiCmvD/zLmyo96jx/LZXd7zOfI+UI6wnYeiO0gWj1TEY611GbORlLMljR0IP2ftjYsQv
Kdjkrr+UrEIJf0q+Qkrc4/pf+bz6fAflIkjdhUbhtVy0fQ9YV9+2sNF2nHDq9k36N++LlQTeJ4GS
1kSxReumNgB+LlFOLNFa9sQbb2d5g9Kl8YXkBYeNSSB20jOJEe68Os5dZmA3+RaFgbVrddJy1c8Q
kULpgugOVGf/Ibc2PyLqejdeugOOBLlsUw1DWu0M/NV1dvJELZidH4g9fJSVKKuSc2OE+O+GDkb2
aMxGrRXR3TGltMmCwtbDIN9WgKpDzPBA8mLIVTSSlkX0ucuCzzrpN/gQwxtYp0yhDMShGzDwlx3t
0rXa2WJp7RBcjZiJa8garEIuwr7/7h3hRwgCFSk8SH+l/SAyPUV1/zX8gqxYJArMEfx9VWcDfo3Z
szG3rz1VjDGQVzjmSdQKJshG80QPjtYqpFVA/JRHTfLqZ6yDrjpNf8rsq+bNvAxOyKt5ywqvFqnm
Vm9b4XyvGgKRWW4rO8uytcTcea3YgpE1K2o2LYmQrG7M1DMvp7JCUnb8DCSIDvemIEvsDW/Edj8x
YuCJq0cUbnJPr9hVtwEwjw55XMFoYLk4CUSfnQCllreSLg3srMo2BQGc5dp1IbXcmB6Ln92nuhek
E23sN1FB3v4zMXp0DtUolfYJb87kiH6pGnLouV+aWZvZE583p/O8iAAuC+w45Shd7EQJSJu6eOFz
5FlnG2mWQEy1aeNVFVPc1xRBV+0J/v/5/WB8rM/jJweJICd/9vfOCJ0ay44CTNalP0ybGAYG6mcO
Pidw/GPl7CWRu3s1c8qZVomQBzqpG0RPd+Ne6hfol846+DtLvzMJQOokZUAiBQK3rt4vFyDYMOTn
ub05TcWSyAh0AChVFlAzxFe+iecBfpbUBkjm4mmC10VhrDQOEpiFVTkURAraYb6darATAwgka4Fz
j9mvQkvqfaSeA2k+2iODbU0c9fttT6ZG3hljNHQ/CsbMxgnGqAmTECHlqGVc9j9GyUheoCrqXsX1
Dka7iugEtsBg/YaiMz1bRW1tk6Czzd4ceeqxG/tQKxzt5DUYihAnomiVuUsY/nCEmeXn9zJYWZHe
u2cAZw0YNxqOrxnfC/ZTNPSe+7V3FoZNl8NIqjx/4q/StanCB7w+U/a25I5jxWCxcSlFyh7Orye7
n2nM8GkjYGKA47IcqBvS20lABASJOfg4XYyY/MA01wI6BzLnEqLypW25r42WluC6M+whtuVCIPMC
9NA7mD3t4Requrw9H+PY5kr/MZY8/0YUrjVVcDt5VuyrfgFUBDpwUjWQqaWNIA006GEpJ7TIHdGd
hnqdUoSujPJ9cHVmP3XH05pQRjmTcq86VhcBh6oXhN6duWjDsCg2uXEYY4G7rCiRLi4au3tLTqH4
7tub8oxStRotkTgGD/D/lVWV/BujnfrhhPw/FFfRz7vAvGFRa67+Vne/zJs7+o4rGQ+MNzdOSYy6
88agPttjXve3eBHj3aApV/Q4cebHlBDYbLNd4lOIaW7PdFggbP9eAgz358pVfQVU0XXvyM+coBQ0
YxT6mhG3MaEZvBsTmC/SvcG9CH2g2Iz8rq7L2jIpVKHaZ/ozdVOIJOkVyHD/7gWx13dXtww6k/ic
Am8LecUDcpGW/cA4WujezznEswBITHmxiwX73xEHeNmXrwcVAMK5UELKQHCw4tkswlPDSY/j/jiz
LzF75MHcrnRqZBpxtBPjrqkkU3B8HvVik6rKtZylOPJTXRMNW+ac9Hmt6en2qMFpuL5zn+ODgCVi
n/wHvcKk1j4+o7CnhkRU5m6/MymjjcaJ/DayAepSHCOY3qGGeLA64gNlyWtuqltvnuiENybyxRBc
F+gcIAcSHT3MTde9voyiSPmQ/oDL8CYDOCwOI3IBBkCjLzEjKuQi5OUoLbBFFDYkrmDj3MLEhv+o
gZtYFVNgBWWlD279XJ5h9MNYC2O/1K+xgaYEIFSej6kK7YZpJR9dJTDeocRoq1WIxQJ3TVpQPZt0
zqT/mOFZR6YugR/eMXIgzYJRIo+cEESYrUQlzFw0oDHfhFn9dEia8bmS4GEXaSuAUdjUDc3C3dNA
h1r7xUwR6QCtu83T8VCz7bMBYco4rMUiwesvnt3J/x4bz9l3xOiNEguCOOnZcFlS4mIEEBZiKiuX
dcheMH9h2gqjJcRzPRflLti9XKnw2R/+1/zi5C4ACVOeYhj/CMFZ2aig7Bq52W2fArf3pyuu6p22
AAQ9eexqC0yvJfnlNnKYzVVYGANmh9e4oUsKMkLwGvSw4bFpXYMLoQr03n7YGswTPyqFfK7b3vF/
WE2fb8iplSTAJFD8/gnD0zXEibO7xVKQWBfcVIn+SCOj9Px1YOM0hNt2u9K6Hii2pYAyeJIAIA72
bzA7sShRhSu6ho06q1Ad99e4blxITXenCIdZlo7V+6QG3fqMb23SJjDR6oJ13K5afmLhhmjPkvVz
t8Qob1XrWS5iy66f9C2+saLdjZ+2norI7ZRrRCz+zdx5kmVOpLFPvmzT3ETm8i5VgGaS8cgsEQJj
ygi2f1tJ5c7e9MwGu+pJhpfM8fkNkIPq7tBV7yqk2a9MS8y6vYJXtNOIZihXGPEoKW+/jSY+ysrx
pMzcA4+a65+MJU4g1x2F7HhnIXrZ/DYjvErdfw8BWSoeuhNcyAW5V/RI5HKqpGNBlbbX5SAHaOcb
3b9iYo1TXhv7Ka3hXhh2yOqmpLRLRZxgKqIpoqnCgzExvf1oYqjq7TNg2EfUUyO+wOpnCSc9HoRQ
honYU8u1Ng1Y3KDnXT8Hv88EX+PHY3UPdju/aE9OHPJyrVLK4jGuloi65tTG3yVweOzkGdbJcmQ4
CfcwrUvBuWzMZAEgrSjEYwVdoQGOETKSr0ZNd8sLDMWDrhHPq01sLi81ooH9SNNyq4JADY4WT8XL
XLGUDp+vTVuM9tXbgpRfJkfvddMCpxDs7llJEZZNo0Q3YRXzWIOkU+fUqszXJHxkQ4DQP0RsuFrs
tRLleNhHe0DYH6rp3eJN09qQdjlS3VYzZqcFcLY9VpuPWw0a5uYEwq3CxumbcBW2zcGepRYbUXjY
sCn5g0VCGPd13WxinJ0kFuwz3wIou6QfFhWWS5nd6TM/BGjMdHoQoAoVQa6w6417/4qs1c2Aq2N6
J4/rLq2ZnRM3pz7SA1EcSZRqvFtrA3MfPF2TswMSxtT5jyNm6ynleJB7F7XwVnnteAUtTdqYd7z/
KciEBMG4L2Au7ZpVcf2QSOOPNSmzHLd+35MpUjJc9jAh20Th7hGBNRPhfsclKXNPMPQDbtVJLlMe
75rO4EZ7FQAHx0h4MXxblhZOYwiYMAfl2pZv/q7nWQEhEeY5621YbYOrTLdO3cWez89f/0t8+M8g
Yd+q133LhPiDFK9VPx8jiUqbmSXf4mT/5ukFi3pBxiPGhYov+8OWOUQ4vSjX+ntR4vDmCLjpTbQy
Fhasaz9UZB1FzNt/muN88gjHJBpwLpiJ9TirWyLRIfhEUuTN4HgWTLHB7MvvL5JYo1iRQLUlP2Ci
mUtcFaCbc/xpkHLRHd9kEECvCR9Xb3fI9pPe3OCxxtCuEvv4tNQ+ohl5Da7MNtiG6E1yPgoieUMd
58EHujwxkuhlvJJDaiHx7drqKggkTakyr3mQCqnZLLOTN/OB0VexUpKv9mLdQbdY4HijqVM+Wmpi
inY71orQ5JqePWP4IudwntlqBgVH09s15WqHLvar+C0XCIWHBsjKhXKNv2/7y7nfzBOlZ3B8TJKw
Kj0T+UecqrIO6659FDstvZSwYHVtlUNphvGZgxpyNic2EqYj5e8Sarl9KJX4OPnE5UiWKpV5uUuN
9MfR+vgLx4spK4a2NTbfr+gG8MbW1uYDuQ8RS47QyP8YP/M3+S5ywrW5dbmtZ27evBSo6T2hqz6k
d8GuD3EYxz0MKG2KzsYtVAbgAaXk4g5XTMzSc164t+AssBo9SsAiiedlE78RdjbsTJB6NY4LZubU
lu6Xij0vDu/D5y6rnoNyOYdispTZ0zJTAh15UAuKp15SRwzEuTEqRTHx/lGj5wld63Uuzorni/7h
8bjDm5fO09zfwag75tpt62VFKUVd5oIOqYuv3Lb2BFM6+Tla+QTWWwr/81i2cPvUUe1GPRtwZJE5
SByfCh6PrE48v93tTKWOQ6W+YoOm0vLy6kN+kgiDRp1feUbn1QQLvuKwpo8O1vnT1HaW6ZgASmig
1OfSQeq4P+5BN/IwdB10/fMF8I6L6pyesaY4Jz6acPd5EHh+xRP+DceSF0KAIwq41GuGBh2Qaj77
59InVV7SJB22ixyarIW0w7Lb8gdvT8+h48PT6wQ8JBzNLbb7m99yojlElMNwMzeSFzqwmnt4PsF2
4bvf+IrMVxg2fnkCHjwK/tzaR/Dwn3ljR1aDuUtvcKfzeS2cYeKjDRjwlYFQ1V2BUaAzcC/ITKrR
ogPivh/qTolMYJqJ6iLYehAPs094VWGsKghlt7TTv7dPFNDq1E19//uaOwwYF9dF0xfL7XT+Br/P
BVM0EMDevxX7LYumo+lKN8mUugorxzen4hkQzPGFW7pENeJmZdj2zl/zjeWMOzScOqctqz4pxPzj
S96FWra25cpRXA6UDIR7KtejMzpmhWiZxF0ZsyHtzqawdLMNkCldFD0oihVlwvoaFhkkNmMIA5Uy
Ujev2L4UBbeppVbcShTmARv4KHgg50JgAnldLEUqxrPz3qZvDT/TGtiwr7Ed//AHsZRAloiTka+p
FiDuhMvKHFrDt85hNDFQs8/5Xq+oZgnL94t9pui7zcKm9qvvqrBRMRWb9/JdSsWY1F+Y8zmu3xpt
sdtez0M/x3ts16R7QN3q56/kRc3iLcHLzUN+0Mcc/9BKCq6oP8tcla2bMEsl4KfZy5yPTVCwkmXM
mtdOBZQx0tGKCezxH8mCMLZDT7zHCYlbLT/OwprOhSfoQ9ngwdsvzcT0YDiyYuWP2EddjJT2SRw9
TudoJERJqiUuL6e2hL7m/zr35LAl+HXldFzK96NxAr+vIdU9ll4j2sAcQI4ZkFAhOqS+xXfhHscs
NeoPLZ4gIqsqqxXpFy51RLskQcNnfteBdM3/aOfrZpgcx20Lrqv2ziNBFB/zhfZuUj+5noPn4F22
gclvsf7WHjgS5HDLfLAr3CNu+Psq0hZN7dR42fvihLCOjpTJrbTqlMXURlmNUiw5iXq4l0QqfLlN
GwK2qSZ71Wn7hIc97Uqj3mCgIIBPqvPC+jDw1kJSaDxxNj43ork6iE6QIGDz9nhTWRGHEOMBkAnC
FXSjtmkX4WrD8XYQYTg/fziBSbqKZmnjQHZ0NXKKKYZQhgn0imYMxqPpWmV4+1JBxYJnvVEsZ594
xGYP9rA/zxw9vg4/GQARFrJmIOOr3IoBZFiAWeXK4UKB0g0hSFjOxLteARH2DbjgstLJw5MnhvEA
zhyxKl4qHJ0/QCK3SPNZOa8FbIAfeYD1yMY9B1T7nY6F8brPsA5DcOyKaLMxOB9tdQV/Glmd7wLy
wcx3wTnymKq0cIFxyjLanPP20waWbRLheEm6LEUPYytIL8PxMaZDlbkTcrJjGHcFxGIceHqIu9s2
NQ1PGKPtdvEWOV5LH4oeM/RjnEdBZLQpGgkvxL08foAapK03IpZEJlvQ8J0hcbhKP0woD/MPNpab
dp4E5GSlkIWjrrKSSP0F5wA8fmyjeO1G+CUWuBAfNNIztp/GEP5soNHbeDGJ1Eu7HsQPeJJJRhjL
34Bi6xFBd7b7qfdu/ScRTyGdOZwKTEsmdJWmqpLrX3gtU1Tz0L8c3BjeKUaD0mLO8iVYyxVrKm7I
0Z25N5dkEbGO+Bm77kN0WDCcK5E3D2YGF4PKFyIMcGF2HTHvP73hqu2Vn9D6NSRBimOh8bWgJvMo
a7Uh74fxNFHq4nONt4kVXfFXPrWOMHz5cdlifOFWkqru0bHPzH4ubE8cONFHu3uQac7fyAUTdvhH
f/8lDAVBd43U3t5MWh10dhmAE+6l9fHSpRnyWPVnqKX6KtsqaH6+SfMOnbWJ+pblso15rWmkwB1y
JthfH4M7cXerRT5G0oaVPmmQiGj3xZdOx9aooR63D6OAwJWE47f5DTUm5jG37MV7iY3FVa9Xdhwu
cZH3FqgshKGNO48l1xXHJX8hTCjhFkb1EiSYUe7OR00IB1ngnyzR6VREMnodOMS3S3uyW2o9Fv8H
mT/McNbDepKUnPr3WVy3bQmZCnC/+6B3NqrMRrNukWQ6oyqxVdCSiNUAZfCUYHqJ3huZhpdI60Bx
g09HwfP1tm3d1BP4QTvdvLE5p3ZLULj4XJRr3obTnG75DdToodyP11eqABFTEWr3oL9VfE3tAsRt
iFLKYkU46IXOtLTSOwO/UXaws9MJRK21D+okx2A2gpHlgdxz/aRglnm09vkAZb72emyuIRGKOrH4
ck7iDt+7D97A64j23ru7Vno/Ri3D8+54QAnSOhdoiRN0Y6pd4t1N4JcNscw0MlJ4T8y9UvoK6ePl
bYm+fxyrTy77qTv7QeZVxpBezrKqDXuX/PahitrGcZsn3mMDktdH7sUmw2G//rZHeoe3Fwwhfq75
T14skCGNhrDaqwCXTfEiAOTa8N01qAU4QUeVqnJvCoFhTUf7qoAdOBV93ojSGR8u0paX/nrsKR3Z
akyL2BdSHy+jXnSktKj1waoec+whJOdxfxgeLiLeebf3SoIaiIfgbgwYQ5NGMDUxWLAFqQXdNiYm
TaHN9W/sx0f15HnpyS1m9F3R+aJ8MMVydY5b8WMfO1ROv73ZdhBaRpWUCs5uKcMZkMV6uHqymMeU
3Z5vp+6l9D2W86go8wS9HKtjQV4RUHp14TBkr2Z7ks88JxqGPWss/z0bRNjwt+iYCnK1jmC78R48
5MmCFxldh8xeJyaSq5AtoUn7ONmxz/8Rgi5VZ1A5HAf6ut0E/xkqSWMGbMC+7Njq0RFh9wMHpUxQ
E7EC+wjUfYZM4E3qm9w8ALdfZsWMUCsNp1exw9T9umTnUwD3JfPG5+BGnV3IleuGqF1TmqrU3HDY
tJ9YvNyYODkhKFXP+rk/hxcjoBm4BypTL+v/BAnKElfOBflIgKHfuN1UzQZRLFLlPvH6cao75hA2
Hvjyd2bTLFHRuNbXysqEn0B462vEpBXvVG5mOwQlNZpZ0ZmmD6R1yBrjUUFX45Q+rdreP1f6UKot
mtxYW9NKxLP+THzJjl63NyT0xs0F4/uwjoz/Wm0Z8lln8J9s3NOAwLo011mbmDXzYv7xcnFht9iB
Per4iva4lMnnuX+YjfhW2uCG8ujC+RlFedyAJxt7NhAkCklSsJRcsMT8vzHrmW1n7vURPZfckoDM
LaAyhxNqO6vYKZ5kBMer2TAg1xBzqpnonmUC490Ps/IRsR5uBcB30ZxL5IzhK/QbgqagJRHyhZRg
b48Y3RYC3J7fsJmuKHaVeNEu90fuMEBCexEmB035DHSU12sC6eu7Ty9XMzeOkP8hkZixQZjw2hs9
Rs3c68m7Jil+syy3hnZnbsc71jEhIeFFGGnMvERVCNnjUIzRA1HAFD8HFSe0usUFg+lVncp+D6L/
PuH37k0eb9+WVP7IYtK/wBhmyJGMHCheB8OKpjgDoclBA5k1W1iXUhCIl1CL40XeNt7wWQX1UflT
qFJSO1SRvAGxQq3akhTdfYNeT4TJtIwUYeHKI1IJnOE6koCHYCyad0yldqBylehny0srulATioos
13u4I9CphZElo8+sCy11B9xfV47aRO+i8jmAsfR2+v5ebt19BdDKQdg4XWJx+CXld9vDtLNu3wxQ
HfIcLAaTgcsC27pdtxcUMbadlIysqU4mEKOmk+r6LuuLDMi5vCfdLRV7jAWtnp/3PL1mVg1fBbvC
Nws9Mt+jmI77elFg+yrEc9A6hxTiTPqfpvBDPhgQaPoro95Xmf5ZON1ebskTwLNvIQ1J513nRYHe
yAoZuOenxi3vMR5jY7YEmKWSTJsnEf+jdMVqZx6dEIl7ZZFD1i9c8PkYWBK551VylTIL8f4xaiY8
yaSrECEi+/HRe7xgw/SLt2RjmIaiPFBSewiHm75odadlnyQKuYumu+T09apdWQ8TO5tAmlbk6nvd
9UcaPbLKXfnVOxiSm82PrtpYgWUIoDHuWvOM2JEdUssLO/wxfBFlcbhUG41wfDtmEJgKRsSttIIJ
RNBrzQPK0vsQELEiFhxqGaK3pXJ9MDKLZ2U1/z8t03LYFrpoV3Lvs15XNzCvw4X2phqvVu1RpwPq
RrrHNuLbuUouHe5rfOP4E9VEBlS3SOJE2bctq8GkTgutBZ2iZCYjlTzsXUcA4tucMj/8uQCur1EJ
XyYR2ShALTvJkwH2tGvzSP4cKbnXIR7ypTozbuJ6+SO+sj7OJgODG3RrZDXMfV1f0S+2EHmoMEFm
jwOGCQ0665v8fmY9hiFi6Vxzo7YyRIU9nXKJoYthKYSZkTC+DmCmUdLfR1Q1DU/YGPEYENn9pa6f
xG5pnroAsBYr7R70wAiMEFoUQm6p141foUlnaUaci+ZqAP4UpP/+s3zi7I+DwR3Egbh8p6LjDzUE
WU48GePPbvP4X83T9XHSwdK8G1TfXEhhFwkRrEtvkpr/oebwP/iFwXk8G+TJucJ0hyq6K/m5OFdR
FoYPm36KLzpzKDSLhJMljSFOfIYy9bwrDwjO2S+FEjlimEBUx3qoifw+3NswLjwc491hNG32IIQJ
eDQpzPVp0cuRK8rt9a4rfILljSj3pP/hzTuzs/Isy+SuOTkIKiMBk7Oor+rqS6HgtIDCpLYlwku2
8EK4hnFrAa5DQY7w5577aK7hOAGGqljDeFkd8aHzIh3QYNO8qajbRSTBnA6xytGRka08sfQtGy6O
nh2AAdedHgjqGb+S4e4OweH/oUCaWAWxgRuGGhA/8yAnLMLSJfrirXMECbdFE8ADPxbSerRSmKQg
M9p6uy8/IBOMfpqu8Ixt3JfxUC0+3iSfDKFjR5zbvRXNRbouCONXr3Ow8GlLubHIONGJ4bmKyQ8t
mUEFr4Nf42RWVKdiEr0gvPaU7EPHO7u5GNakaauCORtA2bnly5aBKVW51QLr742nq8E/fxI0pLvx
TUhphbEozRxcQk/nIveOELIR4ImnWL6RHI5CVqta22xPzOu155COXzqbfF4hqyCD2A8u000KDoO8
LyBZy0ckvuuU3v7VBMN3oe4QhwoD18fbECLJlM/VvKdYwtyj+ZYkVPj4ssZj29f+yywRZQGc9vNA
L0n3hB9tlCCIgu4ObCEtou6GPGE1cjHo1VKRpVEKm/wsYLuqMqSa7bJnLvEGv2BVljlFY9Z2GqMC
BF243AWaM7bNfXCZ+Ek/plRzkG45pQco/MjWfLaLN3H0SScBQGifCge/PZGkf2ikLnJsxaXfi6e+
ik7fJ9sakRKTz45o3+wds13qU57TmMs+6F1y+tlbHeeSaJqMZ26rkojb4m49BOev/+7QKutAftQB
mrQQ1SJfeFqkVwVaTc6PzVkGB3SNG9I+e6A8aVdCmKLXroDaexmay5bJhNPRrzxY92HrlcWEz686
ZtB92pTkIQcjbSxcxJL46E5ksWfca4OiW2B6f8OjaZNqccX/gaR9xDI12nqYg/AuOiKi+AASm4ux
uGVjOjnB3j3WK0uJVJv687UYT0gvn8xrZMe+iOcOPbFNJuIffQBIji4dpqy/yXOJ5bQuyU8s6ubz
MVMTmlFaf/abONU3If2GaCTAsTX4rYgIzPBuH2HJsySNkF9YdZVa9YGGJzgkptIJuFwXDuYWJahE
11IZ47NuhUPlkHqSCi2k5JnESz8xQAnO1xG/phwBQ7Vu14bk2diWcZWUJkTRAbvGA1lHGSQM4cBc
NEl9W6r7jNTuzUmBHbPcbyODT3gQyZOCN1zmB8NrXkrJJl0k1dtBlMhPAN4iyXzEiK5mTeWWg17y
lV8dO/1MVAtZXsBXWTp6neVjHxQYV8yVCi8ic1OEh/H9N//nIKPSgO1S4Q9gOApK8eFAYd5v/Vut
OTzLJ3kpOOvcVvp/kEcLe3f/wgSgoNIQJ+eqG5QOCTymsmf8WsQlLU6KpSNqsa7t6z/NhCXUtdpS
8CK5Xzyo+AGl7dnUu3sJRTOw2OiaQjdsQhV4cY+XgmFF9HBtcAwMfA+aZq0y9Zdud380aEHA3eIG
IrZf8EB61KnXLscpFt/3rUyz96J6R2HG9ATD+IzucUPObZRpkZpLZykx07W1YZ4e9l4dNmWRZkS7
q6GRnkdXbIX1Sls1sLuB8BI81N8mRdE2a1joo3VOSlnM3ia3ONYdbvQYZq8S9+BbdgShvLWQ0SMC
GBin5mueoxkGQmhM/Pqu5bjaXz5dxqGQ993yhuJ796fMBPKDi5uIolMCjFdzLunPRD/rgD5cuIym
Mh9eBKaGUsbeiUaPCmah8MjT+8cPAwhVhs9PxDoZ0x7VXvB4+yqlitaGnocN60r7UiJn0PJu04Zp
tprcHG+7V3d8fa98LpUaRZgDjfkdBouyJv2Yms8N0w7/NyhcP06waah/QPuIGBq61xBApoKvT1uO
zHi8lhjtPI/UkeFEcQEEcIiiitoWjUKjvqu61HeTPhkIbKYTeskDWHqD9a4RQaPFCxX/o/zKYeRS
bUgk1wx88k5okvbPOZt12iE6ZhgkKZ52XPHZKV5CaThqp2BEHYXI1vDXj4hUDUmKY1ygvPlWkETg
2UgAz7IFkF8amqotn4YD19kFDm4JTdB69wOKkW0r/INfUaCXBDlKVHljjMsc7C2a2wnd8ZytQeQ5
18/Y7WzLQccZcotr5lf9ucsC8aGnubuGg8ah0tdcMXK05g3Y6Xaic9iVTZEIooub+5+RFWnQbRJ5
3WbXVOG89RnYUAeCrfYiVb8bpMC8V1neplsmuj9f6OF7uq+ROUvJdyKQBbNE3dYs0TIhJASNk5o8
z5imLKm3dxfJFeis7i+9c9avGYFsKDi6NcFyNY9L+glqYQJpo4lAMEpkpRgswqt/zCJ86u6IRxkx
m39hQAucBRPhgZZzkH41Ad742j/ONx12Itt90UafAwep085CdSjQDyg8s0+TDo7p7/6wY8vrB7Tc
t64qPcRFyg764km+7QqG3gV0Nh8sdfC6lJA+J1vORjxBZ4t6NtbILZEKmuWuZ4KLoaN7QaelLtzp
wF1ejm3dCbUTzI3cTu6EFP81ylug8y7jTr1PfXOk5ZlhzuOEew93Y3OrkATjLQ0I6tj18vC35r+d
4/oYHHpx6pJydJdN+OmrUxYGSYgBIjBTYd/OhFX1RW53eSmd6HcnkO4pvZRZpuKm7cNWElUmHdLh
R7yiTLiUIpb9qbJNdAyCEOlcVyNiwn9ksbuEy937/jjzwao2yCbkYPnUohWsPAi7uUT7ZE3gJR62
zj+I1sKZ2nKEG/4M/9FdZaqdn7ri5bix11Wf3VPv09DGY+OHWdb07AtSwX7GDWbXVrR0EVYhzfww
9Ea5dFvfSsfs7LczHWTIQNrQPv9tZ/k7B2oKGfk/5ihR73XRc8IDJPZSg6ZJ5nk2Rdr9uZ9eTr2z
K9MkOPaR5oIGO0GFHOZtY3NPK1FDjnnaWelCuGPqSYMT70rDEivlEKkx7wY06VqHv7+NkFzJZpVn
u5VdmubdkrnxnWF8kWf2LNtXD2m2qdNjvdfBGthqzJWpRV58B+P2ZESiCgPCC7OgDteS3gffuV/x
NFKF2C3OCVmo7jmi7ausHQXxrYH27Few3BPVSbWZNxRE7F0DFRStYsi2L7C1D9WfAiHCrpI0V4AE
GjD+R0gPo7liR4KizQ7PLOODylIHt/izhiKqvLx8Ev0P3r+Phxhdcw5j08jCSahvwdjgBif7PTQB
1+k64/1SopMGREV2pZp2Z+CLEyvgrXrogDtoa5MwIWgMHe4lEHh7IZG12+C93qcrpwhCa2s7OSwq
IdykvcW5NYFC85rWk3smrCWXCupzuO4ZDdUyTuuXF8ZnPAGRRma4ZMy4dX/n3myUceU/BK4yp4O6
3AudfW4Gl1DMGMYg0u94S14pyNjG8tj9kIvbWX19NsfzdHJBOzSC2hjnnq6v8buyHMyJpzzKb8WJ
kuMAdLyBFcR39AIcb1clP5gGOchsc6YNtVVGE5qNpEUzxGIFSQXt99/AICq2XpWNg+DJFHz/+D6e
eUQzNSrdox0Zv4HqDhiqLA9NdLDtmF2Y41f4vD7wJ4R0YHYVvN12r1RzJy4sW6DYBgT0Q9UD+1xz
sYUJG6llTR3xdZtohKzMv+I3pi/V/HI+0Lc3CmsDGwwsZHGZ2Kxfw2zdVPpYXVQgOorbraV02t64
U/CT6H4VD6NzcFRm+EuLRQVv8Rz6/vGCqUWZCLzV0XP0Cn7yMQkW/6VZcwyLj9RW5tzb23mjIR5x
B3DK5xArP1OFnQhmj0laBYvCdhGmGI/e1PIU6fAplYNcrUAqHdxz+xzYv/1vYJBoOBwXcPJ26sXb
bpGBQrd04QTzEWuHYtLjM7hygh7LvLBoPEG9aQ2m+ufy8asbWg3+SEymF6Avv4cd2sQK5ZWfPrPD
xKWLVGEkfVJ3XNyJvY1HvgJP0wVRIKxW8hm30//pETw/tl7Imnz6q4XCpHRHgX2b8kdQJJwhZSgS
avYtCOXAbT8UR7PGaiR8QPSo+BTBnsBJa0K0qFafwiZ7gJhj91sU67ZyWEtoxHDKmnT5lVXOU7Oo
z8YgSpplixt7e/of7ZWdzdyFJcUb1qzuYrD8srTP/ICJCuCVYenagr3SPtsZ3hNN1EVlbISDHlGD
BsFBUu/lf0qwrXvS3TeIXuXaQ3uzWetHTCjDeuTPTd8CULunlExeRvqLKQVTT/uKW6k1AjSTNDrv
kKJKcESRx6jDHxbXYCnoJ1Vc+glMarewSGrTftwR4wxIiy4mb9BhxavHcwwoO4wYBHgGZaQnAtX6
zi6X2kc0ot+whly3pAlyp4B3qtcfvwLE/ewjNzBK0sOZ0jFZ26rVHvv9OYcXg00TjCVfVtQXZire
W4u2325rBPBSfiRBD7DxPNsQuDz7q7z4+EN/gtbGqRbDX0UoyRcbPlSfncb1QYiotn/3pDEXuasS
xEhhhSXDfjkdjpzApFmgd99TFemf2/lbr287EGLGa+4Sgy8i1zCSQ0qmTDcA1of643yfWfbd7FSZ
nv2KagPdlUF3qJOnc0KdGXllFZUHaVA7h8MUrsllG7oQZpvHDNW6SmjkQXWL+DyoucH67Wxy88M+
ksWHTz5vaBUDkyZ+wLFz5IuuqEJoxrXemCiQtzD9ynM+8QbI2swjZpi4wzb85BZlSrfhqT7VEKAr
kbIjuZ1G4ZTCKNnJl1v6AXh4Ul4GMZUqKVAKSHQF50KU+QPRE6CodK00QlKbrpmAwu5oYVstIFGP
tEGq7XjNfvExBSa3HDUNGoV/0qQsJ6wrj1FLYYEcKf0eFa8Vpa7V6eW+Qy/ULYE9vMkTD1qp8Jyu
S2SJ63IfOX9nIpeVw2VNv0xEsBx6eP03Oo1Tb4MaC2fUC/jNWNjYx6Bh8h5OVccJeKUu98ToaVgh
X/JmoLu3NhvQ6zw695vVR25Sa27bqdjtTbEbIxOVYV9OzepTRbAsIZaioz2Ge5T2AS0GskBhzITe
82ENeWQzNMAVO66eWfmnOTY9EB4EtLigGzLfHJB6wrL2j9F1eKnvGW7huEZRoGgknTVitkVuibm5
dNZnsZJWQd+M61Zyaht4r5oezT8+K7Wksl5Aup5amJXwZu7R/8iH2W2cNdy6nqSC4A2viAfuDdfg
E9Tk9dfqclee1GSVAEandN8gQ/V0Dx/3B/mlAcklFseFgorrAX3/Ww8FTgfnCR2IioYya5HQo+hY
LDghZ/IlqcemPX9Gp936JARe7iUyVkqUWl/ANxkFvZutzYKG50BWPFpMwGqYfMmYEL1isO+oW5t7
YEYR+6n7T6vlF88sjqaVFwzBzMyIPX9fonD2KYYvh/+sCTPK6RKWwQPX5vaQfNyJg6XIR0AxCXEe
BppYKOxQR8pLVLWqg9YVfzaHN4DVkTAOX8IT0KqXvYjSFc+QAFGbIPIsTKNWvt+UxaLNyBlEk6p8
TV/4bo8Gqz7JL/C74v0mLtXCR6QP21M7PQlvo120wN8Iq1+F7HycFBkeFhyYjAG8AzZh6l3mzGZ+
Qby3561ymzy2ahC64yOFQB9YsP7cnB4qtrOB/0GojUvseM3cXQzFOipfXRy/dRdbVUMoYnVylvXy
6/QtSD/EqEtWvJeJ3Scsal/zg8/lkKmtFk6q1OwYKY/cn3frninA4wGIVjcA6RHqTbgROfgg6nFN
tldka+tM5opZCjiAoRaCWzmEyVBMKGfHmNFucU99iBNhNO6psteoYQzDIc8AbPCOTJ9LXTtr1Q+Q
38WX86u9L7xpBDKr6vc+9ttnPHq76FW+ikoR+leOU8wRIfe8S7ZpeDlwHFBPXI7nW2ah3LLeRHck
5EyvaoROw9hyGdF7Lyue4VNyDAlXqtHf9Xpg7q9NCtZ7n5Grp3DIxNL3dnmP5XIVqHtCPA4KIet5
zIE8aNGBDqFwq2qLopYFmD8gs84kNLhW1zHTKF8oDbuBhP1cFpmroL36vhJ1ZAfpHAKfp3WmFd5s
l1uuAFbaXIn+mgVmaD+CxDhcVPec5FhLqEywQmDUroU7D1JuyipLY+nxkOBEicma3ZpdC67Qsbwm
/DyqiSwskkjcEODwhI0VB4u/z8aaU8vZl8JxB7YBdCsjBrSA84yH2mDy38AHCrQbOlLzkrd92pCc
tRtAauREnib4f7LGiA4weDrVsaLTXYmIJSLpQnjIJY2u88MRqwDxKKSCr0gGn8UQkq5PekEfojhH
mxbSTkn//EDJDr9/gpB/yfiLpE0utHgwF5FATozUgpLsFxslfIG9uhjpghqPp2Zc//eq2Tbx9d/j
toskdCK7mBNmbXn0QbHpeoyKnBgQ+BBbvQYzreisi35E16woGszbgwTa/mIZ7CewCnYDnMzNsWKC
ktmCqaD2A+pRDuXW4tKWZUaRp+fgVMbhC5i/HsNCPiN+81IpX57mhuDwVF4oRhH1phMxiyWv2jF5
n2A65ocx/hAm6cUfcKYSACvh0rb/BTzMDZi0s0hgBvirVLR0ARQZskVR+8zVNjBHbG60smwbh0d0
PrzVBy3ZmkMnQVSmP8DlpHTT0dU6c7wmEFeuFETkTAlQfTRgMR5A85uW8+XI47gRIuXOjdm//cHn
X8CUliYFqVwJe0AmWBDuRmzZE5w661X38kk0PxSxaekkALG4cP+vljLagea19psAdGBJo7Un/tFN
EJqkL3yAhmhbOakuP+gEp5rtjKZDv1C21Cl23rEx5YCwY0cyv82xxJNoiFaZgxJ+/H2pdvK9+4v4
rTgnzT8ehf1AxQvrlJNMKMDThIKJq05pJpSd6XIJI/HCcygebVb4i3iz+M4GgSOYteCzR2fmBuMd
x0HgCPbEIuc8WECw0Xxhk2X8tZ0FTLxkSX/s44eWPRVZ8y0JHC1VFgRtU6ZiVavgORrBOwboHJg8
LQp3kqELUQZVkofN70/u/rbV2KC7BkuzhdEEuzx6rxZUqF7QRaR61fGbCNHEqw1AMBNQXGqEpzq2
Z1o9cfHwp0ScxZ0Eq9PqhU9EHNwF024EnniJ0x2mZhvV/hVoaIQQhmzUbFnqwn7UTPSo8iwzLOGN
/XeKaDYxCFeVBZGi5kvFQYm2ygDOEkFlyCoRY9ynsDzcco1FWlUIh0bc/tpbuEoOzivMGM/m+XtM
o2HROcbeMxS9cNuA7b8aHvria5rjNziEk2OWPLCTTPteOUbBS+qpkVl4JwgFGd8d9lD/3p2yh+Sw
ATecQRw4Qpg/f7jOVsrq4lNA9iNM31hUulVUPSUiTyi7GDF5S+2RRJi6RyTk2drKV5UXqQkQ5kKl
PRnR36JspEzANuN8AVt+R1UcHXgHo6hKDkyMM6iFHv3BzC7AaH37P5btwOC2n5AAws2+s+xiX5y9
bIiXuOJslZeiu3Y8hX6a+lWXtiSXGyouEj4Ro8r8vB72Ys0LJRBT5g001bnh1j4rhrIWrgyDYIf6
WEDqtEhnTRPSryxbp6qw69hGG1Qh4i29xX38CFgOE/+rPSPC4rcePVlmBJ3ckxWcv9WgMt0h3/bK
gicq7yjuPz4VzFerUiu1397MOvdeC8FiwPK4oalqCXZ9KVR8Hv82D+Wfz/8UjpGcKCgbZUAyqAam
hOJ5pfstCUoosznKhzn+emX7wtpuH6S5/n0lOCsn2LitGI+6KliiLOaGK8nZ62vf0XAzY2S4mEH4
8omaVSTjLF1xJQgRQ7/dvs50CbQcgq9Eaatnci2x4P30lQpr5YbwdyUZPu14TjCfdJtq7r81uRvn
RVapRAUUiCUXdMBE7/0lYdiV7TFR1ApSp4x64RKCN88c/XTLuKkyYyPuY+99WVK8pQ0639Ucijff
eaa7m6kFni087occWKACsa2jhmc0PqNryKf57re/tYxF+eoloHYBTp8bl80WIEqCS4CNmcBwI+FQ
moo6bDyFl8f1eKKiG1xn/OAUkVvVZQrpsE6LdSmFopLPMuEpBFkJ0G+cdUHJwJ8jr85vfr7kcvkT
fgpJ8Nw2M+hK8XcwvjAtOeGIKox5Fz8y8SkuOO00eZ3Fy+PSWCK1xU5ZoQ9bkcTF+Fs8f536ddMv
BZvgOgUeTzN/+SqvWJHEn2QaEYoNe9zOoegM1nrotLNVxmy7WOloU73xiEU170yw1/herm9AhxXk
Zh4T/4EsEzKcptp2HxeT0fLGFiv1hOuV00CCOrTgmIbxWiKSgLgUN/rVbPZp+7oJxUp8u3CT5D47
ePWLkR4wJGjNAflM0tROaqpQjJOvSybArfcLqhp0AnF26iqR9hwe/AX09kBEByfgpXzXz4sT4YIz
KhoP0Lv7bo6qmilGnblF9y/oYHAbBG87qyEgHDYclVRfsaixYsvUejqKM/kxpiIc+wUmomvbCUdK
NyS6IR1UWhxaXC1AMcNo95FxPsZA6yRb0fKVtYUZu1Os+z6AgzWR7bd/QwwyBo6CZ8tBig4h42zs
9At+vLyODA5V+eyqXqp5EUJ4CUCQFBa5b59g78EDhpb0MJ2UHApMAGRFU0CYjtG/Y2rUKUYtmmOD
gHPpjRhXEKIO/AyWY2nzls0zC4jPIYqp7KPFygrcdLTgSDtYE2Oo+MqpoGGtwl+BS2gs4RS/BJKF
gL1X3/v3EQ0Kg63Uy9Ept23eD/TGJp+CLWpTgAJPJDpMNkhqhTOccJh80CagsG7coZW9MEsJZidr
X3vYhHSe23PrToboNlLTe8/DFerCyquLVceO+2WOt8BCJOZvZsXHjFv76zJ4R/N4+byDjiP+B/RC
TnjN9j6EJGp2Rkvsjjui4tcqFv4bVTyGS2wCfCYJ6lW0iEPbXEGTsqioHYey54ocAWSw7Y2eWP8H
NPRZRpFW8WHcIPzu8pxRE4y+GmS1nCqYagESm3Ca6LAADwKDU8YwVVgfXpMVuy+vA4ogYsr1Rhy3
ZuBNgI6LGeXdKP/Skl8pDsOgl7O259s51/a7DgWuMv3pyUpIZuSj4GiWJz03u1bVpj2Ya39jIWCk
qMn2OC1S5hGKDDHA6XvQfNXjNTsfY3Y3QlqZZsD7oHU1n9A6v67CDfOWsUq3YStXLUPAW3b151ga
FTlu7HsH5KKa/T9zIShFW7lACfUvLlf9vKIr5jIOzJYNROIyUU/AJgfZUAnxE300L1o9AT+nojzg
dHXJqy1bkahx+Bk2CiSJLUvVEfHPeiWRsWrBdgI43115gsrTA+n4eYBayNHB34Dz4IlFYVgakgLj
Ii8uMZhFlOOwkuWx/BxcjyWOMJePTKkWGDzFHt+ufDbwnKlRx3G8JXogWhW9jKfpi6Jj++JGvSDX
WtQZrTyyfP8HZzeC+LNRKZ32rJ2gkvt1onK7BTGiQq/kSMgNqqQ57ioxIcuQXSgGIVtt+RN5M7Hr
exZGp84thuiMYl8VhEz9ZcJvFSK8QHXF4xuKna/Q4d9RaVYIljqgZb0DyGbKGcf4xuBsLITUjeGr
UokOdhfPoKxQWNmqX1eRER7LD/0ynRc5oVVVqEXQ3S1HvlBbZty7EUW4pSSaEEGGF2TXAKwQHm4W
RWpzrFdHbf4Z/0FGk7HM5YopsuaymoEoriAep13urXWZd13pNPvcsWWRq/tMWIddaQ+RtRGir/C5
0Mea/Rzvmwp1r8Tp+kqyiD8iKG14Lb3npsHRUu9QOE9qjOpcp/3H0Zw3LSsiirACyikpmtnhJo1t
p+YNUjDECyf5vV4j06+TaIDFn5QSwHyNyxjUktQyPx+z7OOjNbhgnJrIrswrmL9h52IwuIkPOzDE
Kl5aNW/CCu0nvXxQyng8yezvbqZZj65hr53BxXsqGNsrNbCf6lTB+upJbJrf6nDv5G0Vs8G1D9As
pRyLCFz+um10reneFOiUUXL6P3dEFSyB5AqvXRjTZru9ixSabk3dTQq4P0dgv2OMtR9Y8n8o/heb
jj5ILDEZea57dngq+wDe8ojwpAjyxWABuvcvq7VAUOdcCA0oer8Zl/cCFjEpJ5vWIlTD5IfE7T5f
mR0fDTAMUMsT4Y9mpyn0lL7Dy8pD3+HIO5oJs8OBy/PxjgOF0YPd5xqqIhmfA4dHwrFx2sygttmP
H4DzR2REnSMs8cIbEis2SUT5gXigbPBJdCsP4kUxypsFI937gh8LozaT0ZNn+PpS3zBw3TIZrPL5
W46Y/zvQWV5gSoE9Z/wTTbq+Fc+EIp9UxBh5X96GTLp6S1dALy4OVP/7htp9IB0unfxPxnO1NG/z
DE+3UZu/6nehElw1xJ1DgqGbx3yWSVPnWJRlHgRqRlFdv4IyFYem/ZIQvWm1NN5g3SWTdeRCyFKO
8Ij6wvnQGQr12XH0RaIvR6d9EldrurG77XiIOSr4mW9X7bMP1XNOB6v3wtBfZ871H06+1fLFTM9T
fYMWX2KxH/QC1QcoHJkavcVWbeohAmCRBLyb+v3hbUtVf7glN59NC7bAYOBB9UhQA0S7Rl84a9j3
H2OY+PNAx6aQ0uxDNLfQQ1UY30W4QEZ4xhIrjk8QpyB5870rTMIhiidXs0qLujd+wup2JyvMvfiR
lzuH5/hJbV+znY+vYh/Y37Y9QmYXtMTGLpLloaKpR1J9C5xg+jDZ0jkUUpyIA/xrLCB6SFgRgTfm
sestPL5mfFw4+SBWWUizTMb/pt0MFtaPu6bBUjdS0DcXxcc8TSUJufRKMK02VGtLGU6hDm2ftPro
h5z/c+2kLznF+vWuiDuozI22HCqcWb5RYDTsbKjyWjo6ft+1cDAnwNuxoKX7XpAe+56XjkIVBlYh
ltNyXURyFxFObGb/Tbgs9n7g60S6qM5+EoKBTxhVn6QSb641JQ9mfktKCmXR7JjVRxGrvMGWhbp/
d4FYTiYoxXOtTl8jz5vgGHpjjvSz9XDXDob3vNabtvyAihtVgpDL1FMGA2r7Wa7txLjDGYMeCzL6
PDGANQXUho7lVRO2AH4Zq1r/Od5CQSDWKfAyBrUfCI/00T1954Upgk57GXiuWgdaQz7C6wjgxX8c
EOLaECldLfLL1bVth4JmTVgc/3JDygGojm90JKhlQ9FCO4HWJR5/1SiiYkT1Lym+gPdoydDMvWvP
RHQabMh310sJuCNw4ZX1dzm5mvWYAw41ZyusqQnxfL+zI/LNDEO3wzjScfo2+vfnJ2eM9NOqECY7
zuzY6zkWT+seJtFGEyY2Tw+kJiypkuhn+5nhzrz+iPlc6qJXFv2t2/0j7HXbVmFVqnHEGfhKRkmD
Y0E9pNK3bQY27ty8gfWwVCK/7WnHrQmZqepfD/sCYvOoMeX4TocOzcHlBH8M8iKA4eqyKp15X/eO
YcFf5WwFyvqveg9nqTSj7K1XCuuoEcJg4pMaK6xToz4BwxsKyxVvJbHSKLH3cskzFRoV0+VEq362
Ls9yILJRweNukAgEUw2y9+cJSLHgb061sBYg5vGP6vfsmbkg4XjNPV5rkOjEIOK4RwBimFlKPNFV
lZ73zKtPq4PPT+zSoFuU6U91kxGwjOYC7xJmmaK7Wibwk/v6q/dRV08YqmnjykrYESotImq/Crm/
Mtkv7NY9vZiEtJtwfp04VKLD4aamD7xNzKYfAuG1gUy62sFfOEhNPIoGFXz7vhrsNAzMK/Owjr8W
yaZkAyP4A/jur18pzYKHMqLOtMg141xcKpKUM5FQMecyK6Wu01xjgGJB2gwkT5gfRopYFDyEGsk0
itQYcAKnagDdjKf3A3c7jVk64dYVzZYz7MVXteMXIv+S0RjTAoKHbnuBq9+lWpoDnWAmTRk4PHBx
ZJU8vhViB7zxbgRkRAIjhz6n88UcKWe+LmlyD+q3hV+N7eNCNskygv0sXsk2+oc/ZI4pG7/3r514
sprTOqU1kuyXVjFtCd//aZX0KWkXcSZ3P1ph9GxUDe0uuXK9J7eSTJsa7FpV7/cfzPOkmuhPD8ra
7VgBxfEC7kUX4bWd/bS9veVw00/EP7DZz82jRH/9uTiEcfUuoslpD/WyVtzOrFuT/ljJMxSAL+v/
Vw2e86SHHeVzBmmmaIqebCB/MXnYS5uWV64Ay9/wyDTIk+TF1Z7ZCd1s0z2gMzuonO2Mm7U13Vuk
IOibJnunl0/oeYjm3w3uC9gxgC+r4CH3FHoioZWoSvd14axBFbPUmUfGYQ0Yx/eRHR4ynA7gU6kw
vzuDUKRriUe2Ap/BnMPYkovMm5rE9K7AIflV2cPhk4+sqK8X6NDvYJ0OwNRqCayyJG3tcdNJ6ziv
AJ3W2cs2aAWWaQLpeHMDBLritdErnAYn6VMoInQ/IzCHRT5OfEbxzDjxc08/Ohd7EdtXbe5WQYXO
0+IXta4vsMJIcWJakjij57dsGANmcfnVB1iUGtumzOXYhLNJmlfqHQiyFiEuWqUERdaU+d07fLZa
IjRQOeIfpAcVqX/2wRzs6CmIZCf40l6k8QfmHCZloQYgjoBQ9CgHaAH556tnUsale75SSMBDVpAK
rRjBQ/kf/2m2lno77bQUA/bPE8ITrkWHpdi2s+D2dNsuy9gMTZFeTcpUXkfbJsh5fBLnnihy+QoH
DURhNEj3QfN88X++ivOSZv068/QZmhIc19AjHfyO54vX0UZo/vAqHIE+CMNmij3zef9NhkeYi/vN
Oyw5M5hvx3BBoHh69ewGD5Tqyq8tJaGK+UrmUWJ+NaPNwzK2RhBiuGXqTECWnoHBLCAsDUPxJUpG
j2IquSevChUZnmi2G0J+U01OEH6eij1LDcBzCvb+cH02xnsVH1bjreLHKjBVCfoMP0EHz+SqScWV
eIoHLyMXS7o5uV2/0cmMlNsgRLrzn7XsL/f2jTjqfQ2MIJsvIwACHsZE6GEF2YrEndTrrW8nUshl
aqbOTzj91YW/aSHidXtBtkbG30bwJcV3Xo3Qo0yr9HvjOepmJ725Z/MIRml9CNeN0tNFT7l7W7el
blQ8K3zQTxQZ+Ofo8bGWlcz6M8NAZ1muEsjI8yAUwxLOuO0bAG6dXEuto98sIHhN7PDyDFUO3CTC
dPacVDzdj5kW6NbkqYN2wsvCeB58Q7aADjRGnLWSbxlR8D2mFvfCs973li1d2Lfk5P96fKQxjfnl
yjqPA1Q0/TmBY/ahPKfcDeToV49BOWxx0GzYMRIRYIPmY4TwV+HY79r9X6sbpl4mc3Chhiph1yQJ
uqOCBZToN5Stkiuh7UjggSiMyKzr+8RC65fbwWYo/93q15iMhZ2jd9O8v6sBNzZgQnWz3/4PfLoA
i9lk5FJHC00u6Bnr3aui8IWbRTJ1WEuWgYMczrOccixW98h8rQhE99c0DQobHRkrmEnqKK0lYanJ
pm96kPnfR8AQeE2qwNz926mXrVVznu1IiuaN33dTFQ85IZZgybX7aCzZA99faCWSh70f9uVAZ/xa
8qAxflQdnaSM7NP/WeTQLlKLCzh/QiiqTL65IpM5AmiO1nlkfn23yQbg3rtUmwSPCj5uJc2ILPZM
N9To12HS0lk6rtPLdrinKq7i0hACyjkdNsaNnVHMiKgM02JiNv5JzhCS6+MUKZsyVUWoZ/vcjlnS
ikYuEaDjhucszpud6Fe7jr9EsOGs9xs/mBeeJOse5aBnZdhusFehRYWhOth7EaHcIZDxFvbhp0hV
eAO4jzdq2LDe7YKfx2q1bcSrRyzi/Ej/9Ib9ImmMcfnaHO73ZYnDz8pAKwhH09DEi5hUW+qZ8jQg
UYoa4gRE2/i+0jiMhcXUNFFnhr4+AHjGMSDACUdjgJa7VMdzRNvCzHjFtmQnmaRg5M6v3nsk+Dg+
zaI4wW/a82nECLzqGx6r4Eeo9mF3eNP81KeRlq2tnmOmqEg6Mupkcp06Ie1H118Jvr9fgUZWagDI
+h6XaEHh5x6R6L3S8O5gGpy1EJ4oMkcniNln4EQDa8mfpbFC/Lgz03wLetX/gypOSFuy0hlANZjt
+/wUZ8VUU22SsivjKGwvc9taphmtXRIrk2iIHw3GQTKLNkE1Kafr68PzgppNbiW8Zn2BUlDt+a1m
gyUV7k4lWznIs8tfMJtYhKv3KbWYe+yQL/ywmp6bJDOBgNG0fAmEsvjePn60P2ZW2jebfaQZpkhe
L2PbzTKWVHFrQtRlaOc4lBAdv5HH3cbMaznOtSkmlnMvQ2uM9BkHAxO6JwP8e8PwM66rkymgZ7Rn
CE6TkWnlGqDA+nN9aWHlkVYbnkRhLP51m/SQFqzlJLJfcwSdz0NjJByCqKObOlbXLV35HLSGqHNS
cufG/TrOP4h4G5U904yQqxS6+bGWcLNnOl/VB1LRn8JZ4UZqHII1PAjUvJ47cNIGc1mMiyVuXDxk
wRQaiyZY0zJV+4J4S0HB0r7S2PjZ6RETDhYbuYRY3WYPN+G1nJzqfZgkIZ4q1uEicB2SCY5RETGt
2qS19Y6BqcnK+KhbZkCJeBjuFuaGrBI1s0XDtoKaA5GwsfMQnJ3v75Sztsi7+rw9jfRrsw+gKoE7
RUpuQhrQiT7H85XHNsv82dBHQPlWY/sqEjYPBJLOy258k1R3kZfTovYrTEgfIBWKIYbXWj+tn4eu
vSXK/pQJUO/sM8XgTp6B6gHyQe7aqvYTLv1UEKOGMeKTxsdmxmqTswkMFzUppUg9LqhZUrT5cx8y
N8cTng3ahvptaqFJO2CGPSNhwE74lgBhusfsqi7GML+twCPaA4AqMyjPgAQATFfVpnF5l5/fL7V1
hg0HIq/x6EhRU6KhY9AgE53wHin4ku/H6RvS4GxTDh6v0s9cv5fDV3VbjK8qVPggKS6J2+AJrY4s
YVgwYb7IXhVhh8cKyB3E5uFhS2VNHcIlfrkyLJ8DA3RVyqjGFWHVpH/hczd8iV/QbLxoOTqc0mF4
12JKhBPZ0W3hu4CJUWcMLzg5R/SnDuJvdZUB1ygSahZswbI5McfIq6XOonPSWnhg3mu4Ba17e5yF
xTxbh3no7yu2UPu7+PObRXO7dYn4PyOLYkc6nLvbAztezI+z3fNqYhdbXpm5/39V1y3z3fotEYEO
gtdnoSrMiag8kctG5myxRMnkH9eSBMbKZ4wfbslJCW+qXpGmd7rdVVKEnB3iqzSHQYQ+HVdeh29m
4HNe2/TkvB59AdZ3lzAipY5QRqnJgUONnxkr66NRqmEjSFb0Kdz9w8rojgZa6i89kTyFnYSMojx6
zcPQRhLNqGWLfjNkuw3Vnp4LFoUSn+F30dr0DPIsbshO6QaOBcvdfD59FCIWulmMvRdONAvXkgX5
GUxIdiPZgFyB/u3iDiBpD0w7JyzFwfrlfpt/jjnX8iajiypMNT5iBkA2Ll9P/2AWDkiNVVCdJJzV
t5L44eUry5/L1Z80HcnwctKr6a0GqTJLSOw1yKbxPbWdb283bv8PV74P2LXVDJG19bvpHlTAYqS6
Fklpeh1bolHKj1yQ7dd27zm4gcoqzp2yubJbF+9yKSN/tYzZaVJs026i8pmz+FULjCWYwmAkgXUs
YWMsXmdF1EeVW14kUS3fSb7aieb8CjHsKRquXfnbWA2gMjXmOJS5rHF0iZpwObTpUNnpuv/YWWua
fe7lfM0b5JYjg/ICbKXb0QkvDfMP2mbquR6k+6fciAv9naw+uVKciSUvK+AQ/ukqQGUYEfssrNfM
+mjnqQNj/QTXClMhzuO2yNyKvlPWxNm1iSudJD+xhZmg1CsahYjy0f4ojxu11S2dSbvdkdDjMkZo
3Yrv7uTXlQStyJWSx2U8Ii3u85ayS6VfCyZ8BjKuc19hLnBep+XmImbhvlF74kdmwHLhfSXuoK7Q
fAM/YHvbC/99bUt9UrovcEXJFLDCxRbdWqJp/H9O8VP4tjY2VkPiUBvKLIH1HTqhu9jmRy8dL9U6
Z7DaDzc7ZHqlT7Z4WIE+paac/CoE+KRVa/QD6NyZYuGMvHAevyJeuwFFZ6k4B3E/dYDaAO+9GiSm
omcUCUfyW7WgEQ/z8lS2URFHLrsTnx5PLBDZxcoBKYfO0Xfxiu9wSdxwc5vZ8L31mBO03er9DivG
PypZiCLTpkVpXXV5voQur9Y4+6ClMAMFNdUrwJmLawqWJkPfP868/2c2jpsQ8CZII233VivTpA8J
hgpnl1yOhiZhPjPucUlApOYJRMGdXde1HbBBcv0Ex/lxHLVaujoD0X/tCaNOXGedvV3idPb5+viQ
GmgTWTlCBQ7wubGl/Dk8BnliNNVK0emdS9bRlvvyFfop9DsSIAgtfuYCEpF0kLcobSO9trZPgkbC
rYKrRkNY7oeVLkwp7oxLvmfBUWHMuonGiAktL2SI4OE71H+NrfUy/d6IFVud7o5v28bOWMZU0xG1
zZM1sylfQfBhE0Zp70JJRxUJ3Cqvzy4vOmzlx47SY0hLExtks3lrr3NjRJ+IoyjeooPdZFcR3K53
LqRTfSeyHK840aGkXhUlk1lUs5guavoE0lr8pevRxOu9t+fDxy19S67Ml4JleMsGLsyNGyBhUkPu
ctJaj7IWGtF3icyFKdkK0JUBLIwikzDO1VtMBsgijg1XgHuIHAXJCaudLu2bVYctKUFn06K1GBqw
XCR6dI/1E4sO/i/MO+A18j5QrmKKrOgjLM/z3BaaMTm9lOUoq6XgGsSlaWeJo6vjQU66baPs2RQe
eReZpN1b7FsFjoQoPab7BqKRg59PgtE6X5H69TQz4Bc50ULELqFO3BOK+bg3g21DcVfhtO74q1BE
4nwhiMARdLI3hNWTrqZExxaQ3dLH2kMBXg2ppbk26hMm88PdEKnnCXeffGtuuOXrnGx16DHExPSI
j3tQTXA35yUaEIo0bSfO5mg4mzUJW/SjLO0MKYWL7aa8ryOHGWPrGnAERLybIJRWltWOVPSG1VDc
NNyyOe0hjjvNXvfkEkscLn5mdLx2NW92b2V+TUPw+U4vDWsKRLD48a1tgRljn+K4oVWMyKDe4OP4
ihJAPo02NvP6CrCzBCF+D6gMOfrdK5h1ZhP31mq5BEtWiH/FVEvoetTqs+UF0dHKmZRYS9TdwHqH
CjOZ7EWAq7QJqpGNqJBUVAM+bH3tbo8dVicHOIGfaBCaHygTpwLBx5+Co6EF1sIUPNvlHQANfBcv
3LrxTalqQ63o4zGRtoGbP6NkU/WiCHw4OMp8NvCechi4k7TLcNJG9Oi2AjC69HcI1AnkCZ61SVKS
YTIOzka4AnLkrGqI26q6V38ENzTsecx+FQIQnX1mx1dV+C/5N+M0US77OSy3e1NG+ccI/I6nzIEi
0bL/SJsfTn3sMHHmr8sioALPRrVPR3NEgAivkSnz66E0paMuHksdpMUyH0ina9UdAqgWE32EQJlx
SSSIFgOWTNxXg3m9RVWogrp7bxfAtejqURDGuxtdi5G6EcLNKUj6atdlAphHqCS8MtWPVh/+u6Y2
vr3oJTBlDqA0A3+VxxbLpZLqQ6Yn8OTxqlnqwnHm+1va6W05Zw6jrhhyr7le6Zm7uNxo8cjH2Syp
bwUjVC4iD1GlwgA0NWgj9pCHpfOG48EuGDnZ5W7/5X/BhjI6K9NKnsXaN5wlSnPfCqHmHi2Fpkmx
19TuO0763Ln2k+f7g502BLglwt3PVc1jFsVuo5QhK9ao5aAaOlRv4GW14j5tVly4cXPjkfHZkrOa
ImObzRBs1uCwM8dbcY065tuBNP3OKSU8vzb9oAX8ruJ+U+hiZUvfWvqvOVoBpHysNh8/GFDStIwm
xdO7VmrbZhaQm18EF40FKlgq5f9GgBf9B22ZD7qYP6tfZTif5nFzjhL3Do4HQPMhB7xAxyNMDna3
mvQBAi9m6LeDvj6XF6Dy7in+hRwNn+vKg7kqNAv4Yu64o1bk0hkUW8z+N7TtNn1GIaGQNlJEP0my
nNVFxtyI+4ONhpxcMFlDyLXchNTD36B8lntvDBWcDK2YQ6dkO1/GhHmy1DzOee/kIB45m34ARPhk
T+izj89NQg9vc0Oim2jnt8uD5DoueD9S3fS8USiJTwj+mA1fXjthte8i1dtzNW+VprNmAKWHhbw4
VnBDc38p8IbfEY9gR3+6cVG8GeXsejUdQ3GoDi7xnjtVyND+DCNHs+epp+A/Kl4rvCkCtQSPaik0
NYzAw5OewVgqmIb3ex6ALlC+dt1OEnw5lqQLFbORaJgp6XjIctBJNT5awD+6msRvzGGUnVRGcAYL
d6eSB5+xyT8uknpfuxMYdBAwUTWgsFPkN33v+BRxgGvL0b+6rJdQWHDZXk1cHU5HS8P33C98RX8f
LYkGq6Lbw49VwJ053e5hea4h14EfKdj+hLnFawVPmP1gOORuXI9Z+z+eZTDmW8CK/2gABp7egvXE
KR466mgtQR9tJHPRVcSnm+c/Du200KT8xMjPmB8e7jYJXEwu26wBnCgwfan4Gj//GVTYno7J7lsV
+ijRlrngWANpnvtTns6Zgzy96tHtbl8+CBytfaLffwYE+lBxb8eBLdPtvSmJiree1flFfUfVdZF6
poYB0zi+7XSaACfUKx+ZWY6s6JdTNj2sNl+jDdKFWcOReEqDPooG9/Etjh1PeTF+rcjwlOm/+ui7
CSAaz+7yh5PJ7wfbJntYHisPnmlI5svGzzQoTklxXulXM1KNAKeI0/sLWHCA0eafcpYUKyncZGn3
DkJrFAVSHzoWJatzwu9XLx9UpZw5RoNelANrcylRj376Ne6csRX+xxJ+wrJJ6BQh0oD9WV+2V1WH
cy5oFp9RFxvQKWk9WMqclRmukhkA+X4zrLQl1DQQytPH1dBELswwCRDsPn39RrBrrD8KMj5trFYZ
MRUptkW9XwSAg5omPqU7RPQ6ugzbbbIjNVIpGsrR4Ng0GvugfDJ4zTBawxtyZcOhdMkYvGaS4Xy8
d2guA/LY59r3I+ljkryCLRqNY9Ee2XsnToLs6Ys6PBopz0N1KkglmLiG6d8fcPfWRj3/uPpT3Pns
r908XCgk2AQ9gJvyGltym0Jotoh79g0X2rFe0XOhF+x++i8W0eeDt8l6eSVWE/YeOgADOdc2OGz3
EpdPqGaUPEndef8x8IxUb+sIoJ4P0/jFjwW/4+3Pndxae7Eea374x0QNaJopWBJ4Mn6dzF6Op7/D
xSWqqdQnFn/hlZbeqrZPnztBqvC4EYrVnu+MFZ1FW4KuV3JNBOiKhSIa9EQMNPvqVJ7m7SeZOn+L
4lE7Z21wUjA5YTRObQ3kzEm3FKIo1WwjzI+0wE5ReeRzufIRK313Ji+JkigCHPixfkrd9mAQ9OZl
Bjin2stpZo5eIW1n0ii1qyxb9e11n/nfgyYRYgQoQS0nCxZihpoXIzhBnu6TBHBY0uH/MpKoW188
0G/1h2xjoLZ6jdWB4czyWzw0u5UzAALFHXYaXw8IvIS+UxZN53H/bZYDg0+ScQPj1193w7CTdv0p
2H3+w1/R/bqWtvtJgN1bB/lDbzKyPD0RIY4ginQO01eUVJcbXFSkygF0y4BfmaxL76VdIEyphDmd
gzFS/QCwNkNmIdBTDpZqZaAdM7nOEkcag4xptdKnCrW+6xj8yQUdzuMrbsfZUtEK/JRzq9kj4mwZ
ki2SU4sVbaswgYYFYtK6Y6doKOfSfN0LPlrm1aPwoplKk79DlzsEM4/NmfWZojF4eDMnQvq0U1Mw
cy2lrQ/O4KkeSOpppoKSiURnIgtCANUYOcqOlBpUPiKuqUYlA5mu3yX595y1Q3rhvwG+zSEMdrww
sPUPXzzpyd4HI4Cry4jE25ASM3zk1/O2nK/a7b/PjS+3fjCE42uZLkegnj3/CHa3DfP7ExwRI/HG
fe3+rmYJgBsBS4TCIzzdji7fLz3JsEAE7TedKsSTXxeVHScpBNWboMDMkVkLhkUdDj17EjsqTGJL
ZEtY1pliKit5LxemF8P8Chhx22kCTrT3H6Rp7NqiB4V1yK/PccZMUkopWaX9AUHAORxKxqqDOkR+
VNR01+XoHwHQ1lUcKQwJPEZjD4LBJ5nJqhnWYOJJBiFBhzwcvkf/2nVXJJZzV4PmFEyHQ4CVPOuP
f+tlE2U4XP5B+HN/VEV3OHefdhkSHA28jdd3AbF8XqKQ+FSAPA96g+hxmfcElO5VVCVAMdfNZS+H
PPBFRqGS2kMr5t8Oeick+UMqq5uWzawf3clceXI/LI2uSwZWiJqqXcMSKTWhNcfSTs0ck8AtTEA6
GHDA7bJexG7bf99t9nCs1s/4w4mTz6fIqvrGQqK4IID4Rvr0hGzFner6fgO0WIggRKJbMObMIrCL
71Buh23mSjnEJJbeTAFtAzKeL10yTU2uCHKU5HeZYF0RFDB4PNtYMQESGM/T8d7IQcl1rGoxiWRe
M/OzjBno8D7AF+X25YF9B/sOTZ1DXDtZtZoQnlvCmcyxwjAESudRXd5kyuHWbnC5MJwJOxcFrHgx
lB2tb1Ue7xPJ1tpgLR3+xUemNWnw3zqfQIxtuqPi6yAh7gqp1g6HQb7DiHjkBWxq+O59/zw9WGRd
xcO05845A2Sol72dSLEBQhbz6qCGZSGvKbYxVwYGdt24C1LA6iSwWbworiBJZOSyk/qMDyXlkcNO
VOpMkOz1dgiPfn1nxKcKqnUrqZqvxBiZnESOfQoAn5PQ4j2kqe9CAsg2TQItsdokY6UszMmJWCuq
jpaDfZln/vAU4ap8VZeThM5aijDrGGozl2wFIYXoxmtFY7KNakjZb5Y9kxOdwrISPPEnJZ4VFzO9
4bsqQEbwBLmFoQm/oCtZpoLMbk8wM6XGKgo0aoLuChN1UOFum6XpgBPi9Jt1qa0DL1DE946LHDNf
f7R5Zzln3Z4KI3G7Fs+1fr4T9JBBo/Bsnl9mRZ4OJMel06mUYkDQUUK9ZBcvmi7O+dhh8rjRsZRB
9Uz+lRMYw6LPwTsdRjXtEOGLwEOtEYn1RF1QbDSDSaAz0AtIXrvQ0mb+5gvXevyhnl8J4boKrDPF
KDtnnB3DzvnIE1B7hj7dbBpoC1HWA02L0CafYQqmAMLCx8H3oWckdBrJ2LOEbHzCKFGxX6WZI0af
laZIvrMcZzH7W/j+JOfV392B0mDBlE9Pc5zq5CMGJDrI8gR5SFI9Qv+MOakC51CfNnqCSFcedgbs
gyHOq1d/PE/hZM2Xn1x7ym+HwQllPe2L021ZDmwN/ut9yE9KuNYR0JYTS1atNTlNFBMYu89c6Tck
NrvBKECJq/Sox583yXGpnleXmFycg02IaVRD/h9nC8gzmy0b6Rd37IRPgkLJsDfideztXMQBqK96
Arj+pGuybe+dTCqrM3wSwf0pwsGfyVJUHQwPS19v5VOGUDBAnngH6lJcS3aGQgBU5Dt4j0d8XgqF
Vsr8ruZniowOBJpMbVVqYZTR2QsK4fysiOxhT4Rilb6lW2lCt9XM5/qNx0+crfFCoEsg98ag0DuX
sHbCpxEZKE8mcRno0TbTlc0O8D5PoNXRe6QsuJ3oE8px2iMUsleZp3w7IjM0Z7WT62pf569qDUvr
fA+xZQtIiOiMSjCSjtRN/cmX+KthQ4ssCc29Oe+QBd564vTXVJWAt5+MWCxaTn32hE5ogavETGf5
Vw3m/AyAqhp5ziNfAGHaxMTc/Ou4E4zlmCRxqGRVo2XRsHN4PQpPElfXCwYxACO9Yr+s5diYZz1I
P771xThFWIB7YUWJHaCj6GC//d7IopXi6v3MawsOr5lq9jjszeeOP3yXsRK22meBKCThGJ9tosPH
pUbWHVG2/u0iFnwo0qj3MAwbVKIoMYjlfHyj0NtT2IodSZaZoinIK3Ur8dd9c1loeAMb7ny6Kz0A
Qkfe98Qd5AjxGii1SLOS438mz8I7PyeWGwdEbF2ENZBsXxoAiVbELEc9G+ffrznBnTdNvUa+y9UK
ajObJx+p50xs2YJ2Nck2BrHa60BtCZJXaHWLmHmMdO+vFfFOiCCI2n36M3lkABPFXnxgUYBjhuuW
kOPhUzc6HqPKRp7x3kdyzDkAkCprcexlY8cSS6GCBB1u0vwtTLOuhP02EwkztiAlmklR5e8vAYzS
ubjCmGHNprrDuiCRQZk/uGNYdakcrRIRYosC4rE0Zxrsp6h39HCgaDpB+VtkkpjK0iuHdGhybe5P
WXKrxKlCHaQ0Z7zogsj8L3vFO3GYkZ/rzuSHt3gGi1bRzu++75FttwDvjxTEnSZvA78VXteGEoSs
/ctv5gxNQbexTzT0eeoLcqNjrm8bshCP6aMHWyEZTiKk+h9jbhQmaU2vsZW7BHeGeDquRlEgSbtn
/ZCWMVn9a7758ITUVSmPhBXqPKSn44QFtORFXo1ctQsBddDQliRz+mR6kgKHv/BscfciSWdoGcwg
85Sm0tb8VJfW/neuU+XggPLzXR5JEbeASFABaubWMBqjt6taEjvLE0QxUtkT+zl8IeBmSRELtb6Q
jS9iZwbPcfT9Y96wvd/c1R8yOXF4fTfKlZYC0PLWxwQuZXUSgPPcUUb/aKrwobkhKgVmYM8Cs3jS
jFSeHiPd8mJgyIbwC8l/iQn0HD8EGTibUE2d555BE4MurnV9XJETzjqXohP1Ikj23PDZbGwmqPKI
Xaaaxmy0h53q7s7ebj03mSgTXQlAJtvI4ksvWygbKfLv8a/zPcnO/99OTFnNEMJBxt7gC2LwwK/3
K2Sdpq1ILtsM3JVD6ZTg6RndJy2Y9wSul7VqtIVMrTjd+wqhO7LgnAvUCfXBpRO3kM4uc26ql0kE
zkSfpVkShnwu18xVSws5Z8DfeOq5nXFuQghBdicwPTJ6DudLShLxxXzgUN7pV3tExHlJyAucbWdE
MV8k/Mn17bhzhXaJMZgRu3shium0vKOzppEIXs6yn3I6cvLJUG1dzfIyxQzbLlZnERIL7dFm7DV4
hRYIDihRPvlO08XYG/Xx0ORqYzCfCVivSdOj3HZa/rFBo3IthodULrAuPnyXctfAz13DHG2WRww+
fRFtvxOUHrW72dAogdzv7SE4ZaZsH+ju18N5CddwBrbZHdYjMYM4ACgJHdCPPOmqgDafLOntxN0N
JSzjPDgHAPf0huMr7aGBS7MW1zwG0w52FNo+L4Pe1paX5s/Uw0cnI9WsM+otzXReuuoTVjj9SPiI
XEdE9lM62au9DXWXOXy87zWmp/EY+eU8TWZPQeu0TGIUslQApQp/MsqfL2o2+eTtYECpOp5BXSQD
gCL3uw/Z971T9dDAWwlrpAyfKcQAzFJ10VjQdoTTNJwBmGpwViIm3OVK1iR++v7kLpMLT3GFX1gk
PbdtTS5MXq0bmlYI6L9O6G+B3yDYQE+eM+1sYfbF1K+72f35Ccjio1+TQW7ouFVqgOwzP6BJujTK
Z+G5FpJr45e2P2dTEKs2EHoLFrWQokKy0psM6FBOyFoF9CNR2YvGg05I/XpGO5tP93XFrCGJsVl0
ryKZzAFbhy/zMA0mQ2MiL2bXjPKw+75WeM4VoWMXkpTilo/VHg2I7sRuAceX/q2NtgHnVdkSxSRD
bD/FN1mlrgw+SzeQmUVc9XlK6sBIiRM2kXtqNgHV7HbbHqNCZFzPrddsU3Q3RdtLxb7gZM/sLIpo
S5DaPht0jn8AQ0ukFpwlZ0UXoa8OALzV6KR3cMwe8DcvPylx5hPLO/FdUh5bwxjLEMC/f6TlwvZT
hxENWn21+JwLJ5blfAmfGr5B95le5SnmTGu8pFZNhmzIPYGqZzn+Vlvu1r3MKqydy3UdM7/3iJ5q
FHrxhQDEDWelJr1H6sW5ANWSp+mhlhG3NJeNdo0M1r33+KHnB+GcF3RHgmpTuvHxn9HfPFPdYWqH
GTAkjnC0r8Neb8Rmyz3IhByCgHWkJC2VpjU1QuFbuYTie6FdM8O+ZiO5o1ou0JhJK8c79Zsq/ZDe
7rSOsxtHCoyBKW2vCYqmsxm6GEbgOdh+FRNrucfZn9rKtLsENHSS9ZSs99OGFE9bLnwiltfADCgn
G4NoCWMI6tP5+BInp9rvUf03o1Ky6mtk10K/StP7SVBXrG6BRoYg5ajYbsKCOGE0uoBb2NRv5Grn
16PEXdDXXVam2CdoID7NpDGHOdbwmAR2w988zyJOltYIo/ksmD+5qLQWO0SixRoG0xR5toTPwamd
ThPoRuUbY7TlUbT9EdZARDEA/eJkveqtKlbnRQ/m9qfpmh9pDzykdOasurxZ0zWEUbD1YUUDdgjo
3+oIB+smqjQkSOseIvnQIbitax48xR4OlmjLFwQ2LJ1Nx8VRFTMF5KfR/fn81R6ZcP9/mbZS7HJc
F9NR/YQtWQw1bI4Fy1r4Qu1djJBSS8lsjgDEulsb+W9seO8/rp4x5acQmPgaCESKEX2O+U7H2kHc
HjJOugj+Z8oN7xlSUoxHuYU59Z+0fteC+8Ay25tFjBpHZKUBpkyMUWRlGSo5eiVKvYS3CYvNgTl0
S9OLOGrd0vZQgfByIm4rewKyzgv2Vki8mopqYEUNDJaCjJ/uKemA0pEIAgZrjMhNTNB9nbJnwHnC
c6eybt7Eff9patSvuFWgKcOsjxEyuKvwOf+Y4tTNMC9ql7LgII35KVWPZKn479Qrup2cxFjwNf4U
VrYQX6V+QYwH9NKxKBnC+J2/VV2uvo5MyOJDSBa/S4Kps6dsrViUbBbLYa5hjQkUiHG92KeMLVJ0
pM8u+EvFecpwqAtd94AtoFPGggnpTdtZXfzE2eUSsEpAYr+zpgM4z9KvmKBOZMkKxSUBluZATSJk
UkAns5xH1C0ckg6nK/84tgBQrdrfkKdvxN43xZVCXwrHqmF+5fV0kPiWujd+gMwIeydhJTKpHMZf
aMDx96hNkUmrLydLQi7L2v1bvxTD9SGZkP4YFmHzoGc6+ORm/HPSY8Agk/TGnd4G4aglMy55afaV
c9q86fxKk4jJB10fOw8dZfEJcdDZNsXDn6ZlS/XaN7+9uH0lEaJyuENKPjeVwL0SOnh7va8nAjs6
1pq8e6NSGntSOkPqAsTq0U7IWBP49bRB6hgwpRN0oEfFFBziJLfMM+5DKXvahqf39jRROximnBq5
RVeT/cKjN92naUwRojIrDPD6B9KacClvjdnj3Lq6HcxLKeVgwnunX9VlA7NKZFo1UtGHSf1EnLPf
+wdOh8lO32fE+vg/tEcBOmAVeFAlgSEA7M/aK5X56r0lSt1TvtycY9LRlRYphdNxNUCXKqxLMHUM
S1KnlbwZk4fQGYT6hb8Z6PrLL4FW6ELtGn5Pl1i7W5JSgjhLkoBkXgO+lOYPqrRM7u0w0tLgdfW8
DfY4OEUxWoduVCfEIWvSES9R9oWK0Y8x0TGXx/agcpCqpHtHEtesjrrghj8RMch9fBEcqBB9vuVp
AzE7ggIFjNxT8z2nzYCiSwpGqKxIGme928+8dDFDf+ZQ8xlsuWArxuVzG9xaHWyquE9pRJZcsit/
atbZcHfDKGFcTqDCbDZZ0m+qQnivcPJHQPV1JBrXgo9ahL3+PXKk6k2zFyZ1Y92WFxNpkOu21dcI
Tuq9c/t4cnyaKOB9Y4NxdyORdlCNT0OMo09W1uMM8CcZz9uMWOpro9Ia8HZHGjfzB5IaPCWYEy3B
zhzMDFHTkhCA7aP0kQPdPNbksPILd6FcoW7lcZJCp26JjYr8m37mMKo/N9FIPRJPOeZDP+C8DWSI
hePKhCHpldKRNJRmVWFa34u059aAAz4/Ia3qmtD5FAWV7gX9J69oe2ZPTVoErDwKmUiuz88DXu5Q
JJkbFoR+l2YkrwzfGWgFC05TwMSamXDkT5iNm3dovj6gCnwWV9VFrB7UBM4tCVuZUXmcxAWkkjyF
AB/cZcY+W8L2XQPyWtOPrQVhakLspwV+TxnCqKBaKO7el6voik9gN7vUaG2GPhLY9aRlzk1Vf9jp
ZVE3VoJboUKM7gaI5sd9gu6GG0hbKCEDEHQ1n+H+4yHQmsrzwPpfu232JeSLOP6YacXGycaHR4y/
mdfURNxbddoBUcs7Lva+Ayh+F4WWEL3NUlHq7CCDuwt41NpYapnQn3TPZ8GR3NFjfRemMaYYBxjT
NoqZkzYRqizxDPnWkuKtmgkzOXPxw/CdRzBDCRTWRPWKwXtYVmKr40X5e6Yck/8opohF9RilZuuP
JosJ9LSiJ1tOgk/tNW9WhCs04/6XWMSJbVNgwaFhg2+O4gecTASeN5AgxMde1/pScxN+NEsNZKdI
FUC1uW0bIabDpkibAh4Zgc/O1sbePv1E/HQ2tuTabsyc0MQsU5Q/rW2Z/yLqiWKq/nNRKAHW1lIy
JSDzNiGKCY0ZBPLC3Y8SGAq1Le8TDr2oCzljl4NH9cUFL+Os2nPqZZhPUMZppC4fnUmkgnm7AcB9
oWKwPwKGmuWDPaLPUr6Hy9ZtumymWBP5mFoJTA7q6El9+7RQhknAtw1WppTPPIV9LvB2hORW49AM
3YaygGmBWyzNmMunUdS3VmxSSFKsYipK9qAilji6lPMYNSTt/t/pcvxBz5o7wYw3FFilgagdpdOi
0Lno5PQ0hB+1KWPZKXOReT3O9Gr99TYQQ6HLoD9olA1CeC9RqABrhkZCm+oDT8KRpteBL8atcYUF
TtPRrcIodyhUFvmAI4+U6zYJkVUb2r5X3P7G0eA78mKZh8tecTsdYneuVh30vaybY40aqPOuWnIT
jlq/Ff0Vhm0CwvAjKlgeF9DJUKSk4bwjGmnBUygqc5Yoai20q1VkgVb85+ygFcBOPr9vH2OaOyRd
iHCGzjd0hyb6O7s4bSx9ylI2Co9/RePqTzhY1Y77GryNxFJMm0ROT1FcdVhVwX+ZeNulA9fWkL7f
Sumhg5nuWpEylrO4MiCrdgc/J+k4FeKPzbVtZKUVZgiFI8fI1pAR3dvGpb0GNlTIAPaljn6nEWtx
MSZwfxPkAGRN60/HCg55QZV4qWsX7GOlaulFTWSAsA5Uz3urytF5EyZJy/aBpJFCRkHUyiX8hd/K
M/76dYzzG11ltjpTDaEdK40h8g8+qt5X8eLW6B+TvNW/rd0Pq1M2zwuEiFHqeVWri/28ppDLmsQQ
80IASjZFg+ohP8n4ipTUbVkEin4yv1srqqOeN2twFZA3ADAdLGjp1pik9X5Hk2BZoNVuErua4qxN
LlkMN9IDE83SVVwRnB+sgxIQTz0c9CqYzu5IhkDaGPnRYNlbhE8VCFTYiTY2zfcN4mvVbcvuWqSN
OrKWOl7XkMjX+GbcTN1s23zsm6SoeEMnGh2us8fx0hxANT9B7ktTWiV7sp4K5Wr8RfPRPZqjGjYM
AbFVG9qkmJm0m5wDKL5S2tKedGk1BLDlQbD1xpUiOOXraZazA+p8Y63b68HRheaGTmcH+iJB98gp
NMZ4shsNFNHeGUpLfgMjGBvkbXQtOifBuRSMCT8p0vyQBLQJpd5HNAwgEwWLgSbH4++jC1RwXug0
1XQKJ8M5D6+0wNryftixmn/fDMsYgeLeV+aBGYQL9n/fEVwcKviN6QnBiC/khOOLjok8mfPkYNuC
Q7+yjYX17CdwL8JTNlvWLE3U0tb0QquhacxbCBqlGfsWMRP4WIxBXFgonYlSE6xJEwynREvJ1riO
dHLNbifXzsRQd8RNWBNZDn2wJ1QuXQuEURGW24KxQKRhJ8Lxua8LdtInU8Gfs8fn5/HN/PKjhBJO
sSDrpG+ywQGFIah+1BoYQUmbQC7/gC4p8SzITT4niyYs+OdnEc8zWTIA2nUkthpCND5P0qy4cK+R
82K44qbbS2OjIJzgtAEgHL0cRwVdsA39wG2yN/ee3yGiuVUpSBNiiZNDM/KD945JAq61tUlZFCMp
ThzttHtLhvhanJ28BBiUisLc6mUk0Ahdsxyl7RgeElgZ1/JF3qjK+KfJcG1cUo/OhijlVufzF3x3
s3qsYVQfVXAWfzAA0CuRiA4nGxBBfcMFO5bGVXw2l4crBntwxezZkUmG7KFQtrsuJWSb8crGGb7U
XIzxKHCkcUHMT2GhLv2UYK9RCGwnqZqDO6pZb1vpqRkr0vwyvxf3gcWTPSZaa2oVXHlTjZbOsgAL
O2SVoES4isAMHPMOCT+MNX++imbITFFBgkQCE74jPwchrn2Dz4UDdLUKHvrCsb+AVoTxJo9lAG3m
Y1t1AYR+5TvvVOFMKbOVFbN1peaazmvGKl06G/haneuToS0b+UYR1krJX5o6wGoN85X5IPCpx5gY
fxi0iwsZIlYWKGeePlSCVVO77PDOXMxV8OcQR3/nKx82HUzUAM2QIw+HTkzSqFsBnzxKh9MXfX3k
h+qxey1jw9sbaEnbyL2jiAvX9C2F8zl4aP9V4p1Vvs6PademLSOw6KAQyK/4fBaol3uK+71ufHi3
cyi2Th0K3B04kiFNlssAOauETo6KwtOOEY/5dsjQDydR6S+lrxjEqCCgSXgWQyKopX2Nj7EQLy7/
Hp0qg7wG3NYaLHyWPgbrIFqcE0uVTHqa7LA05uMba6ZGKN3LHAIwjif+JUQc7UdMYtjMyplEh022
2y7L3IkS/6d2VTI9yZpUM8m9BS37UHRUKW6bmjuMty6GIRpjf+equlh5AWcK1VCTHsZZtbI1Vb05
viDSzLCnqRJdT2WlNMQSl4xCrFif1TvUmz1WmBGo7mknH1wKNrsPy0yqcEgBpcbsuFMhp6CVYdht
HeSTg0JTqQsieYj6OhOmMwYnC/UIj7IZFbmDpwfH6hVDxJG8aR3nlQbl4axW4xi5q4+0aSrmc4zD
eh77KYLz46n8gm4+gTzIPuJpbRLpxO59VDWuO5s3siSjEdP2DT2l5h/62zQvi7HjDYw1yu5P+Ocq
iRSWEmubMl0LVCKFcQqKTgT3EmB3AWGdHltjrYj5hG2IZo6wgP1MZE/BKq3i4JOYU9mPpCf0tvwX
NooGRFo+W3ERwUU/BwKN7UwO4vO77l2eerJ/4OgpVdIKOCNbUEheZAejCHF7effNpUoRR+0xYnVw
8WWqM8Hi5plH60NFSzkFsO3i/CAKETiFCe3LRkUqrmVQSDyO+NZXSE/eIUzRGbf3NZur94DZLpIt
EARIG2nF9Z1vjegqCqgCHq3UNnzqfrmcX5cOrGjUw+O21jLrDOjHpq6XW/707juIB1wa9Kx1J5DQ
OVQ5kgSVbBtg5dXakOdWE07rjkKzWWskxUsmP/R4D4PpuWLZeWtMy5lea2RerQKM88SCohSIixiu
d+6dd86/ZFV9RDz/ksDLw07MdnXZtBScnLmULbrdlb0WFQuhWR3H2o8U/nMDzwQ3VEOWBteUynZc
bhfPi1hXImGaeHMR6AimVLP0YywdTpl8CyA2oWrj7/TUKB2AgoVXR2/1V0HgQPyJI5sD77A4uK/p
WM0lBvjCVsrrZsSWGhRk/yiGHKh0fnBJ/d/Bo7oB4NdXXef/ToYDtjeanBBbLdKA+2CbLC7eX4tE
6LvfN20WDoF0k6oLIyvpEAAnw8ZTWfqjnxzhxEdSkrSJg3kvBiA+dv+Zp83wU/mw+F0nrYP4QKkY
6485AcOaQE0RvATfzPPu+/992b4ywsN7f4l2O+/tbN9vllmP97k3FrlsVyxVThdebjmra9ebG0VV
S4bDHy0AWfFcV5Sv8pHoM6R+l58JX5HkD/dyHJF8EF1FmFn/7JgxmuottF5hz6dBHk0z9OnU9L9y
q2BKHfjbbJn7IE0tCfDnpjlRYXuCJuZDjxb4OIGD/3H8ZfbKoqr0l0VWyBxp4Ja8WS4ozRufbnRr
tyAp6n7v/nTdVFHiz0qmBW5473xcgDKHexXIqUPNzlj+p1oDi8Evw4tJrgYIlanLV6PXvlUxdQXO
f3hRhX9LmDiouP4jHfzjKSXAkWwcWd+zDaCoXYwwlH+VEQi6pGJKCBTqpnnsWevv4NWb4AVFp+IY
eqe7Ele02qQ+QS+GeXmPT53+W1y8pmU3tO9PZxkl6l0QihiKKFisMWnwqdteEj2wM4agE2bScfjD
Kh7L2zdR7OUWX3JnPOcYVL9JSWvwr6Ev5+BR4BNUJnl6kNorzb/kkNdkobMxUVf+pZXNLb02ue/m
zAPMBq5Expwsjehrjfy9xY8CVYvTtfJ83DXKFcSviAxEgXixiV+GaJ+UlADqw7ICdE1I3DBwQ+TF
JQyVu4wIhQiwv9kOtSMTKRxIRThxlaf/BONVfmmMiNEyjL8JuZGZQiByYWdcOc1yYC7c5nKtJceg
sgxjv4l08Tdvhaaj1v9mHSe2yek6HPKgDbOBzZZYUsGlEbkLsS2cdk0ZmUtuLpQPSfq2S7GSAaXT
t7NqMd/eeKdUvzWghlanV7uJg2R1cyxysUcDZ9lE5m4lQh5J39HEZhE+63l7U0lzfYIFIWmvYaXn
9Bw8IlVNKqEakbARZ3SFkF/efQhIxcxtT00PBuhiXjCWTwonFSfTDjadeIZ3MwPwMSW5aFRmlNgP
tIpRN7eFWYyDMk73nKl3azUGC/TEuFK2I4QG3Tmnun+4wJ5oRdWBIgAE534FAw7T8I3VHVnPwgev
bkIlZhQOKTDJaTpbOKtP9ldJwoC7ooob2jqFTXJeYkVfkJ3oaMJ7fFV0hWx+5mq/9n7eRmcZZp2G
59jC/n6AdZNehofQuOT1CxWqu1bnrKBN/Qs+kqNdGnNHEqMpN3DFZq062fCoKNGVOzrbz6t/IX6U
Oh3Tm9hQufUMwLCFGbeBEVwcqCLHpLU8bbq8TQO0k8CQGNRTSKv2/ZAmmn9TM+CiytVb4v8n8dZg
cV2Al8sGKAWMrreeFfxRyx5xI80qkXjoDaja139Kx72zlnNNJumTL0bb2yleWl4OZCxVRSX9bYze
A2Y6/XsJ6ljRWLRfQX61uK1lrkL6OskrymIXcTO1HDBluzz+20IAcGEhbcIPL98EXIPVBhhlC1w6
9Fjz/j/ZwwuOKop+BY2G4n18RihRDuzeq/HntJlkwYJvcSdHlTXOY8pnUNT5VKIfKB4P8iNL8o7N
32IunHjyyk3OgFropkZ6WYOVPfplkUfClIV4vPmqTXYL7Lu6AlcCokBU2jeFHsRVnyvJx42naWN3
rA7njn5Nub1Esz+28s0pYY+HBd9d+JakflZO810zklqdA6W+sLvz+DY2x1CP/56V1Aug26d2yHNB
8Yv7qcWOtHbPM9D/j1Vpu8EOInseR0JpmYD8ERKdNThsU77+h8AVdr/tRfpxH9PsmPVGrLaBigK+
vgH4GukDisTa4YowIJ96sePd7/JoNJx0JZUGO22CiFGpxO5z1J1LHORjrmgntK3qR5kBjun2TUyj
9OWz8dFt9UMvFz8qksJr4Uwgc9xJNrqQrEpt0og9PpfQic6cogRrdM2dWjaM8w4+RvPMyo4waY+W
wO7rIkB1WBUhR8svzEOCtx5SZFKGP+zbtgxqjjBD7/lvUYzs6Ajr7A6y830mxkVrDCr//bxPzl6Q
OYlP6jKl309KlrUeUAnhCwL+Ol8W6YjssqTwcLFwVQjx8VZaTKSpv0ireQZ8jKjp+q7sdxKA9hAb
evqGtzhgYNoxL75PMa908qYEZp9zlS3WmVGqPqaohYoWPJ0yQphX/4yZDkWKC4RW9LcjAYdVSwuN
HTF9Z1IHqA2w9Ed74QJcWY4CrlXeVVoFBmNy2eQY0gKKhDuh8ReN5l80OOJbRoxrnDPYGB3txp5g
k7qGl8kU3rU4xrLEy8CYr8zJ9RVvSzYIE5idpg0svmgX9J8Tw8mzb9OPkKQZM4Q3BReKcuBNQb4Q
WeMZBd2b74azq9Xl5oafbE9FPek0P8g61+PhRjfMvz4AoIRTdqs4U6mSMu0Z5+gXHC2Pv+S2HydT
p+dXHykpAKK+wI3l2AH27X3iqZR5fuGFzSYMSubN3dlZXZ6wLfWiYetrVOcilwkhJhDqkNCHmzq6
V8551A3jfljYFWcd90tXJF9jfFCZDwQAwtqZH3HYR2/sZCgxMB2lO80PaJUJRdEsrAE4hf4DiMRw
Txp0pubfnjp6zjY4gAfEYAqxHJJUaYTPIdtgkvYcPHrqW0VdrVOiMgZHPaCFS9PE1s8xIvevgH0v
Af7mMCPiCOykGeLregVV0DW8cycC74SQlNMoDewnwmjTCCM3VWmrz6CQ6+NSp/zXoZxlRb5ufR//
aPMY99ZwxfbTyL4rSJ7zAu5s6KeGXbeelZ1BiRqQkdQ7EJ33oBsQ8oGbsvZA5GIQrxl186vLNyUp
ljIG2QS+5JReQYk3nwivOjyC6rDrRivF2gmeDVDIsZ5Cp1ICfG0AKrXjIeHEV3vg3zQ612j/CJop
oHpUGkEF+TsQflDpCyZdPYvr3b9Eu45yEFZRFVjfzqj07wrQSfVu4ZUoydvkBObJU/BeJa1pLc+c
TOPTQs4HUR2+45JdxViEOLN9rhpQvzMGmT3hxZgwzwvkQmBjPDWKEcojM6EO5IfTiniqr7ufSayj
V+sDESzqTKQCwwaDGwx5wUrTKxhZNhIZZdyEt/hZwu16ayXOro+WarN1GaGedKa85qmwr2ZU5hh3
9W9ESNtsRBOtVgGoYf/FKdi+WS/WnyDJrNKbtGoOZQxliWYyUp0r7i/5Db8xmSEJG2ecU4uITAaH
87UlAK+XdYBWUuzvqzcra9jAFr2irlRcD9yaidsdoi0ivkwUUb7ktpuMoTBttxQx9FmYLuULcBM1
EnlOcKUBYmaOhH9x8H9vq5vLpIrGF6J83r4knBvDK6F9ELO9YG7SJbj4en1HPXA5CnVOUxuka/vp
Sci1kH2W5Imn27FI77IsXUvwkQo/hsoebsQSWKozAqMWIRikVkYDs3wZoy3M7PV2t8UOMCVhKek7
k2trqSPYKl8ryPBvibyFZV8riXAWRZQU36FQKMvWZO8RhZtpIaQKVoa7VTxfsQ2AjsThEzsOy7gj
zqjjhumizncQcc8LkRtVLd+DT8tH6ZDODvImP89l7DJO6TQ7ppnCtiSs8DaESHI3cQv8bvNYPo91
9gw8YIXpjWLOXJgJ7jIibo9wIYvJDuXwrH2K3uz/Bcb8WWXChSLZjERpm2c9LXNsWfjVH0xw36FD
WTUnJnhpPqN3cOnDVFhkIZr60JIKYh2FCJ5I7GvYegCubrV74yI3YJNzRtOTA39v7D4ypgyikhqR
Qw0r0QLzFPIjpwHqX62NqhzBXAbUtYl4sRmJUYutr0XeYhhPg1KVnQme2cTnussn3yNRRO+4duX6
/z1oPG7snIMm2QgqKJVXt90oZcDbSRVJPewfNs9ufCu6gljLlEZk6wymCnzpuObi229fYpAqSoIp
ldhlNxhFDsDKZwsyeCAQqka1GnEtYOaTUea/cl5erFZm/+1yGm4jCy329OXSPYTiFgNzKdK8Txus
gLPLv8eXetodLzBS1IM5BqXYEuJP2/KyZPppHR42nzuWZ3x4AaAbgAWzRg63Z9J2bOzOrIe1nqW2
CzdurMhe7HgjxRCHTdUIqGg7RgSWyT2wbTGiPsaGuviaTx1M0vyRgP+8QrYYd/8Rc/rdO814lrLI
3dw27YHhG0i0q0MoLKTGb5Jbpax0Z+E5lPUWwQsWGSJhkZ50RNyVX1SV/D2Vw9VI06ylyCcAuKls
x/gB7MGHustOSMsdqz2NYbDxVPkxk0qDZqpMRv+l0D/uWRd+sRqHMDzSwbmjd0Lw+m/Enl9DqBbd
wdVRnnVCXGKQq7Lu4nRApGTUlQr+JLX643Y5ki6Wom7MHmk2N1h/jhrpeLNhtaY66xFNrYQGAZjO
d2GyecAW2bxvsjWcZ2fZ8VNnlM5xY7Wx76MVdTWLICmwEryLpz5ELlmiTV4XZozwKXwyAK7WdEAU
pX6nbCCi8hqPOcnKy/rv7HpiX/hdb+6KWwYPGULqc1/ToCIk5iU4RTjMGab/WusTLhtumXLoBd5S
CTg8fK/d5JxzGYyGvMcvsKmvkNPaQMU3bpj9jkgw7KQmjiexvgII8EuLWOsxXOD9/hacp//8YCex
yXLqQ6ppL7b4BmJjBi72yOIu8syH/hFj+e9VHLupWaff2cGPDTwmFay6r+KeLWay/im4cq0ZVDXd
v4c0lTPyvUgD13RXkVQtH9FP4rzv9TXnDjF1tf1TA2H6yoZOOAAMi2DM9IwpIa0yywQOri3T7CD/
2JE1yBjz36F5Zl9ZU0z+Ig0rF2kuR5QhUgiKdNutPftE65tZObNHzgEDuz7h4EcyRYb5nltRHVyS
u6Vm17fcDdYQeYw94RcmBw6cIHDvamoqYjMHWkgXUgFapfeMFQo3DizKvwviUDU5j/zT9YJDsJMi
Yuq0nR7gYXvFi9dGTdIdiS5LYs562pqGw3jBrtXyf6C7OJUjrkwb15xEP7b3xcFQo6aV13kjewyh
fZxi3vNdU2efb2RH1REZUYsIj9xxxp9m+LKvDO3RfOpX7XSZ25jacfb3BCjpPN0NxIVvJbvVM/Cb
zMB3DZLzMmnzK2/NCjwv0ctSXdBSi6grPj3ni44OqqApjWfqOTtCmn78FGyWGCqEqP9gE8jFc+mr
mUUGh5f+EyrX2eXvSZDMczrq3SusJgW4DGJkiS4DnJGi8XvBbIko0LFfFeTIcVZB6UrpEW7NxXTt
iQ/1rT12uHppZqPeHV/7QIFBlZBewwCCDJghhM65PU9OCvNh7GyAmW6w3cb27Z6Ilskq2XWwUYWJ
sWwXQv34m6Yv+bLB2gMZKF1o3GRpaXy61DaaCNBWiC95cmcpxxbCN6G5vS709eMtdE55iFhJqymi
nk1zrZsZqpp2PUri8GBc2TC6j3ENmJXhkRrP6WPNMY1GmsODrVGLVXUot25TSGtw0705xunGnC4L
oD5vKkgq4Ao0JEhTmGVG27nK9ARpdJK+m1DkrYqxAfZuSsjZTM8maRz6BSV9eX/Cv/fN0KntLCsH
lngWk8XyiaT2uROJxK6eVwTPqCg4Zj1c5WMJw2Gaj6nXPlFSZPOYmltO6G0T/k1FZoLxo0IEuGxl
gD2BYt5kKLNcFI+s34HYWYHFEzNliZiAcgcSUs3xfYm+SDxP3p5JI1VFQpFIH4IbaX5jZBFJloK1
LZYMA7ds+HH1sxHO+YgMOMyM5Fp1soMxrosUTvOn3+FUSlcBHgYH8hQvYj6nbi44iCbMUaQIkf9s
TEBzoJkIZ2pfHLlvznh7t+k1BZo8TqEk+p4UnpJLmiSOa3hmB2g/EQop/ayTOF6dOMgfEeHFLj9d
PCywGTo3yhiCnH2dPvDf9rgAhs/dWADugD12+lj9oZXQ+pVxvQyal/wvTZPd9yBpqj8w7+fwACaQ
QmKCgJfEzmqOfv1De9t5MdgvIEiXkUmCuMV9Mf9jRO2V27GW5bKJRjdR7+Qb3zrKsd//3ztfvmOz
fYraVdP75LAAuotToaDrxRFf+KUZwLBVPPtMRVh3kbxIVxHUkzKmQOMrYJnlVsw9nxTtfGOHAk6c
29ANyNtwgfDJmvHH2PbyKRISJpPy1J0FgAEWYpJz3NY/5lytjQsgxUohxQlGS4oeUQEM5zxIJBrk
Qxs9porIX3Ddtbstru7QZ8zyhshUXb4O0mVdFEOGu0gHEUPm9Kd/Ox7ITXGMIJNkmiog3mANMNA0
a88v4Ess51mH1+B7riykBUSMvM5wVRRcF+gkBIlD/jHCZduVUCP4YE7UEu+MXAnfd+dqgD0ZUs3v
OAjS1Z0UmR1HBwySYA1UM1whFa6V23MX/f4CTheTR/pUQMtIpOG2edcvgxC3HRWbQ74obmIardmt
bKiq1yngepz6+/VWG27aZ8/GP4Z+asVeUIG0EzxO1x9R1fV7jKtiL7PP8vCnA+TdsQrH4YSblMM4
41xezwtRZunByVtoc/K0qWyHi+PIn10EFOoI337UaqystB05Zf8PYY8t0iJlhF5dSmkqo0ecTO6j
FcJB2mbJR1ssWlu9DAPThe1G30QXzxBYTTiZyNFKjAkUamrHmQvTI897EL8c4gn2C4/xq+iLBAam
Uu8Dg+qI1Y/iF5F4hNzXzURa5+wCaYOrByiL342CMoDCt6lbP/DuGG8g69Ml+CZNZTLheDPGJOsO
WwU0OP5FMBk5HgSfKPHvP8/ZnKPmpNov0LFFaffPswqlAt4Fl9aZIyZbl0Li+kOuU5zcndP4Gaw0
9OpFr08+SZT+JrKqVfIoYom4V9ttvg78kdhRIFeQpGpzpZOsPg+U8dGDi/RtBw6tL/K1VirpYfLP
n2c1bvvDnj/Pfg89A35ytm0up/H7Pp0KtLobl0Vuyu9/kPyd0/Ub+pXCI8WCSB7wZ4w4U6ACXYzc
Zhiuayv7k2zYzb29fYaBoyTkf9n8Vf6Ts/vqoShiY7B3gp/h/fnJUF2/P9IQCzTga1TLD/RIQkw+
N0ZkSUHBblm4FtZiVFxiwimVEVfAIMkdL5wgjjmx0tJ+zhLTfJ5mQtEY9A7XpNHC0TDQuTVq8lbK
a5MBJrbTNXQAwDMLSN+FlXRi80MoXBohzpws2gGLFoRO4daMzWzlnYz/tCl3+O9U6pwowt3Kvv8Q
f4hzMcIz9nZpKmyQVD3xFFJ3Na6PHGg7ZoaPoLJNOGxsz0E8qe57wguOAXMljk/tITRDXlsKeCVV
ESxB5c8KRDPjYYwpQu13mgdgkaHw83N23sfaVF8UClY6QakTM1vr3tEJ5DXztKs3ew9r1bw082bf
xTZ4Ur+6pH7WxBm1Fu51ENJ7YG5uMW1lJj5LOtiinv/rKYCScxNUco6a+QZKHok42Cbx0PYBnEax
JL+verDn83y44ctZcJ5YkUkP/402X/0J6HaodQ+gK4w56EqfkZOGbCmczg7sUbp2Iez5EckIz27H
c0mpwBqZzCW04dlYDKbF/u8blYLOH4Vagm2OeEV0p6fQilGIu66AtY0G7jZeVJaH4wSAs+QJzHwc
m1szA7VBlpKr8UlZaUYEyYWi6eAcOgInMhh97hMytuEj2ZDsX4Il3fX48kf9JkozyVqoqyRUe9FI
JmmxNH0zcw8kcOqRMBPPXpAMbn1UrqGNqVITI7+5qCfBySWKDTqPH8aVX8TNhEFgW85RrA3Z5iOp
2Z3znSg9yH/rgcRUp6akWdMS6bnGPzm4Uo1bxrseftDMkIVOfCoqeJJwy2GtP3jMfNxZZ+wroAZp
/fJEiKvwBwu4X3SNbv1jVBg3Lgn/Balonkrb6v8DO9iTt/DiX1flJhNCfgyrWKLvdzzyFnFEARrl
ecDg9wV1r5d4q0HXRrjtxToEWpAH9IDJZn8zPJOTqd4IfyDyOxteOSbs5FHKgdVIiGyo49skZMIm
c4RH/hpkUkrIdcgYnbu96OduJu418E7ihMlEkiPot5JmK360jB7PDzrtXphPpPpSv6TYqkOLcXVv
57/E60V8KDKFcODR1Ifx8OjlQLnyRiKJunilZL1L1/9+2V93zjSYyf1NGCtnlS8pU6n/h5A+i/ov
yPiS36o36bJyMNiYrtu1ldqxZ3YZJc9iu5c0q2n7ORrVM4IV5jTco+0JmoMf4yPvQdzD2uKBMUxu
wu4krsWoQ6PXRswpdL69BlZnv3Z58N7H1Z6kz7h9SGuQgTAwaM3J7r/MSPceL0AZoQWeNf8BdgP0
lbh+yRUa7EArGyS7ZE/Z07yrXc5KY0M2XaN9rOWYga7xxDJlMruQQESOyG270LRR7CLhBJv8oB8g
Tjn12ZZWScHu0qmucG4dQTEkc1BXtsEGfTxweJ4ibZfBQ1BwlwLSoyUHJnT+pqEpw61Ny3+wWVqr
zrRRH6faCaaiAie4IMRNUH5N/Qt4sFDqs95pd9zdUdwqhkJYHUujbEBM5futrtihiNUvyoww9Yq+
vz7ayFVI+FQSx8efSnb7MMiNHp6/9d/VmX4eaut2TSYRhzfB/mcxxM3Qb3+V0/lrI/L3zFEuFq8K
Ksw9zBTD63vnN7Wd2n24lRUpmsjS4l8521S1Yby6YRbQirEjUxeeubw7OiZs3P4WpCrKxsQZsHKJ
PcQ8qT4LSAlVvxYpNzxtvBkWXktBt+/uu+daHK7BsZ+hhSgwALzLwXv+lqCaj57hUI86CQAX4fCK
irz0Z7l/folcErZIStAtC+DvoiMDx8FORgJfd7YLuQX17DqZsoGPWud7oJ2vJURjva7chCpt1XBt
AcYlkLhdsKF07hF7ljWEBLclQuBgLW9P0EYv6bEy3/z/0lvTo0+Zar9CaFufmcbpVdUv0oZceMfM
LmhHGj7feQiEepGnUDZ1/Cqu1rH2ZILhUTAXa7x3+dzQ+EnMww8OefLaT66HtdTCF03thNV3sNQV
J58tZGdcYu17eS9JyVm8WXnWLIrGo55q+fkXzncR5O2E00eMQsJjmKIW4EqthvbFOcap2KMqsO1l
WYO7E/swLcSO+7fedZUj4cUkWHkgxPkfKG1z/Kg9hl+aiUm/Aw/F/qUr8oW0Lwgk9ezO13R2DD+4
RXkt3SGEK8iEZduUdxM8afQ1hBEsi0Dx8U53XShNpo7KRHjarL4QbJVsck0vtfV4LPzwvI2c99ey
JhdOJXqbVeFi4Zvs3xEJMx7SFtFV41iY4RZqbTsE7N1lnock1N4VXe9lEaj3o1Rp6nQ8AZkT/xc+
NNgaIcSrDiHW/z1nGR1iuUqUv0OwmqmVdxvZU7kmQBpQ8vwc7BuJVkLLjLjnZBa/Bqnc373DJCqV
hsQXiZiwgCNTyeE1eLK/Gln3Ycabj178fGWbFFuhu4V+DYsyj1kKlusYHMwNGBxDXEA6m8FEvYCy
LLKDX+teYi6hoA0Pel0KhxFe8hjyUOgz6F+FViSlLvN0nokOvuUZ0UCkiF4/POJlgUSmQj2t/DM4
A02KxSMhjkxuADGU7/gIhxNAIg6AVQQ5ss6WtaNTNH09w6rCyWM4p5IDsl7ibzrESofTAyEcfIPO
/sR4SKxj+bTHpn261WafT0R14FMNzkLif9g20EJf1FEZVTPyh8B0sf4rNP70u/BpfgX7A7MBb6nn
6EauTxwYLi8Lz+pdgprqPqVCJkIIMSH57X1cw6Qy81cavnBE5Pk56qSfCssclEbev/pkaPTO0nV7
p6MH9DDbV7YM6Xzz0l1JSMWhxvNTfGXbnmUA/oaxEKBahv71+4NTZPKOAuPO2XcVANSGL8jlomvI
ObkYYMH0QQeAykPPekVDPhEDThLR0qhM/kqsAVdKTR0JBXkPEf0Xy9HaY2XrhVPI2rtXDKvQQIbI
fpffF6VlI0vRY/z0G7uq6VeFlEDbj8CtpQSF6YDwYNiKyh8PjbVHp2a3W58zrdzn2LeVHudgOI6X
61hLpIywApbqXCu4tAcoUgiuT8iApFGo2d4vp/AuUuuYNU1Z5NFLbqYeekWJQjCDqaDgdJ89xW3S
J4hWSqiCx1GG+SSvE6bqAX/7K0466kCSnVd2BavHvNZpf5M8n+shmK6fMUQKEAt4G+2VmUs5p6hk
J0wEGRNeCy24DyFBct/YJ/9UFLwl3TM/bovA/HHe1Y3BlYmktO4BULBqwcAgkmrs1vM0jemVBf3o
+Np8PxK0I3HaOOT9DHBl4ED7KMWV3lUmy2nUPVYg+A8dv3M02mk6nlUNXQ8/hPChLapHj8Vdb23A
D81EV8eCk9eQ+gDvmUORR7FKaU0JkF46pgXUf4yWnSpITkmBR6VOoj7EXaQ6Jb7ddnJr9zdT8x/d
KJ4n3Z3RNL82DOJ0+Hoj9SHyazSudORvHUkvUA/uEkpM2fkoc5ujz69x2xaJ4yf+3AJIP0oFC3G7
/I5pUVIuHWGu0VZJ/0mFJ2ObQcAwPkkht9xH3kOb+v0ccx/q5isUVDnBvN4pJwm4QtcIANJSzIbY
O/70EJxZnU2/y7sDtUVvhoV8qSFzWQW1eXBKlc6jsAUJtNYpqC+K4OuQfljnjyDN8fpMgPQDQOjf
aDhI5nHe2im7CjRe8AI5eJ17jredjS7tgxbbHEcGCba03/BITPmUY/UUQXuGbc3Nk7vDKimznl7Y
XqQ2vvOn419WZSbhTXpFJFSu+lWYt8co7JVt5i2KnpVE1+jp53MXyKlNe0+do/rZ/AeO1eQNYWa4
6gCHYjy487Q9m9ue6aWwMk8T93sdtcyNRgbdREYVbILiNP28nh4djr03wtKC8+uJwXJf+i2JeAY/
RMDTXhdl1baneHrepQ4C5Gu5+6Vz3lN5xb1+A/5qCFC/bTt7/38q1rW2pBftsoRimBOJKyXJYpN5
9w4QeyoHFpHhSbu5XKUnv3aXC/ZRqsm+JzMMMKZePlHJkqGiNyIIUDa9WgeserRv18LuoELWNvCa
1L19cGVkNQFxsWKm4FFFA7R3NsLDOMrFhwo/1Z5pJdK3wqnJzbmwFcLLX2PWkBBe/9FesYHB+PGm
WyoV57Zr93tRrvJiTqPCQjqJnFIf5/opdls0WbC8GW2Rsa9ZvMlYuGO06B71GxB2nXkMlkxhDoBa
ntyQPiUEfxlinuDGF9KZMDq7WUmVa8V9/YovE5cuZIsOm1oQDIvvkHyumnOPQ3svReLmraJjkQoB
Waz8xHcYS9B1Yy4ykbqqlsg3dCmKI4bLTm8wlN9+FtZmGv7azste4LGJXvssGa/7RGi+aqeuLGjN
jqfA+T017Eymv1hlzf+NOd3F4Y3Q/jcnLxNRt1X/HIXP7Co9IqhNZ88f95krmKWZpaJcJFCbMwL3
CViLUjFkUwoNiOeQofyuw2Mec4tXI666jQ6cfMoHRGAz7c6HEanXwZD2ejuHAxeOQelDPU0LnMGH
HvI6aQgjLqumJ7GUoD0iWWy+OAtCvdBG9tuSPKy1plH7sELKVaeY85aEoj5hDc3fFu2oktVd0h2H
mEB5KcKQnoJCsK/HIpa9J67DLXviU8bjcO5TE9mdNdqSCwOynXyTNpj5Y+Ft5eAhhSzc9E1b89sk
T6zlPZ5XGnW2NWATmId5qXaYRPqkKE1f3qL9gZ2K8NftdVMO/v436KCikz9bOHnpIlSQv1KUfVxb
bQGUSKuaM3EYf57ijfG3vQeT6WsD5rvL7JvGGcSVDdGuowIr48HVoOeqTgUYmDUPBk+h1gIpApUr
P9MCET55Fqq0Fmr+PYHTTeY2nmTYN6WDmzKDVn/t8yqwfVvff45TKJS0bXlmxvJ9UVhUkzdQ7Hha
pfGw5qBOJkdTr2MZmzGzcqodcaSqXdcz0bF7tQ9u/YwLgze/R2nWGM74b31SHMVcog+ZdFUnhxz7
Rr3NVbfweF0H0Gem/Fin59P5r1orbl4w39h8fbGRRyoam/rlFTYRSvOP22p2Nt3T5cN9wdRbG1TA
dJd7HMUhsCLiLx5TjKGA7kZivldh+Q5zcBB6un434DM3F1lgQ8Rn/hREHuKzvXp8/Nr01YcuYVEI
p93uYc5oxs15+3KTQ9260ZLWK84GosOywcHw9Eag0Tza6zq5OpMli7Vq6gcSiNxe718gZ30uqaOY
xLx4KI1Zzmd0Jd2Ws3/Vn8+o4bctREMmrsEDel3DvQtwlVujkIlfl9yxKCztfuKRtGxxZHVN69Bg
/hP6zLJN7HDCS/P2AJjAZNaQxIkl6qskyrVUn8qET20Rvy2UGM4OKNo38GkHv+n5rt9NvJ7q0HmH
5nMHLXa3OXxmzqQdIzM9x+IKXzYl5C8mzeTVV2WqtqxRQDtXh40a9FGKHIlM7aop0ICrg4pNGUbm
rB48dlagSV/zmaBWbxTLmQ7Fg+SmjlqL+fUClVCv4e5HgjJ+xi+wAmi0vdSDj+LuBAJ+raCJAK0n
RYixy/7k2VA0/HX9qax0qH2kJOt8gEF/Ac280Z8H2KU7SyYj5/xLhOEGupKj+tr90aKBlGGl9QqT
I6prQLUhHav/9yUr1pKYpcDp8Jf428bXtsF2nZ5c5YP8JyMuuACDzw1rc/RcpIkmVckstM6cPz0s
ET1rT27Z+POrXzyjmE57SicLCjOggY/b7PGS+HKc3hZeHv2ylzUUb/ywGzPdYXsFdbHBl1y4TrGo
CvCvfEHD9BNFMvP2bN+l6D6tsPpDWPM8IX1HoCs2qfM0ST8IMzhvpjBJ6zRIfyWlX+tdCL8k9m0A
0Lc14getLSjKTV+K7pRjddF4ptOT7IhlWDOTEP3VFPaZdZc1NMxqME46o8KbpbnnTsXHEUQSY2Tq
J5Dmcgp4F4rEpCfntxStOguBIbVd/VxO9JuPoJwquuBH+HIi1H1zYtYr3sFUnDSUpUpdO4c0WoUW
aXJiH8nyBOnLAE29xvXjmUGwxSDmxq11aT7WyE7ULQQM25UOXFTuBqBE6jA0FidamOixI7FbRC6E
6Bak/N9eKCllia4eYmQ05F34e6kPHOz0uS7AIczb53PN32L7ri6XbzNrgYpCfwq88PVHYHQDv1+b
Ag9pBNbpMIVFCxFIaB8Zl1I8LRFYW9IGZSDl2CI3X2yZ7vCGVm8i/s2q/4i0kJb4WlvOtrnloKLh
WQF8Ne2duN6zGsO5IEvwtT6YoUB9+HnyDqnrsCRsGe0rham/nSYXhKDXCgWv280WA5332MI+u8qU
+LS+OrzkKiNGGKcDyxmktDqMzOtGRqkrvNJEp7fcVThQ4/VIOAICJ9JwnWY4khX8xybt7K+8s8rM
jgt/fdtAPZTgIxYbEgfdApJkKj+HJYKpWxhGDdthfTpqwo1oCqypve3Ns/wt1l/IugO/NaaWqTrD
qYMoui1cdPTJAADN2R0vKhvLcQHZ3Pvc5/8K5xwYoKpPj3Ww1ygprmR6/fclEIzwq/2g8BZBJ+QC
oM3J98Eudmod/ilotyBA8nxA1oP9xPTwmSayCFD1NeHwsXxlAlES2BaiLsThGEnchWwQOL+TODFF
4pFoCW+ZfZnJzSLPt0yAjkThOQgtC68HZ/IkuBm6dBaCAoDVFbS3BhICW+Sa+optjONmxbhtZk5o
ktRYq4nGEMA3HCqyHQNU3uQiKlw9prFQYQRmmgzAzFRi4qiwjHbgfuFwLk8LlnMJyf9y2PcEuRfU
hh7BlPM2Ylkx2x/AvDcPtwU9NSXwSndN+gvY3j6lXWoxkvk99bhlMxLidxIf3pjT2z4NIHXbLKsW
/Kdgvd/y40TUxNH0tIEKnDhsHIFJQqwB+gsRJTBOW3bYg93gu0c7lL/RTfRBunnq8t5X2eOJQKaR
WjBYcX/qVxJar9L83pFe0L/co5cIIhplDcDeLXCnJg04WmVF1ubuxkWlDBmlm8GTcVf2NyDSnjor
nZGOABV7UL6fpNIwDCz5POxBV+Pr5644z/9mLAL32VS62+HKFUARaMZMuZk9/8kB9degvGxtqUSi
JMQ7/p+B0fbhcV1w9nMUWk3sPSJIzoKV6YvnatD+nkDasd7fM6G/G6KF9uC+05KzHLVBch9YfzVR
SErCbJ16D8hiH2Q28j3qw3aV3uP7dkEwS5Y0KLdbZybqlVXlNlJWO6rG5cTYpXNPmHJzFM2B2yei
e7A75IbCvnziEbdK3PZQmn7DrS8vO391fG0vY5TmwSwbza0mqX4XauBhPcZWkd8PPjFwVTH+lVV5
P1Jn233R6pgoIhX1VEhZ/JW9wVmX7P1I+WJBnFJQuwnp9Qm/yxXby0bunSL9FQP8bhqLkAIjqLx8
jgAUH0RpeMopYzdNIKbWmWW2Tr+P6NwS6rVzKlmRgJffmVwPxB6e2gwR1D34vIWUECa6bu9VP7Aj
l+nkyRHLoAdzHgdvbnjMbXeyr9f3lnvV/yrGquMrWkneL1WwUBBjE9Rj9tk7E9ObdHAjKwpXGjJr
XGVt3vEfRK3Sg55FHK66qVwGHgBCFloULt2JmK+WiJIH9VvH5LnnehMrfUKNQRh0bxcS1Pdc55sp
vPupvKg5WkglEshhPRJy7nGdpPnp3C2CAW1/quPKfS0e+TNm3bLGe9EyxEx263ww8QH1G+EuzqKB
5kgnpBpdD0g+c1i/C49F7NJ1o11z6KkPgjkCyDFMUoJy1ik34C4YkKbUWYuiV4l9YflP1NFPIgNL
m+NGOeEvpOZZOtrb5xKMHoVodBresGoHoPhvniiUxWU/eqpCissbmAjF9X5zh/4kT6uVmmRQLVo2
2PHTxsvQc7C1ue904Ve08XnRKOwV+TjMNPB3p8L5OsQSo060QZaNouRCuFLwKjPXCozQjjnRYUcO
OUoGqNKfZYr/f5whViHNlTURAqTy+jmjogY10fh5cp6HGpbMh5IXvQXp4EDTARVI6sejTUaJAYUQ
+4BddPCxZSp5zE7Y/JC2On7+QMBtHlSE7JhRtaLf+lqH+Odyt+Mguy02Pl00mSoPKVjEis13ieOJ
TgcXW88kRManA9nY41qslxtMxSu1xJ2pvFYHyasFiSp3uFpv/n0L/eaLW50qex8xO656tWZASIuD
oiDfZ20mRfvXcWzvEz7f5qQcV9TiEklMcfqy2D727HtVRghwNWa1tqL/tSkHSrLhyJXXLydkFWd2
Bg5c27SQhrmaWlFNO+Cf17Mh9kvldsWid4uZ7iq/uAGBtIqp5UyI/oghw+Rz2S4OQCHM9HjkaTWQ
R+nElXAOCV3LvSrIDEHkVaervNwbg0CBWYVVX67by1nacApS3/zHPPC+1ISUvQ8nH/o5Nw9zaEgk
z4cxSV/uH0NLtp4MbN6Iznnye+Lty1IJIMG+3I1DFMRJFzBkMY5plaI30YaTiLNKUJqk++S3HckU
1mo6KhnNLchjgQGmlq0aO/1/RJaY/sM9r+fnQtr6lk1XQVm6ZLbk00xR6OkFGPWApuIO3llWymX4
syS8rdsk6dwMD4Iv/wMXZN6HasF+hL0u0NW9giiRF8WLeUUXFyL3Ft2tDMztt6vJu3F/gFLD2zaQ
NGXUNE7Hi3LTLLT1I5EYE3YBP5LrJYD4MWycDRv9HLAzBfFXnVoCPY26LO8G1E7RH36sGafGHeOW
9rCiChFnNVopaJ2s94pNJdAvaU2IrRmu7kz4g3iSiIl0zKHv8g4SRMkEdan15OGQD/kb/hux45zF
SJzjrCHP0DuFrNlm/U5nvJQMfY8X64MLik/6lvkaGiVVHR5yWwhiOBWMp/2moKc1FtDZNtoObUi5
RRTbUgCDavi8EA8+Zwijck4AI8wtrIuG65pY9SLn68v+vqE6ZzFUTXb4DMd0+T4p2iamBgsSsKTG
94ICNIm0ndH6q5hsA86Rj/jVFxtdVGxCYsMk5vEWe+v2RZJ8iHuweiVhb/IyVQzXhQ4HeCpOeN3L
0Gdx0QNX85eWOkmM+/qGsxDLl3uhqZeXVNTTr2cNUyKw+PbRgPpcuxczVNEZfXXijDdsfF83gj+v
pW7fexdRtLpnZajocaR0wgVYduEN8H8vAl4XOsp1EPPw89INhFovVzSY3ykrI2vFNWTMBh7MGPaN
jlum6ljksOAK9Gt3jm5rqaiOlzft+wgbjy08FEc5AAIIIz0QZIYppqlZX7X44YpORPQpXju6KPr+
MJRPdc+14DxB5jdsTIEYHXgbexb79iHjP5HcPLMyjONt67KHReLX6zIudqabdwZK7UCLjYo4QTj0
a3LoLizv9GGPpeorae+J3NfMzVTFedq1iy2gDPwEclRznHrfJYETcEBEprRmF0Ogk9njUnsVevJ6
/OK86Rl4Yr5aU8duSl+Vlzm/ExJVyCXK0A2PFBgMxXAKWhHNYEPsxH7XLc1CxfAIkhmBQVNcSCYB
q/oRLhS7zn6td+ZQMSWbnvFLM1yj6oDrM6ryMVj9rahs4ohnH6FFXBhDIAXbaIe/+r/8E9/+vcp5
/P3AoU3IVekiljGXfzs43Vkqu8zK1nPCSA3vd1r/+weBTXKdIlrwrpH5+GEA6fUan1LgEAEDditX
wJM2w9pn1RSE/5Q34usQ+ZoIotglpNtzh1QAc+wvyRXAg+hMIZHXmiv3EMTnI8E7ct14PKJ+fdWw
8H2vgNmPhvEZs29NOPe0m55s+zh1zg/9UvcLHytJSo6tNGOtT8HiB3W82Wq3WtjkWKEaW5aaC3Ao
wU/uc/kfAzy5BHnzKX2fv9qK2eNHA0gQqTh8w92F3LcSkLzh6be2j5l5L9gKRVxa67V/btX42UdB
Idcla8j5yl4neJDzUSrAqgV72sO8BPHlaKbqWOrbzdhhAS6AjaTjY4Ku8g1wIrpcLQ+vAZjZOUQI
YkJkgjjNQ50hkvLaqEKf+ATUbuubngPmcpanihkhHRuHWhdcx2AnE691O7ah4EhIIIc7HgKtvETX
7PYxNWmZ4hsUGRsYUCIBPM0uKNgSaSMEhKeaI1bCHkxCvypnqNiaCccMAihMqHeLOgiXcKUbAvtH
k9uy8XCNawGYipguHZ681DwVfkshsoMMzOEPsgO26Qh/lIhXN6NNKgzqhOoIZZLVbQ6bYWA2O2FL
ixFwylxIvs8jcSAN3sxcX85yUeFQZe+H08QAaho0tX1Vu4I01dIUURrcD8eiiG76xbtwkOmK8FUl
bAsnS0xjIaTGYC/OV8BqOPbUogkjvSUGqZLQq66zWS2ARAddXmD2VUT0IIhZPE9xCX10K8/QxJQR
ns7wI++BYRXP6tS+9FRVLpRHOk2CJOjEeIFcq33l1+nzR/emIzStU/VV1t7S50HZtZMffd2T7KQH
fd4aCHhn38tDs8819D5iUZF7513bpz6OpKQ/WESnK5JFcq37WGlL2evCR+os2/Nmm3y1ZWfIHV3E
CREzOH/WfZC3B9m5G8AaE8sxCpJz26gzafTaJHMNciJ+kAnBaR/6B4z7uxzqXWr/ASM6gdCSumIs
bylYutguiTwsOqhpHgFhnUMY23jt4CGIvrGkuO4hE/f7nOrY3g1r1ZFsIDKEXRgN2j7MyNJj6+CC
xc1MWh+se+Tnj1EW49sn1hIxFnhdIpkfCm+GrgdEoQyi+uOVBl3kBpdlovUQ7iG8MVZ6mLF/jF2l
kS5QBk/MFF8m6H1V5Lcq8BlOFAei1PEyljXIdsMG60dM4Be4YQQ95aCI/Oon/LYywbvbRmzil7Zv
kCacojkxseRo8GQ9a4UqYaR+X18XCLY4zbVW15S2JvMWzFDkww6J5BzLhWlz1PHAnbUBs6aaaitg
T27ZHIEP7KwxsTs5ST3HmLlwAQmSIi8dBT87Vp8ckJ66VW+3ikBZRzv0ESzb5e7fLVUUzXGsa7Kf
sgp5DYw9NyJuPS/Go6j0jvZUf8+XpVbFAFIkv3QgxXWQEljjlMjKsAA1YZqOmO/ecflYIHnfwUCQ
Dv8wo5qnqB8KLaruL/KlbdVRvkXWt708+vzv68/IbtuTvQfkQNNZhNvYHOpP3jTjQPu2azUVoiDg
BOmxyySxwrYR8vobs+DR94+kPSmVNI6A/ViNNY9NfIf6HqMIu2b4TI6MSNa37XuEK/5in9uSS5Jv
BwgT9F4IczHa1F5oysIgLFbSeA9ai5B/iYDOeJxvykK863vYDxlEDAzV+T2xl4rpjGnEbH7KTJzc
qDTUYukhLkt29W2t1IQSeiqxzJjku8QMcm0eIhWeWJI3wQLiLP/uSET5YEs95iXd8LaMPeWqoH7q
31zAOF8Fu/Bp/uZsVzSwBSP1YCxrrKKKsMXAx1Y5M8nGNtKjpmiPAlsqXv3ZVbgnQe7anjm+zMCw
x9RkftdSWE8Hv2DOa42al7Pg++urwYPHIo+KW2+rAxPgnWMHA+/eMhmKu3vJ9NO5sBRJwNw0nc/L
1PeLqJjbYRj5IUTVTi++1gr/N9jvX76JSXBmjkXrpZmf92z8GwO/0g2407ix13ydyOmucYmSgDFP
y0giCY1mKbfW6mQMh5svsQqjkfsnyXPQMszCsQUB/STXBSuxJ5LPwsxQH9UqA/nwqcBGlsbRdy53
yqnt7kGPbHdxkqeBGn1mrEsDrLanaC8ifkCBzdWorleKNSfDPiwVpIfStp/SK6+kO0/g9xPkaOcu
vvK0nm1EPN3mO6pDqybChoWjE1d7CgivSbMyfhSrXGIJqBmbzuWMT0NnDrmBglZU085zKclenASv
/s3fElLOy6z0SulICHGExzC0sIRljK51NHjsNkcLLDDcvr+2FZt8sSdxVUVmx0aStXnI4GxaIhDG
p/VKOqPGzJ3UbKL61JqwKYeVYFIop2PjZRH/w9KqcC2a15d7phtrzvj+EF4X0ntUIAr+Jz8KWC4O
CuW/lA5BkiXh1EYHFPJUotaqwmoCiN3xF/FxeR3ZKtbgZk2L42lLSKi530JkoBrZbei+pXHuH+pK
GkMGlda1BrO+7FCxgjwTTgr9a3k8K6Lxgr5ghEMfdpCgLH5g4R06RwrO0IFL21azEDk0CdaCmkaN
xzyGXf9cecZ+txR8rrftwLpBSkkWX4xFl420CpBydqzjEm4KUlE72jGqqWvufoLnol7DrCGY+OlJ
YQsVcew7d0G2DY+vg7N9yaNXD6/P2yYIcT3dWg696YW8DacaXdXIhcTjWSFFk5lCXCPH7lZb6Pxe
NaDxdvF0mllVitD76UFzR0o4cMcYKaMDrM9cVlhsYmycu1bqtOWFW59VHyUBvtnvTRvyb1s0y1EH
cy8UkwmJL85LoqylmtpFa6aeCZCaCprTsdCfClUTna4GeMN7sfobOmoOe6EC8k3DCxkZ3aNZa1nc
PTo8dkUyFCprYowGI+1WAjAwUf3Fj8o+kKZvXvJeaFgbQF5zDrQ4vgnJ3luBjOoepSooL/mi88Tt
YgXXJG3dBzfOQwAItOvKxLFH+JjqwSqJAzAiQ602CH2eRrh6dTG6iCiPz/Q838cEABbtJFLrx5U4
KHw6oac288u11mcOw/wU6f0Hl4/WxALHjWdRGI2ztRco8r766eBDeWcCPfczENIMTN6T3cm/g2mI
gLQqOzwlq9O33QzI8QIkhpR/96B2EPePU8rXMTVgaOIbq+s3PgyAtEq5XZpRTlZXZmEOI3WBERgY
QW/pCSg2lEEaHgfu6sGnwyLmtyZfz4VEibuh9G7BC2MIDHCmDbRqW55cYoxsrjMfEWk1/X0MKbKp
Pf1jteMQNLRUkOHTcKcfojAX230MGKpccUvQRvoZa5HD7zmfY7Jxy63UPIrZ4Sk7A5YtkmN8FTMY
WpPBpTuspM5/ags6Rf31UmBr6keNAIYi2vqohbn+a52nHjM3osbiea3kpUsYB1zArBRiqFZLh3Qb
Yo8+l5ExCkvPPr9TcwqOkYUcSmxQ0TdBJP7g1z0P9mPRXOw2jDSoQtHsTqLltQolBOG90ehKAqRL
Ilk8mQ32wgKkARhcv3IwXyhJ/akq99m9ktDbMItmLsj6ptYpQTvQmt6EZWMWJt/JR0e+ApNss01w
cBD9NcLgoEFAUNAE2Y29MFxlAV+vHQZUq2ma+v1n6jmbMqsoXVyZzNpBA3SDDwakQ0ErgI9ducD6
DHUE5dFNUD3L+DFCC1SrRJS3qzYszya/DLqprZ4d9C1bXp72R2alB8eUIShypQftYi1M80rCG+tL
2kBAt9uIvj7Hz64bmbzxMACeKieGt3iOyPRmYUNnNT6bNqeCJV03Lr8JEi4V1m7WwWNijIr1sHfn
YSCRFMQBkkCff6xH+0iBVT1CGiF55t2hcFYWJXZzSV1oGEYmXLCd7mDDKmWrU2uGnCEdJxXQtXXh
8B4TuxuIifS5q8cGhltiAHy35Sur+9sqRNC4zEiJfUUYtGDwL1K0qEtkHU23NuoyXVbZ019sv6bq
E9XF1rKY0eyAa/4xp+zTSBlDseGxMoXmdlMe2vb8QBn4fRwr94Iem0yzlOJ/MhbMzgnPXXXxiNF4
v3YnKd/zJGDctc/fmZAQ1AQMXwIHS97I7d2MQaS0DCwq2TxiL5qh6isOFStcI3yiOIf2PsOkr5CJ
eMW8UNHj8eXuH3AseqiqXf+KEsuXwfPcgW6ae8Oa9e0c2c57LaFroyLnQ0xVEZ2CWogV7AOXSgHt
QmjY1tut+hsVERb/x/pRmsScQSR8Xa80LDEgr/FiyqMgu2jeVKor6KXOt5HvRuyDR9DV2VsKuRzn
xZYhaRBSxoygBMdG5X1BJAfW6d2N5wl4KelIO3DbGxy5kP8XCE3qzw2L1lopRTJE68lRA1YWcF3E
soczLumKgsDWRwj13rgXUUDy3WpWunPyaa8kn7jXtGHteIA9xRtlLOmhrG4zRjQb1HKuTlHPmux6
7jP/gtP1Mvt5AfYT6OAOvadS7gqXgwu5z8to3LN5l21QIwRqI4+dE7C8bbCyh9Tr0uHzstIzz3zR
I+9r2sP5YUQ+dP8EaR+sx1Adj5DV13LELKrniEvRI42vsR3hTdn4lwJgZ1rj37FfGPCTxin9ZT65
7z1jOZYh4MsQqR6v1X+stfhVpodTgsEFCZM1tbn/P55YkWlRVhF1N3LO1lUPPz8M4W5J+WrI7d4b
9hxBK7Kmq7X1zZ9dyCJxaqJPmhVqrZWqxyVtmEATcHQ7qaVAA3xs+fmpRezd/mX3lAXMg3zLNMi8
WfevFl33nV20pLEcE404IM9hN94sBYY7+Mu3GqRPXQUC2it890pwKclReNNnaPFO130Tu+UYrlwU
3Pi08rUHSJuuQUeTQovSKR2WSIq9Q3Mbv6wQtZ5Dc02cdpJz4isv29Y6xnQSBfN7E7q2k5TnK1xu
PNHPkZ4DnWUIN3RMBxRbKRI1xOLfO/+KMw0wACVcAMvmXNbe+J1prc8J/CngwjtritVfixB08p/1
8gKF+1qo88twMP6KMo0aiNhDH5zS1DZR7KXkhD+4q1C7LT6XV0F0i46z5bunZUbsBtxGYL2FWakt
qDzj6wpRM4AZQujTIb0XU7xRqp/lIKFysHpAXqKUZcPOGOAq110EwHdrH9VKWRBjJxwyGWIKYCdO
cAwvxX/F1TaTk0/pYnXVOfSEkvt/cw2PjMw4LnU4WhMmnAqozEn/f5tbnPyQaMrw1/uciiaISPFy
AEFxYs9QN4DatbjB5Y4DrjNAiPfMUNytG2o8aQwVfI7ODnokNQMCqUrFQ8zH2UR12d99iIBGc7PD
6y9EzdjK0iqlFkfTzaaV6felu+Qs0tvTlbd5px8n38+MjRrk0T/eNXO0ARGJ9u6TQWT77w54WtJ9
XVzlKY4aWFNKHx2WC6M74XVzIEo9NfqAB0t3VGt12Cao2hPuiokVAOpZQAT4AcsT1/Bk0o2/KVPr
aIOSkRbCQO4CGsw8lSgM9TB9TWDHoLE2/oMSY2hZV5wiiufqH+4B8nUzfgbCtQdDksgOBhnPV/tv
C2MmsCg10lORRRHCnGjevDF4ZhdyDFEba7vv2czLI/8VzJwB77VxpN1UqTTjh1Ri4cojzhJoXUNK
aO9A60WBdx12EMHb7fHH/TeoC0sV8r/JVoSFWSVePh+eS/y4NrCIAv+0p6y5j1Ay1V4vbOxKNGOL
/GLhesK+kz7mcXIOs+yrraLk1bYtUQ46DeNwpRW7h1MW1owXBNhZ6Xf8PWJP+1fclyXWm21NuKg2
k64zlvq4hSQJTRa9RT5BaZ6sKSCPFW8vfjakTUng1ZWDGz7x26xnVTXgo71uf+7i0J+3llLRkJKF
r4oq83LFjs4yAnSUhsp9wINvsgYbLOwQ14pkjvhDqdr+iZsQlrayzCy1VYue+cdAoDaikupUd8oM
4ioOXGkWTvJz7sX/Wy4ykm72rVV/rrXzcdPlexA0O+KcDHJUxhMrDAcXE73J6r3h5xRV+zAVswrn
e0zhyD0gtpAUEr9/NZ5rjnlx4ITm29PppPF1rTk3DmYrLJZwk6oqNz4yaROaBRMu36WaAozIEPAO
T3/LoWaR0TPH4obJ7976wHjXttDjJXDV/Rq8SYbgHqdq8APRI0Dlm2SYLUYciOO/38dKXXA9lhlp
tekJUsABvoUMWiMBBexcaxNByuUlt7kEJxOwYWCB9jgOZSvw70W5FQ0AYfMQ4fpnY1FG6BLy+SFA
IunQhbqnUAvyA9E8k9xOUPrvkNKE9gIW9xH70V3IefzZoHaP0VVnuSYmirxkQEeSuh5+y1xX5br+
ZN9MJLIzC71LqwkB1lyEyfhBnvEgS9q4FlwcPUX2RIgSPUykn9oYvdbobiuAhnON1b07UMZRGM4L
s+U7Lp4m7RzXnCv+aroG3qHSKdolVUCdrNT6lYEqt7EUnXTTr0zEKlKjyKXec6U3xPOgxxJiOIkx
7ecHK6kPpfeNBnBfE+DiV6GgARbcf5DTFNvXA4jwJIv/7e8/tpaZw4v0AFPF/IJfR/W31wgnrZju
NY+F9Gt2JsMgcUQLARmG2jGr+kfwWpuKeG8HJ0llp2XhR0aAIq24ug8bTFwFoXgcJc+4RwQ1eDei
LI58fZyab2m7DZeJIGT3C/yXimkMmxnfJZe+Kz/S3959k/TZyzpUKR1hkesW5yHscPMTv48/QPpH
96VBF9/sb+ts5YUs9M7VlWs7/gMQ85bYAxjyfz/E0zCMg4EkkAZBGfkrON0jfZ5WicsGQzK7+Wz9
KXU6mFVv1Rl5BGVPZeSk07GA2RCKSMz73OIietmc082Kb45NSQWlLxKh/Pv+1cFrSulcFUw6F6rG
GbU0mSMWHWWHL4Mny57uL8TteZRi9K8YTjP7OLJaJkf/JqMixwXnxZhsl8qv9jPv8oQkim84IHql
ieWCFpW4sKLoW3ygmeE9m4d95o1cyjBZ+k1Lf00su5I3ONXfzMlHky4brXhUbTTJdb4DfVTnDZWr
8BdT34HiPB0Q4gcYypy1VpA+ueHz6n6U6FvoFlz2wTW/hHIVTyoKZLTUUxx1GWXaANWJi2HYLZuK
9YcPX8FM0f8q2JbrlMHNEl1huyn7LKNW+9GVGy3P6w4APIuofpOD8cuxRVIosEzSieaoNDYkA4Lp
pz6OGIiJfSUKu8+B4apFyELmqvv0whjXhWWUcJp2ynXxMs0rua4XOaRel73rOI0OLhKx3atD9FJa
jH00RzjIGfzCq8Onqa8rWlZLxx4xiFIbIACH6C4TVEFQPr3i543EKnkk9t3kotIbxT0i3blCUSVV
nFhMSjhCsokR0GM9tx5C4yD0LEqotqBAzcuxJ9nUoXrMoNs3wAR6pCXbSxB/R0+3ia8LwE7Ml0uq
u1gZ4S98FC01gu3DmleNgMQkjDQb+dyh0NYZ9BxhTUDg1pw5b+3+xxQfJ8J4j/xCtrbiq4xfMuxd
8g6O3jBMnrwsTrcv3aiI6xLLJomqiLed5zI5IAzX0gsvIiZZeFB8CyMpN+5yr6CuzcUW/pfyGuFf
WHiY2naeL9CrulRZVEN9ZQ68djBeQ40Iap3vbRhqfFsNjg4PDGMhbhPi3ZlND90gqDVE7RdKkA5w
u1S5+Kw6GWF1MTXU9y8v+9uMXDUMCB3FzFPgN9r8wxqZsifRYEkuSy6i2T4HWnyrRSe9tBVf0U14
fSyeE8zpdVCnJ7xptXhoN8xQHzn+YVHUAmBf2bJGBlOI0nLH2K5Pan7QrTRQSQf7/UEdPpUY3Xjv
+40E2a7U8uIOM83DhIZ9H5baNiNsQ+DLRmpogNdfGhkpHVSJ8ge+6HwtAAHTKSY5cc5dzE99Osb9
1eQa8lygEEOQl2/HJnJPiSUO/SB6509iZ4/EEa01xWpM4WHcMjUd+1nJ2kmLWxVO93L0B63uXHQU
HNIIkBu+IrjFWz1jZivI+v9NoNGA46ef3toXjbxFu5jm5fSzQ1aIwZmRc2HWsBrB7KXlIpDmdvfn
eNYoaZz2iBsEi9RpoS4r6gfdrR+cFrqvkzcZ046jNdWgzqJVhL79nTin+22AZQRrUJqdNHh10HL6
aTMOa6IZGtpTfD5E5Az42ph+gOzhFrJssoorFJn2JJkdBTOBmalt3010hAcdm63x9fm2RSjOtutN
ui+KAsj2d4xMGECAUOwao83PS7P7zJzHtuTLqbl1MVuEWAEV17RDhrm9bvX9lrnQQE4Q+7jmPJDa
Iod9YVTfb56lEWcp5Lcw9b4Wj27eccFG7Nm1A8GHaDEZhk1gvgnOr0pUkrimOJVqwgWEpMw6zlnj
RTREnpuAdRFisgU7QFv7H3JHs9QOkKXC52jAszXL3cHvNQJNiIes8eC9AcFsWfFfzH923zkLMyHs
136F37wzXPQ58gaU17B6pxuJ17OHOtn02zCKxmJP/ow86xUF9r+dNRh7oiq5KYnOsu9ELnlI3XNn
WSF7Lz0+vfetVtVemGcrPUYO/Riu58O+TzGeCz315QxZ7Xz8Os6YkAN/iaPfXxjBJpf6yo8JYsFt
qqK3ECPq5ouaRhLBhmMq7LwhxGg0kjTHhek720EJ0D0v4Qa/j70VkMU1WUIS2VPUhyyLTmBP+KkO
jNLFJQM8MjysrSVxzZzupK4EMx8pPMLMNo77dv2DDY5EAMMd5zg/nn50BYgDcOTRKi+dm8uvR2g3
IV8H0i16qbSrpkFCChAdBxVdtO63ugGPLKXLi27Mezbl9axuZUPP4FBt/TVABKQ8QcqmIUbvCb6p
YoG92tE6x9bKDslpL4SgxRCuTcF84sFC3xRDiRyyCjE+Emunw4kdmGl2xsR9i4bwmcsIHC7bdEVD
44Tzvp9KO/+2CdXsDeh95BPqHBvmNeY6amCE5BqAVl0Z0htVEf20xy9MFsTXFMYt5+Okb78QdGfT
N57o3y3jjSWfl3GFZxkhgiR9Bi73dK2wCCCt07PPQrFVP5QVeUZYiOR+a76tSyShlFzmNzfppZ2g
sT14+fSKbVG1MqoJjYIkV+q4s+RODiaxPWhizYHCvbdZ9R5IdqvvBTsT4O66Br2Cj55WsVjUDIhj
tsICg59qVNAZGMm/XDH61XXU58/KvLwt463F4IoC94jO+MzY26drZrljuCdY/L+5V2C5WieCmT9e
pV0FGSQfkGm26LItBcIPAc9RsUg9699n+PB+le5um31DVbcmggA4huXX1X5ro457P+EsxfYGHjO0
+Xdq6BTjgsQLeLHHvqml5nm5+u19S0azzjiWYG41cBp9AGb2+yu6H01Q0rIVsbDP5Cj0cCggeQrz
lP9p3UWu3iMN9yEzaRIIHayOhFz1OQMMM1M4Mb/DTTSvmZO59o+zHJLfUO6OPUYbo5FdepbyUF8b
Q3MM4c4cMXhxwYpEO2E27fTfNm9GV7HzTJHb1YRVzLmEIAt/tgAYf3QwsvhPyRdY5d352anWdw70
AYgKdX5eFpLg72PAG6daaY3MBN3uSAqwSpi8gaQ9xodJEFRVgCKNCiQ8pxkKo6ACJZxUNf3DT14L
EBeReKFZCHbcrAyMj5cRnQCIN4cHJpxWhQDW79SXAuy4pwUt6f8huxS83FgluIgFPX2tUtIdZUKO
kRL1wWamvobTWQegEHD7YwZL8rg6Rb/brz6tqoMZWJPeQQhaDMhzO3dS1Qc7vMuyKZ9qf+lcJ74F
e47qyOD1KaipYP1JQXfIzdPOKB4azGxpWo9KtsZLPfOMMaMMneAuTQHaVf/aeT4/MpqXVIo4TH0K
pvReke0ZuP79lpsCczSoY6PvBrBqnPmEJs5HRAS2mgpI/w9NlK36fi8EFDa+C8a6gTuivyi1asKh
26rO7RER2ZTRyXr/A+Kq6myjH+hAx9UvpvXdoaiC++LNdXSkPDaMQM1tbhwdtwMkMlhjsVxaIIBS
ITtAYp6AsxVTfVOHgwRrNx69IetrUYwdTTkXBtsu3tmKh4nbLGD+nvhYl+DCwEVWRfk28BW5V+Pe
2fD7AUUNoB9C9mc/yrjHJBww/7JVxw8gi+cvn9wlO54G98ySY1etQN1ctdqo5e4Ckt4ZzvASd1RV
Orx4zn6TD2MD0HphSd8tHokhfI/vFJX5zqJ2YQjh9pErRifdrhWcoGfVlTnpk8JXePIR0c5pAS0t
KteWQcW7Ns44so+SuiwYJ/fbMQezuvVDyGqtpQDRLHp0/iIdcZlx54SqRtgOx+QRBQtU4ulBkUHi
giVDloDpHpEzXpcHXPlELsPNYmK/EMf1k3vPfow6g7XrJi9ya5dTIStx1n1KiLhN1mWpt39obRZI
+IbYnfoottr/RVzAi+FsrPWsRLN6nVADW49ebemUztge6+pupSFAP9lQBbzzbGJRvEBiDQ++DpGb
nL2sIK/xp48JESGSkem61Jq+K62O733asnFFgf/bk4l1K87cNUrvCxKboZYHDOaGHIPBgg8gM9yr
Xn3BwBkERjzB//aVR4PLoiOAXOPfW9lKNzE5V6yaPMPTXzIa5yfWjzRzPtar3taH+/zFxgqgmS0B
0nR3mnFDEo7pbRMvEbWEykNgFsE58K9Xf5Xc1BlruFIoeiKsCsEVLddkejg66oVHdodXdMN78WKy
duap/9UF0xr9MrHBrvdPopMuWJu6QlKK1qDbMCvursZBimehsCCV6lrWV6dAj5Y720xUIErPBiep
v+1z4D5WNOeP9CuAvRhc3eW3g2Y8Zcm4VBKbTH3kqcIwPsrEEdvbiYqcoXrb0r/kYpCDFNEoXgp8
nxR7OQ4X7vNiTQ+uDcJxLER2NQYvituC7QNtJK/GWsEf0m0UoSH4mlMNDpB2AKgX8wn9DfDnr0Dv
opm0UICr+a+08S4HLt4uB9WauyKGceW7IP29Q+0pYN7jUnXjNUD4Ga9mPOZsWlerQtsuYMkGUwiC
211qdFotfiVWszENwwObnxIlRyiY1JVAWp0OhpqEApyufHpTCcPUjdwps9GjbG/nbeSvVf3yMQDD
nQhyAySko6QjvBw06K7fLkr3hJcSnTE62mwtaCsCPukkjC+CU807GeZvm9kgV6i8VMmPu5jqLmie
mB7L3Kb4okB4DtLf3b0hwG11QMaNbMum0yoWrfLAaZZSp7M/kTJe5pkXD4cM8pFFh3okvptXxwOC
HKrWpw5Ak5ketizyNuOzW1m+5N3k7KHWeWeMdO30yCO1dNNc/qy4apoYvWMJWt7h3ZzxvnQyEXiu
mjyQNOSuBhB8ZB02v7aPHomqjkXhjXUJZS3yqVp95ikTr73fRlQ3AxT31b/3MmioIMOKX3HR7QBZ
C6fYG8bZzGJUhXsUgYBXfksVMOLl6z7UaHh8uVN2VCeA3E+OZL+k5SlUguOVXNCQqlKNI2k7rj75
/yXyzUtHsD+z0F4IrPsbKbU1DtbuG9CmpkRE3VV0BDbYRGHeJ8KZLnKYs8Y59FUZBFkBE21L1Cvy
XGDJRVjXnk3KQGQwcJUO4Gst/vKgKyfR3hTSxSDbVdUJU51duxqeXHxD29+ZEftCh+vIP5alRTBl
ppJA+nrdaCxGhswksmA5StvhZdj5LuTt0WV44C9jOSpJg9ncPDOKzF9hl89yqpZJN/uaC+WImkFG
5ePf3Wc58NO/470AeMLSMNyXebNnMe2wQ8z+MB7XleLKS685W5Q3wgF6RrRkf06n6NWADP8+RsNX
CWHzlxFS0imGVBHFRZoxBj6RCkkX8i32CKtedkvE10q5Dpwo4Uxc5cwlPPK0T5Sgmz1/GESYaa25
vLBadnmFoWiTMypKwZzSad7oW2vwX2cLRcXa3dzIwPMCIPy5//5Yi50n1cn1eREVQgEPGDec1JxZ
OFo4lLF7hHMoxtG6O+v1PxDsBc8Ia3nKCWhhMWoeGxutsuf5MF57GafKEDdGNHJnSfGcq8C7tyoe
4s7U30Nzv3VJzGXcWlN78XlqeQ36z9yDBLCKsfzJ0d3iHWcX0tEtx59Ahy9zt3zng5USdckJkQd+
2rphjAFC91IVKp4BsEhqSMJw1IC7yH5fs3GXDgiQ6yqT5tAhULXyuBwlBveSzLAKy36WFsKIVPp3
DFXUQJtQkkePvRZmrDrsgmD+3XsmRxqDWLurBb2w7akLmFgvRXfCnpdjVxu8A7hJ+vHtS1gNhTN3
eljTRaUooizZOpfo22U37FMTGr0ed05zZmDYWXaVGLDwIgNd78Cw/xehlxe6rDdzIV8918VCs+/I
GOnO3bQf8fNjyhHJitbmG5Fbz4BcskNn+AWP2eqOE25t+mQnZncUzAvPSq5+Wui4TErqAIZ6CdVG
fVu3QAIBCrtQik5cMWgJHcAu2pdlx2HT+8ub4iiceMvGpPjs9KbYNrhCOpZ3B97+E5b62JVbkFCL
WFXCiBWtL0fv1Al2zwOmNaFzDPnu6+LXVdhtU9qr3j1plSSHR2D1RILEABoZR2CJjkn/VW+SRRpj
m26U+AzjTc5IXIoT4XJ4ldHxdD4OSEDZdDqDeRAWWr2H8jz3hMNVZZJvRZibLz+p9cFCchvAV4SX
UXNzggdJevdzgulPKuMKPNr8K+IIn8ZGVBYeHqFvrrn4wrtw+Iq1RvHrofk+Z5V7WUHoym912jN1
AdYhi83B1CQEb5S+GZhOFDgvroMJ+Zpdorq5xIoHw+1gKYUePkq9UMCCgDem81KxTIRZs4nH3hZW
pnN7VZmDsBxDxIEDnnTmTYQtHbFXyaBplTAo2Inf2gPRm7Z372+KbCiFcJXS2u/jZJnvAQJ6Fa4T
fBn5ZF27CUTJhIM5ful4xSm3DVSQHh0hY6nqoUWZiK2EyuYYoll6oQV5BNi7xEfB+OXDlMXZszig
f24LFV01ES+WHX4eA71c8uLC3/ZXwr54NhgUErr69lHrl4qv20s2BHzt+FyaB3wPz/rUFLPrtL7p
mtHXB8yFTSiqC5gRDbSdUMfCelShjgBbr32zOgcGxPme/8Xuw0fgTtBhs+V3vRP9La539KlZNaBU
loAnLxb6lhZREGiacDiQ6nMOKET3tYU66BHZ1Xt5PMtjcWrjc5nWt6wbeOJGHtgl2f4wcSTGs/QF
9ylozHmEnSlKzekVbhe/h4qL6w1nG6e7eHV4uL8LXBaBqcLtx/VC0FIvk+s4Cndw42FnIXCt66rr
2cibCaYCEFt2ujEa/kfVW2shwQ/0eXwIo1id650LSteODZDNKp6ydqIfiPtAWyjE6njEvjLzSgdA
dm/4FbSkMCkLUYLS6gU9BtuIbkbxd0TgaT7zEgfXmXeCq7Ku2zVIqmytA1WcdUKYRm25G6oQis5M
A/E78qZQRO09D1MXFXOZkppZy9MPL9MEL4IeJAPhU2CyOSOh+Q4AWa2B5ccoTXRs3aVy6xjBMwcO
ayuJzQrwAnNY+uM7ZasIUD/eQWPH7pr5nLgvRij2fFDKa1YoS1Ih/PmOwImpKbtglX0d3JHcDz5i
FJJ1dyeT6Y6UfuGcQX2sKmgEJahoxgCnWR7j3W6xEo2YzpBTRQwgG4Ph016D8/GsAUmtRNnRiSdT
RLx5J2hVcTJwgvcS14PLtfX6AJF4IM2CRPihWOJ6a8D1wYtrMqYV7tdaiL3ln8pwAHOaUPxmcotr
pEDJh+3yr2a7JUS58htup+1zeD8SndHkGV5fHi5kfOsfZHnThqC9xWHpD6rpz2407aoJER+29Dm5
y8UP3fLyn2kkC6GiFTaqWK/pIgug2BJbQcEGY2kvp2L3sW4983Oypae3KVLEZRGm7jMnqwZPOyxM
BvaX5sHt4mrjAgWwrY3dCgTNwPyikC1ZPhzsEv1OwAkXj+hqEOH9BTYbONpNbJRP15/ViqtUqt6H
AXYRQRhl+IBBPvBs6vv3MjyG/VSL4jsrM3qsJ+l1NdBXtxnq2WIdmqb9pA+WjSyxJkdD11bzkOVL
W78whz9D5gOTzipv3RwM7mvgihPBdbrSPi8ThkamC60c6S5piYH1NI/Hy/pRRMEm8zmBSxfYdixc
7udlZX1gbRbHneKb9/4rRC7tOoz9RZI2vL8pDuqDjeSjAXwjLhBv9aWwDgaE5j4BRsIx6N2RCaKa
jsdWDbLTslRJ164UxvVQQ1WrtdMIHlUCVMPgWuzAItmupTPuz7zS6aVFoYsqK7O/Kgm4qGqaVdGa
uo6g4L//t/OF7sDK9EWVTRy/mV4aOjYB3buhFblOXlaMIlCmkqKkoz4R5hWATDIq1hLRD/ZpshtQ
/SrdzG5YhuOO8fMkM3gmdQYsFhkYZlGhfbjzlpR3Y4r2RsXOHls5dQN2m+7niV3IVaP75OQAOF6f
yGfcBKMjize4cmH9QpnJfktBAU/YxAUd4F7xJM0VJk1Hlw6S4OyUgAGvMfcBB0X+QMbQj5WZCZY0
nMGdlVswxl71Bnfr7t0+V4LGvQe2D43G/vPg8XSmVj89C+zTo5XzIg6QJFuhOOF7cXz3UiXFvwVz
zlcKg1rFy/Kd3SyAlp+aG+6vNwhwKGfa5uAMblF37hVqyWpMhkGpkxVT0es0CazTsEBhUZhUgxXa
gKuAkn/CC7W7AzYWrYEqTwXcvu+DmTbdHoZzyHUR6aOO5uSgzgTcTwXgWAADm0tX384bMsHfKnfE
xdZzVrYTy7oehfUnQ4XUP9PUoUIOVu7mzmNWUDW9JONOW2MhoQyEZ+kYLFPXT6vf855eXBg7YUFu
uLyga7B3+7adwXK0wi+mrXT298KDInb3JKQlzj0CVlv1WK8/s7Y3b3lRNWoZZLWFCoEGrB5Eib00
rTrjS+DrArsw3wKwn/w4vSH2pZ5kuMFNRxVuq2HJBWbTKjsz2jLbDXwh5Y0sK4lvUvBs66VVdQA6
JIFpgXp9opBa/lrV0Cys850FRjUKM+s+SbIqfyqbB8/tyW1DxW6SiR6+OyuM5YRvqgnjGvFwfadt
/KDwK3+b/Eqtep7Oo1fwF3QLjRNUb/YJ3P6Tbm0iyjC2jxkGRf6ttGABIsRptM6vFJ46gjulsgs3
CAL9S6m60kh3LVW2h8iI1pVlKajalZErWJJLeu7WSqn5eapnc3rW9ihpLhV9gNfALb2SPbci5NPK
UtHejdLJQBbF6S5MbeYVu+r/adc5wUg/uiWvTcr3ZUvkc/6sMkYDUFn+ZQfVWAfaAS48qnq/Jqnu
xCSfXFJiK/sNqNv8i5Hp19KhRmOAws2a3ondSKE0a/mk/UaQe8y1YnJaaMPpgeIB/8Dx7b/ibM69
RBHxKnaTNPTVS0wsEYajGLI8X+0rMStcuk19UGJLwFrnwEwQcVRW3hs4Ycsycrz/3qMXCU3hh73+
Y1gLm47NVL6GeUiWsSj4D7S8EiEFmH8KZUI2Q0+lkHPSunox9ZkxCHAXI2MligB+ktjcOi2dqqDz
XcoFTKgAGf8/VO/yjMvhepoR9YjeZZubh4lyKoUAGlgBCYy1kzenbD6ceRLhz518yyVBhcEof4fA
WjHzFeQWZLs7X0JxiBFGIMaxr/9I/Ww6lcQyR3C247LQLGXyYxaLHX4V/SNlhHqbBO7OVqzUIqP6
l0UDTO2BszAHmMXAgkYG8ZprOnniRYpmZFvSmg2B9WtTnJKWVu8tFEwAlcE9VyzdgcKqOxSOHYM0
mupAajtC+2XjIc+3534xO2WGIb2e0CBG+QE8/I3q3aeyIu3QpiU+ix8+7cxuzdBCWDfXz4H4uT9R
axro4ugP5MEOGp5St9Vc/nj082CjNb5LAMk37kDahvdhsqUYKV9FjPdKeED0ijFMhb1kL7zH3TkF
bBp7Iptav0S8FwABL+9tehnndj9GYUKRSigWFs/Xh3SjPbgb9dzm5hZkmOfWB7HiyJ9jwZF5o+kQ
abFc7XMDuiiqak96O5efJD1GGRTx2kJ1R4HYBYot3kRuq0EsLMZRMhvIs/TcDbga7qVSbx+XdVev
qvj2oP6xopkqzYbbXm6BHiPA4CKYhvtSBNh+RQVQCn5sVrxt6tIl48fVY1VEJWp/3F0AFgL+EnR1
kinTerwHJbk0OT8F2YMBybTns6blyxsr7qzIrHqXLLly229rwaf/+1jAVkZNAHMS0f6Sz3Ej6cIm
kiEJSkyqDlvGBtlg3MM2ESDb/DcSYpqlvYr6sYLm4oQEMHkXcuxms5niosEFs2pKHS9NhwLvaV6M
qaUD5kQEaGhbuCQ7+diD3H+HTsC7UKV5rKY/ge+1w0T6St8OLN0+2WZExgBHLfT5x2VkZnjxZKV1
vjXAlPo6yfF3pF21OrWTID+0sPjubB56ri84Y56AfI7Cq0k/9tWKdGl6mk6MVAoFGWNrglAGy8i/
NXDVcyq+xcy5t6phRJInT15lwzCDsub4qdYgSM314Vq0wWG4ZtMNjHxR/zdCc9WtrsneWhINbY4z
b4wmeTXUQvUqE4ub4G2ek7c2t7OlMiCGRzZSdKlGyvxu/8GlBVxEKpf28J2QoyXhEY82Qu3caMax
xyc+mxDJPQSZSgdq95NweGAzrlJfiLKjDleBrXmSTA6R4G5QhKb0jEVNSv0FT1AeIqiSHC8auRlq
vF+g8ZOn1txR4YXSfTilZWcQuFdW4UsPQ6mZrdfOo/2VW5aRAhYduRZeMpQZO+vc+T+ugyPpQjdx
D8sYv1Jq0dosF7W5kLODR1kg5XZAY5KzpNElTQ4jRmnZtnzBGb+UAYrB7ENaptwzKvApCHzEMgFI
6UPxs+l1YGuRZI7q8DxMfaV1iaTOrYyI4hrrcRb7ZdBSDnRsJHP7gTgjTUDO0u/Xndqj255zNC5z
x0/6ylTE4sQuMNfMlQM+Q0kit3gNea8H3TMWFGIrQn7p0VMnhpZdVJHGJyu1hLbAXtrhv+DRIETE
uGOYZ5NX11DvWZkF96xPn/MYynbrJw+yKBcLyERK9MJ39avL4ng/imhWoIgmpucQtMulK8hs/YfS
JQDu1EuWtwLxaFU7R71quohe0/fUFyfxNNf8GVwaOhChZx/awO3sSCIq+LAeEvZIHiZ6R3uG5QG5
WxIQ7iyJAVfKk1GS8XbzmsK6gKf3Xwl/hWyl9KI4BxDbf9ZZCgjiAt+DTbKfg4cwtEDafmKHjgwL
EtXULfHWWAUL5oO4XJidihPwLj1O13dBJFEiLoFWbLW2HhTNX64SoINXvfzPinGmZCiCPTOHxLn4
3T7mDfQamYMp1rlDvDes56+r9pe4VZKBZeoAsc1gupWHBRFGiQMujvGseVXlrlWPFkSyTfAwipXR
IhWeR1ZyCMMR2RAVSGZqsS01u3NdK3foHvS34rdQNwRppIpgRUI9oYtHZAcouzwEI4bEc1YliVG7
oVwafvvpTElgYrzoa9p7sVozdsJVSx369BpI8Kq6CmNCzMDiGJGMzEAKwtzlvRa3ql+zYo9dGyZf
n8Q9kJbTUL7BlYbomhKbqmcMDwLJTHpSC2JRUPUOZ2Y3DMiPo8lVg4ou7sba5k/WIOxWOubaz0e4
75jy/4AZHeNrEa7OwmgSy13luboKW0YrU4pU9jhx+ypRO+NC9G6hvS391zkwVHMYnvCMFnujOK/z
B5NklnTDwJlg/1QO3QKas57moKJHcJDwT2IzGDPfmx9zemv9bhppPWxie3hd0rr/PuoSsOqF+PT3
dNtCEibLtXKcxK2stxJUB1ZeF8PVxLoN6an+swMv1/jbpFBkwmsuDG8430bE11W3DtURtrzeg83K
uz7/FTKKcGspnI/VvYOjcZ79wOI4ufDHhbJVujyyLm7v6b1tTCduMcfBtIHM9L8yz+T/fR+dmTBT
kFSVkCT/Kld8gIn/T5axQ6/aOjgVG3dtfLJaWUP4zDzfdxrF9QqUYhO4UErzw5gtNNDJs+BiCJZl
48yCPlYo10z7QgxU4lutz/EaDwJsMhlCDGzcIpameVR26XoYNWgPqH5lrD9LDAV7Op5jCoki8fGj
LGy+4sNo+yTfsbAc9oC84vpiL1xP7VIKlbGp6uz2cRkGV8OgOUpKoMOeuzsJAAun4Ha4Y0PPp/3G
mcDw715dfqRzpoBgxJ9sjEQiAqQA5ERnW/iDmDk4nTgneV9cGnRKwaiIo8TL5N/WRBJy1QKRDygl
txabCVx7JpPdP4dGo5cVj+uxFTUnQ81GTInD0ePMCZE1xtyx8VKqrwLPGjIbl58biq/WaH0vm91v
Hfofjl+aqJ/Ze/F4BbJrHwdKwnt6MVq68wtGfVnSLSh4aFNOCO1hy8++OpqPd7QjNX3WpcHn4dS2
4suSR11F2D82xN5WLL/6B1u8cPht5uIK08hL8gPvbsoT/LkEKhK0lBKFn2Q4KlhX2wBzkSHg6tEo
TrooPd2bkGhVGhGTV+hBq6CoaQuKqf7m2kHZd5hot/2MG5GMxEQ0QdFTUCxRAS0jA1JATyDKpE51
/UFf85XkZkR8Ol9DDXnYQ9ogmK8UK/GZN5GtpDbN/KLKGWgVsxaXg9FgUBO1Dd+ilM8wt9PwWJia
sp2wUV4V0BTMGiFYhO/E2FuA7TPVgPx9+ol8FtzJOnG3ApwQCFXZQJ/Zz/62u92PPr6kmdVmmy/Z
p/tUWccTi02nEbZTil3Q+1K8kBl/3Ll1k752E63qhsfDstugC/7DzCQJ3UiC7tVHU/StnRNwsA42
4yP6TapTgrb6PhWRLLZkbnSI/KZVwDZFh5ym9wxvJQ3JEEsg42L48MAEQwkVVjURAJu/B0nGvWYC
ncbcjnaBVkZmMV/2LR651bS0UfrlhgbgO7pI8Ron5JLU70phrcGcUPcMeq3sMtWuaWk2kIc9XmxX
uD200TSNagl9btSp3/vokf2/2zweoIGb1R1C94QEpLjTmjHK+pCui75xGkdNkp1XZwA/9/IU57Da
koR3Yl8Zip3n4Lw8WJ790y8X4FYfABxBxXsaydfXJzu1AxZfJwry3r6mk82gHSxuxVZy/I8OuVk+
E/LeNkb9NZqCf/SAZ8uAkZO+pzc14MudHVgDSPIOaPySuBK08IIfX1/EyREE8+ubRMC42Whns51H
+8qJEqEBcqKbRf7oc0sj0v5jglW9llZSjLp2m596hSpZ3oIIGjd3fB1OLo0KB+xBJHstsfzmBr3z
M8/+I7LbyoDqUgvHmqfReox3XVjKsbxpTLRtnYmpNKKyMa8zDfqe7d4e8rGPAYFGHMzzHIKYjqqJ
16RDW1ffyaWwgEMhZ9rM6rIrs9Bg0pgjW+FmDIa145RkPxqJoE9FX1OrCV+aFK9tKgFxAmY/sq39
YD7FatHHgmwxgByDRBUbBYsxFhLZMrDRBa/SXrbX3DD1MgYwyb8r/1sNpTAUEzH3wMam6sAutBl2
87Ayn2OW6YQoQJJ10FWNg7zBCsjAOjdYVCTUzxidH1VqwPylduHZV3lSeJd4TNLPJjDxpAsisYQy
t2pHYKgbwAcNZOumBuoo4KZKzukZ2UOKZW8tOmyAo9wWRaGg7+oQmgJxAuIBxSDNP0k6wlPX+K+H
0syERtgALw+P0MZBZ3H2z+7mVG0toi3LYyIvJk/thiZFLjlu/J5saf4upxtiIhIExTE2jgbuPlys
La13F6rg1nKjaHJpcRIM27QjTr5vo4uTTBq0fyfklLHj2+rOLxgQd4RCTif3qDiehQuc6XzkEcvr
gO4h+IckZA8cLEPaa36BJN7GjT7P1yEfIAZmfOy1F+5ST3pBvG8iKlRNO+Vrl50aQcZy5g8q9gcK
IZqb96rjSFNt2wEmDRuaRgAUYbLuDoqHnxPnyRhm0LUWZ4ADC874GnM1ZEuwXXF59eS3ngFnXbfv
KP1TUUGevHT3C69uhkvl67DZjyLR2haCIzvmJTJtgIcukKHNAR5cix14QuipN46Yx/nDDaaxxpnH
sxrodiK+7gZopC3X38gpONARfUmZoAKwa3aTa7fDRuG75w4yPqivRIyiyXP87OflqOEuaJRbYVjG
BablIKCC/ru/QsVGyjiZWGeohSyo+o2cbpuL7w82WHSepveUMPd2PcSEqp5IWZxNLh8uZqwbxSxs
j/D3tC4w0v8N3ljIJKdpg+V3fB9mxsU1I2ceLsl5gRFoLyhhi42TA+Alyt8ViNTRc9DmG5mqPAE6
SzstVOrT/Lt4ZDZqarmZ7MZAHH01dL3yzSx/84hstSHKcAqtOVjQKEIX3o23d/nP8Zv5O2fnD86Z
IGaQvS/Y0gg6UeIozWvea/8FzKOpVAUUffyU7IA7E0mXfoWG3dIv0fZctnxevQ4yZr+n9VgVjJBe
lQ+JVUYuz0tp/WZNQrxbpYInzi4sSem3saoSeSSQnBvGHdeftQNKc2RWYY+Skz+nTijFbXJDvegW
cT/1g223GYRletrmA2mdxEZxjxMHtofzDF2BQYqhsqnGJra1/WkTqFTBYqBxViVQA3zmcrQIF5VE
w9yBS8AP8wAypkRvbPQN+GnCbxvByYbp8f9FkcopCVQcHaftVY9muW17DkwnRkCKNb18pZoMdrVK
C+WM0rl2IuctZ5afFHedVG8kBNsF3EXelYHGIIVR0ZyQjdE2tc+0mGvWtZP3Gt6oyklz9bYkswVZ
NrQUr5z2fJrlcK4Kg7saAvFF/Yu1RBM1wK+jT4pBlUUKLe0rrVijYUHBLW7VOowqkwoRHdpJhFVE
koWrAJ1q4tptwp0AjcX5KhSXs2mws25g2uwLBbFVeGE/gd1ADCY/tOMiqNRkHccpR7ZBK8U+TiZW
ATOhhimco5UzxD2DuD8optfLtMqQ0qZYLv9Y4BrwizSTD0GiLmYv4vknGkoMpPF9qHrOhxhYYfda
AL5DPDoZREZjTLDXw6T1WxoEbggAJU4U5ODmSdh1lm2868P617cEbYJVdr34BraSq3kLBhym/GYG
oFHmqlt7wxXR9pymIUkiROm2E33RouT51MHAVKEHvOsJQR4RSq7m47iuvhFAFJiPHwmThXlQe8vI
nly3V5iyXYJLeu6TUJoeDfYoYw17bgRc++YitsL3IhPTca1UiBQPS7tdVupkaAdaDm6MYQNYw2jY
95fImYmpIoYO3xtCdWGhtAcoHodojVq0pQgM49+DdPPwO/Kb5JaDvYAZUyBGiDaa7V2Yw1GxTBI6
JpYgLp7EgIscCaTz3AkZDTVcf0J5/LSpkOWgISpuaVGMHV/KcSarpdPkZh/Ww2KvHhvVytLnXhY1
pg50qJuNwM3Bm2FU9f+1gvestaCyiZhp1omPX7HDHx9eRZcLScXKac2uRp/ajRnl43hKHv2gEw2N
+lKJENif7pVJKEPWUvqAipxN/8KYzm1Cwy39m2UW9k1dGjkgtEIAwC/4zDMHjKu+Oet4De/Xl++W
yefX0ULE7d9YElW6QiB5bkgbjLhrO6wdKbe/kX+eMvzAVTWHwpg4JssM9FljUAugB0IgtMG6dKvw
Ws0s7WW6NDTP/MAOmgOe+JMEeK9Oy+YO7DuLiOBqXyR+SN2d5EUsLI/xQogQEeDRTQv88wmhK1ii
aReitZnLO7kTCVbm+SVksfKq2vdjG4XnawWNMGsmaDbj7HrMqBDFd4uVBNcQ0HVJCm4oCxOw+wDl
dppnXCMqqk+pRPe/CIaGiMyYdwAQLJHQ5lodQHrlzi+bAjGbFAwXwl/pQP47cX9IRXNCgBaNZ/sS
Mq31itRImoCLJCfTOON6K8LBkv8xMu+NDKRfnJAtehiCJ8TJPvdyX3Nkcu0H/b0NSZbm86U3sZUf
WO+hs2wdC+Om72xOD5Uop4wPtJ5RNVUpg30J2E7o4IZy6J3AnPyGIYM+VpRZ5DVecTJQ6zoYlkHC
VBH1SIdfNDcRtmXU+ihBlhcjmDVsRMAjHRQjSvjStVcJP1NX4eoaA/AIfmoidDQwdkdAH5yvuf0F
RupjBZXosWlBFYXLgQGJ6HbYqlVi2zT6FOwnBH9ko6yH1SsZ2Sd7swGCDqCHa2oLq9+eKZ+ZQRcx
QFGwaQdtFxL2KK2cFTmcTv/zvJveNYnXmMKOko9liZraAKea1/O6jGUXz/+BDIgNLo3zVqihBb5e
VPYZmgyn5W4jFYSYrKNfQxiJR2dCEA9UZoVhF1/Wbbu4JxaVGs982KzdrHOPgrgoACkng+Ww0jYl
4ZnaRmDefC+4PhTtY8DeWmcw+ZRczEdBwQMCrLdmmFLxDNbgLE5kcTM3cQf2ScDDVbwOiw+qndgT
mQl+GcliVJzH8KNplkPQZG37cKMwtlB8mhPBQ2wq/0R2YBHIHJM8K8FlzhSoFx1DEOBnTnqEIHv6
B9Us9NdFViB/ioS+qoZzX4g21PRKWG0hnIV2Bs3IH2nEBo21dUex9xPneSFi7uWHiPeHKnlqHgGR
Xz/ifShcBSF26YnbF98osbQ2x1Trb3NHKS6nXRxxYqhfZbDj83zjXJregaHzAqxzj22DQfYx4FB4
zAKmXOuXS+z/z8PN8e4L4gBBOBlkCke5h5lXkmybjnvjT7RnEnQJMRfZFBuGos9/Rj3JcSMqsAjO
SP7qsVg/3BD5MkXBQ8PM0WK91UAW5avSHAJKY/Ry02vfakZ0ySPB7wujAJLk05MfDtrjYr90+z7c
q5cynun2O7KNwNG6nu9Pff9i+XpolQFEnvKr9s4BzqpcgIxH0an8qy3arjvAp5TNtAPig7JANm0+
ist2rPofZFSydVXtFKafRz3sZ3CItP9y/GcFVy/gQssso8nAZ5s2gpSgB01mIIEtSBsDSqEa8yXD
BrLezOhbzcKsyTtGLTx0YjbcKzrW6eb+Nb6Lxbvh3L13/h9vWeRzcibUk7qS9Jcx4I3mmt5cx0YY
GIG0AvkFEkTgjbu8+C1RsclcmwpQ/XWpl2XKzw68ERYLLn9SxQ9oTxJX9pFJTQHRK+bt0YBGYQtD
4acHFbhzxeJheUOOYFZhOUQGuAefiBwU58hyRiqWyZGMYUee3yXWjcuTfTlRHakvIu2JdCMZyg4O
rooS57V+RmiKlja523Vn6g8Kt38I38h8QMUiymWrU5yNYRaDZ6q4Qf4U5LYzohHt2OGDelGrzr/Z
mwoDWrGtDoLZ94wkrMoS+vVjhUudwJCOZI+e3F4MBUtqYoMwYEbFf7D9loRCx0nXYPaIy1E86hzV
4JqTz7cMV1THGhsVzKcJ4RZbkJkzq/1fYIYJYLTW8EW11Fg4r/f9Q+V0n/7e8pdIlTRsaYRZtO9G
RcHF4OEOeMdJmj50KpPJkXWIg1PfBGBnPsdfNvWNRJJmDsQBfkyvNCbwoj8jTJVgs8spdlgUrIKs
kES1wExyj4GD+3jv1gLOm/NaOnH3wBHmqXq2yjulyPl1IYltfCo4FhdynCxe9eNDx1RJylQzpVw3
OkoVBZq8oaR9QPrLVsGyeiXFbQvhcZyPMqCzY0ZsPD6/kifUQgLIQbQIEAgZX80k5ZMQN35MVzsa
6i5qNspuQzEj3ApEe6bdLehJDQQ+kWGNs6MggbZ6F5OpDkIq8sLkhNnxbIQx45AOvxNp8C1Ko3J/
jtVKTd6ArAUV4ERctnSjqHUZZnKhAWHC5GJQm+m1MzUwn6Xc4vCJ5wMTJ6psqR/nY5isnmA3L9J/
O16H9LHEwTN5eLs8eL86+N9magJjm/5nGroMxI5DwT+0qABepTeVcTPNnSgqrls86xvakyD0YmoI
nQGMUls5GZ3wsafFPl8pgj7KQikFOlX1J7TNNj3mGWOT6uQRhy/FD/dTTFflbv37fwUx6fY3vBlT
0X42EYg7txxMW512eq+q1tXgPlpL8C1qfJdU7DGGDEfGygom0rHKIlSbY8Y9psyS+DU0p7FXn4bM
dXzaoOFPFP6WmuRY5HlXiiJuWiued+7JM1AzdCn7UXRj9Olj6Gn7FGjUTNmd+QhfahwYstdxqNpY
R/N5x5DIhfDm8OGXI0KGJonva16ZFw8i9VW069DCO7MgbmiCv5dj2YGyfomkUupkmNvvxoLMfXxf
E5rXp8IDxGiW7ft/tvCsstCKHTw1Mq8izfALlwGIPLiQxrB5t22jVQelBJoIY8WjSfGzVf85OwHe
E+r2UwSRDvfB1f107c6xaTg4MEWK51KGRCap07jN9FVWT2KrGIRrd/I9LJGAs+m6xFMk+lC1OfkV
m/XVlrApuUDmX5VfCkUZnZHJGU0knwzFiNSmsFtg0g3p6NH4ET66znqPbt6tfLJPDwFL79k/FZMs
9xT0kVUUTjJcb8YmFOMOffPuxUnbG7D17QsKCVzwC7G/ZLdPoLargovoq4gNPwC+g0xzTutdayxS
UNNwsTGypfks8VmwWSfRNKXY4p1Y448etWNYlZd8C/EMSSjXObX72w+lxqZJgSXkuKA2LTwsMPNR
k5g8Vy+WwD/qKduF61LC7CdIA/KrZKWF/x0mTCEjDUttkzzmxM1+4z+Qz6+s3m0JkTEn0YAjBza1
cFaI9TdFoLIO2xFS5dhT3qAbc+LNcCPMzT8FxNxcPYeUcMyrnILj9D9f1HcY1zhtETzc1JzAR9qr
trOBBQAL+rLHX4gZUQOxEcgAw6+2xqmfvWYZOXEwY1pMZNJr/KbWB6VbhU5V/s1jGYPHeh8TQDpd
NzWf9JD1LAFcTj4ASq94aU1Tcimudke/5nQV0mxkL822PxWLH6uqwCB2QVmnqmtAqjAJltIErBEp
23Rm8jz9P9Hcu5b/Q4kVeWDYEXbPMrQQ4DEHlnIAGuY7bMkvhNpAvvK40Xakp2pV2SlZyRAUj8Z/
jAVeo43aOvhjtALli/Ui/8RPvSr9jAZldIjF5IgBnWEigCYNUlSOS9XoJcM2PiZlsozX4N8dDJbC
hVvokEXHVWpGhVPXjn07cGEfApuoynO5oGebImReRXjZCCtceuN2UweiOHJ2lZZ369bpvGNdhtlA
HsrZN2Px0qPoKwwJ9nXO6Oyi2ZxiSJDMJWGJpn13Gc2ByCVECnckZlcxu+72LJVdj1scaXFn1FZB
GZkMX3F1YFetDeKwXA/26TDwq289gqMHPe2CAXtn/+ZzCMEZ9BKZ5KKc6CyjiP/69noD5RLAEWHK
VaOAM1OY/7gzXQVjOd6jLtZ1fZ3M1AToJRCXJOET0aT+akdBr6CRKq5x569VSY0qG6nbKL7q/ChZ
QpBvi3K48806POXLVJcaHB5c8SqNCpJzOi0X25qY5T/eySqAGSjfTMIxRZW0C1uY12MgmVJP3IAa
KfPtr+Mdl5SG3VfedC7Kx1wJcoLaWBx/VUHACSDiwOzgjoZjJ7aXpQD8zs6OyR6cIjngL5fH66AI
noNVuUqbGAUql8H6pWDV0wilChxp5QaHbYESRxK4SaO7Mj8EIlEI6mesBX6kHOBdGnbOd1Zt+cha
V1V/yd/f8Jql+xwcwSlJl0nb9x+x/wX0EN3PG3b/ghZBJ/WL4yfmVHcnlMpFAXW+Jvm0dZZfaOOD
S2Be1a1ghTRGvcrrMr5rRteCuPFPoH64//+uLOYt4hKegxsgVdab9hfklynDJqDQawt2N8k38psI
edc2y7QGQ3oKSlBt0Z21G+QmpI7WgGhQMtJJLvlNZSxtqpt6TlMzXVr1Svg3IUFT5juBHXXzDV6C
ihtN/5CGRzOOjBRSm0I8yiV4vaS3HQvXwNw+zZs9r45tSMbo2AaYWqnZMk4bfbzUm0D6URp9VOsn
ZR9knW5uB0q98qyDyFEFnXrQ3zmu6x/O4ix+OohavfkIRvkM6U8SfzFUwGJ1A8LaAOhS0+ie4MmA
BiLCwNBDQ6KrLVb2Q00Mk7/wE6XKr+rYW8LbdhPETOrvQgGOHNN1vdiyqoL73tK+GbQsiF6C7ehl
aTL2RqDXbf4ffLkFTWUAx2W0iyW2kK/+nw8b1mEUpv34r8vPV1rvtrkbQaxJUUjTQqm87qIKU1cA
9ew7yTAxqHHBPRlTkq2q0ZLwfoO4GcM3QsEfnIl3GSgNWNpQi/WJapkvZDLAW7Taf3N5WOXTvmON
EDWsjyGdGHgHJCrhfK4CAqedNKVpKhtIUo3EL7D26DHCqxm0DIyguJIXVG4LqX5Q5VKVoP+x9FWn
mX1VyFg/GQ4oKsDpuaDHCFIIgfU5lNBjJKCn9NzbMGI3+46eBDgbFgcT+es5+dBd+iXzXyR3haYz
faj0izoFm+ZNCbPHGfdA7RUI5bIfpujEjoAjONGG2RNAUx3URa9thlyAACFmlGGYozdia0ORz8AG
fxFJ0jKnTETt7urwKMAA5QL2rgBbIgTrm1y4b2VeW1HK/YVhjvFoethOKkavl5pFYbnQqH/Vg2s5
cteR/r0xOeYGxzkVfbx1RcT9prFwNQekwuW3vneq1Js4EhDftmf27CvZjTfKkJuoKYF92Mf4R3HS
nNfYlmYBWt/ns5XTJH0EGwWbSaXuMbMIM9rJJBovwIiso5QEMOK76cCQ0RlcsBx/bR/D0sueZZza
exjQeS36jcGvB5umZmG0Y2d5fdCe/CSJ/69Z5L8WNU7XnTidZX/V8Af4Z8HlEuKAWyQsB2/6OTnU
C1BoZxQTFrvz50Kfz9C1QXq6WjLmU0oJw200QaPk0YAaOdxTTLMP/6UOzdGTAvGG2t+fUiczxcsj
TEgAORCboP90/hoDdds1jKNY3xlYIRh07tW7HcQxwXc5Ee0YOXwzpzy1oLZQWdl9y2dL7K+vEFzR
X6HRIbpr7tofiSP40QSOuLSRRtqvXq1rnZDIBVEklzuI8SFdLIAsTPNFbYsBHLMoeWh2+CkmdK/s
zXvIigPU+lA7jiJxfFfYA/rVh0sy8SwieIlTr7XTSzdlzRpElrSgfos7pIw6fjlvt2NxiKPUljN5
CYZd1grFJuODv7x0EAKfiGUUlHRTTk4tHFts3d09Yh4d75PqjeP6dEf9pQskQpjV1mrOf1UI1XT/
b80WfwUXonUIRNlwzuA14a7ksJlcB0MgfEMLoKJ2qVrXrmq5VEc7EDo1XvC7LpE2J/5ZxskooXYL
//fXhBqJnFcebOFgpJVXylNLXZ2uWJktenNIoySCwB9q1dklYvk4d/HrwaO1dnCU47cGiEoMfPzg
G+Rl/9WI7PnFDSRDrnNfAcaaa25vECROctQawTs6vgRNR+qHdRTNX/9Mi6BB3XMXp59nMzUwh0dY
tdpIkVTTHZnkdo7Sm1han5TqFUhdE6PqiHtmYiJrFghUo2ZQFridIoBuaLzQ5JNBo3IpeodEl2eN
G5kzex5tLlrvmDfvZ0RkgawWPfDf7yUTeujpQXp0t5VzWW9eu5gR9dyC5qicVXVwA+mqQngMjG3A
ilTXZlVFEIryKuh1TDgwRoniUmBVw0tyrKP3PcAkZYWPZGCebchyk0auuX6BRN3+g51GZ92/gNGY
XNGlpkcKxPNcYS0ul9CQDbYwD/3Ik4dbkAHDnUMlSmUdzQHwRZ+anhlVxof0g5OPWZ4wFcRUL2cK
gkTaNnBs5GCal+0bsTZTrZ6IKIES/5pWmANMMbHqGrbnaYsku2pB2lBiqkI0XqspOMjlkYs3bB0N
QVigPkvFPffTlPHxa+4O+HZV0y0Hw1IxoPojm6nVh6Ua42QnM+kVzkIZNNUkcmYU92tdqDiPCjdc
Q4imJLrse70J2wx8Rxw/nyKryyVKSLZR+MoACvlwIu1yAg7LzLpwPH+hv/d7oEPPh2FRYPp4a4Fk
zD60LCAzEe0Efz+INpFGc/oaTq4H3zlb4l3s3y8Kfi2vbQUUQjfDfOqlnqhFQUm+GSHXZlkIt0ow
gFphuIDKZr/2U8WJ1d8l7oKB7FjWjnXB7e9RpFflWh36AN+NDsdxpmbFSauLk3HbHExa3GGeOpl3
aPg/0YXsNxV/JgkJO2GELmgKQvJjM39voFCPmItPVkDFxUtUrQW2igLZm/pK6d5eNOMI3qNypUyo
Lb2zAOmFsKQPNqXRAvZy2hjP28n2+HHMTHXSaz5qmA/7QV5+5sc2EMeFPyDVJmWEW0gLuRWrW4u7
ewKt2zs8RHn+yvxxFxIvXxTxRWy2XgkdemC8vlXZo77/NFT+STzynysxn4KiS/oj0/yM+cuVom33
Dx26jTEVfOTvnWsZWH9c5H6qdM9oUYWW/sK+nPSAt5wMISw3sW94/QN1jdy7X+xZWoTdtiLWFY/+
BENlcZcs9AiQCTkBtTgM0O4KTlOLEa1+NqC2GFBfu00NDd1hqfVxkzV1Iub9JizJX0IozSzf+gPH
PvGQIa3xDqpM/BkAxX6mzIp/oHJgXbSz41SbhnQ7HPAah2fJUb8DpOe+7vDEZ4TUbf9HZx1AyWml
UZIGyRnsP4vbxbe/VOW/Rpo0+5yd38rkseEFhL1vFt1a41A+cjUXeDxRZSzt8EqRBP8s6YlN4cl1
wtgi+zqj8Wn5hfjJLVPMATw/K9MEa6dykqYSTLONWyrGFP5u3eD32XvBEnoUTFL5hdJyrAtipNd8
WE7nqOpCGQCnOcEl7a/g5LxBiHlptkDQJrOYMgKL3FwLxmLdHGvWXRDC3fuXxqdH4aB8nJEn9Eb7
Ynxx3pxGZbkG7u0cm6UKzXGDd+ksSJuekN9zOGZHoKr4rdz7oyA/0FiBRQRJqBR+w0wG4oE8k7OR
yEJFYS6dWOhJx6LQ6Gih/L5T18MwhY5hgophWXfrGjlX04AYAz4NHNtoPEaXnwslr9WbAfzxT6GD
Gwr+/+7r44bofIA91iuanxAB24zK9vCCHCejbErG32YDa1DScyKg9nZNqM55QMNmbVqpytkmjd6j
kBQkpYzWZQlrX/doSW6uAeiGMxcTVuug55tZvhySaN1wh7mjg8WSo6tLkbR/aNCvXl3UOBDBGvK2
sLHFXqz94W9kTJfDhnz8ZCNer+UHP5oeDPFEyNhy0wbARmAASn5Fad9jXJ7/y9iKAdTa2Guey4x6
fv6gITa7vJY1bk+69jmjnc/Fyz2rGMVtVhAub7yF+aZ/QTm792Knc2+X2melazwQkZYmP8NftnkU
1QxKwo1FDENWTnJjgOajRQstz/DOP9quR0xfMuT3kBEsNQLO6D6IcFosThIrIjsmYzZf+eYTlXu6
JUKWSEHvCQRWxtLWMq1WNSqBiaI4qTOBMnQ1S0VD2K7XbFpMAekel/1Ys6pZ9158AUGb2ZCdK+5S
6u70TnBWQWcD+78ummJEgCeGSe8q7PuX/nJsyGLFNrzUGuNLd4SEJkrtG6ZZMXiCeeNjHn9YzuDb
Hb4g1ojGb57M8YielrKQUtfvMs6vWJKnR8mJ4EZu7qafKXGkskCjisYCrHja68VArg+eHnUcIAmI
QP/XKwyX1rf2WwqmI7TVBCgsHKSp8cHt/EKBgRXlZn3NC9q8Mf70lBIUHNcl25pXM/pcIVJZxUH5
ei6jS0a8U22fQIZutlSVMw/MK1eh9d7Gggm4ShCB3CkZ7qUtaCI7NVgvKOzbCKqAnf6FyVeI0pq1
T76GKcRvw8hMG+aw3DYCuz0o9ur6qKUbbMMTNPJMp7DitGLOChcL0VnsH6PYY3Kn4OyVBCj/qxQp
e16zBdQq0MqyBo/bqaTM70OU05j+rNPWzYsSiQMch+g1mC5l68cdLmhLBuhSlpfGu12qReZQKROF
JTxgUaRo8nggKRts6C8FexWrVTT5pWmK13NciY/vbf6ajOAi7fE2m1O4qo9rTC+2DC+7UH2S7SCg
G0Py0VgW7S0CaRYEZWjoSQ9B8OSLgPtREVUFE1QPJXFb4hZTHJFBjhA4FiEi8J55gTtksYjXBHgp
IGtmGEL5H7990HaByUC//9HiKr3lAHnhN+1Tge/8eN8U1VyGoDMu/tTj2H8QCosNY3ZrzL9chQuU
IFCrFBfM7F3xDy2yud0IgVvg7WYxmpSI3jfDfA0zY8h5Eo0kV0481WGyvsht2ONz9+1kYbvDjhc5
nPn3HXEFotILV0BJnwlCcTGOFM6tm6onPc9dyVvK0Gkc5n65S7x3gCCVhP0HjgcJYf+aBxNiB2Ya
Ehyxb8IVP3N5cvw0u0wXmwTyycURoNRQH9cDFe9d+t0MYS38FgrfWwtlz+/eD6YRkluKM9/brWwG
ubajkXCZ6qh22OCSUPoX/0uDCE34x2j6pkvK1Fk3yqj5YkxIt+hHtSAAXrBYOTBpaJPAw5XYZOMS
iH2RE6UFzk2MilRRs1abKoIcUzdyVwaE3cBQSq3KB+9+tiXNVikz0k1xhrZbSzajfpJuD2FI0EL6
yMehn42VIFj53+DW2huhkyJiIq/DWW0mM869A/dE2Gp2G+sBCGWyIWghq2kvmwFN/JOiF2oLESby
t/MjCMNKRfgl7ux1GPRC+QTTqXHDh0i6nKaCataSqgZcCt8wNLrr5XTchtAUDUcl41iIIqKibjKR
XN17zBRXsPV7O2oRr0ZOspZ50RzP/TzyU8+cN2zGDrvsmZ9d79zlcYMOx1eTznKPsc5W/7dA7ShM
E6Hb0nrC0qXkBAqDy60Bo6Yt77Pj9/KFRvJil/C1CwFOMLCZ0xF7k2791VHgKcd6aKD0QPlABbb0
QDslqp1ug6BRQyDFdvMJBecG7JGDkFLRmjXAa/sCOoNMovHwAWyhiNDmbCfnjpRabhGFm8Kjw+Q8
UEYphWNIbpOnvtYf5mUuejSL9bFWhVTv1tsTkE8y4wq2gmwhhrLUtVcqXpc6GzibCTHA15ovOxRB
ZzMWWDd/Qez7MhtjmyV1pP1d6H3AYhMCvjPksB3ZfqkpZVkUXTob/VlqNnpUiE77+zEe7vZ3ZGjT
549xKQTuvwqhoIyhZ5jLTNP5Y5G+Kn/iXvuTC9nNkID0wY0rx+Xx+jlbndfiZPqvXbwQaQL/GdcJ
2yqtXAYHhOJa0W3CsJj0Y+r/MhQd5kyUJ76f+MHOwXQ3i5O6egIISaJfwmW+W6GA+o/ECbMaxMKv
u0uVC9Yn15iQtzTUQQH5Vg7l7dfdgh+zP7lIA2wX+PGE9YLzdUBnreQ86RhguyRXjs/UkiDCzUnG
G0vUZTxHvAG3GP313yiZElSMTbEFJW4y41NhGRhWLsP5mC7YvdMFhsRdEZL/Mnrb5XCCtkgzkZ4s
bAj8EqFPuim1xSB8nThJ4KdycC3A3AANjvhaFXYZlwN8J7a6rwmkONfKryn1puGCzsLbdlwrJv8H
ehGgyCpcM7iJPNqYak54hv7h0eXZxaW5ZSR63OpxsvrRGwEtTmnoaWSat5e7Rr0ZJbJaZ3yrUo81
zv9Qh7salPaauCQ0Ly81mHeJbbjZO6z3mTOKcrE6bIzwp+kUjsCUnYJ0OR0wP5YfKZ0E3uJkszGv
y6+uZXMmDwsG2W/xQMIvD15lGU8g4F8e1hUlxzxGxNeADMfZqndNcsedUuA38ZZDZFHyN2vkryrq
BjeBTxsL3viPfEvOK/nf5c3T1jZG2tPJws+TGecCqcmNIY8e6d8HXThUr3tkhx0IfudKwwluzciy
aUbwbMw31HSxwVxUramwadqj8GXdPzjeRanY7czRwyVXtWRx12Z3ruw2EFv1RWnPlyKN0NJdnTJZ
U+7khqGz/Q7jtkFNWO1Sh7bGQfyOBiLp78+Pfiej3sb8ElTpHZXzfHXlKACRIwoHHg7E4MfVM5jS
zpDoGMOrpYZ8Rco3NHWH/efvCejgbUiPQkjCxngsWk9a45V/SS2xYxTbee31T1P/cSEgBMri1Lz4
wXZgdka8IfkUBWrbUQnr5XEkc3vMAKEVNOBu3isz3zsuE25a1jtwRy8KbFO9iW33HdWMyPhMd2X8
t2zDK7ySkm0EJiw7ijflIyVwR4E7hbjML7LirnwU9AdFvNqsWy7ZO9YgzzSTV+B0AODY0Wlp2F5Z
vBLlf97UumyNGXyqjyDZ/DWwAW2oXrY6yjs/gQ1Bc0oht8GLLnVS9QQ6hp7LdiC0qnH2SeGR7REK
vzSzPC+/mdNmQJxC3ajdOepe0447J56rvFtHUbyETnfns+bbXolta8/cq2bWvead3ivk6ZXPS0vh
QRGhgcXstlsMuPDdMcZqyOVm5FSPK5+bWdT/nXJWiFXrSoXiwUxB+gCz3rCuYKJafRWtst64+CF8
pKH7LPke6etLS/dOhxrqqYU7uvqg5Rc4/uIwGeqb5ynG7gvXmgYwked1dGTecW5UNDcPDQrH/H9a
kf0qa4h8Yb6O7rFoeO7TMUhfKYWARZ8iJPX+Y9fA2A+mAr7DYhd1O+NB34e8XYXmxJNGkYgyIfpt
PiuKd1TNflEReq1ac8K867eDc5DFAu9cIf6LOdLgoTLkVuq4HpsiYnekV4y2GeZNoBAprX5ka3H7
SA0Fnv1hm2pdM2fleYf9on9jTZibzdre/RE5EQF+WSBlYUnQFWk2AjVdbStptQOWDmn5MjPAHSIV
6cYI5KNRermWaARGYF2F8VtAcxi5rGcBAgCkJYOprJ8mScXo6L0n4ezx/ieb4qCpGqUrNLh0f0Fg
wB33g/P/Pke17qJX2idCRsfkWNO01CEZKIjfOnUh7jRZTphZf61/d3rNmBekH77GqdITZ8M+ShFE
Dfhz2csqQPmbJYup/5+JclBgHm4IukvDIvFjnutf5HgZ1N4GBWwTAgzz1czctzDSe2TLzALcJCEg
DNLbZopXl46jIMmRO3kq8rVDyph8vjpGwbuDNsU+DWJ3A0N107Fql6pwJFfrdLxbO6dcFRnpksTC
3JsRF22LBiJGXypmEF4qRAXwWgNnQJPV4jUSUducX9JUq859RO0XZBEunLErOOJk+y0o3wD37C24
tliamPwnqJlSbEN3V08XVIyd5mbxKgEq9ZDb6cfNOfTR1+CzUCukcELJp9/P4k0gynwW2Hwfd00y
F6FaSviW6g250Sn3efKzvmmoMsucs1HGQHu6B17nIgewXEI252wJBlzJVUNjb4n4znVM22JBzhcA
PPagsADxRHm7M03gWl6wncHlPI+iLnt0tAqr2+7Mtf+TIeTNdwc//odaMuwGPMZWNVyZoRM6SxJL
c0Q9WygK1iphl+PFbq3H9n4pBR7W8OctTp60z1XvlQEhmANzeJB3zDcnMZfPT8YozSoiBJacWuWI
DCVIBRcXcaJZKaQk6XL4X1BoeQoiPapLZFro5ORlHetaTvcj50a3lWet9AbBejTMD9I5qi4xZ8sT
smsEdYppmh5AN7Iv0EbGpwAg/KglG7cR/JuNoqC/e1m8C1CblDPomUycO0RaC+es0JhddNTdGbW6
nAzhFLRvxwLG3OGEHSjfsjnWgRwfYDCTYcUQZ+3uSFe6FUiqjSqlYFsHggvltHK+KcwTPRxbKSdD
EGQzPOGAhoIUw5GbfOuMWA71Izp+WZWJQmXOM/N5vUBV+x7hNMkkuzqLvohkBzx37VevQkjcM1XP
6GwSCWc6STZh2IM1jqzngtOm1yZABRHBkM7zY7NOqBYDQsFuvXE9Qxr/nKQ1wo1KtmgSnjyBEcIW
25b+v4qcYMqVVGW47wa5ixP+27SvvUwEzNpJkAia+sTRQ9CzWeagCDVdfqCFYPH3Xu8RKMXyTrUJ
HG87HqOQQKR/GXJBMKYcWBDovrnCueQZOEdOGN4qkr4Gg3pDdS5HOw7KWE2NyqbRwYoUL54e5pLh
049qV/g+baA20c44FK9S99cUoh7966PeX8JEi3Rg2iOy2tJh98/2QBrQtFXZtyLqPdLFF15bPskQ
Ys6jyEC7x0SisXOvUjyKWB5ls5tyn97XVBpkwf7zUr3C3S7dFyM2zziDZte17uM/x98oZS9Z6JR0
l6tDZS2Yv96fofSyVLMgPEKmmeoAjXzcxEG9lUDxaI5aw08ujo3ySGkJ8qczuachJfJHQOOYrVqt
Om2zFt3K6kI5IrHMeWXoxJhyJ5ohxkpo+XEgvpq0O53rhcj8aSp1N0jb529T0VdbyWvBjtGms8CE
J+W6emcSz5fEcE+vpdXTG4CL0/5OEbubtJByJj+zO/uZ3cNLhnzmLW2mSEibl4PbHANl0aEvCvx7
vxe0xVgUnKgzPZxpeQF9fWN8ypZZ2o9UQnFGxy5Wytsg1fAutJ082mEGVbLoIcWMVXuGyPLr+hkn
JlyCP6HZQJ7uzu0Dy5o+tDNWQuAOftHhbCV6fdqSDkBt2GZkIikebFW2BVQqzYJjYVMobVux9+Fo
y6j6S5o036GL4pbRGDy+sXLzyJb0/HSuaS9oOALti+q17ME5cp59XU1vH1XzJ3+P2tKBUPJzICRv
1ftBqw+TPTXUYezf4DgSFvK+7HEyQwltjNhZdSrAs6lt8631nNSWZabcoptrO8s/rsZWgIitYRxb
g1agMrfxIgCHBd6Z4gB5v2ah0g/vOExQJXi0RTswGxUR5Ph/TqxadjjEVFoAjsPOoxkZKFDQTEO8
fKzze3LlyTX1dGfbzX7ml91ChlT958b/tfnVpfiJH+kWl90eMTxs245SAknlnIia+1cd84npDrks
dy8zVhrR3PFnJQ/CP/0ih7mu4WIYIJsyASvrzBOOiTCuD9S+vbsgkOa0nxFwBwD4U3ZNzyBtloRl
RRE+3aD7V4/e7Ktm6pm0dMR8I0j4/C6/QeV4XWHERwiWaWJ8O91+0BxeUJ+8jzc3odwfrJeDrD8n
U0HyiKenuD0XFFq5tUiWm4XVVzLMqaNKmPuzN4slC/NJwbJRJ9hl02q65kf6q09O9bs46vzO3vZX
Be6NMCUD0E6iou+iGmZ+jGPwGnd3OtcGAAdmO9z2JB8Ah7rH25gla3uEjVH+GkkjqunGGUP+mwhV
eNeDuoonOR4DluIcLmJUX0JC/LZo8Lr/67cCRmNx8zElmGitfaX3HCRputRgu++HMPt2CRjxCjX4
7k2zEGzea/s/nlxHcMEz/5/i8pC1dDzOM7eU1oRK7ouu7GlHnvXi9QJr1vrbi6uT1hLaKk+4ElV/
UOF622RipC1M29WXLgdUDLLahFr2MqAW8CbN6qZeAUhyiEfxRf005Ok4QNmg8w736d6X7MApd2qj
KVPp/EqPtVBKEsiQmd51++Z+q6jNKzm3EMdwN7QTc5Nf+H3FeST+79YnGmlWn4ys6qycejDDHTG8
wTcCxk3ntwwQlOXc2UHqMe2LBl2G1r4x91YD8ErdYQ6ASHo2f0h9Z50/VprG8RPNK7tHcKwBbnAx
HDiAQwrqoATPIRWD4voNczSPq21ko+mqneMYT8Pmn8jnQAGX5K9/Xpd2i5UHcbB/NXKGlF4q09pH
mznrkBl2Y+jTZPPPDB+Kt9VaCkhp2HR3yP5X1XkyQ92L8lHfXAjSUXozVdApshn4PWd4DDWr4UM3
ShumJKdrDyPpM+NsQPGwe494BbEfofD/1vjk41zOTwtHCJy9EZrcuTATm/cp/+Y05i+Bg73BCg8F
R3V8i3MGSfpeVM57k16JXOqGEdDZx/a9mByIa2b5YHLQfNULyTmrfCIfFuBP0XbQVY54InF5E0Ib
VPhd0Poul8uB3/VjVyNrJZUhdqvZmDHn0gsttbaW2dF5otkJyaUQPnA7pOY0HZU9PAX7yWxWwZjg
Po6kSUp+E0MZEQwwCSdc310kxaRK31oaFsBVubyc/KlG03xDASeGqhXmZaxaeCLt8qPC7hYNhXbn
WfYBu2JzjQvlDDefCC0Fp6N09HsOwjt0f+z9CRyB1w9x3tMNNnMou7yq5Q67Zhlenvv/JvV7SUvY
1C3DZ+EiqhAXk8xvwGJNgObzxi2CsK0NFjXs3Ad18AGJvvAPue0FRa0IpvbDyfpa8CaaEzNwawVp
nvOh/5GLlHiVmudr98s8d5tb1QT9SLNHh4KS+P0APY87WPtjowzFokFKur54EqfJkSMFf/Bsiu9X
ZMIoZ7IQHs2Q3lndy7R8l4CvPRNXH237/mHt02cV0YoTB8wHraWP4EY48IRPTcjefDTo1PmZsQN5
0Oma4+WXLW+VdGKqbAXbpbeFfgqqQ8wWRnvzKLz+0VTEucpOgb2UezFgHD8crNeb4VWHnE9r1iwp
e+goqmVp83/yRbSysrslgmXbu26bX1VEwpH06+xlcx/5mgOR0QG4u16sVfITHgxVXoap0BBZq49P
+rJmKiSdgiTyXAAYEpu8bI7PEKdHgkrlVrnweq/uX3SSmC59VwfINgw2O4B+yPUhXnWg1o0U1kjW
N33FcJG88RO10T7/aLCDQ40aL3e1BNhjmbshETw5qS2uwA4YkAJJ8w65BMTGBVhVIVhd9mrYxtmj
NRn1nT0pAbot998AyTDhjSgEwRH+sSLltH/14hMWZO9LJwsoj0nAuDLgDWsSWV7TRXTLl4w7FbDk
JXJyfcT/9yDxq+gidP1WOWgjJOOdlABmSnrtPOrHlEkSIUXH51DSnogdmgzmfJbaDIhFX/fFzyjs
MFUCQS43kYcymLR6BMd+sAlx+4MgxGFU6jgP/7aZvYOCdmfTLW9grRnbbI0cfgMrch1hMq1oTgxu
a8O8V959FUotf/eNuXdv7eKkI5ZwT1gx7/4W4HrJbSmc6FCK0wNiaI+HtVKQnL+vIq+7JtSN4L0J
mqW5XNgePnE7ycdz3v6dAN8Xd/RxCq3jU+8cp6mAtAREY8Yoob2vSfOkXy2oT6DRRlycTURLKLT5
lnTf4bN5PHaNCVKYtcVRpPdmSiBVqP+STT6oSLJMmzb+JxKdDvxdr5ZEk/uht6a0vIjewBK7SSfj
oDrD1nevMlw9vCD+9WWxDCbxjhzkBoR9kymGjsZI1VRv/6HIUXe9xrm+p0Q720CSjP/Xp1yemzSQ
yoYx3Alq8i9CAOqVFOVZ8o/14xacES62SSHlqZZrexNwXVxcJa78Z/v9DIrKDa6/a4diQK1cl535
9Pl+auDtH247NBQpUlLU7iD9VbNGWabIGS7nTIS5nLnDDWJp1hMA0nri9fDen6vlqta5JARPrvmT
0GLgTCGWojtRp9kgFizSMxDm5mqZUKzS8mkITPORj79awUghbOx9b7UxqKQBzauunt8vPgV9otJh
eriB36TQ5RHHN00TnUy0YKCz2IODfi5t9GTCOoPz9VBzaPlSNPIaHlHrGIibivQtqxUj7U2mQOtF
GxgbWzrdeDF6hfefr8LWls1TeJZfqGFG7Pe2dmRHBh4aO4WQ4q/fmuX2GlvjGipbRVqgdbrt+l9d
h0wEWxDelymDreMHvGUwFDif1/fbeD99Iq/rW2tIlXGHdbMBjTRCe1V00eoiPX5USPIOAuId0MLz
MdCbFkt06ha7vgzp+KfVDdY8D04W8FbjCQmAICwSkQqxhRbBVTScp55U4OnX5LAwU8xm2X4k7MGg
tWNWlein0GkJULwZCfZD8SIy4riBhZlqvqZQer5apKxYISgtOjcFI2CahaM1Y125IQ1qJlylfgCg
10bWanzdfdOVKJQCFQGmEh+0HPSg891TX7UmblOw282fQdBLsYWSNlPHjIjVb9uBqHzmOzliA6SS
4o7aZLWdBXmhtFFY5hYtMEtstvQ3F+/Hf/zFjLATWaTSH18sCogAda5UOeZGbTTV75YTxJwBxfmX
f9eLQoHY6Yb8OoC447ZuISTozssIcFfHwFpmgHQcIjOg3vgS7Hhna8XaxT80ntshAz83a2rdJoEK
Yx9HhwP01VjHlWN9SnGG65X5bhexFwjWoTuDnzHfHiO7phb/yiyLfmfymLXNEo0FU2zMg90yb41V
lV2ZaxWFAfS6hfcyK5auqxuT6JBAz8RYUizPiuNJmubA1MbYPKeVwnL9TtXDQZIL6ZEQoH6L0i+v
LBNdopS0Orse1c78TT5YnTxWbZpaw9hSYMFC5nxecSxgmdHqiLCwvH7R87X5mjASy23C9S8Dt1su
RoywJsvT2w4ZZS5UitcUMqdD/jfxkbGoTsPfCJxrZbWL8ovGqp1mAfxzFKpjDl6pWTJAt5KHsU8v
LhEZXbDWEUxWzQz0buEUX7hro1lzeKpH9XlohdG6xHG+4jIalEPmTYNfeOnBqjoAGkeIrf9jOnPz
5OmP2UbyMU+/z6NCOkGOEYuc72awSNEz6JDVrxgjpXl/2s4xsKArAisx2nFNVC1F708wwKZ6ylbw
d8M0lHrIa523E25qx+M/C2+1ATimVgCGI0jBD+fNUAtQB3hVKnwEmaegg+TBtCNrt8OsPRIZzvWy
MuN6Tn9kiz7vjHhJoH3htBAwnR+29su04NEegLqAV7ccaa2uxLtW/qY0bvljwCTRyYYWTBeGD/CO
6eEfM9xbzU4pUeAtdWXWRUj36gCQfR4w+tYBiXra4887jAvXAuoEa72HNNo58dXh5N7iZ3j3xIes
umKLN5jx/9CDOpunCbXVI07u/r5whbPqjBE4mrW4f78NgFJ5YNImEMnqTWgy11WZuZ+SdQNhuHSE
f2hnU2L++d1RNLkGmJLGT0EPAHpz4j4G3Y680jkbMfTmbSSp9sIEvPSvwkFwNwD7/nsiwubbZaq1
Licj5DFWnYrqzGhTruiKU+jRnPH0eBlLwBwPeV//g5fjpw9gQW2EYBYxzR6GGFl+uw3zQeeBnbN0
p4EoBUPsqcmYlCRxn/pWKqfIGH+NB6dFqeFjvDHLxIdGhwtwddXsuZV7O0kxG7Z9a43LxKWMFccX
uE8lSw1rcB4M5xCdKga0lumiGkZqr8SWgwYUC7FOk6uTsJdR7XpBl5aHOoGRiHRTOOMCnw/dP1kQ
Byz1aubJZ2NJQXsivff8CjxYdNYqprWQbIFU6njU264kotig0wVc7kiz2R/OlzHfnSAr+r25yPsT
PxoeBcksle1vTUuQ33qv4MAOUNcj/KfAn53jDLrYGJSBLrdMT3SV9UiGYBocDIOBEsxHqUtNwwZe
nDw0xRon1PZEvacQnzLH0PBK36OxIbO039GmTN0FuigqGpB3C6IlhC1IF3TQDYJgksj9cAB7oyU7
hrZ3NfgO0Mjy7jNq3/dud+6K4MCuoyIFIapPHEqrzaxyw+fnbdOUlzumIBDHEsrsLBbZr8uNIIdV
/da24hdjjfxVqVqiOrPfMyclAvba8/N9WMlDJTuUy77LxapWCC/N/UZIEJLEylZTWkX2d6eEkeOq
AFUvKOlPCY/zLBNmcqEhnSy7ArurpLPgGSAnlScNRdl2a0jifl3VGGNHOYNm3DmQGCb13OibLmIw
AQCsWltyT9x8wumK8hsceWWfVr3EfhIPPuKPSx871JiXSKP3WCLmZ2Pyo+erdK8tq+tKucjuaxHV
mRitLxu2hoVAw3MaKFY3mFmhcwCZptikA12pIFCIiJUt3N5XWgrPTXcirz0EsA8BMUv5yHLR6Qhe
QhKOP2Yp9GrnZnZ0O3JOtXaFv51dSaYiITg3ve+bfVxEcRYFQQO6OvrqK4GKYLojDkCaS/h6ESwJ
aK/dlyPsfUTAygm8sqbBSpORXEZOoqWalX4AgHg8k8/hmGiFru71oJMoCI44pR7FmYo0a4Ms6Bsi
C9sK+LhJpRtmH5rNPLnF8kRm1KPoG0c+kcXAiNS0vIhQvLtc1f0ngErHWvPtfTmZu3q1aestDCHt
2V7srI6Xay9b7YYOGbTjpM8gtxRITAzq7GYr7OpBZSpZBKi0Vnnj1K+gFPRJoaUyk5f0p07JCC08
mXCLas/LuPea1hNQA8d/0r3O7b/ZmpRtxKovOPy5OD21GSCfngLDl3vSm43zfDaw+wlidSxRgaxo
KpWn87idCTekf14918s14Dp3+OGo+COl/HQWetMsF/TszO7iQ6c67CrL573la760Vx4K37u9XS1I
1CZ6z7TgKuMlFrXp01Mdnl0aQhQZd2EU14Q6tY7Zcn2rIGOkNFL99d+08B1TrTsIuyuADX+qKzWp
Q1cVN5YtmMQQ3W9iWgud0FIcr5FYz57sOZN2v8n6B2HmLPBOhhgHrYm4bB5eP6TWfLt3VJsLs10g
hc7J4HVgPltwtzR1JxrdfYLJxlz/H0utQQg/tC1208pToK0rbZ8mtS0/W+N/iVJF8e0fY0KJG3vP
JK/QiMJU7ED0bvEThi1AqGwmp+EcsvosNRjQqLK6i68Czwb4hQYivA/e8Oz6pgG3qxrfJvaNsmjZ
Rjt2Oia8O6Ji4cMs5MUp6YGdbG0jzDtpV4OiOk+yxP4KQETI2qro+L7MlU19obk9ANNVt5WQCap3
3sYQu2pNE6ZAKE4LJtljnQ0d/hyMvKkm6wJFAivKp9CzKaz0JeeW5OThCA3TeSk1R/EThw5JCwF8
zJruIyUgQBWqfQmP7kP8+/EkUgJxpJMGs6a1vzRaH5F83bAumxOtgljsgZVA+KVyA3CCPDowac1M
DLJs943suD2hgn6GTwQ3MBUskStUiFCx9X/fL+NaRvtNjoj3GTHwM3x5YVA3BuNPSWC19wz+Wyec
1GnJt97JlgLeq63ShHlpitSix594Gp076Y6SXm0Hr/RY408BaJjg+SMmBveOKYlhrAnHqnD53Lkb
y1pW5vpo/JsWozoNGIszxhFPnPM++rug5npIGmKHVwldRdKVGji/XvsDQqfA9TLyJsahrY2aeE0X
Y7bFUKbZRztK+IyNGWolkE2EiqsKQlKKUUl0CgM+I4ki7ertbTjd4HNs352dVEny7kAMjKMbP6Fm
y7QrxebYd7nlRqCeAS6jysm0NWi6HocImb4msTEo5xKetefyB0yAqlmkNneONi3ZPc2wBMefRsKN
5xGKQ7gPn8MJ8Irm13wWl/QGchlSjRkG1YJTT0TOKKHxWFW2oRzPpmFa2y99TvPrCSZHFsBOyVkr
aodHd2VkJxdm7aXQh5NpWbIJnG6G3ZotNgFSv7v4Des/Oma5S5wFxwnWBeiqJi+43Zzt/d74MErO
r4ZREhKQ3onT/45KdsellRL7uDMw+8JIACwYL/hoQU68gUmYhyqRDWtwStUI4s6UrwKUxk37T6An
otzP/Nv6OIAUiKCM968Cu7ZeBGDEN/qwzkg/N6oW0axFGZcBlGGDXL6CxY4hZtQqpjXMa+tSSti8
VOa/IGYBDhakKcsUyIlB0L9ydgnn2IrV0+qDh9bruxS2pJ817BQFv67/Klm969YyrnMkuUHcC/i+
llNDQ9ReUk/Xp3qMDW0+HNWYwUPK2vnUr4O76Av962Pwe9cgsXQQj516788eYj5X4r4tqOlq6Ygx
R+Uw7vj6ReqXzuZJCx7p6fDHfEVPIZkOuJzqdfojDC5S0eSNyYH5rMs/cB2ninPq1opuMxU3YeJL
lODRgrIyiuzaR6Re7XUOOwO1N9IxnrLfVribEWH9teEnhCEsfNEFERmtbl0yGJ+5myEEST0vdhnM
2yXosJmw/QD5w6aAq/El1Nft6np0wiiZu0mhzuLVnJq11+CTwK8FfxDwLPCZfNY5Te47BnDmy65O
MB5YfX3w/N4sb0UVJxusOK5z3+KXpyh/0gMY65sJD98dxOFM9ENmg5/URqTyvhVWNZhELEPJQHkp
XPJ3Z4NRF8d+zWU7K50o6SUZBw6uVu5Gt/XfGGOx9eBISDIRn5fBlo4ouhfRbeG0jgS2NJhZ14g5
yANLbz5ZC5UZOtCeF5Wb5dcIl2gejGpngJhOSSZTcjl7h1ro3IE42jC4diimT3AIGO02r7/KfPYT
yV8bqSx0OpK1rhf4voJFLHDpId7wVdPAk4l1QCkIqF7YhzDEZIGYBuh/cOmvWpYWssp9Qdfmq8W8
w1fyYyBO/WeWjZDWdPU6KzDf6qM1vOITEq6BRoqsF6Fiy50ysMkXYZZBDNbF4HPWBD6jeCKiqPBm
UACMJOTbamRCCS0/3td34cyckMy6+/BN+OmA9oIEGwfa6cGKoPD7fc3E2C/YOWF/pOGs1YnN8G6j
QSHp4OXx0FkI/EkFAniJdbpyL1gJeFGYLXpv9lTSvsiP8pIXODc8XubwdGoDQlRlZpj9YTaydgcX
j9T9iNYqNqJ2ua0u/gUNM09wV++ji2K89JPM+X94IklyOTOUjhQ293wzZqCxbXM5qvdm9yJHeRiN
PGt91C01utU4SOscah7lJBOhQKAI6CjFDQrTE2NPUq/pFKd7RjHuKIA5x93A8e4EvYabNX1Xtd2d
5CGuPDqgiWbzB0YJbFZonR2oGqlHUB35loYgZ0cBA3BIC/9PmpTJ4qGebRwEn4RQT0qNU06jaW2B
96f4PyugWomH20aVsNLUFwjrFui01GACBEWudcr+Hlc6Jza+3c6/xmyeLopi3p4x6CuPlJIdVpop
D6y2Q4RmzOWjMqjrtDB535BKcP2VRSgHRy+t1PK5QJS/XRo+RD4UR+/ivQRuuhI08uMfZv188ilw
w6Thzv1DXz+RVD12fYFDQiT39qbinGb0jsh/hHHPGktjoozpnaja/vtqq+EijFp6+mi5pKWbcBZS
D6tirK+OogLPztdHIEZh15cUS/0sPJTru2XPlyCfvrj7hxf5YfmMHKUV6OlKTPsNK4EUGmMQfIJV
YljcLXdwlWhcBr4SaNA+dBMJJ/4xmHfuA08kDY/yo3mDhiFRRZgqJIjSme8s485nhJgwduWQ/e1z
RXdAhak1zPmj9IyfriY6LRVm+gfJphKf1ArLr189cG66J7dWsdiRi/vkSl5ikw14t39/oHrLqMvG
62JYKGcQoWbQOIvw3DA6ZbxrzWg/LBccJtGL4U+WLnqwQgHxlEaeUF1sAKbN+H5JIl7YSEoB/y6p
xeXSn18DQOa8dQdxL41vFRDYSHcZdTFAZ9LAYb1fBL53JM9PdHld9N+Ipz9gCtxnDdhqr0t572ez
esKfUNDenADP3UvK9pi11LUdWipY2+/5/zKw2OTApCTWz6b6YhQ4nZJTUGYK8KWyJeI3Hl7MPXF7
3qOwrQb3T9bdNWUkfPOHjqVPYR1y9DcTJE8gmXGyIoRpAIWG+MkofWM96IjQJTPkymT1P76ZQ0j4
u5H5faEb9mGcRa1pPiVKNH4h/ezz6X0dxTZWzgSgikQZDocoQUH70ztL+1EeMB3m/5ILDvT+oBaG
PflONJuNGIdDks6sUe+GKgveWh7u58achumZXjyirwxQSweqSC4MPcNRdnEu2fa5Y9n9CTlmODbq
Ut/iwkkkmw7qnzYfch3jrqa7Sjr9CmkXySJnSlMeQO71a+cH0WTlIzUMZBI3tfN5jtgmL1LiOkRZ
+tUoAfNdgc5/KA2Mi5UFMCK/LZ6cGB28RSXe7SpObnJJpY+pXb4P9WI/dyX6RM8s6BIZbbS5sr6K
njJP1IAFzBm7r2taZcVuCAW0A+tW0Szpg6txjskVBb1BdHoZ23RP4cKY4uqqWWEJQ5QhJUo86aKL
YHDlVyG3x4SOKSdvhN4/FjbW/rHZT08UnBb/ZefM+wawRowdGmOLStGDZMvODc/I9R8XcodgTKpC
QWwAR2Zu46FgVCU5f1aRLLspTnecmxIsfBq9gf/l8qgHEuCHOv+7xOusVvykVsEGw6nRpAfbkUhN
qSjmwxCb4ApHbes1EwJrU9sE4yc+SQCIBDBP9Wom5zxoWTINqJ3k3T7GxYvmHXgJIjoq3Z5rectx
Sc0BLFZ9UhcMEODTz+dyVPCjXznN7AQcEQmSmlNX7De4j68XELXOxqlmtuHLVEgQhZIfpv6esUBV
1P04cm0Ub0OSu0DkXpcVwghxI6ZN0Kgqxpb4ckanLPjKqY+2G+OkMB0rrNkaHqQlVah50ylSnUQL
uebkVIZwR2P4SNWmfSJ1QDRU8zk+ucjTyQ+HRIK9CTUZygnkgpznybRXNb4u+yLzGjD+jcL0MvXY
4I1Fla7dmCH+hERRv21aNuYQBfqukeCCP+gsU2Ci8FCkyUx9TL43qDjY6Z3RgXnMtD++1/DsTy0Z
7kZMFZeEuWMC3NddbR/ED3O20G3bR4BDV3kFbbcR1z4mGnZ9fv5Gjo0kSx6HVZYiUG+KDHpGNJpi
qz79D62I7yodUp1Ax7AErMZyE1kf8Wx6Za7lHE50/d8n85bUaOeqX1P6rXHA0xNB6EvvaDakUF0x
Ym1c2f26rj+SDxGz9dq3faWiodc0FK9nz+BHnbzfMEN6XDt4yjKiUxS9DlvnS6OHa5CThulJeFB1
+okdIXYCq6OKqidYi8e6frlvwkGNK4TXtTT5x7IEJFgiRLvA2LJoZkTByN9UCbWxJp5ziYC3/vyU
Iblo+ghy58PZmcN5Hj85pcIjGZUFMZlFPDnePhCDFso3IrRYl6+msJc8AkFEXYIqRnvUzl1ANV+U
dL4V+musUi+aWIxr4c19mihLtD58flzw77rvSJZu0kq6bA45nj/Xc+H+s2T4kgDdwtqe5zm1B+i5
ZZgLkiEp0vghIrRxL4A2CqtfaP76OuShQ82OoByxCi3ZLYwB1BRberVkcAqGsoEl8D4kwjCAaKnf
AMb0G9UcL019S7aVsRf9/HbBjpPBanpUZnyTBL+dshpMmeVT5IE4T4PC323i4tPF6h815boGUfFF
wJNp/9/rICX1rqceBXkRp+w0hf9xcJtYLrlVJoa1FLXhsZLDdACSjCqK9dxWmgZ8TjvYZ99pmn83
wdbPbXOyd1xOOo7bTEOAeFz/dScRjBhneoTPb+yRAfMN1uUpMeKaE1Y9GTrND3thOlhj4NN/jMJa
7FEOwSpbF+WVPDi3rGqRTsjCltAt44GToiTcs579jan8/6Lrotzz2mW1c/uIV20xMckj/83YAT1G
5rouD9ZKIPnDnIWTDQkKFXB8ulzS56akDgRn74eFv5YMnKQl+0ZFefUvSdMwd5OTVVxHfqiAgpEe
1mXZGvcLHvyuUhd7YZ4EgQXic+7d1AZzFxkMsGNjtw+gS1Mt7z8sMuOHxBjgtyOrOk8OLcMnf+Rw
DiTXhsuMcCvdv3P8w5hmzabkgk/g4/9PnQjOQmziJFRQgKFTsxH0UKn3tuZX6AYY1OvCYUOUhz5o
8M1Ky94qqlJMxRxkjLnUfBVIKSl6IT61ReizAcKGX0P0vmgdDqG1FmLPsFswapl+f5QY7Mowcj76
IWAj0aOGSHuPchTjkIifvHlFAt0WGQFzwmd2uQwQz5TZtsLJ8zwPw0BRFa4iB18K7LHgst+Cnpnt
Ck7fFs8JVpCvfsM1Upz49zuyLHIfs/Nmli9KfbsQoJWxqFu3CAXPtQqMODFe6wcYYEN7qIXbTUSe
H09KqK1D/zpkn+SrRwyGXynfATN25+AXNac65kgb9qZPN8BNb+RYJfHIsVb/CDhIVGI31ZNT8HQb
2/InS+te6pdNeSdR+jMtUrVJm6bdf/tbzy4RfLpc/BNhlRy7/zZ+ksaLKd59Kt8tJlnf/Ca6pToo
r5uyLfV98Sa7UvJN6pVW57a+fRUe5N7I5uAlH/29mCdWeKG1zgWIrgP689e2JjZYGALjbmJHeJgP
XcFJrxIVZgxDLEhHGeBIv7K6Amkwly3IcdZHJKX4mEbTiR9CijQpZ4jrrk2yxZIsbKVFndljtuJO
NO8cTlSsgNckGCJf1YL+MzhG8HlIJSSlkjwM8XGEuitKSdDjZHiy63eNVDMontqJX6iuIUCcpAfe
fcPQib5MTZP/7q3mWySU+Q1Vg+jmHnH4ZS3Dlv3BFmwiAZOL5jEkBmMVbif9WhEiNeJuX6iNYHJO
q+g/W0wsn440pxSz8YHdmaMqBnF82toYfG6hZrk871TltvcPWH1z+8temA4e+SKiUCtL+sptCjMW
Hp62APSnuKxxafQ3OUwAdmc1javeUQBqRYvkS82SPK7EoSlRgr0fiJ8PV1YKZFQcZlLVhPo1m0Oh
mUmo5kfCtDG8L6CM15huv3J42fLsINhVRC/lwnLbvFZHWLluUDW27/+4VjvJ2te5fa75PoAKxPVz
GK0/XlKOgMgRVfkLo8dlEKQh9LtZN3KPGUaer+YZP4Jj8JVrb2+gLEA2EvXEMJnOZ4mvSKMoSWxj
9jiKpdge6hS0yKGw87uhtV6JliwbYDvmn6erJiDP5PvBGdVeIAPM8rQP5pFs3uXCE66SuKu76Mp3
rxL6bg6b92eq2X0x4Zo24urVK/fRrEOuEZRbrbZz6FpDmoTvlEopsl5Ow3r6fF2VcQfPjM/l3EdC
ZlJhDCrWizv3BGUzx3oYnFD20UQ9AGp9JB+t2OJLaTtNjqJ8kDYdGj/GbUlJty7/Ctz5wKH6Y36l
evVus/O6/xjwTvg5P6mGqW+sbdpXBHUxafomRfM1t3ggedfZiInMdS/QO1j7+WDjtTpy9RSGxbl1
ziJyRNVOHc1lHN1/RLaxhl7822BgzS99dbVAbVf6AbvQtcbaMH/+GZUnzpDv4MA906nnJE/EBufu
PTqOWmbVRB6tOd19dZepAVjL1dq3AVYQhDF45Co+Q5U6Y/pkAi/ugIU7WQ+FLmOHLbWYhaKUrhS2
iQTKAwBCixjNOg8lMbuaAEyV3Oqo+XASi/OcD9RfFZal/6Umc2/vSISd2gkhrrx5sYckoCXVgU7m
tOq1F1Um9QpakWvxwHHmUYzfCBIxzMjY3pDiZpUBN+N40xj/XE0WjZEbMj0XLb2wYUPZlIyXZzxm
mXu7QPSkTWWPNesTklz69tKnZIKvuyIjj6xsCCWXNK4FZ5Gerjei8u17e7VdHwC+JET130jF3jHz
0cWmz9aM6OADuQRAw00DJn17ynm+dK3y6/NWOoon1FYUUY92/msfDlZBEKKOx47UkZ9KZ4DwwPw7
MJCGJsfGF0jwRVKTM5x18YjtnXcwVB26YRWx6pRg/XGbOtcp0Sn5rIEU1k+/RWoK2gqNcMVuBZDR
D3iHCXN3fo6FkbrDIy2GzVkcGdmXt3LlqvLCmq2Hx2SCMWQHrcKLG46eDIAAo9/RIj23cpB8IB4I
gnSjvDDzUicTHtkZVONXbCslAplGRFr2w4gYq26kZIcDXooGcAtRo/UYXQSvX2ULemqN/CbX3pG+
W+C9lJ2wbKXOL2JEVrHICTsKxha+R9ju9BTCqfenQcfpRunueSywVzQQQRjaR2gpMZeDp1fJY69+
W0HdHZceh1khs1E1vt2NsdGFPg6Q021REfrrPbBItJMn3FR+ZGHSoXzKSB+607IbT+uy3K1Iiq2w
tIIPR5pSufmZJbYf0kX8NZgC6tGGKhxm/VlRlh+jfRueOVR5R6i3DFMOX3MbsRj1MDO5MDTPkH17
5OGFQq9KE+3tpDYs7efMTWJSs/4B8Fch+0btVZTe1thAhPgTWN3Olk1u6XIP5RCFHkc7OrFf07QY
3RngvRJ2BzeA2KLfVjE3R+CeWqB5CB3RxraH90QXfOVRl2OC80KyRR3ZLtQcjKD244T/zrXKRFCk
xkxF1ujpk23VrZdieb1JpT9sNdNGpAmhDdKvXFZajJfQ+rDAfzB81f4tXZhMnXE/XRWT1Y4LLHkL
9a7QOom+QfYHOj+fnw2kwwgKerb5a29CFGm6kc+TI4TM/fF0Jr+33pJ2vC7DUNaGNvnJscYsb5Wn
BLiYx9o+cg7Hv/iaErtsu4lCREZd6LtSlA9db9qBBmEp8h5ucFvKcavPVwX8znmVp+QQzJS9Dmp+
oLbu1fFKRY/zqJvc62dlwyLXK7n3YSMHUmCgi1YlLMIuDV0fnlD8M7GaTuP27bwDkHYPFvVDq4/G
7iJ1M7+4XINMjWYBNjFsK/QoHulMgFL3bHy7FQykLNAA0n1foW8yvsbYIbz09JK9vPo84gfQqot/
mp01G76Nqy8RKum2JIEdJDf26pzbOMr26t3R7YBjrl/nslQ9DKoYHXMBsRdxFSXJdlIO6iz8iltG
VnbdzHOP2eJGmWPhE/XcugSJzJ4R14OxtUOOVrqeXbeqg2BqmVKDAbSodHXW0nZ0pa41P/yNAnkH
ldXsGdftViT9CmFxbDmuySeiVWjfOYjqIzmWcxAwRNyGV8Tb/Wn2gO4o3MT9QTZD6rHpp6gf3jts
NVT+qzm26XbtfVQ6LHuhiR3xcbkwplX07O8wKGpes8eMPLLAyafSpkdc/1NV6hh6lzKUy+WGEGSL
7ihU23tkv+G7/2AsHrIrznRaHrdmnMtt8NicXw4hTgdekcR2osh1O+eyChK+FfIqOQ6W6/B4x2ok
u/P3TyYapxLRz+aj7Xwm0ALH2ENMcGd4RpldH1pdMXLY/wL8qrUaMTiwbpISPym+W0EIkWSR9Ltg
+b5+ezhm7qq+lSvDnW5IpAcP6UHdugAlSHAhULm+E71jTKVQ9NAp4435exhUkZDGxu2N/uSdz5RP
mEa7g2+gdCZ5wN3zkoykKdrYVxtk6Sx1pJo1UayPGbqFcIIO3KdTyWTx/rckLT7MgxkUClH1p81h
0wrMNzg3jma+UYMgaOpUrQUY/+8XFpqNb99UU25iw/f1IbVCmppzaHxymqxsT6nGRT44i+ZfFthm
fEwmRvsPuxO0kzlo7v2hSQgLVE8TBqclS+sx8boFVhw2WMUyXzp2XvMklS9zMJGZ8J0Td0VaiWNM
EwdczFQMWeDNProNq0bT/XYLburj4dg/fN1sZakuxwvmhrRGinf7ZxTfrxYGVlPbBRuNrRQ3MlZO
eUcRbVj3FrIexSjbpV+nTgCrczD37+UGEzqiFO9o8Pu46z0ANszYUnaf5ZhRdhX0rrAmYR9dfMAh
wJZnkEwP4Wz3MyPK5J3O5Qyalh6tMdE159pPKNRsxQEavCCThRLC01LeRxyWT4rTJedm2IfvWrPB
etJElqb2SuxcV7elCMk1Wf/mKe9yNwgaXFFH/nCJn4fLF3mP8F2CVFvnXRcdMeYE34dNsLQEifM0
3+iFanU1cqOr2ugiFf8zJ870C+N6/qBQVKvQPZHghNndnZD1z3oves5rNRE+06NoKwRRIvsWxMP4
V4rBrLE4TG0Dzje8xKGZECoMbizdC/vSDTfBF7G7DCDf5PxA1e9Ma/84i41Wn0ITwWHNDG1qUBkT
Hokj3HC9CZurtkPmMWtJH4G1dtK3dVBwyTA/CyYokoqgLqy21AFzxwM5s+byhCVzQ7shViqiW10V
XLSHZ/nW2pyc8+HFjFlVTY5EcFcTPJDD2UeBugNPgoJoNbDsD5vEKf2/b6vdxEnElaPO8ObHTl7D
YVLKwjh2yb04prKSPfW5hW8CjpdNHbwv3l5OUXopH0WZghHBHUUjujA3kvEpUunjLmbGLjoKns8Z
ZnbxLwGgWcYgw+OkWmlJsDp9UWrWqe96gsqt/Di2qamYhwNQmY2fh/bRgIskqevNn3KCQZi8biLO
pzkiiKqTtIVxBygBbEkigNxZ/Om1nSzGNhMbfD3HqU/j0IJhw1IIm5Lad99EKg8P0JvJnsEfqRwn
mPO5qvFAnu50DadctB2GupGven2GF+eNF6y2y2LTxFTCmIZnlZ+CbQG5SFKETA+Tv4PCcYqLmYeQ
rsW+j2L133BSc9dGyLiqreh+IxAHL2jqvF25p7kS7/ulLqr/iyGUyJmbs9RuT8HW3sJBs+MBjUYM
kboQ7wRqwwoZ/QBdNPawcbTdvGyvSTg6IIqrhkISJOZpN19jbdLJ+r5eJkmxrjOhc8mVYXtEVHvz
ONaCWQZMehZmhTfy+tg4EaONIhJnscmEv1YbgUs+TXKYXbMipw1I528ZXvjqZ09c8Rb0uUeNmyvh
LqgYsu0sMCzvUWi4Cd4qFlmKLpPwb/Rri4Fx7JtEJ6fILiHEeBFwncupGXLwJDCgAR2KOnF4mkAt
FV3rNg0SVmRrJgW4W0vKKgrlcD9Bd6y72+0jfwBAfiiow1fVFQ+byKIjUUWoghz0kX1PNzWrdyTm
EdeTR18s1sxYS/y10dBXR3nsPcsrq7wGiT/mYFilv7hlNv94hn/OZBJBIKTDLAZTfFuybkHxIjuz
dlmGZGKKE6OFoeu8RsOX5uT405GIwdppSyY7JnwbGZIx4Zh+ODlW0caNI4a1G/tnMFZEcPnsWnOr
Kyrk3tyq9leUCLorDi/LbckOQYqVEZK3uHuO3Nbf9mheM3V+dgw8voiFzoKCUe3SErz494SosPA2
OP6ZXU63Y4LCUhbxnrHamCBeuKMh0AxZad2GoAZHW3eALTwcJw99GZF2ajctANKEj5rxcWzGrvpN
G4KQOUQ7VAECTCCNZduBHOC8zaB7jc+5eovgbRSP34CEhoO2w0gsevV0xHgxlVji0d57MridpCVf
F4S7j1mbft5BTX6dQmadb225lCtE8IFYfryr/bPZeD4VkaE/pWLS48u38HivXJYmMc+qlRcQrsug
IfYiwWcx1bGtf/9Sdaxw/zk7fD8Mph0YwzQC54fm6QMzyzIGPfUo78WSEII4kbFowzl7WwymuBOC
owekXsWrlJ86GQkP96BDHcnzYa86850RtHkH38bQ+EZkj3aBKyJGZQsJZeUEtP5n+XmKZMko7Gui
4nG3+WZK8EM4wjV44iCK6wfvcTmnG88LxP1+1Gtqune5qYnbhdT4XVBe+upyW1C/KtiSiIp5/6tF
n2ERqMIC+ww/tL+taeWTdYWNsKJS1zigF9HSfyOEzIUmXJMckkXRYbsNBV727CtEJGnggJa+YSrQ
wTJfrd+xFaVgP5RFufm+fJD99/Lx4GytEQge+s9uWye6XszMaU4CIdbgKozT34bbOLCsMVaUq1xH
na9pYD+zh/i0LpNcYlOF0Lcfquk8oexCgCxn2pE19i4OqCOuf8ClasKxYaTF5Q0VCZVGSOsj2fcl
gS3rQTVJPVpzuK3IK6kAoosTsdg2yAxTgwnLmJwpvZE+nMbeIo29q49mLB5/JGFmP00hFAzzeXMR
1bqbbaN3CQ60J/mNokBsfwagHgkNGr1wkAkH+tKiamtZ1sBwhMAPM0wvqlRdJeYMTEmMrXjhcUV/
8cWcBVAxNwVXtwXySdV3ecMxnCr3sbWnn4cE6d3q9j4v4qEXZ/45+Ic2v4s8Wh03/0J26+haJU7k
G4n/14nENQrh2rMEoCmUcQQJDPMaUWk5wEA3eeH7g2cYogViO7fbP+jj9z2D6TnF1hEJ6DBvlJ3D
uo4Sh1RRuCpnS8SeZif+dM4Mh0tiwR2Eubn1eHMdlxgpuU4kR/87lwcuQsBW5c6E15rdQuB4m9/L
3BsVKcON771/CGi/FHi5A4NJZTskJnEvSLcsyD28LKDg/OGnUEVBZT+YjujtgPhEyHZbRsi70O3y
oUb7WvROGw+6J4h7+6Klk3JT2PQRiYiWlhPMnaYaP0IUxlbAC1HEhZCvTysrz1Shp0z5rExJgg+d
nqRoDSYRON0J8QlE0nLOc7WE8FC/P8Q1uFGnepCnlpCya5gfy7Y4XZemwD+tNdkbFq1ShgID3prc
ajmVJRLw6gPknOatNjMrNPU25aM3uRSTlfwdsvMwaGyltqeQmtGWMhaqmnndZQVQkwNygQ0Fv9Cv
4FFvSvbtdrGI14dk9hpuQpk5+XI1YBLz98ulF2roahWhAKIMHS1+JF3SL4o8tIovOW29KVRM9E29
/w310klO22jqWgutBpaq6XOzUxj3ZloAFPYftnzKzr4VMcYyXmWujnXwX51ecxE8IRPkBp0BRQoY
1ma2rtMYV+8R81WALD/6sx9DApzPbN9/L8LSTucBArlNlWtD+fAxDsYi1adKWzUMVwFO91J3M+13
xS6vGhvIo5A9hFEDhCXA7E5spBc+/zDJGOCFJUzD/ooBbRR6Ppk8UUjkzErh3PTAa4xwuYFAvqBv
CZT3Z/3tew1EAuQ1fxobv6te56++VqUGQtBiHFYcYrPfHkDt9yInZ42zR4eGYpYqeE9yeD/PudOH
1dQErJszAcJHCx3Bq1118m4HfdKRjwE/Omo47LW44feZraR8sGwKgH8XV7IJ2hVk2WiddBejpovc
6B5DKmKls19m+5JLvSUuD4UPsU0wCT5r4u1Dl4pM93uX/OFHgNRBX0m+XoxEnPRCytHQEP6SaCHZ
8igUHoRl/M0bOKAozaGcx/hA2UKFB6QZ/7Tmidm1vHaOPagsCNesHSn6jjR7IaOwqmlghEfO+c6X
waUNG80cjCuHMijFBPd/Mhoz+Quaz2FPGECDWO5JHOU9Hp6zpjjI0d5a3S/OQazUNfJ8UTxdAMIz
ZpEmj5iRn+Qn+cVCrDFik/70zYmVtm1JcVdgawo2vF4HEcdHs1fTyzQ3Wi1d/bOfJ23B2cXCt3kR
iNB/gx4Cp45XYx70YfwTcZzeNTXnBh9mBOXUdY2Ne/3Ufsw8GxJ43ohE6OvNdVZOUi7NpYha0IML
FqNGsv05qI0CQ53oqK3JhrYUzxzxVeNszBGV/dK42jZDib8JKTIM1dXNAeuNxi+vxE3oUBZfiUjB
LyasoasPpnOL+M1fvWEyfBUMf77jR4psqvq/Wh3pzXn+i6xpPv1Xf5Che1xIZmvv9lHwMhBjZnAc
QuV6VQAx2dBW4uCWITPZ0G3FTMHZQF6zse5ZOVNhKXcSfXCFHbFZ6ayPIG7mQ5CepFCeFHwxHPgu
R5r+JvKIXanm3O4QD1SA8HVGK+ekyXQUdypAZJIDNCH/LMw3YYbgfF7yL8JGKy+BHJBilgqsfq4n
K7MPPEjc9J1uMqAc6Z45tM25RffAEIgL3GfoahBg3loxL2DueENoU8ELD7w+YcUY3bgUhs9oRldH
FgFTK8S5DNODHeQm1sYFC6UMijtRrfqv75luhA98MIboSzoFdMEemL62JlmVWqYpzrzi1A9M2Ua1
EWlJbwEn9eEp4y6JpBA0lGlslQUXNPUZgRjfPH+MYzEKfwPHA9xIrQbpzYD5/tHshUF/rvv3giqe
yP7FpXH3KX+sbykKdBAa+k36CdAcaKSXLNYJYrZ89kSPNWNc3K3siDZ1fUdRm9Z3Gx/xUtB7dsGY
QVmcbWSk/Ne9exfrvVhqQhllgTz/wE94skkyr3JNlMweTJeZE+fZpy3FT116+Bzq1UR+GrQuz8a5
RKuqHZ3nRvQ5yu/x73wj/5qvhy1aWityOkulrQmX25z1/zCf2h7PIHeGS4owWtwn+nDMJkdge45j
OAUdiK98hjov0o66CHanm27tVXkfriiBEkDON9vBu6MZHTPzHWMkGRkzif0p9RzjFCAgdTOj+umJ
D9LPojoW0m5Uo8G8A1H/XQK82fCkdVaFxqb2/FvKOO4rJ2jollfGexmGeISi9TRSSYvDw0eS1mPt
MQrCD2pX26b6peLibdVsydNJV1Hrl7Qefcs1Yj9Ie5Z3+FVyqfN1BiTbSWvCC9xXHf+jrd/mHSR1
8E9/EcjY1e69CXLtaE+uizsH+a7GEOdJGrcSUfoMR1bIxGIrONuVG/OHecVQfyds2Axh52QFVjB6
WOEfY5NGyOrOffLipm53cXwNXSO7MUarpgXylrsWptxDiIiVwCKJB+OxKxQA6PPdQaNVtMhkmH8h
QwlfZv7d5wSHM6qgFX8pBhmEPQN3bGSJOrylZScEQkAxVtXsqb+d2XajLtlHsMlFBpo8LSzQwMac
Z+I9Xg2gPbiWk7DUmwV95YRshO1Y/A2e6AsVXgRTRxrfFOdf8Q3aFowNveAdw4BmePhKIH+XdzPW
iOsGn3400SObgUZq9KRfnDoaLk3iIkCLclOYvaSxKRc8k/9KxG5zvaMXrV0P7cCSmK3XqJooT80F
PgQPE3EJkwRCp0kay1WOujmcI2bVmWnbJNAO9JNtUpH5tM9IUUXggaCtvyCt1+lF/odvVixw92uy
xIfAK/26bLV16knUnsa0OrYB4GEY0KICjS64vKDZ0zaSdj96o3xF90E6wizNm8bnFhYm4qHAzJky
Vtx7SHtbzli5WLH2sb7Ggs8drudUQ1Qvypp9WHGFmVjesjQQS6balhHEurnY3OOaX2uYWvrkbqY8
XHxrQ9RzeLrOvC0h80MzRY/xQ9eyVQkgmhqrEGS02ZCrH001iguvkZH4tBrJp+80NjhRNx0eo69T
BnZv9opPPGC5JchPUlS3hStsA+Ud484UcSn+QsfKiXapYNjJcgCzoqptNdcQX3rmD83LsmqXQc7X
MGOPsieNZS++wHy0gJ9hsQIBpKZURn1yMf6ktTFRo723r/qSTZNwH5ai1i6yjIB6a8qOnc9fESx2
go374mxIbU3nL8etjR5c5ct2SswWfP3QvmNI//KiZBKrdTEv4ZySHE4rs9TMyg60e4tdI31D/m3j
o0dAD5zP+8Dqqkljw0gne6xxOnnhqD+6BwK40frYTYgyjmeggQPBLhmNnT3c5HD2Er9nemyWDaQ2
JsLnUeTYz/nRvCOvKPNxtvxd1v1GXsnqOFIJ+/M9FF3KRZW6fdjHFtyJ2t+wwfeQRQu7FoJiSCR7
3zFWo+u/+P1/Ani2nc8eEtMhWbsd3T+EbWYdLr1oDyYSbctPx7SpSL+9pIUwOSad4Scdqcl5xoRo
+C9dE8uv5nLikKMEOFFSJC8O27MTu2nrrpizxM7S1YpGjxjdF1YS9xF3gidLVVmp022UHCGnJKQE
FCW+5KOu9N8ipmNehIzubkI6LymSBPCrzoyM6zwdaNi6rIhJMcNwSzNemo7iuSxRhAFd6ALfvV8x
k/lEYqg57CZ0RQ7nSWGaVRbJuhfmYSDq74r8q5ILyP37Vv1PDznlkG+QbrI9N/uGD/pt0s3pEBcv
KtkPYzZX+NfHyVtMrF5edCfd9DHmd7hNRENbQIEFj9iUiI7MRdIewhPe78NRk46lvPV5OjYU62BY
dYuBg2Gk3l6YMDe8vlEtNDEn2MxdU7iow6JDKaRdcQtAcx14rEOx/SHqm3F30Bmazn7oV9HGsZZA
0XbQXnGD3RmRQWYSHarBiCSrzeA+ald7o62MiwQr3Qrr+/N4higaCztyZ/wa1fZEurVqiv/EWPor
towkF8AJ2D2A+mxgsdi3xzgy/ksk1tLe2OjZ+97zzUKXnnL2EM/Xxyu3mtH96+qNWYwOWDdNzfcy
POPsOWhb7RxqPKObVftM87oLXlp40GRtOvWaSdhgj08hBE+bpBoci6QB59wPcOIAynWV41oBQue2
hV33Rd6LFY90jbZvjW8gez80Ky+3IB1eK/EJhtWx0PqDO1TEm/KLtIa8zlaxQf+IztYnsJiGdstN
60aa2m+MVQwRir0TBhwsWqpO9ETP/SMUt4GHqodtMDrhGWWht9/10RI3UxV4A6LerBa4XFKSJWt8
2VhZK/PgABqW3du84d5uqLKVvOemEXrHtx1ly1EoWyt+k3l0z1GrPk70f/ERmm/dFzXaI+uhYlJu
ENwhGQ9ORh85Vs1VXL0QP9u+/s7ueXCHCE4rSZJ6zbrIioMnKSj44rabxCtNbpG34mlEgmFoBmh4
ML5yrjpn6TjJyaImGOSCszwo2IqT+ntlkMbThxWa7xs+9OftlCIizVj1d26Zv4HIMXY7pHZsyiqK
siReAQeh5mFpuz6ldRmFfdf+bpWRT1YfJqO3T3MlEdsKv5EeUn9LVA5BYPqxDcvCq15LEOPI4CQ+
D6IAfcCjdVaS+wWbnY5aPHBPLx5yZZy4wahnOLgAq9B5Q0NsMyfgBejDWBMYZziZVAZp11XTOi3u
s/d4DirwrMadD417dTQd9bQUJA5OC1R7muSrgbkVTk3Nw8on7qDqdcqSb2XCpNUxCZQ1ir09jsxy
whp3CIBrJFVbCTvSFpn+AOZi6BfLjLs2SfXaWeVN5qOTfIJ6/2F6DyGbFJUL/bUqN8fTlDc1yf+P
Z9nI2xWgtAPU+FdnXp48baU5S0Nj+HldzyAY+vhdJyq/Z8jb1zwCgKOOuqn7hjCloEYgoOINLtS1
fmsM5abrDZLVvwt5V4xlbslA9MB2ASIYMx/znQEIGOkFLnlZtr7ik/uw36NwiXXqdodtCuQYWJBe
D9fdSjwn+Ys6mPaXs5vBrJh+9QpH6iMWemBRIJ6QbbncmIAtCL3XKi09HcEqW/ssaggvONyYQla/
t9SvNSzusH+d6v4i5sG44CnqB9WWiiesiXR3GyhqB679K+EC6x2z895SKQDln2whmg0buH324wG9
HfU7q6U+EMz6O8yOCmEfm1ctLQnz/06wwnUn8vQls1rel818PxaKUnjb8c3qfYZy9/mSNlT1fU+4
Gb/FdjsTlhIUKrNBO8KtXbt5NHRlAPWc7Wkka92EufYLjt1iRCc5fC7CmzUlaIVgoZPhcA6Nf0RC
CxS9TUjJoTKI9apCbEITBj8wLpm2FG7UHk6RERueVmz4ofkanFKud5YPs7I/7yu+NPE7QCZdP7/j
uz3zFhxJw9lL5EP4lG+cqy2lffrRLvWkSfeOTcDEUlrQMbPygMa4jGLHkjGNS2t9S5JKQdyW+ZrY
GL24biW/aWf3EHfl8hEqtItnThOg+HPISRDy2ZT8oNHx3xm+NiJTh6n6UlqaQTt0cJle4F/tYQ9l
V1lqIImVE+PccKKs7jjjm8SzsdbYmPkeg/kPYlXMx1YhHqOaNfz7KBUx33bZDLYXhDKzZhYFzJT1
FKCv6gJfSCrOuNLJa4uTDKhRZGKfPjk+r5KvCGSnV3K4h22ry6DUpKUmnjEPkAvmh9kjtcHBr+A/
tp+LvmW1MfeHF4HaNEYQfCBWNSWmK0oo6xTTvIqSM4K06na6UHN7paLfPmR5By7lAE2mXl5y4MaZ
4VoNKAN1Mf0jRMe3ZYvDCcJiPw2/cpBaZvnU7gbzktK8spcPpYmEuq/zsynKlvDVx+3GP6qT1v0t
5FotDEAoSWTwVmJXC7/D/FostsVmBA1xuc0EocEpk1xlhtvJvOyh7+1hddYQxokA8QRwBjtxg4i/
j1MqX/Q0V+lqw/jo+3rT4b6xJ4KkVbN4MpXuKh00+P1Re8eARMYi9s8eUkrYNSoRTXjIpAyKGjzj
xGvriUKgZr8fy4vQ/i5X6KKylrU+dhzRSDrAzoYO7k7B7p75xetk1X6gaV9L3le8h45HX1gb0Hrt
6U+7chKv4CfdHWhonnxg09pkaUKHnjOA0SFjjQ1Ytv83lJy1LtUHPsjdZTrnaKDUbX5cPIu90Qn+
phT7GW9FPMohdcMwliSi1Ie/KKXAghmRhf/MrySe0kTxrmOnh8fV4QmHeUo6rMHUVeKcHJYeaPHe
/qFLeyMUqCpHutKHxFQxuOv8oXTUA6cAdntDxFX8JaD3peOjTC1D1/63d8d06zpfBd6hcTd7MvWU
hL0VLVBC1zdCtFY8EizysLKuZYLWEGe8etgs9KlZicudvWkdkr+re57F9o4QzjrnH5ttk8PTZKnH
8da3pOZN/A7vjSsPAJ10b0nTUFkX/KB6et/WB6gjek/BoWFYRvkpRXGXW831WiiRe1flGGcq5DD/
gWztbgWLg0DDqu3pAp06TnnVelOakWjogonNB+ZvzhQLFcB4IeuKsA8C4jukgqIDk3GMFv65AjMY
ky+nx+Z+lT3CmX+FMHX9zMsFpgLpp2wDQ1PNJTwlYAPA/hhdgVpoqOaAHNbm34wAUTxwAMWElOgV
mQpk9Q+Vexwgec53CZJMthtX9FkRuwBUeBG2SxoV7uYllz/APNjgbKO/L+5qGpwCSL3DxEIRoUjZ
ZGCTq8+L1JoXAe8QY/2LJ+EIz6MrHIwfDdce7XatlVssoqU+O56buz98ae4b2SQ+NoNUnKoU1kRf
qBIaDytfx5TTsqbWqzsZceylsMOYaMmo4n+h8tzrgPM04ybWYJsB+u4ICFpWWPSuTJkU+tZJEkkq
nEQS+9s5viIDt4q4TNFLKLvbPNkLDBTa2Z19mA7kSsn53atBHlQZ01SXH750d3fyjtZF9yKx3L4v
XSPY2kda3c67nZLk9BPUZ8UBMwAtjE9Nn9+U8vRyrWeAvvsxG7NUMeGHi+VozvUyIRvxUny4c1la
bamggTuf8GNBYc1fv0P8QSCDLmQwrFxZin92kG7eShSQjAAMgCqtSYr7RodRacj496TEE4C2eAzK
gKkXStSIaGTxCOeZzXcE1kCjuzKlHr2H8V0u4UAqfXHlwc04V9fxliSD103LwP6AkUZiZYN845MR
ZlbCKBF6a5/u13r+0VCJMscw7hvwdtreiUcwRKU/hP1QKnkjQuKtRsuCw1YSVwAFxRT6JQNZPapa
D9CNlIpjU2Cy+IN3shIR/WPsxaY8mkAVKiRZcTrwL1EpNhicEbvgl4l0UaP2JfFzRPWTE9yl0LgY
L7z2vIg89DRhVyhDRFHzCHYXuFHigX2ETiL3xcCMV7pk2xgT5/3xwEQrf5XUA8oByXTf85hud+GW
qtO4LxK5B65m/yk2iB/U+LUDmnjFQrHpfNS9L3WhkZbU6qwPfb4eC65kCwlhUioFdIKrjV40Vo1r
4dYi973QhJBEw2rStnj8UdwxqdBOdFxIIGO6gDx2SnFwT/XU832sN3NOlRJTgOpOTdhhGC0N8Ztv
4/VFCtnpQjQ1S0V6F2cI3Gf5io9kRlJXzwxmkLUWyBorbRmD8vN6jRufwxyYiylPQl3wf1Y9yf18
lylnLw927u9Cv/FcHzgHOo04O0mnGpHEGZVqXNq8k5uCAIkyd4iD7r4CGQFzyUm8Q3S1di7rJko8
wKDaZK7TIQjWFixwYBySo6736CYT4dVH0HTwcahu4nhb7izXtefCfWLn5XGSK7wfXs9AINcCMyWW
XTkqPEuPuVtGLn8B5atP+yrb7PDmOaN7ITsDNiUcbK+z5N/b4p6jRno9n+qwVos7hkORmljPGZj2
VbADYlB/aJxxjOSFc7+pcVDimhK7e2UbDXMpwxq+oik7xcLyG2Sav9MPcQ6ji7UXMQJkStkBi9/Q
Blib2i1fGdzG2L4gHfByuZ5MK1+S13VrgR8YrBw6rFUJOxDpwnmFuz/S42XrI0Fp7zchGq1NjOAI
O3/CgJO32UBdNvqUBY1JYaXxkAKSybpNb7L4PJ5buvaUYt77ROfrEvRCc7KEexhAeO/jE1HJ0iJ4
pColnMzw4tll+0BWDir6RFiwex5MFvnZh6/e2Cpp9KpIlVUbW4k0FSamMUEwUpnpXJVTNVD47x/3
3Lau5IfPaUaisLqBI4RWTWOnT8z+lz31GcDXO4HDZVg6kYAHpWX3z+mBtv2yKVprk+NYTYWC9/4F
B1fXY58b3t1h7P+89MKD/y+2U+eY5yu+6+hminSBhM3zNtyDWfnfWSTRxo7faqIkExhInUbuJOdp
ME7c0rxzE+iAFjnOYH40/QJxSucETd3cHvrM4aa7FaEQRPZSsggn7jybasVl6b8BKzT6jl1anHY4
bpsYIX1nwu0Mtk1lt+6D2llpRXDFYFxFiIGctsMvAOi+Wlstd21HNmONZHulrhTvS1a7bLHeQcZs
QzoK3zl4OrSYTD2WHqpNBui5/PzDxYC2ClT097QZWn0ZomC5o3lQFOfQVIXXv7oBF8qJ8Uz5x/2O
JWfwK5eo9+J6IzkMz+PnnTXsUit58MUYIZwcbhk9HUyL9OluhnQ0ykUhpYTXA+VmgqhG2GYqZuLY
JxJG+O1o3SJ8CpxjdkwXOgBmxlcj/Gyzic+j53zZmsfsdW1R4Zvul0eBceL0W2xiAHd0jhpItJCZ
7o80DAGLiWkh4dElyoZ736EOF10drsW5aiSZV6iR57R2TQvWRTQGuIFboOd1liulJ1V3jLYDdcTP
DU38q3Wsdw/y+fqTXqwAsErC1SNytDLg/BUqJ1nqkDaJJ4PjynrDUS2Pm+uw67o0002bkHnI7fsF
Jr0BsN+fx8EWx2HNOWo98KRiuIr2oIM2wVfe+woX3JwDdqexEyjmiwe80MxC3LgrjF9vU+Ybjk47
NY5t80x8bNdRPX7StEozovzqoFL3XHS8AsihjXXwdvm/YJsHCoE1OTexeJvt9hPr621O9YYSPvPr
mFBJcvLUw4UOvDjD0bCfqlYBot8pkMyilZQ3FH/QbxXViHLs1+NtpW1F6F1n9KEUC1q9RkRR9Nq9
BBxrwf5vp93WWFVhX6BwApQyF7xJPrRFBnr7yXnAg9nCDFvTBi96k6uhDhD1GWhIIrA5v7kudxiF
pp+g+XQXCPWTN6cZxO1M9MrjnEELFElHO4w7XbvJvFUaB1JIRR0PdjYfcQI2WEhZyxaumnUuFxBd
so6JaZ+5WHXtXC2+Ub0bW2HTtb1UM64m3ECNLj/eGoXj7Uli4jem7MHJtq02lhTGfzaPwsZQNdOR
Z/7jLaxT2ujoU2BZ7CS6KiMJzcqCNexv5/WwhgE//d+N6Hcx/8d4knFTNPN5lGKk1vvq8bOASsNh
NCHjUrIO6e+h7BL0oa5iCtE6cq4pLgBtFA40GVBr3W0UZkjvUBrOy30QkH8AeZi2j7cf/IXlKr6c
D6PwL8/JnXr11yCYvngcpimd8X9rgPq7C7XB1cZLzzjCRBwWhSyMrN1bSSkR0PxK64PiAn2V9466
4He1AQe67OEwLY2X/tyXjgPP898XE+3vAFKyA8o60xBWG06+KdGFUT695q+ZsfcwsaKXrkV9RZ9v
me6v277Xao5VHsF8MXp0YnrD84M9NL3ceaqw+JEwp0n2G1GkZ9dNrIM/UAzGVUdCOZCu+TZOrIL5
X3oEfKS5VyD3r/0ACV7nL9C+kyQ//GwG8cuFysRxBWqTT/RrgdDRU33+bu0kYkO8OMSYS5Q+mb3h
24E6AXrUGVp8LyJlwiawdyHwmvpYmVp6+HTsZzo8NldCRo8edWXbLTpZy3fL3EuGeZQ1WILvdZlc
HUJHU+oncM1y6pALOD008y1n7/3DQtX0nX3lyq94blPclPW8dr8mLClAPD8EC6z95l8/m/s/EVD6
43hI/9A499buCDtz9TlgVugnh0yCUzjlL3UZd4GIgUSKzEK/fmh/Di9CsFwHc/k/BqSJfEKCFzsZ
j/Rd1Z+A6z9OztZRp+QSk7NKlY7u1eUp3zxpsv6lWd4mMIukwKDhDpvSa93oMrMsJHGD4oHzvpQT
P98Aq5ZzYGXbwRXUuvcU8oFkwAa2d8FUkM3gb7PGabmgtA6Z5eXQOJk+/j83hX451b7IeNWNVERO
zQLqWqL1+Kkak1/BwQxJVtpSmtEjMzoQ1cWYGZ3frAWxQV6iDLpFbE1YjPcpXMp6sB1yPBBsEiWz
aNxLPISi6lvyCyfEjsfLtpWz2qQLfOMaG9FS60RBHTj/SHrOJXdznnf65pnBvEJLhClqKPdGjzgP
iAdTwdvxuiuIPcrgSuh6t6RDNQzP7O0IdZ3zwsMRwaM691Huz7wgd0Pstd1jBz1UwKHggp0NC2NL
R0t4i/NVXR1843WjTZbGp9xSlqZBdPb8FUMmB0cT33Vc2NGCOLgtroiOK/GbViTU+yDQLJJudZZC
yAmqWPZF+WxKM49WwDZ6wzdee4rMMBCYhbzZDKHrkvo7W8jwEP4a/YbaND235kKO7I7EcvCXNHCp
B9dXkl292baXWdu55DFBQ0RJBZaPiGgd6YHb53OFfUO1qNYwpgvVO2GIkSnk8ikYGyAhIZU+2iv5
brjlThzwQGbDIimBm0RMa/xszDNLtywPtiGSpBJr8DBAhzh9vXxX8C1iG6N+o1hJVsX8AEppmnve
Nxf3B4HgOaG+tDTXd4W7Csw8P2BnmaGz/EPQp/iCkO7ks2L366PeBLVaWoDWJrJfHTU4HmYEADgZ
G8gwJY/NGur26bwktClMPHi86sOSDDQm0eHOHf7P7Sqt+L7lCPmJyscpMjYxnIEmn+A4+uwQ/wmQ
K6fi1GIfXFgRgR2oQmdZRZ3Ng28Qc+VEQEhzLjNnAew7+LIt5P/Erv95VxRgGxB/9Pv6tDl7mQ+v
zCtGPlEYsPgrR53QbC8lfa3Us5LO0+qMBQq1XQ8tfKIAz/C1zvsCD4KPPc6b7cTAeQFUwcmlWME3
FyDruO5jiDhqnayxHWkzacqKEyZd210rdPSB9hBDS48OuYY1n7yMz/bNEtVf1oZC1m7buuNAXGk8
gQn0qJHrLg1e34ZpaEuLl+kIsI/ma9M4LVQNGSFy8VxN7dOMuuH4wY+iSsGiuKRExFBQvy40zgXv
8mm0pc2iUiKNs7S2wTx3ByrTc15Jx7Anf/2S8QorSGRl7FokxT1rog31tHYbDW4hEdKgbOwUW6Vy
P9gRbOLC+VgBge15VNxG/f+p9jc+oY9YV7LHAU14tNThsbvK1TbkTOQqJmPXILL1RAf4xWr2Y5K3
9JM9AyqLnERhms6/O+BajO99AzI2T0p0aKJN0ZaCyOjFeWU870Cqc+0a7CWETTZHO6mbxYusUbYP
4J6052XodzOC85tLU+hBNZHklNYaT1yn67UiaoKx5iagdFPtknqK4m3V8uYU8nTZAh58LFvb+y6c
EiQyDLRSPaao9KfBQnteN7xeacNq8wr4yB9PyoqLcgoAth7pYDYF8csglvH/AuKnWDrBmbmnr+Ic
eFGHESDlwfRKC+Tx9Oijv+6IKjIpV1zP611+xUlrQvIJaW1iMOdEtPeRB5KRyXhToRHNbPsPJHYA
D//zEU4Vw48GVisNH3jj53FJTDDN4WRWpNDs7z4Jp+v6XV2ImeOhR2jeoUcX80Z5c1JtK88aL98o
vctNFZhVsxCadatBaU+iG9JEllun3TTwMzsjYxnbmtIGF3v3Xl5b+yZCPeBxZ/hU4+vphDD08OLX
4ZjK8l7D+77+bx7u6zUynflesILDM/+0ijhyjNDRXgGCsDmZq0CSNdnwbVsM5xajHVTCPT+/ooEA
AUlOaX2tZh7etAJ6SaPyIrg3dK7xxD3Yu+a+ROC+mN1H/hxRXwZCA6jdIWK7iWJbS9s+lY5qsUKY
xjRWIQvAwMGI1Sw58GYJHkuWg7Isr8BY7H8dXJuOn6l+LfV0WXZ5+dW+nZ4e8wKI5iFObBHY0b3B
uRZsR7haDQ//01mTvNy/xPJ8GX98FL+yDd8AjNxP7g0PH8rMFUmcj2H2txxO41ixdGOnJePvP6m0
9ke0GmhH9RSU7rT6a8qP4GDr5EJtiDvHtaHVqaLEitaWKCuF0YMb6yR9c66O/ywVdr3MLtTSwcFh
8C5YXct/PtPNze7NMwpWAF7S6ARiy6jBVdVKTdhmddTLFUysolav7HJxIq+/0YVbIRatdiIDIl4H
cxnGztQBJGkEGSc6FWtIY1xroWpNS6HFm25Y8XfF6X6zzEdpVmo1y90XzAclYUnNsSlWmLQvK4nL
pF428UkACdGZev2uDmda1rRDHlUx9Yr0lYPbfL9q3RWTqG/0b9vdaT6P7SaEMxgx/hO+NJtATnux
nWtpMWM4r5S6ZflHF0BAhns0p05ttXJLcd2Ec9ztB0IFpiVgNedFGgiE4M4feA/ZQzutb672PR8u
6uX2YI6AQUxFaD/Lv4uhlmNY5V2bCN+yl12JZKFGbzQsqdfuCjV+IGIAwEoB++ClQMEQh28U7AYU
7/Kw/SCRJrpslEayrKz5Tdp3YUnXzVq/GnfZs7D6mBaANzMO5rjLG/9VClULrwPUnlZAHCWt+ZlV
bWWbTVVCn96kRuHnh618xizEpbN9PBRfRAdLasEIHG65vN80V+hSIxTdfGf4qEYVxx2bTqiGXsPD
jIEufk3Qjp5nUxiBJCO44WQtTwX7O2dza9NLVH9OZR8TuuFiBXd7a9UDypuNafU/oA0KWBdOg0VD
EQoHyvdE5J3EAKtM7kNP+f4VUT/Wd2/IhAV1ldnDF2GaOvgotHEmAQSzjuf71MMfD9yBgzINF8bH
MlFi3+z25uHGmQHq7riZLEU/Ja1sutoUn6LtwOhsploYCk/NSCqlA7gFhdKpshnrzEqilacxcdWE
6AMDXxGVBtWsHE52Tp8KbcKFZjVWYYtCLWe4JWUW3zI0oN5rK/DFm5IexPGnnfbkanb/MmhC8a0Z
hOxiPvLcuE+JE8A9T6yf8TT/jtYZR3MYdrm3mHSRbKrTLjBRq3nvLKuy/oWNHwVEagFK44unzJyl
2Io78A1jFdrYgyQK0Vp/7xpoHvxKMeptTFD6ZMlQN2rN/VvvVnI9HjqA2UGQj9TJT2leK+t2cj5j
5d7qobOSMGpIhbGKMmfMCFxbvf/lKOf3wPAniBTuFHagqXLgF7vMdW/8ZAsVFd6hkjZ6umXKZ1VD
aYe3SLbotukKifhl9RlTeQz9OH4hBBknDB0mNvk02le64pQg/7vXzT0rzcyJqEIRN+m6lo0Sf7dS
58SgF4i3+rQG8juYwOoVAwhuQO7Kb7LcIaKn1hwJ+CkNsDJvFqBYa+ZYtCQ2RyAjqb/A7npLIngR
i8GuzvVwva6kKD9mUsuTqEwGzPo5Kd+i+RUbUkhDRhsTXi/lFPI9QT0wT4vBD5e3sUYcrVxVgxM4
wPZGCdHlyOjinuoi3LLtVDazWKoHdWN1MVOubQ1e7dA6RQXP0NoRyqb0WwT38hhi3oDfnNmqhuJJ
1W/RoMYgZXZ/Q1l+AZnFPyJDFBRVaSUXw65TU8w80wq6ppGRkrY56uCpnoLcV5E3N8qnXRjtu9CG
G5in1+e74TLbrPLsaIBP/SeGgfVddDZglECbD61ofNVfG8qbM4GjDHfU2scRmCi8LqLE8KI+jQ+9
J6DUtXQOPht+mDeRhR6lycaiapetZyJKPoObax/ISbFpmZxGIhZrfRsf4V1NAmS2ih1M+vtHZNYq
Ppz/PXvp498TrIGpARLI+9XCYURGWTdxVjzfFzXJ9j6g62Ck7o+CfKKHu1mABxPLnH4WQGb1xhMP
+wCJS3loA+/OofkC+D5BWaZY61NtwEev4HO2Gz+/1GCzZuzWOZa1EpAuaknDoPE7Pz1rh1E8x8ib
lcwlo4WkcRHDgdSDzYJqSD8JXtx7e9zjSpzjKVUpw1Hsz/pcVfdlSh2qoKIW/ywQ2El3QNieDukR
MnOfNUtkYq8GYot97OUPuizTWfRAxxVm7kX4FuRdvf5j5T8fk+NB27VilyGbFjoklh0eStW36KUK
8SCrasvAbwr9DyqikyqGuMz8nH+iQRiLJWtB3WbLe7VBzVZH4TjQEIsCYM6fQhTPMqUDZeih8WFO
0NI994BOtApZRjCpmWhrbTEn5kz9IUcerDD4t1P+VqKcqFA5zs5BWDP4vCaDQG0QgNJfPugAj/d0
YdgXVCLEzeISH/KqV4S4bzBkrIeTV1PKa37pOS6Lf/7gDOF9LLdUD23YE2MuqlaDWQBZ7FDDO8BT
z0O/Rr6aGvtW8slv9QxRMaZ1pHAJxEtm0E0nij9x8enMnWA/dIQBOF5395aavMKKfLG6Z93C+AzR
NmrWH8eoDZs0L5bTPvupqkafUa9ulK9IrpoCqUueheOIm9JEdn2Tal4+JhvFwK6U+Ht7IXjyEsB+
P91rC6VMO1ryy58OnimjydbcrnKu2PtsKyc/+WLFktBpE5ROzksvTBL+ZPR1e9qbsn4RV/Z17Y5p
sEyuZHZcUy46vDGFDGDZKclzLXjctRPaRoiN5W79LVIplfzYj+EdYK3xQbf4WW3WS78qbKFRYqLg
dzxNAti94hz5+JLZVqhlRgZzVzjoCU4MyYstx2VnNNzohtFVkwC+S+HODXYHfhj/4Kz7xHaSwyWB
l0bFibJTjbH8XUa5xpuFBSPv86RM5TbMP3Wjh1Uiz5Sjvro7mS14f4qeXzZtjWDt3ZHHZF0uwZRe
fYw0D1e4j+ZcGtzQwvjjll2kjL010OukSAYbwr1DDmD97t/DFnXUcpbaYPcywjrloPETP+ccDLe4
iYgnrLpFd7SOj7GQWDEEFtlZuEUXzeCT6vDqShnovSB9flYSj/zmw1mD63GdSyd5t0BJ7Ype/Ujd
HrxYIh7bkJAkBngwae758jiiOWcNumEHrNHo79qVnQnWquCPxprZ25cd7FqsDBSYLr/l+tAO3Qbw
CpqNenLAUfLhtwVuccrJCANa/3wQ6qTW85yjjzgazX883/nOYN9xnvg4FvcNHjQ1vhJcHRuYAAf0
TYizu91hti7LrjFXf8ORYsAqrlJ607HvOQLmMOwmI/aDoH2rkJk08lQKs0Xbqq3i+941m7v1j8TF
hkYV3v9eN/KaN1CQ+YAj9MYBU2r/2SVgZ4RlEOHh+8NIvjgrlce+wgj4q5pCrVaIljkJzGQySDrY
geKaAziWr2zJhghn0fo6lLmzOGcD8r7HKbjR6Po6S1zhkwVT/uKmCC9LDBcU4sz62hrD2c7/9qOD
wWdec7kSxXqKr3+9WeaMzH0DijGh1UR4dIWj3RHyg8/YhLaGFd4Rd2JiHHMCxLYrE01CGK+mSu/A
zTU0TmhsewZIswT/dMynOLpp7f24lx3RJGTz1ZBmWXcpmx8AczBmQzJ/lvi3n2sIFTlcLszjLzZY
49tuUdVyBu12Uo131tzWrBSj7J06Bdc5bP3dQs6pE8ABhApVrNZp2hDGTC7qrBej+c1rCVeKmpIP
cW1VeXWm3nRtADW7oDBMeyuVuCdYf0EIs7X5ImWE1S/33DpRtK6xwf5GW6VlXBvzp/24DQUz0QdS
PflmJzcD5r0lkDiwud/Kt3QEMxcsFbpQdiilCac2JecVXT+9Y2kUpTdU6o19ugCkjzKfZjIqcASh
FZWa+pA3EJ9kik9wkEPkG+ANrht4/U8GPWg/4AI1DVRahdphBqZF3XfvMMXdfegBc/g/APfcmkTd
Ddurg1isII6qMeTMnmRVyMKsQd8qT/CYHJm4ORirEefZoBvAB8s22xZdZIv1QjDjIxsqzJhh7XZj
9BZ9c+A69ZZMH0vnhc6tR3KwuQz2N+cM/ubsiM4xLxcVNUAiqJIxFd2Yt2BaoYM44eQvnttgsJCv
hnJ7C5/sEbNcS4bZBdi+EDY7WbG4KdkCXY+ZrB7q9x5ZOf3Ld8FVMBibrU8BMdG/Sx77Kp5AgBTe
DdEt6dLBD6RtHQrAUO/qTaZfLwnHZDOFqRAi1ISlcz0ojlnx6N+v51Pib9fn+xrYQNUkZsi7JMKb
jqDUy9o8N4K3D5D0BQWnRELitT12jZiu8Rx1jIapOY0lxs7uv8wB7RHRVR/FpT9X9hBva1LIpdZI
NWR8Fh4nsBd/lB4O1pD2VDx+RVLtltq2R9pDgOG2v+OhWiqXN7tSE4nOU5ohqLDpROXRSPGW9cou
bcwS37uEiwwxiEM30DuakvcIw47A4A/P/khOoaWI/zbsQ7W4vPe6xVPHhdN6XAnN6Y/MplY2AyX4
9NggoJNwF5rn/JxzvSE+P4CPVJcVdyJ8NsM4+T7OPW1c96Fs/Gct5Lxgap55NIPh82BDJO09mPmF
RcCYWTrU04wIlAqb62OOQaOymwCW4m6qIuedUjcyOYKn42FTMlKXy2tFItD0wS021IWWMGZbHWCh
GrDhYg8rAngG9O6d0bzs9sPjXZ38Y0tbQ2A+WLvSfIHNL47jDJCzP0CGqaBt8IS1L9r6Oo3VwoKm
nRO/jNekb3WQZpLaAMKDk3NZNzRZb7DIMwJIJjmcP5xbGyAxqIHKNw9sDo94F68nQRoXcDf0OG42
QT8FEJO+7V2OjxOATcH89Gy3nvwFUSNfQc2TmaBnKmU3aFgfpVJgBMR/gTGKbcGa78J8mFS/jLdF
YAY5EAxuFWNAcJA+hPkBXHcELiBbLB4udjKcNwWkocVGd4IoMk1t0k/Ix3hVs71fathsaphghe/E
DsyjD3G11tlBJRHAPh1HcxLmKB1Sd95KQeNESHTNufTu/OsjMJwmOI9p4Q0STwystq+A/ZxUMr8a
/oD+L7ezfuTobpXOJ44hsRW4EPG4q/ctVzStjzkkyGAn1k+ikf9JxH24vWGEeIfoLPgfpZWUm/fB
O/qOjiHiz9nBL44YGnHkDV/B/EWLiJBzaO4j4xMlIunYlkPGYL1M5AZlbsmue0kG9rQqHx4rv8PC
WD8cCoQgMrTilteN+BTraUfwejVw8isA4Gei3wNTQa0mpm96262IDOfSpAj5MvlT3+/N6sBwH3CF
kK0+nKKiKey7kymjTM29X6ypYDyKHR/9FN6S+5Sh2uBwo0+JaYvSLPHYHBQyeiPRJ/SWLrBt/LTq
mlSBHk25onAi9ONbXtlQCrUQ5rKEH+n4BtsF0AxjnEpBfvavOPIztLkYjGPC0gMMk3mv/VE9blYY
0sMxP43H0zfIJ3WuZ0LFQU+eE8KdcOG1japgSZ1Oi3eoS8Ft0z+FHJJdtQdNhAsdsrjRq4JUuWJ9
II9Z+0SO+W2xxBr5Jql28tS4o3kgUrn3Y6MrKTBc/8BolfK2DXlRoAMQDGVwnC7PvOIrJFCz/ZOu
ONvAby0xJZMYuwtczENHpH1buwz7FAxXAMDCldmDC0O1yHnWHTq09vLrXRaTjSmK7B+sSC81UnJL
D4GdaNkRMLvUY34maVpLm5pfJJ9fXxmy4NHAdrfiJeUuVHJTdvUuPfgOlgaD4/6+DcSyrt8PmRpN
sxmYZVBa7jo5qUWlBgdR41AuqdfGoGxmpgRbairioOeO9WiVDgMOf+VtSSW36S9kcp+Hdy6GdXrq
4WbQ7qhIDBZSU3fAkY05VpsOx4a1x4OmFPK0Lm+qfNOh5mplR/Gy2r5qd6f8cKGDJg0OJUbXLz1B
wLCwdb9XzL15AtAoegZTRyaLNh0MMxCRws3SpN8bPFE794iVc8doHoR9V8rruXthCezgzk/NzW9K
6UqUrQDl4CfuHotJR01ziAyNTg/fiRFBuGjO7hp/LP+f76FxYNWW/TPPDGKbj+C4CMiZlz7ci6Za
AGgziSrE2n8ehOjuXRM24SJr95wGPBScquhEAeEv6Yt6Vhn7ByznqFwYJCwMcGahxNyQBWCcxpOW
3YKjcHP6lUjJOzfWvK4EJQE8iMl/W0jdbgpYhAGYESZf28QKXEZbpeyEYKXDUjpKyDrP5dBf4Wuz
Wn2DadWhVuKcK1F0B1HdaYC8iqzE3MwzmR1O9fpGmi9qTtLGNZ4JmIcm/Qe+0F7z+TBqKEA1LPmF
wRxnSJ1i3Uig9Zbi9/Esbi3NOjhDCwRKSYLnNCElMUk0gaC9y44XziD4aEKnGfI0Gb6M2w68l7CG
Lg3zYEAyad8jrqElAzizlOdJA66CdZHhph9boRHMO1Md/kyjO8ewf449Cu6F/HaCwChmpPlxKAhn
xhTGD0Fa6YcR1buvVl5toGfJ+eMYwJrDPKnTZxqMJy9Zm2Gi4++wtc+r9EYAjniT+m8AOXPUW+7t
qhdJR860DSy+s9FyjYKvLgbxHbHPv9TjHxpJd+iSv//tEmJbKmi0bqZzt4gGW2tWO9kbcqD5hN4j
UzMGahWSa/uAV1rJfUtmSKSv45G4ia5nfyi+0iUXO670f3McbK1MpMhSkOMlvsC94lkvyPO8ltna
u/5LcaocI4CUjquct2E7KqcpzkOXLItyCIP+RldNy9jtEfHjL1TzwiKwcMv0BUB00A5UVbx2AW0g
sm8RCsQpMKv5DZDpMXVueg0fI1l+O2RoXcWKNN2kJMf74jarG/tp37WCNbFKvhwebWZmRC5l76C/
vYeZgmZB+/Mpeww+r3T+sVcET07DRTiSq3bCA1ICR3LuOpxWE5KCC6WrvsuITycVJxE/ob5d/187
hRmgLOg8WOyO8QwfGkJbmPBo/RnUYSjHdnDyzB525f52nnsZhw4cKs1eP+Ss35G3R6bb5W704YRK
unD9kffQFYnGKVDYmqupzOifrnWxOY+wdcA54Cel1MeFfBGg7xonbV475dISYMYsP6LH+L98YFeK
lBMNkDF7u8kBzt+Mc0EYqSK8wuE1pibBunWlIQVlB5w8X0Tv2P1Dnq3zMsD4rgFKJklDH7uwcxym
0/HysS+Y33uWJar7NpCE1+ub0HXgHgb14BMtx/wooBYdyBLRPNRbVKqSNjUxI/di0Rw5A+pQhJ4D
y1odgEtwJFsD5mHWxNGeojRmprK9pnK2vAJA+AxCqwSx/pb+81C8wlUTe+eHaC/1WbKJ78PqqYkj
Nr/SS/mo1UbiSRkG4K89THHXapdA9qVvV8ZjoMy0NxObVYHxhgBrEhTHMSZhmGRb3DD3xpcu99hl
5JP2EAgqF5r5gwDiGNG8K1Z6oDc7GnF0y5lCu4KPisDDt6Gozi4dIPXTQCNfb6rg8XngnKlLOiOE
yiIbryp8xHRZ2R1OZNWihAJgFiSB/QRznut4s9eJDGLwBbI4f8gywsKFodu2GnEKdFxEkZ9JLpGh
F49qyS4GK5fC13AGP1rhcf6FtNpD/4E65HgiHoXfF9r7Wa3SQkyDzN5FoNdbdWrrhjqbfXg1qocJ
fI1ImjMlfjQQre+nco2jT+sNkLMeX0pXtZO+olGThnXKx9+6zBPsNuvxIFIlU3bqpEXjCcmY3fDf
QVfW739PX/j5O/K7UMi6HLDUuQqVmxhAdJPj/IY70XSsDS8DuNR1Q1YEbmIo5JA1g29XeoJfJj+s
lsUMX7rD4H4zYovRaWy4X0NXBO2eDb8g/i57GxMmI84xUBoqY9N33Jv0ovR+QNdW9pvdd4YZjM6D
UHoSJ7jmQO0qTVRDF+rBZU2QMbAfkWMByBX573umYE7toGkB2eY09HQ/O0wBBEMCPGoYTa7Jt59U
0VJXk+uxz6gtpRLdmoNmgm/oDWVtErVJC0KT74C8Vm6dvis+zBv3sPi98tcYQ/VHaiJr4KDmFNcW
tKDiR4UHtzF8JTtvFGe7KS3Qss+Ft8QloS5BXwv5BaY/IeCcTLWb8xr+w71e+nqC1OQD9XTbpVT8
G6Vn8Z4Bh7w65QO2NBy4SxbkwUZpHKq8aN0+2zfO8OFWvZeP5JYw/w+FRhPfF+A+k1P08Mf4o6Hp
okZiQWj2QzWo/v3/G6N05aHQgfp15eJtfZ2bMvYuDjblDRXWP7gIGUbxl9m0Zp7gVSVhMGTHPEgU
2eAKl3YqAw1rX2cFL+bvrf6dDhFDWMwKmOj/1enkIpIk+m+m8u/I3xBT6HBMtbEOQRH5W2aj1E5g
F03zeWl+kPqyvNfjisP3dcuvZYqgeUNO1n3NaHKUkgxzJyzd5o9HxM9ofmBf8cOkK7QQAS7t6Tqi
g9KdsESQpVLcTNMNNyJbGArpxyot+FxKLGVPVF9a8mylzxUm0+DN1DdlcuLiN+hQbCnfEahz0Whu
VVanv8eo3frT2z5Y1ZKORKWmtw9T7yxSiAlSTh1h83x1W8S8MKiEOzY4D5TKu3+UehGPSHk+yFyU
9flh5m9XLRM3RZjAZaObsjyyQT4tulPkOMLMFgEltZ6ipZEmowq704eJkO3nZ/y3TdDIggXGyaCl
zV8LviFvGEzqlBcxxvy4JpmaHKKvAxcewCDk0LUe8gWk3nfpfxUqidTHvQnJRGCSGCo4W/gBlRb3
B3efkWTnwGY4lSVULaWL9NcXcL5xqaOfKR5vItas9cSaIGxhvD/yLK4tQbSuYsWuBLwXgPF97Av4
BZDaR1jitbRDRfYQhEvNk/j2ZRJffcjYRVeCs7b17uPqMiC1WWUWngQebUpP1323EYYMJ3SNWkUt
W2h3ZsKP6QdqfPjdKpPQ6WGwwDGpntgtzkndaZOGB1/SpMzBkgkz9QKtMzd+b4K+5KCpIHnxYanK
E44AMPJ1yrQnBO1pj+HbZULM8x8a7pEUGqEBMagQ62d4Mfhxn9WqYeMryatsdiDK+ANj3EzVrCee
Q2AhafuI6ek6+yAwzMANQXD7j9YiAtffxLcYuKyRwQoS8k0IXEoaYTO0WKHgqAZMPhCGdXt0EltI
AVI7OYVa1d5iALLpRJJ4g/NlQnYHct2Sui4SdAHRTYqW+UyfuAZTbRvE/wiWij11LCO36cjh1OdW
Vls62OCHdyumCAE8rUCF8I3zzsOgYMazTfajvg916KzxgE3SU5Pf40OvxVtsHlH7AGufwRG8Q4/S
A0lYlR2qL4k0uwkvHf+66wJjrIl1ww+/gnETrb9LDFsqWneBGzAm9elwWl6bw2Ahep2CbAmJZGjM
Eqc1wXh77saCuEl6P/ztaZvKweI1A/gFliS7H8RSGZ+Ch3MefJsUdB8nlMXCGUYwczy/5izfwbY8
HGLeUN4oFOttVbHk6HXGhW4aeQKmWYial3HDdBGRxHjBPs7dgqAu5JRHNmJ9eal5Au9bp+SGbuXQ
Tz6YhBc5bzKhrDvmFYP+Lyj0bC3LEdU79VKrWsIZ+2k6tKEtQotXCqHcR2RPvE285hD4/Xha3qCj
2NP6aOIdE3cVDUiup9+yJuabOKGGQwVohE3C382PSTq//bcNS2sjZ7vGU4O46n0bRkxLmg9YldF4
/TpyPS/ULXBv0M6nZqwijdkHKwX1z3/dG28h3zhP5gGUNBCSLlD13jjLhzguVGjsasQHu/u4ohVG
fc6gXq1CC9PrKjhszCybBMGudW7Uv0omcfqxbwCBeGMfkasZxncVGKZv2HXkY5kCIB0YTqhqmv39
NohpR8on+tN+WnWHeunPCgLnYfJBFe8loJQUQuH1aYSjjaHg98xhSu8aNjoNv3ZtQKoBLMSfMtEj
9AbDO7LoDNmMlbWprwUvWhZyV5XuP1eewtteyIaHHrJiPjWxiVb5RPvPVX5Q878WUTMb/zy6C50a
E0BVtFfRcKjTHg1wrOqTjC8I5bYjQz75md5nWXG/1ZHSgJvSzg1hnBkoQYdnGzKI5bkhz8oiXLHW
WTp83i7ZrmZ3nCix4Whk2PO2vBLtS5au5rL1d31t41/IAFIiOlPA2NMYe0xsaJvWM0fpHfPq/mHc
z/R1nCLaEw8JM5s9X5KqHe2nLpDEJky/0LGVLG4CCUZjfzue2s1FissBZkAD/BMwJmV5GXbr8Jr/
LyrWjXyDfapFv1LFTI9DIWWdz1tH65k7KiioIuebkegrE+2mJQZJ9HwZQVIXng6yzITRMbHGs65q
nyQ0WdSY47OXN783RmVq/n4aWxrHlbxWiRYX91nSl1sxi/66aa9Zy8fr6X9eZM3DXHzns75Ws/Eh
fu52aFw1bsSJURqysGLzptZXUulmmqMDtBntO+VCnpWLPny3f6YbiGQP3OWhaVobIyNQcT+G4dYz
uH52xfVKxmo2KopTuLc+5RK0tNj3S+D1Q8QqlT0LY6v7VqFPsKdZOW3mdg/ZDzMeHsarENZ7vmfo
sipXIR5d3NT4kBOQmKcD24B/UKCYs2RiJVVPju/PBOP85rJMIZdtUTwnoqhGeIZTL07hNMeG9tCL
0Nbikp7nm6EJuqW/QOP5kqKdqvef7DHNBG+pi6mKzZDDHaNeYsfUViouggAM9XzfIA3e0KoQ1wop
KR0xlQUHGHnvlF8rNhRaLIP6Phe3OWnQgqds/SN3YoP0vgMqCijjcCvPLxOsAeelBKbglPNO4Keh
qsmbZYbkrHxIXeOuyUoGQZtcSHCKZb0sD4Sb2O5y+Wgwx++8YX5YL13Sev7hqGj5Nf/0PHEZrdve
N855UwycYkT/3VmBjAkrpZ/gVuOQbDrx49eDXvwg+8zBovGfTDPpYR+cn4aJRz4U2ekyBMb7lsDQ
I3JGu59H0rIx9d1FcnJJcoHcofFQxf/lxpPgM4fYS6HuoHzWJJuKncL5J033q8SO0V/caNh+72L5
NOiBQHbBuoafVLyybvkZJHFUKmzcIAkvux+npLDMdakYu+xTWHZNxvG9fg9LkURx4Igz6P/sLhAm
qYX5GfDXdbyjuIleznFThO7T4WtB1esJXgGMAcN9s0qiLupDTj7C7ch2fB81gDrul57yVs+Rxqfp
ygeS/ToZ/9oINyzFrCmxTj6ioowf+eo6mmbFaNud3IL87NLRzErcZTi9S2Rc27T6NUYlETlYcwOi
Aox8m6kCeYNrEiyoRHmxsKPriTWdHf/n7X6HpZdN72xPPH7uBL0AukrmZvuFZ9maWu2YDgKf7bp9
09oxdZC0ZtBm+aeTISrGif4XhjIJLgM5wLIS+hvB4PiLpIv/PDjKPYgnuRm/apCwNGhSgNTzbnTw
TepJG1Wyriu4Vxtr2l8xNvRAPacyHg9xu+O6JHew7bH2JYPBVUbayc3vSC/NLscsr0DGta4E0+Og
rimQ+1Q5tlvkFe6YxZSbSZOHqRsKUgIyirRC/xjH5lBm2xsrKuMsRutGXc1O8RYzkvGnKmV9q9UM
zgtPQBbs39RYce+jf5d33cFM/pVAPWncUGUeyi48xob7cR9XbA/Uh5CcAkpXDatrRJq+UUTuM1WS
5uYFfceqWV8ME31G+zFninxmYv5EOgy5IB/Yllpoj7ZomlMLsUKkGUbO37cJgt1oIww5e9/BJDSQ
Dq3S3ctvLxU3P99rfSwnG48LnStIYSRYMMDjDSlo217cFrgulutZDEk3irXVzhHLNZ5vOxcqQO2H
84VdiAjK+j9lV5+MGPhEL42t/pGayMdFoVkfEUCYGZlItNKtz6QBtXDv49BHPFkUMaRDg7pqr6zq
2N6zUZ+bBrS0P8gf5bFZgZJiuOg/MfU3wXn57ToleeIuNnO2Y5AZf5Dn542UKcyf6jwdKfw3Npek
+aNvkPuI7fxICjuDtvjBOxzRy8hWDPRsdFv03LnkBY/QStJgYkY1x8BTkGYgqtfhLW91szB3B2EQ
y+T5kTy9EE90nZkrYiw5gEr0xr/K+0CIqn2uedLYnw5BxvaHMeKfxW8miPhcWv4dFuJ//Nb0aUhO
VUGveEkHZANsRlkfCfUurrsb858zVkL1ccO2Qc4YhHhqARTeua14xAuM0vhfxdlnE1d+kwNrTdyc
aqQ7MtKBVtJ+bGIJewAvgXAcZ99r7XKGTHJ6vCuVzu3HSMewjwfOoFiIePLTE6xeq8is11e51VQ2
Wk0j8zmKYkGqj51PVW/0GAVhjztMzQK0vnBiSIWurTQ2KBVYMdk0NX/9AB6Jif9VXFpfF7MB+jbb
msgnz4yx0IEL54lf8h1B4dVrOCN0vWYNebkxowOP+WKZwKri/jZCZJviEiCtPFkDwJCWEuTo3fCA
qhU+Tcbxa+NBJN0FlmggVT3CXGbhbVlnwjNjAZRD4q9cUofSPscMWNbJ7uTrqt6vAzSQztgHSerQ
VZ1hSbSSGUb91lvcumtrkI3dUHZJnhVXW7o5B2cioZTK/bpVanXjqN7P6tTvbwj/FWIwpfaMpQcq
v8khh3ZW5RZHNcJEReEXqbfu4PeqnrOmiJQFCpwUWyTOfV1PCPDh9DLRA9h51dmpZ7avf3ldMeEi
B0lGQlglSbHgQlD9RNpcuSbLF2XvrhGVPyeuMObp3jsg+5ZiVprp7mIdjPr52y5Se0GgqPTnabm4
QSQLYi/Zb1WO29Wix6dZt+6nW8TfZi5WVTUIDHA+67r9Nbgtzuzn8aRNqNRzLQzEcbSracLVvVOg
M+cE0dgQ5dujCXzOlL2XWVTrM8VYFfgn0ntY/shcibXz+naygB0fpD9pGxh+/YNpF4l5h2VDe+Gs
hEs07gLL/WMtawtFqjMAsUgUwL9vla66f8YehUXvjIUDpcuvYETgqUYdRzTYTIymlNoO2pnnHYdP
syFKEPlqw4wXS+uuG980hYAqC35WRYw2I7jiEwNO3p2iFtf+s3RwGQ1SeR80Dp8F+OsN6NmXozPr
7ya4orAi0HZWbnblwAsWLdgZg6ZVKLyjHTQCHa4/WHDBe52+aPp2TELWXu9bkvjRc8v08tBehe/J
Eu/gloyArHfjgq9v5wskAe2cRyNG+Vh0sBAjRwe0z8JLi+6KUAL0cm4k3rebTfqGbDC09BmyaChb
I7y2CO51YgB2wZnoMFXeuce3FyHBS7m+j/dG+3sbGu6Ok1xOc9ucM2HsAvKVGEc10b4JdAQKdG4j
OuAfRvMyiafe9LipJfvUvNyDs/kd/figll6mh4pZHWJpUZcXjrmi7N9aXrvWHxriyAWhcYePGAsR
jvQ4zl+aCIwcxO08XeDJZXV/HEA892S591DZbYfQZJg/DtQWsb2ndFZX83kU3q4tB2quPkiyyq9M
uIoSRULb/CsDprilIhgV5w4WuN6RF7nEA7sVbgbL4KS3SaTwCp2uhR70bH138sYA/EUeRE96xDzP
vpDbaTaXaa9SMGAiFYUqaIdmmIlXl0NJgtbOCcFiv220QA4pm0j9lZBucfBmTUx6F5NArMh+mhui
Zbj2nrXdm6UY0xnWNV6RdWPa9K5z/OQ4LLzEqHOt4KyY7SreQeKL1J85LgwUvl2zkTEKtpVD7E2K
wdz6X/yRA1yassF51g6Sl82EPQoid7UZ1dmIwW016Koc7WWhH2RPR1BTu2PNsKMxDbePjfJ1/0D/
bVHZhDI3zCPRKt6wpTMrlfKujMmtNHcClrHtqKy/kMmBehsIH6Hc1wkrVC65VUtEUxKhFqdQSRc/
STrWnSK9rTEcUvd+2Pr7UJtHzwkI+WWcgj8xrPmOQIYtvDUDOTJkHKC6vTMgaI8nb8atr3qzZQl+
K7R5GC8WHjy7dL0EMoAFrM1ciKRcRXG8wzmJYtGoTck6JYiGRiSXbC+glRoImsvn83SVFMrdHSH8
ZTsBhPdzYnKppBUTq0jTNh0ycHeA6Kg8A9Qt/zDRl3HMeJA54D3sIN98tnLEnuriqlMVt37XfjF2
8wXYrAFJMu/AEirDvDg2zgrgp0BIlQ91WrumQigdYalusByPRbMY/fE92PpQIDHyqIJbSxpkvUlh
AACHStCTSR2hQwV+io4+YW41r8AO0A/Z+gQ2iGCnAGZIRs6dDErs66TKgPnYi6ijw2ZguvX67DBl
0Om2UkBv3w3WMiSy/iWLZd2mEOxAOotbuOy5ZyjJQBqQ4NHkA629+Tl6sF65/uRtvSyk7pWkEHcX
H6ORaUcgh2xhYZz1q350IHKrNIp8ES+ly4V69wTERWDy9atnwAu5hPFtO9Yxbs7uOzT1FjF00EFb
cv3qooBbl6zGm91uk15BKajbLIBZ86Io1UV3KUeo6RiXr2POL/ulQPXN9xeLKCz2IsH3kuY9CHgI
in+gqUZjzl2mhq1bVIOZ3T2T3SiHCM2YNHFpkqXWJzza7+I74FNQbp2Kl+cuR2DiGeOxUfVY4aNF
Fu9NgRaH6xYldFahYSdQPfX8LG/uzGM+gcVqQUSbaugaXZW9Jwmk+msy+Mnn4Tn88txPL6hu2hQW
+bHMTmNxj4siY0ZcT3yVK5K4PLvROCwndZzIj2arEoLFzsK9qhfDVNGH4Yt+GG3RGgM/JJrLCLAy
f/5jDLkAy8rZgiVBe8ffhxqTV5mfIaxlNZf3QVkYiFQlS8tdeTLefw3j6GP5KZKOyiP8hdFhzfSE
SRx5nmFK20xqpGUKzsE37Ws5BSHDSlbZvbuCa/htptCXEw36Ua1qW83ep4aSz13QUmpAqYUHOmtk
kuEuelYPuk4YHANodirId3py50XM5LjdZ+zYYP1F7tMs19mNlhYOfgzukc01KDmnrYS7vco42i2Z
uxOKkq0HrDMwK0oT4oV2dEUn56iE33Pwn5ksldF1ZeNJJ4fO/IUlGbqvDrA6+uAYz1VLXz7IQz6T
zHU6Bw1tqF+MgzftqmNdEz0qNKsLr4xikb28YIdX6s/zHqbqh+JIfj7Htlo8ARXYK0nX2HQtR38C
kMw3Hr1xevHQFLeVdtvkYnpGb5WU94ixlZanhYJ1JNR3thZ4mOfxptRvwv2smlGEBzyN0sDs6mV6
JeQv6QpyaiBhA/+MyabHgvSnkEh/1CypaippgeOkauTCYJGgZVfielvXkLGGVauzdtY/QNSAPST1
9tgPdpn9nAEa2jDmKwa3NhhE7Lak80fnH542xW7E7YNF3zONBsP1XtITGya+95mHwP1nQa/WpYTL
glhRtZChSdcqqApIj1mb8dqgk4dJB+A1FXe70+AFae5BKL9OOrqjRYdr9/Im7b1gIcrAa5AVvDPH
zvyBUXXyoOg2s4mzouUWvkrhe9ek5YyYphTpc2oNrkqdJXpDJV1WbKUD+VQVAx0825EdC64Xo/TW
n2GxE8vzaKcHb2MDLXZuk54ghJJiKpJ3KJIrw5CGmDtSzENkG/HhiQJ6TtMU4eAdJnvSk+8hPTEB
LD3LCDjmJphERrCFP9fdkGAxKdARqqoRH2dNOsDcmUA0Y8jYcCcVClI4SuuWGzcvEeOhfka3mGMF
KWWXJzPxP7UB/1QSk71HSNq+lmzNrhFHOsMbpDr9CQYQkpi2yASU1lSoxVC0oDuSSFpVzJAb9vBt
3D5tMueSrCZiiQi1gplYZx9OCUw1beJH+n/XfCzFR7rl4/IAkA/HMW4vxXK68wceLXXd3jCi/DNQ
/qbAG970wMLvGjLWOTzb779gY4eoDa2clG0hsYB1tv8Qtv5vUo+WDoXJ5K9rKgj6/pVj7ycbDoRp
6uGIStUhAy31jE65p+kIZwxubCvfzZEsAoFyZiSHVo5o4Ll9b2oaDdICTRpPqjNxJR/7TYqnI0zv
zcLOVFHOK8QEe0mbKpugkBB/av+/PJxyMHp7qUcNeLKpoZP2z1k6PCIK3aBfyI5T+1Eu1oe776RB
c0X1uAzh/iJbek4VFYI4Z3Hby5qROjl/oBZ1G/hu8A2mJ3BmTQrN/pCFVIB0XOItBJUPU0CCLt11
5ma8wwoNDsgCmVqD4DSj1HJWWDu5LfGigy0lQdw2rmO+m+EXfZwfzhLL+Vv2WEzb9OMYFu3STphZ
g5b2ONU6QPQpL/kQJtX/+5DlKBJrFjeamaKP3KJOxegp7n5QvgTQIsMQn4PSxlmGXL/LvxV99k5+
ceATY6djCJDJLcdu1kc2SctPApi3BTlm61oeqMFE3mN2wbYdROBULOv9iLQ/Al6/L9loOIDr/84e
+wR+ANEdN5u+SWjFWMGYKg/p5Me/RGclyyjWiXzY+tYQ+W9zEEFUGztC+WDuPDVEvnqBQDfC3aX0
1V8s5Utr+uuzzpMZHsuJfuzV/hc7rWMac4FLQCawBbaUNgeiegZE0fPzvSvtSRrADuhqMamuSEHP
BJA+z4vpq+rvElYtGcls7M8pnV5UboMkmS/Dxp4eqTIJLwqHirco7+gfsc5p/HKUAB75bOgNfHUq
+xzJ5PUca7KB/+XQ/SUB1YlVkV87cuGiuPZCUOWDu0b+1eAHmmNXVAMkh6sJvw0C1jU6y+gllt15
GD8GuQ6Y5mtgBbdQBT4yy8oE4mSOOlJyaGbIpKIdk1erwyK0mB5+9Jlp5NLizb3+3VXBZpDNsHTZ
xITkXrQWlVegVmodJ9jnUXxtyQvvuxY6Mx0QTKsW7C0K3336xLl7x8DMzSiH4CwDLDRKLYC30/lh
PHIm8tmg4bQnTJ9vA6xtdYG1Pw69CKyn51BgewmFsqIz3icmAAndjuh969zgEEGAbDZdRsZ5TRLr
mwGy4wROrorby/zgN7D8XCtHmtVTy0mplbTua31dBN1lnazsFG6B2f8jjJxbOjLrNnqbBFV7hzCz
nFrqGQKogzft/oVVb3GZfORRqP6/yzpDuZRjNwWXkVKKIo2V/a9j1QZZRe+wR4A4SZYatfHcINW1
h4vqxm6mE3VD0TEjnSodpyASUfrcGdzLQY67JIl9WJw7FH0hU2JgNPL+bVTBMz5r2CDJ66qm3F+C
pmNGpX95xJEGKAM/suogjEvKAwDMU85Waav3T4b1ptHJJ3pGRzBngb1B1XY2b9affXsHVDIHO3p8
N5BlaIpEZmjCLC7WjC88VlR6KoCSI651UMP8q/HYTQ35tRm2WXAIyJbsNyQS+2NLJ7mxN22LFaP1
x0xb+r8aYfycN6TPpXIlfsamu8tCVJwfiGS5CIZrmXi066kTFUgYXDlGfy+4yk4jo2uGYb60ckSM
Db9MCnWgJbGhQrB2I2LzxXSs51LLeRAWmsAgOvqY0qUAsZQYWeOoxiIAHsSdIeT+ue5DCAjIW1rj
RT1nntMHlBs5nmruUMSyO7u+odh8lL6k4Fg+KTDiESRuvWhOHNBl1p0jMJSm9czBGcfpiFmekQwf
F0VvQSRaKvrtAk2FgpoR2XezWhmt6MN3kmrtCIu7vZrkDY4dDoZp73kfBFI/jO0BmtWG7WQaEUls
FR2KVe95GCtwQFK5uytyS4YZz81kFvllO1AzkQKkDmUlTn8/zLU9Y6n/3nm7ax4WZtcTzqh8bey7
Y3Mx8apvZ1JLBLxfiVw0QlEz8qQN3LPA8iowQgJdmKkk5D9Vq8dsl/nDimFYgbRZoJhQzfr47qEy
u3xZ8+Zvp2CsyLaMUPN0W6N8X3e2lMdoJv5SLFbv2WVTSCxhFQ1B+bJD5pajwUhOyjbIHXMfO8Vt
c5yQ6PTKwJXq8D7IBMud971ESI99kMcklknnQXw58e7B4ogBkQEltEz/qtNBTc6PDKJegvo9e8GJ
G634WJEGDs3zJmgDPpOD9Z/xsC7xmoUZGsgcFNsS6fXnVq6n633FPEHj8sVZ28wzu9M/U28kFTVn
HsJfPaIOLTUCVFxnHJOKgPwToBBou8xCSMxt8dIdh3BDrgM5htU+nVI4TzIMAo5HRGZj1B0LxUb1
YxJcWuusKc78sjs8ZQCGuBzYv/NebDLfU/0SbYNMUUO46FqYLg15g0S2u8B7hAcCBR0Vw5BSDada
a77CrGA2iN5zI9PA99A0oKbnsuSnsBw4AtWtGO2zYrMc421fv/x9ihSbVkmqdP5hEi2Qzuxz58Hg
lws3A90zT+kx36Wacg+114LcjJdOgtEs/q9RiSTRjiqohFZzn0PkHwV+mx+iGom7GVyQINUeatyQ
MxYTB5XAM0288cnwOf9qLik87ZONrdeg5mZlj196usLSgTWtFXPQqmkDm+0vEq+GtQ8s+4a4WMEh
A5BxGBe/frdGVB9XY72BHc3fR3oX9rKPhqrSH/GnCVoF+wHztxeWq0adsmi6eUDsQNVNfoi5mQaJ
NBZ4gfcasBQwXIkCWaNgDeFsplxJ3JPTmVA3KjsKvL8DXZ95WWyccZQz133ZYAU9EZbpI80TwsIy
qsXR7ZioMiSzdfRj0VJ4VRRYVTaNk7aVXVgJzkOkdvRSheCuL98mnsyaSXBrUh9XS8uIksSVYr00
tqWMGf2AfJqD/Fkg0PC+vKy/unh/WnWPz0v2gmlCTt+q/ZKjsfO8k7xO07xQTK3RYc2a0tAGVnLz
Aq4u83A4L4Ec0Nsp6s5HHOsJOEFqrOELBk8Cpi8gs7wqkuOUz5Hnjz/6yLLyBmF6mvRBBnRIzUgT
8WokF/+cQEaV17eyejNFmu63mN5oo+NI5SMMZVkTxmy7wj/lxWpM/4Trd8Xig5hdb62QJOhpadZL
jJZIrCB9dpkJgdQVzzBuyI2Lg5PQKjsuPQMQJsrfHbDbnu8/3HlVvXIMYkPGOMuUkNHta6trtqA3
PbZ0sgikYDAS4nViNHKCF60MCQJCpxJNgYbDE1Q7zojm6NcBmZ6GuXIaS55XdWX6Ck78azUXs1x1
b/tUjMjL3NRHqwqKv6QBRh5cuA6qIfQrxryNzHP7hqBuo72ZZB9UXNDRcCa9IkI33khy08lkieal
t8WDqHPx2VlJhwDwGt0R/KOmDxzonq6wpfzJFmRPfFVejNyKsmrG1IqVZJCgrAn57JkDA3tLlHy9
/HiNEJ8AXJZS0qmQk0SD2g308w7Qf8ag1SAPEjuADDNGYQmFcq/vqHmFxusHqu/cvqEsd+MwylrT
9PHEo0U5cPYr7Fnyz9c958xM+x1KliJlJyzeEOykC1bj8vcjZ5AVaMP/tNnTBVOQ26r5zcC2PaP2
oXqTBhEwpLK6Bu6AdSWGokUqkAiVJV08NYTIeNO8AwwvsLQZEpadpyYiVigcXDYjrrT1inYe7FTT
/n3J21b38Lki+fHMyaogYsdh5aM44ZxrfnxWg/QYZ5uDW1onNWjXQGsEO5cFWPC5aRg6wVrs+hdx
rEC18l5IAlg0vAfidT3It3XTWiXzbfMJ92pFcTWUGkRW/Nx9/JyLF6w0/8TxMGtuMPx10bBSN/IY
vL6WgjPDIc7Y73IMfrA2jZb4OdrtzMSekGxb9O92RQHvX7W4C+KuOoFafzQz7+eylmc5jultybDZ
PRU0VtujVtGHXLS/5ymPIlSo7+UlK/wbqVXE6U4em1LcMq1bTFXbIy5zxQZ/Hpyr29+4U9FtA0nS
2B3lIWyGoTe5oPRQCmW5FcuSAvUxyVDbGSt9CormV3Y8DzlzO0rj1mHQO76vPTt7KSuRexTmHYgu
QVb0IFs0WrqLdpa/vA/q4LGJuYPxn7KAINh9+QoNiG9sdLU2Bnq8nciSGIZSo3EUby2mHAlEuS/j
vJ+UYTnmsAQvIp9MCUeC55BiMN0y6ZzYqr/a4pONyhwVOcDG/oMuHT3nsvpGIyvKhzchk9yA907j
Cp1puzxgdLK6kAnck4oOq9BKGwyQ0j8s/CxBTCacwWui/EMPXJ7B1pAQmT5SuE4QbNZVtHsbjFQp
2DH23UkvsaPff2sZmf5Up4PAIc2yU1sBDirDxlT5Y7TK0F/UMxGeH9s2LMR6+fs7eVfmQBmgsE8C
Mf/njjiCiJsosSvrLRHPQInfih6gjFWQhLW4UczcfzTiVG28Ag01Z/HJtX1VHlz4P1VXHBqqyluB
2GAwHITe5MaeiN9g12EGkhvH3vesKNlPgE8vC3eilom/hso9lv7Ygt3nqk8/yvGhgcf4YLbnwX4x
kIMG8bO16cFLn5aFgTfLBotnWGzBXcAxt/1DWHx+pEkeU1Fm2o9ML+czLXSFgG7tlbHDw29/HFql
buCiSJFBp3btJZZSocsWunz7jewX6gttPy/ISx2cOKaYnO0zCmcLaL6T3nHfz8sSib/LiByrAPkS
iZ6ip+0rtpz//E8kMp4594XOC7kAbRVuLeMVrZ9J5u0xJakvCuHD3qoFEIPrF7gv9cTNFtgioM56
T7YC4xbp1pWdY8ICcUyi225uhzNApvdYHZyOXXtzc8GSxNqzYVDxe+NMdRFs3QuIecRnP0sB0vkR
i91jz8uVnTjI/hPG8DObhcJ+Pvd3JHsfIA2PnlWfelMIq/nIU/Nddi6sSLAzR3qhz8pJSeSjmDiO
rotVwH7NlUhwvdrh7aTQyQ7qj2SqshbKNP4W7Q/vNnqdl23wCyp+E8y+OO4bY3EOHwqQfqAU8PSf
jQO+JyzLuJlfc7dE0HMFSJdtAtNf62zmXLr1kkoTVlL38937o79YZX2lDW114Simr4ycKYEiCc6C
KClO5XTAJErSYk10wjwBeF1WYHYOfSzutKUEt/avdvjHWj0wQL4UYPbospQTp1kzdUD+ifWtJ5WQ
Ueq+KRq9Kyj1r0oa/T5TRmkP8t++Hx4AMEQSCY6D4AvHXxVTTqvDcClLUtb0sYfCwyZBUmijHNhx
phNRPVsqATsa1x/YpS4OzB25ufKqFMp34oOh6BWCHM3IeFXg9a4ASaz5WNsWXbcA196M6+ss3wUm
E6C3mwN1Bg/bfNub3e1RiIG30GTRfRYEPGR+foznVOMA7XDcbWOFj28SHSx3wSXflfJepevifdbc
toJReh8e42cIgq23LFcBMEtlHAiDTtCjEZL5cv1dYVPAB/A5qsDjhjoEhJjGxN1/IXhMqB1D20Ta
g2+FAEA9oY7DB5qb+fWPOQdgfNyGwgBSrxq66tme5lqPSf+AQIF3g6g3hBSygaNION3fM4S5nOBp
542r7T6RlUkACVvZYway9sHHqUrnjaTPlTS1gx7OfKXJFojAJE9+DIF2e2TUuYJtmJsyclyQxJrn
P5iNr6aLRVN2lyyaECZZB8D2N8RnysUzK9jtCjarCHlAHhcMS0SiWcikmJwPLksLxzS7qs/keJ4i
7BVoV0Vx1EpzY+T77OlS9Go2ZvLKsTwIQ+4iAj7FDNmFE1Mkf+GbFAe6vmgypH/mDuTCK4kfaWiU
MA8/Q2IOBIq+tEDiNWo5uOvMxBvgW459Hm8F/A9qMwZoG2Hwh44VBqZ5ZSUB23vhSoCg8quLxdZf
idXxjPE+qe9C8FFZaHjXW1UEOBvElHtx3T8Zv7/+WVOVbS8ya/BH3myLrGm/vI61lkUkidOSBr1M
VhWIBfuEkJirt50mm/V/2Hn1PY83adou+eIcfhBqCNKMj7UKX4O8ZAo0C7IG1mfzNl4jpH1Qfcz8
RCKnnH9aOmmGZp6FJDb75q8Leo6EncNPSFceX+Ayz6tJ7zDOYZX2FzrXRzvuGwAL8nDxXtWb6DhU
EOBnOPV0p8jdKIhR7rfliiCprzgwz5/URR51cOPdNmobqWcDEA3WTxh5ikGrkycWhFaJMBHXQO0J
uE4vtJFZlK3UmN3i2ebLsm0/mPKuQOKCn0zQRUV642NvmcpfATeFq/PFYeMf5G/guKKD3HIx3yEl
OqokKsgqKuGe+q3Az7dOpYGgnRORr7nuztgIIRIx2i+L6RhgGxu5Oj/m0rBHLaQNq15KIZKHJkHK
qHgbzc11fgeYi0mg7oDtDP6w0PnUcVoTwR/a7E3C0bjG96YR9AdPigXYNg1/6Aj+geGDb01e9LCS
nG94ejd/GsjpnMAqRoM6EDXu03/r4u+y2F5AE89TiwJ3PAbnbNwqh9hLjFH9SSII3SO/4AOVeskC
XnfXdmAuuNDKrT8wETRpBSsVaqJESv0x1fHUnrOiN4iCPDI7jpDt4XU6pbtqi75FX+XV4t7k3SPV
ZwRGXdhHDe/gg/jLkLzvatWSxuTxeGciDsWcCHadikbAHRQzBJW8JQxTM1CyCzFDBfts9KkwDMpS
+3KoD03l+du6X7Wmxglvjp5jWEybR1PKmStGKE+fyTjpEVGvo9UbEzwRLKGvARbxsQ1i59jHunlz
gGRCYCUve01h7V7QeBKQSDx8hkoo9b2Ghz91MFZgeP9/ZBbgp1p9MbDst0t5/KhrtBS9pI9irw+R
1N0zJCIWQCAdg+pyaO0nBqypttHK5t3DONz4f60of/F7Baa6XVr1GQs4eb+lgXVXS/vaDOa/90U7
3B7fe10aTY7lMxlo2LoW8o9G7d37gfujTHM40QcNcSsISV06qgMP+sodZsqdl6i2M8DiBAqfntoL
DezIKo1ZIAyVIqMtrlnP5Pkoe40f8t9fAbWD+W7It7ZcMWz/4uQDBSxpYNFLaF5E8LmhpRFmV+5q
IWPMN0VSzyiraKrNCQNuwopEvws5Z5/XEKzuVXsVsUpgAqbbFgDyj7whujkiZfksQfEBOoUH+R4P
INTgLZ9LZJv51OPTveYx87gC2F086rrLhuAjEBq6ZBgRSJjPM1eCfCRxa0yvTUvW+J971RDRFkD3
9gzixcm4fKpSQWYijmgO68Z+v0Dz6vxCOw8Nd4sd0ijoa4n0/werRqvofdCgM3qfmy6H4nuhMNoY
O41lCPHwc0w7jG70W1hpylrijs5W6cGBNi6xbx3F447J7bo7URfNBoUlMag3ixtvj/8VSXjQT4bp
tlC0H1MyuHxWK/9T8v8ypiwPk8/UQP+wx0N3VYsGpdW2vBepppmHNtC3mnvtVKVtqQJwFN3lMLbw
oexIUcoV2LM7f8Qg0gniV1JOHdQMRqIqj+pv5vrFl+JEY2QGMD6EnCKpuWTjNwGynsc4Kp7mJuC2
UncW1YoHSn31CCzdtK5/6CPKtY0sMdPqrxGdSDpKgdPvuVdI21AP5T9d+aBVxxoIJY5Sukr0rl78
RyyYjvDtnhF4nUI3rbsXaqWskUOQwWPNzB63rX4eszRhVI4f0tiOSJzdk/VuqbU5FlstKgUqYmve
m0FhefRMXTr5/nw61ozK+4e+PueYrzUSKObr9LXmmOaMSD2rl+bs2lAk75Mq9WKNdO4YCMhxHi4v
EfGoBwgpBDwAohdv7B3D1QXw9uVQyrhWRPEwFPv9tBT9bJemJ0xkTQY2dCXeOQQoEa4NS9abn8m8
mve3GaKh2YxQ7gwN+DYeXKqZ0wxtJoahzVu2dBmIi+279gIZbLnCUJtLufAgguF24EX9Rnkh1+pi
udGrn8l0UIM8nBEwuRLoVa81/2z/Qxg0nsEvCpVHVAwJs2UfrHyZj2+qxzmvp652bEgx8ozzUtw8
MKaBy/sbQbcsJnlYBDGfuqKx5YMuio7akwi/mCbJjv0ag3EG4kK7HJCVL4UNHkltCiU2yV4wEPD0
gBSOTaotVfgPxjxepkL0mfHai07Itn2DKL1PWfzZ2NQeMlXXY8SfLQTdvkbT2ny8kZS8VZN593Xs
3HbwvFkJd+f2YoWOclTL5Oqi4coME4voDuRB46C890gpDf2xFvZpNKCtuueV8jttGXblWhsBtTkV
cheZVnLkOhvzJeSoghtS6GgOKCje4hFJSfY8wigf0+V0bij3x5Wt0fl0XtVvvnp/wM2jaSwyXQeA
+d8U3tPE2ax2142Vfdndpz5Je0XavU8Y0LVmWdjVAB2rs+rmZlghU/FfMb/3B1vKxcwfNbC3JjEt
NI/Pm9KJ85pHsBcYubueW9jPTu9Z2DTZWj1EIb8OleNtUL7FnUE57H9YHET/NJ+qlIi8uS+jWWYs
CknHHJNS4zm5x1NjrhdiC1GAnKwOmcuN1OISepYMwPVhxgrfH37D4P+em0rsvqXeQmPEjRMCOKj8
isCdwKeB2SqUVGSSykwnU4IOStUjLkZISSYWIZTi7H0mSQjtJmki5aNBpFdqu/EuDDooXGWjQvav
gXlwPvHcHJrE1gVUKK6isX8KuDGtiNKps9E9qTH6Uriyrkp9a0VJdkNDLa+dKVYYFvA2XcUir+wz
PxpCVqKT4wNVJ8UOrscFyz7O0WTrtBjydlvNv6EBxRD9YrHXOiYN1FtseSjACKguMZfrh/hasj3x
A/7yZBX4RJ4MEf6Bo/LokbkP4gVLXy+mQU2ftryMimJP/TTZqBOZfVGJwYI+2LXn3ber8F+iX1l+
9a3HcXHc3F1OFMSml1O5NdJtORxrtQkGcwwN5MA0kaw7qSeso5Bm652nwoZ26XDHKkYE/AXTnhDX
908lEWibZiVxxt3kaOjZPBVHVMHDrXc2mkHNue1LEfOpUswj5PJgAso4N6FTNv2scg/axFpyhtGK
+pfnM3av7ttopbSreqfnnSEAPp8eE6SBf7UEYDSTAvz+zwUqUuRemXUE2vUT1ei/kikhYjpJwEma
4I0qoUXkkD3RqCnoakb1Uyupfq5kD+v4RbTYbx5N0ewKkmG5MVj2F5bshNxVW6VsIVlnGdkngUeS
muBdu6tqc552n5aMcUbuK0BoH5CdxMf5DmBIzalwTAXBGFS3+jHHDZcJYAyJUbW/DNZnknuZixYV
T7GDXdAVyOrz7YFWxKat7kdQaL3QPHpFUmuUvs/1AC8pRq3RqeqO3csoIX93Bnr8wZLqzKI3ojrj
IEhrMCjEXLjd0sJfEzxISToEQG/l1+5HaCTGInjA6Bz7DeHMEWmYPRHuff6Qwt8S/wKlgQ6vnNTt
jQMZEdmbRMh2w+PE/t2n4yLEvy8/Glj5/eAajfW3jNxkQsIQF+jjd9nDVmSyux04hr/FeYFnB6uv
b7JQYMz9IMSI7Cml/oNThwKRz5gGj/GJczxkKwQaEgsTOAe+lE2pA2B00sxlXEav3ydJnf/zn02m
2xDjF5r5Vdb7hf+miG0m4VV2TMg92DA96fpOAmk1mgf65mjJdy2ji2oB6NZHeHZorX+4ASi2xRrk
vLDtbAt0GZcM2gaCofB2RXAsSEdOcI7eu4y+/5nT560UYSyCBe94djZHE8f+z0VjU8g/hPB7e/P3
lmhmZ5fHld5QfaICNU4zd5cothK65q63iKqfvbIzPvV9EeaV6RWqGSRc+PP+96tfzp2H59MR22cG
47u2dUjSoqZqua9nZbaAHjQpq8PJkMr0mbMvzQ3sTUD1XlgKhWATS1F4UqF3kKhW22gTayAImNpS
vsb9Nnhj5GPlqdRKRb8QDAn9aM1kr+D3FGHaQ0rm+MWZyvbcSYcSgatY4gbtuMiST0PCDtYkikUh
DE9gBziFoPAT/2D0lYQ9RDYzMSqJSLemZyZvwgATvcvEhLqOgDA7qwEyQ9QTDE7MPZLp8HaBjixs
FkDPLoG6DKo7btuDJYT9kUSJ9xancfIm15FHw8ywVox4kPGQOZRFBDLwQW/ZbMhDZ95IE0evRP44
TgLA4xO3plrhICiP6fP/G9KBoNDrUtAjUyNUiAIFh9SvYU1YoY/LpbXSS7GnP+CD1DfuaCYeTqOT
mNf9jmAZ6NYwDa38x6NGTie6xD28B0+ar16jkf9cy0eLi7sMgyynn3ubK4HmOtv6aTYz92pgdOrq
LkxR6AKav+uGflG5TJzrRmpVVqnZdKGoHlncTOn4bUkEVycgnOuFxJJYQg9zL31zzR0QzrGGLUs4
lkq9paIEX4noZDoDX0aupeGr7f9kkw906PwggolkjVTEm6+Ec98WItv3ZHU9PmngPKRhhhj6Z6ik
iJDGLUikHLF/ZLbArO3xBCFDifm8r13OIk7jvW52LnL/BuumHyXQLZULrHSV1QQ6x5pZe14p3QJM
F72GFhRm8z9BFI0gAz+rzXJ9lE43//l1/jvsvnLdjpYlBNLPmIqKjZvArmexterS3GXhlCfc+nIJ
JW8DFHiMZIeLJnpnhNmdpO0tSoX8Y7hlQrv6qqjhz3VjTcAUYNRJWImnCkXy1AZvIi6hT2KieB/+
obCtJ5vpHYx2NZDpLBYC/j6ewuQIlMEfLqMf9jPFrsbjpH2ujRwLLPRSOY8OV+B/58B5GTY0/Spt
FuYx+ORe4Sz5+LPDPWjr2EZrbAcaR4GSlxG2hBtSlel0B9sUIp92UimJMNsPnlaHTMBiNzoJ/tb7
yE/eUE2vbHFE6rY9BD+G2XGOmIo1f8Gcdw7EwuoycdO4+YtK8vFa7JCi22fE/oeutmBPiZOSm/sg
m8YD/4DbI0T/zVyhTQCHvUj9wZoRvDXGdmDdIo9GIkxG1X3IxEWiHQnqSZiZQNZ2PBIf12STiMTA
RslMbh6XfpNbUNAHMt6+TLmZJvJvxuhUEk9sN7YORjLRGWpoqMEVBc36kVuV98N2Ugmt75X30aXa
KC4N45ysj2HBNuB+Ju/zM4pdAmgylPoUQaznFEJZu3fqH4O7VCDhWDlIvxKNJ90vdslvr+cchS9u
Ho0VhXEDVrWkmk/wi5VYm9OlJcqYWSSe9ZRLyNUrjIekSNb3YN7tqr92/NWVMGXXCobvM0btcsJV
jc7xy2E4dyKKe2vy3eFjfbQG2GVLN2kPTR6Y0WrxBcETLzBtxOXuz/GvdxLhGXR41eftVJgLKJqY
n6peJsW8q5yNj+ObqgQKNGB4kmKIeUh8fqQfBW0qBuXbtwwb3OYpr5vyY/QrWJYEs9EN9YDUSEt2
S56dJCHM/c+/Fvv59LNU8KsNWVwQbNL1zfE8CCinnGr9pTUnrVAvjaMpgz+JykX0UfY+a3HXHkIF
vQQGqewcMF002FLEx79SPfft8F1icoG9KEqYbO9oqiURMu+aaE1hQm3MO/oKX5ScvIq1sTXfP18c
2req1sQJzKQ2OY6tUY1ZQup2uA853LF01kIpBw88PIKdS+vCKHwdN5MkY8zQQbdaYpvxLDPGptq1
4+JiYuugTkZfXIAuv0SxCqpa75IS2P60j9S2b/4rQxt2AdiCWWgZoPNU2pSBKvsjHbLonV/vbo+9
VEDIBxDt6CGdC80DOXKt63AiBQg3obfC5rYuVQmV3WV1jiZHHFzBi9DfjSzkCmb5u6hok3Ccc9gm
19URe1L3IvUUVEMyWJnYpzOUXQs+sKJ7iJKSEKOuQ5OFBcowvurGfOhzH8IqSTuxL1+aAVAsHjlg
rYmLpH2uh0KEEJ+kjrKnSRvLrMyVdjCfpzlUjv7RZAVrPeLv2Q9gnf4NmQW7sWsLxmi/UIuoLDLk
BxgYW4DEwmfvXS5z4W3RjxkVBGXggRk7mvxwVddLCC7wP4upkigFO+U+1vW2K/q3H4s7o/OryvVE
zc2fgcfBapZho/FvOTxHinSLulTnYilbZb/MWnRLDT2hAqoyHijYEXkTahyHTqZxnZt8yXpLbDQT
3ugwnPHxu2Igt9rCuZRrc/ac92us2mhWQWkc+8+uaszUydvkGhGONhqBdttPu2Rqn+SZfiHpuieK
v+sDozzs2ceeMZd/NEs6QEzpn+o7x+1jdNUO6WpYJtc7gCfLGVyKY5ndUOPb7vs0q0+x2gsQJlwx
AnEvZxf3Kp5QyzNDPMUZJ75rAdqhPZ+YcPkTElZJ96hc5vu5GLA7IOytadYCMTbY45V4+tBS6P84
vWUNwsEodoKjGrUQtl2a/k77MNaRzLE+3ImAJNydOYYoP+LxIWjG3Hd6RiXi10gsIHkDTgRDTYjo
Q6tpWk4QxORX9CIWopIZRCItWtwOh9PRDkLBjCvgMnOj4opbTTAP6afZiF2edtFiF0SQdFH+3LjZ
SF7OSR5bh9YMjrk6WehdRfYFYCFeSi0mi/5ZnbWYsjBGM8q9q1lX6UjFRC9PGlfgUZIyF9StF7pP
QxxVCdgJFEcOyBthRwr3IybranBCLWynblroH2r76ar9GBbbhtnkast5R/nbrGxb1kgivVei7IZC
fEdgiLtCUGXKz9ah955NITE4yhGF6CkyLH13mMucqzXKVy7N24RyoeIJJN+PCTiCNFpXaHYTrC+I
ELZrbcMWk2VFq9EwbGNVu0yZxegS0w0wEJftmCBpUV5KzIOVzAhwWzYlBeEe8DtfV0uhHkJzc8di
cU9LCkTj2foJ23oiHv+seMfxVmd0d3veGOQX8avtCymZajAj/kGHQB+uZzxr9u/+lPL2KGxK7U4K
G8aJXnx0xdl98j8axmtvyxrmsK1txikJmN9tmPyhwOjRdvD1sq0dywwqh5Ooa6ICCPUI7cztaEdl
GNI23K7bI65QzrIdPk5wtQyM+VJLP/S1M5Zox72Ng+epTpdt2moxCsybWr8JnRNwQXE4YuaIXAUy
/Azhk7TkiLwSdMdTvgtj2GfW/ZUbuLG01GsYqFTRoN84IPlk61sTiPVULg6fgu4dEaE12IsiQIPv
bY1tKc4aoi+5GPJt+QaOXd1huJuViHqWJVUEx2NkQrz0k6q0syuhAkFX7D1vF8rELE6TNp+M8d9v
opLY0fxxD07TmVcixK56jjpfDp5XIViGbJIe14pbCr9e2dq/y7pNR155GessjUzG/l4gm7IuvUBN
sqgYmfXTrlSsU4sdAOR8bAzECNvXcUpFVkKYES7gdpjqdQshzJp7jRCjSrXlVyM8h3mR9noiTSzN
JZBGxe3EpvQvqGhLuK0f9+NM86UqQqBg3UEPw1E6LnHYknBZv0QjJL3vkITUltHagkm8n1odH4/j
LJQNx88HCAyLkFOEi3/pkZBxue2pfse/OzKsJFuFNrGzFNeVojdnuk6G4+WW9B6RIY0jzUe7imVW
FNV2BUxb+QUgQK5o6qB3urx+Fyd0s6lN+TaiEwH/VC3LjbajfcG+peo3mprjT3Lhp0IfTNSmXPjK
BmIg9SAxuSMwnWco0dGvAxvz8XzL3xLSczLTzVktdZn+MLkc9+b8wEn4jy78YflSkFVlj4jx/8sI
bc5y9Ybw0ULzMruUf5IBcYLDP/Q9Cls1X2ePZyT6GfYWsggxjHso5kB6oGhr4F6R/mE3txSauiMq
JSylh521cl5saYnAqP4LvBe6tU1m/ciZHq94/bWq5L0gjX5t/HARsID3GxRQrovU2TdqSCynSM0l
jwXKTvhiOQbFv4J8PX7hsATkfEhYtq0spELyJT5Q1exLVmNrNtn2DcLUXz9HbiwSw0EAJY9EV++H
LOBTz2BhlEQFzaBFJHXUpnGMeLglHhOQtKUjZemFk/yNVsxQUS1MGBW9/CFG5KA7EOyAFRIkTUM4
+I7XJbj+1ffBeNvXZrEcdKTw126uJjx7i1qFSk1P/c0ORarZtxcbmpdxl7KsX1lcJgIiok8GbGFx
kCzVg23KuwrjOyH1TDV03NWMy0aUK4TfBQy5mYmHcqDyr18blAmfp36v74N9I4OByPBgB6wWTEXR
jxNwhQo47Ii8BoSs6cXXhCKZGpkBIo2D9/mkvkNmGaJTR6gJDIe/pdpIMp/phZMCo11p2YcXT4s3
A9XCSDBgaT47ZjgDAKIpqo2j6QyHOWsxQYMaNSEXzOjj5gKkfv2FhwtNIX19KTtjuJx8mzHCqN32
sT3iss4kg0KhE4ftnXu+L8YLlmHTtdN7YJv4ijWxRie6WCoCWv2bUzk4SCxKPkyrySw0CSBqBktT
/Oy2aHb1PL2vWC6eh9S6YNzKEBq9AgBGM4mAJpDNrNGFvs4DyvFfM/MV6X5SwFkzyC/u9byP/REC
w+dgN8uTPMwtkjCEysgp6C9668mjmuVOfQ48EaAfdncgFtCeLEhvhRkqEhfxZNtr+Pib4eGA2wUt
s3mfofa5dlvyjnxNf4UlwQ+MvAQWUrW9F5EjPCOzQf/JHobhaZRhvYWMvAXve+Je3/7nmRmGZEbU
ohM2o7bSnGIzMtTuFm6Y7WKuIZpIFXY5t9sLsMrflGFEKo/p5gTcSw57es/I2cp2gTHfAT1qQs4v
tAf+im8xL5Hdy4ulzPWeqezTMGAHjjiEd2XuitXrc0vod0h+pkDjiYmLzHbrhYVoqk6TE7FsQQaM
wTiL/7m/wI5P1CuQGbr4C8J5ZHIh7ATOkhmS37onIBexFlwGYKf54KKuMAhMZF0MR/DAL1bcBAC7
QuZ24kq8Jp42G5xslmRY8zZIWloq/IU8fzJYYJeGMy6XSaePik107X1J5JXUY+obUflecce/tgpf
sESKbsG8v1etL6uLXCF65qdqAq6A5ke0WScxSzHn7IZQlQlZGb8zgD6dwaAIoN1oy8jJh2HhHBGN
TdoK7o5MxSoBWhuAzMUIyxcP0qPRVZAgBknkX+7ovd1pdVE3lZhD5KX40Wfl6jQV7XAnu4US3bO7
RnA44SxSwapaoomQ1DxyOw0lZ8koXvBrdGktPwnlXTlkEqFxualjSyg3QiTI0xQWwS2zQe1uP6cM
QF3VkVo3eRWFtGixivz26iQ7s3z4ZMApKarw5P7vGD2yVT5SkOdRUNnosdN7w2tpCmm7lsXU2Yjs
FJXrCEeBso/5b+5VWcBA3OajocsO8gR4XJBth9ndfil/SN2Qnnchm7Gy7WFgQiA9PbujDc+b1aSa
gFWOUoxF6csZecqbn7ilKittFeG5NqEj8tjeSqZ/hajfUW7nKvjaJlZqHwSxiuz7ZgmnWff2PK9+
dcXk9c2N5sV/5Bams0EVQiyRhZwXVQIW0sR+LzntJTsO55MATEq/LsXvmE31m/yNRXZKLHmTntQX
Xq2uybK/nrDe9JuKWJoUQUofZbtWJbBJ/5HmCd48IPGfqQATD8qejMOr5LKQ7hVEIi21uAqLV0qy
cVun7ckFoczNO/TmdOuRzMN/ncFQiuvJhcpWbySP64dwtxWqyRyTYJbt6Q4Obv1UyPAi8Inxms0A
wPOeWg7VnhPe5CQKjfU+OaKndvWSYusMLrbR+F3ogqudyjOd9PED9MdIsdKM1cWkTAVqA3MTzBpY
1bJiXkzZMVBHgVFUu3fxJhyJDpwZ9Rw9dCU8FKSbOTixE+wbD4FLTrIlf4uGNX+Zxws//9nRJW+O
t0YVQI4DI9GgZulHmuS8kY7ueMvKLK04BUIPYNVpMuhGKHrNiulCf48roNclKqfaCGJUDGTSG8WO
7dNlLi4Kc0vhJnsHJWMNG+P4Z3JFILR3Hgj88xSWW4lMBqHFzEA4Cl9CDt2uaD5vwwIu5rg78Yrc
ZjeRphTRBAa3cRngTCVyUF6LkGtmemxNwqS605h4q4qa45JuKngp9NiwkAFw4hlt5vj8GZSfGzer
FwGuxnc2wZxw73YEiijMYdWjQFAhriQFtSEkxxnFQFi+u8CkPzZsG1mbGEin7Hk6bh50WyF0ms74
H5qNUfGveevw5NqhCtftlqtLqCu9JvdPM8gwbX9C4Cw0m6e5N5vvFdJ/aTwQ7/Y6nOddUNa/Bbnw
oZQ9w9j181RTswGKE1JpWcskkKSZ4CtYoUc5Sp5S/BQLg3wLV2vrxkxh4pG5998+Rcnn3a6FboU9
bvZloGAy9cmzDQiM2e82S3OMDZwYnGrndeiQJf6yMy/nHQBj8QU/olsJMYSiGhmfpSNkrm2bCAsq
LX6GsjS3CHPkO8aD3nFSoDHgB33PzTfhlSuCPYOp4Ht3+BvtygQrD/OOIXWUIFtu+CXU2xZO8okY
r3VB/k4O+5hauvEPj3JpBnsjhT9ofc/phX/RamLuUVfXLbyRfXUOsD9AVUX6KXTvO6I82bim2htq
4zcMioqj+2ZOc5kttIREak0XcCgkpexdViorRkwQJHewbYPAcB1p2nwAO+/9U46K9JISgTy632+k
Ct6hlozNRoV/LgetrsOkX2i0ivSGxPMBsfCEllI2Vcu85u9g04dbKn7BQzg0NKHM6kns1ROVazl1
kwJhLKvnXkmihlqKqWkQOx2bJLXtAMcXFeQ4e9gTpd44Hkpuoj3L57cpvFCj4wfT7UL8vqux/m7+
C9x6dg4+wmBlP8bF4DWnC1cCqNIbMLb6Xoxi+/Wa7zhQS0IUfGKjGaaKzFZ4ltdU4VZOWnvFJuUg
+DT+nWRjdgWQBkJ6YPAc60V+glZW8l2Y1CEiscmFFt+Lhy7giM2bih4kPkYaPXKnGtw2n1jBCGlW
ZXmi+dsXl2nD2EM1jMuuTSgNjf6U5kKLV4/JgU1Hhoo+i/0roINHUqaTMvFneEyai1+0DjanmLSU
gZ1mSK6I/UigROZbSZrXrGMfDeoRcHfERXvJK/e1kwIyDbl0tN5eKj69+lfVpj2osrPmB3OgVJtp
kiuAOo/QbCELuALDOaJe2PCDjy2KKW83yWBeHz82Uqp1A+qVnFGoD83XES4L50m1gRTw9A6PQpIz
NSHEeiA0s9Y4/51oA5XBYgh0XjgLMzNp4N9/9o1PEV9RPTVJCxi5VSRlvsvVJnRJlkS8IdJF3sl6
oXNfftNXI1Xt40BHqEKhylYsI2ByZSbSIOT8/q5i8rRRk8QpDfFVS3ZWU6BxN5HSbkzJ4eCUySD5
hOts7y+GnQ92ctR088WdynWGEbMTJltOvktEn1DGf1XhV1HiPWbLKwjzwXtFNGJKSpdPy5mBvS/I
yAB4NGCUuILhUvxM9GjmEbLSgr0Mq8M/c3EBkTG0zXhpnMOmh0vuq6gBk5+M8/xjqan7lgmJHlQt
MBUT/6rfy7kCD9zkE/eZ8OU9+7+zVLXUByTEd4Ao+eO5DfknWtGM5UjB0ySly9j3SZeuiowamMvi
7dloODj6vaUHgFxYG+KdTDOBdJJhcYsbbAgqLxj/7iFqlcG3wcdW0SEyOyBJrj4PVeGZyq9zC3iG
eI7qfkclw9HlHBEHLwHSYYFcMbXKEiq4Y50ZhBOWy6j8NmZvetdT6rBumlipzf1oC53YXMo9+ROI
GoWAHkRwDF8ALhH+iQszw4KvPYDyaPcIBGgVmnSbC0S63DIetz6AXVKheIy48FI55lCUStVn8ZSU
SeLNIvwEBu+n94/n1WDbXdkJ6TPfWsn0eLQi+xBQea1lbgiRp2zNERt4lH1r/tYtkDx2nqulKb9S
C0D6qsTQJsMhEtIexuGz8b2wfQd3kauE1vyzGxaR2hSyaXu0BlWn5N3rOClFQNM1jbNDWTZLtez1
u6r3A0DUORAd8BHBW5eWT9MfSIpLIU+YFtsQ0BacdGTpa7EqeO/dTOPu6xlguGma4jd9tfrv4SJw
cgkgFGzgbEuWAaUa30KYZKXD8f0qapU45rK6zZYxTXfP5n8AQ2tWw9KN/jGB0OlHPcOnnuTqZ9sH
SGF/x87arShheWrB/rf7pAlkpgFUaYgbPKwk23iMSlopXIoMqUGtyk0+fDzL/2xAdnoNPMbfVHDr
SuvLvwoqBT8NRUjHcfrFAljvgte2fx8bZmXUGS/dVco6ZEmvmWEr0ej8J15pAdkzE6tfQdmVoR7r
z4Vsuw/PZ8M5r87wrKhiC1ySuGqEm5ACQXxo98s0qjy5ET5rRfeoR8SHlCw9PrgvZVon4Q39n7Mn
kigULbgMLjrZH56oAQDvCAeoiXUa8ZVfccBdR0SbYhH1xNRNwlPK45fXmirzmaK+lB91OrNG+yVR
S6JkdI9LzMx/EHj7O5Y0UPb5RV/CKsurzo1xXj8lZfDCkL+YDVHId5nm+PomnQwM5x3bVplCx+ls
7GkXGNdDCT0abJ0OdxUadzecw67KRplTu2WmAd/8eqnrn0NEgOdSJ3GYUewt+ZFfWj2AMTgvDxCx
vANhI+UdP5ZLbo1uV1yGH/ubTlUI9PliiQCFdEEvfGhAW25Kf/QQoeNPG0HnJczrogbUxJGPcyL0
txWd+tap3Jcw4vWCava2xyRbEAIVgPZkLy+ToTEcf/23B/J0JTsRzGTSNibAyOSn3ZLIO/iy4Tl0
/OCfP7UDuZvqfszX0CYMypiEMyY2V+L80q99n4HFqfNRBWn31szvM340gEjgTeIQNK9UtTeFtcKE
tRcMTu5nwKn55s5iXOaTXJ/F6dEurcTfe2y/AODkIyzecc9zbzaprpAfqfj3PZvvQABg30GiC8SK
2Mii470+qY8rCKJNm5Xuct8GYVR7z1walDFbE0k5F3RTSb5s4VV4IbW8HWgpc8TkJvzNSMhRQ4SX
cS6zSdP9SfQlCfkoO//a8R3Pk1zA36MaF/M/EbVZL5FA+j1YDEuS+0jo9UNRDRQZV+S0zj8Dge1u
+6UmxJ20C/nHPaAXXUFSAC+Y4ldyuN2rDk86Sc1/ubAUuck1mEWF0Rpqpu6MFjPI6vpTqJA88PEQ
VSr0ahnt0bIVxQgNQELF2KkaztfLCAWiwBSgKYjG5qh017RdJsG9xHZ+YNQXS2NFMdRWNr7tboV6
FOOq7ymnP4GqNrLC0nqbnLbRRhPtjKYATspZK1uA+7ystC0k/79RbjTJj866BaXMrobOD7nYtJAm
2FQA3OBT1MAG5rqrR2fjT+alRcikldkWpioEOXumgjkmLesZD0vpIAcjhhEE3XygeAD79j146TA/
NGlM7ptmTjSNa48zBbRsvRj7P8j9yqMdya+qH0OuL+3M2+gAjn5gyav92NmEFcT//QLgNKiitNF6
YB6048Phkse9S6YsoQ7syXft6WpYQpWoQwulwO8InyXEzA90Ws5eCMR2gNXQhHrwC/8NsQp1+R0b
f8+F8DWAi8pMwL1Or6rmpHPCTRLT8TKf3M3nUaYyyU10DNEKdyqV4w10H9IUxQZJMyd8NQL3mAn9
mkGrVIbb8SjhdSoFzBCqox10/uU2O/NuaejMj2O4zEckOSH2TndciiEg0W2gLhKo8tL+bNeOa7cN
0hGwMhx/owJXqiW1iUMcXD4x+NLbfiHLkXpyDup6tWYCN1Et3X2fFYFaE+3EquH4U7oCRmxiZM2R
XRe8mIvykxegeu1slK2plWOCm47GAU9Hc93zu1+7f9yMtDOXPaItnyIlGS8omRsNoh5WwRInOaY5
T25QnCpotSNILZzyNX06kkvT2I2dh9B025HoKm/LYfeDdRBA1Tt4u1jtt8RmdvYsgFn5cS5bxpah
NZqG1gfhlkJeEPR34lxZT/omahwogGx8LdqiwotEKCTd+ECZ3fmQ0pPvxtyMukgdQi1Tx5kVfUx1
2BYzPp99It07mj+qQXYI0ie8OItzNqhA0YbG8e0v949TVzyVrnTOvDHVJTEzG8wVeMdudXwzb8Ii
/3sHjjzXNzoM+Xpf20xLwnEa/TVeq83Ig+Tl1fcr2V/+5wW45WREKmOt2d18InzXceedKVt0YzZu
mmI4Tqu2mN8c5mSQklHRhyvMA5aNldusbc672jZfrkRQd64NDV9hk27S2bTAd1ZdTsaqYl/8CZ2W
a6o4w+EcdeABlua8HdDaPZqLXObU27FvJthoKAtIrbjuZB07K/wJVKWUE3P+6N9SvNauFu5wHnU6
ocPb60FccVTefeYf4vhPxa6e+VUiEdX67pzEVrpJ8M/PtGp7BbQ4gIT9ddHuvlfTSXphpEZJYsqW
KhXxL+E3wjoUV0orcTEg7yC5xsyzkeOd6ynOCi6D5luQiuBLdQLe5yqkAGfMMv9VqaVlOkmI9pRd
XnIr99VMLIzr9CFoU5I/Qd6uLUt1J/gHwJnFRkwiVLVX5Jj/tkgZhSpbDlHm4B0mTa36SKhXCMAa
4HoWYi8bQgF1U0S6/PyeA84jz3jCe6uj1IbhDV1B0AzkQfFsFYFQSNIn3ObUumyxqyn1xPKzV6Yt
hOaABJxTqg2vh1x8wRT5ElZwa6j3N9bWjP4rZq7s14xP4VZUk0MJ3c64z9P50PewENrDs+8VFmxr
NE8SY1Ab305gOvv6eRP0nF7sFei32Jjw7GqGGkAv0QtZe5oTq7PylwHkheuO+gFPDYK/3p7qTLD+
a6CC0ljDUor1E6AeGjoEZGEtjv2rpph+Xjhmogrl2hsnOQx+0L2jb4hu+3Trg/QezrMS3fpORh2i
fW/Ui4GEknOdwkFQIHVwXsHSYoEAKdXeSBAH16vabg5L2sgaDJV5xRFWilHqy8zry5bbv1Oor/CM
1LM7hsEB3Bx9ODd4hopaExyPWbyxxQS8qZoVk3wtHQHXgeee9e4Zf59zeUYyUf2ep+ehU9iHuNZl
oosUpO65re9YSgMIv9RC+0V79UQK8JgFXcEXyQ9snDjN/FTmijdG9ZiBQ7WrEcvITSwWcA8TtjVk
3qniqC0ZgeuVdcxUBkLuvJalwi8UtU+LkCqny39W+m1icO7/81kgF78NpM4vd0A1I9mDN/rUU5ou
22WbHSCaD8sX8em/Cl2lClMNkVNS1wwgco0zTK9FWW0ena50d4dPLLV2kv0qVlA8WEC3oIBO5b/u
KG9tpIQ8GdCyC+lZFsxwvhte+ZwejPqQy9xxw0R3uLi0pVw4F7nAQddxIZP9zbdeILKKKcbZN0l+
QxMSewLWgDOAvAnTo7mkGH1CKVJUihObk012mJiJAU7eFA2XyZUFDaSmP6vNRbkHT+8cDvV4vlos
HXAmBDcFWPlSMHHiCESZM1sswW0V0+mUdd8MJ+PlC3hlfKzDU/UZ89IjGlMBIBilI/nsleQkY2Gc
EWfU/p9ywjhKCPt+hsPW4VWdcthg1HSdgf952gIVyUYPvTGMKz6zl+BfXsKcse4Zh7VDbZ0IXipT
CD8Kee84q8lK3Yfejhnm0sKqyR2/yYmr2a9X+oBZ+hcIpbqlTKY9x1SSSKiEO8SR8keV/VglE16r
9PNbAw6vTDecPsnQ0v+2y9mQR0SvVNK7BbXZ8deiHh5jyy1BWuWFS+bWe6Ef1qVjCb6Nj6ID8Cuv
kyyIo0+GrCQ58XJn4UVK9g3hDmx7wSfdL3lcV98VeLU2UoA/llt4g5qM7f+su90cEZWbtI5yGu9s
ISKSQf68da0e2j6EM7PCwxQ/ZvyY47ImU5zJhjLz7k8dFWcDHXGryXNeNFqAbdopKBdhB0pQEvJv
nywpvVOIHsOrUIzeBFwkWpWhR1iHVinYMSMo9d2QVLMHaczOhuyF0/A35Oe5//rN0+eUFQvYLQp+
1bQ/KRb3O6vGbXxF1uupal0D7bY0eZ1ps7FCQYNRFQPdYRUdXjUdlfHMN5zag/kwyMlJABbgtH/N
elTeBvvcbI+lQQg0IYLVvWdH1k8+P9ZjEmvcsj6FOM+EBUJR2xNzDiScS1ZHeEmeRfozJJ5A3loq
H6bfvTk9cxQ7jQQhZOP3UdjNE6ZLgk/pOc3TKUG2LYL0NABdN8JWWUdYJCroPslAYxilLJyZb1BX
sqTR0lTIhnYshYbchMWSPdHmJNNCY4b0eLYUAXjBPmfLykihqK9uf+TjctAXAc8c8fE5TkDrs+ZF
8Ki4NF8rNte5uLjFanVmfmHHiLBknR3wROpAaIqNCKzaC0peeU6oJe5yzt+2g+EWZakruiBQ9QbN
ABkk+sBYzCF1weQkOv8YyxOAhMnY5u7VMQByCyaCCcfJywhIhvCOue8rIRgQqO3u2I3YOIwhbLSn
89kyeNSWXnEsVIWfydhocmDApCjNHPADHTwgVQ1ga366MX11uuT2g61gNVolvUkgg/dINZ+JFGik
fkbkPpjYSdIfmuBBEjLIqRki9lj7MsPib8Y0geRQtdZQCacKJdQNw2sRLbfgsALgqcGSz7oVQBbq
Pl5WLjK/UAZR/Rfucxwi4/TL+8c+Qpcs6VbG2SgxjM0mAzwH/INj/l2KwJCBVmjcdOJvbmKYCmjN
nMSscXSS1PmHaQJ6Q2qO+rswGHK4T0FtTV9lITdv1vajImj78vYbofc/K//kVdlM2rRrpPK1r9lk
ut/LWI5BAme8bfZPBZiNqhaDXgUCoOAEt7WRdyCTvKdTMzr/NRKu+gOkZlFBW9JfouHaohB5uSRO
8t0BNJxpVPurAc4Lf1ok/Qk8pF7NMOJvFn6QZ86i2bVYKHojKp+FaeikjbVKqiCsT85Uzolj+YRI
1ekGqvfvAsgCFQRofnlivxMvltiz6OCWp8/sUA29vEN2Pat4cjRjPXXnUutSvXRWEtgKLZZYGoFh
+UUDc4QeH5ZrdpxjGVds8wAmw2LXOjhGUYMqJG5Xh9Mw+WsSe3078a7D2TjZT/5erI/CdAPU2PCr
eFY4i3oxlnVMp+pXvUNb03oToOzrJwNTGq3Nkf3k1mzadTj7BKG2rTU/0HNpKvr5u/o2zREIGiRw
fiIFDNTffdStgKK30h9owG7YyqMb1uqfLWcfRHlTRhL+rsTESknTNR35AQIj0EOlahP+1Bj2x6tu
31z4Dsyk8noNlj50Dc7h/U/fR9Yjn8zm7Y3dPYf2ieS3G80Xl5D+irBFZMsCeNVcz3msNBsKHArn
YCge7NqKKztE51TwXK7mC59dbqsHVxS7Us6K/jjONx5j2ySy3h/FjTr0UDMz5rG3f7u44MO9mS1b
KIJHjnsdRhcdBgVtp7qcOuNtCDptDyRfDtrJX7kPoWoc9k92FJG85Tdb4WE3ZbsZiRrdMXQ5Rojl
US6QZx0fSsSx3IS7do3faV8WUY0sIHaP9zyg8sTWoQSR42bJbazDUBgPU51MmiUwK2BMX6BEwPCG
TYbCb8AA4mfsGEkE1l6oEKqZMd1SRpFCpx+2F7GFV2yI6bArYYZmpChAijSljuAudb904csNAOFd
qYcBCVaV298wjSIx0u5eCoSQDuA81LcO+mTQxDRXpdUcImUrq0yULcGdkisojZ/lIQWis5cXSxIw
2jY2R8yKaTiSNcOuaKg1r/YWmvoXKalhfYeB4OAAepLWRZcGkRiCXLLYhhKp3aGNHahh+klbdQ8r
/jt3WKqPOri5H3o8SrphB6ETJxIHi33K9lK7wfdkB+pw5yX89FOgT9vRpCstoqjPxgSMxdHmEPTA
Pgg2tRjeWJCLOreY9e4vS13HLnqYvBLP6phRyqCql+JgtxvO9Wzz6lDoJDWbji8VVM7ycrWu9PB+
jJ+4bEFFTrr7+fY4dumbdze+qAkAo7kzC3zJ411HnE/1dbO3vUWaGR7fupzoR9cBEWkT2er0wOdt
5D5RxkviTRb+rv2E57MWxS7LFFwPIvA7NuB6DXJUKSRg9RjqKim33Y7bmehRsvazlSb0tRqwUOVr
T+ypSvk6Dj5u6oXfjiLGUf2Sju5ES4Py5qmQz+GDNqHju4ctqhD1NkaE2mEl9IFjwNJ1AS5t2FUq
JFGM2og8ZoyeS23gkgkEbLL8gA1USrxq1qnkRsX8IU82Ibv/oiqNwm4D1iAuihNmZDd7fwoRuZgG
GnMcllZrOx1/7SphdPfb6R/+1uLHPqlcvgUCmPLf77S6g5P68ivOkp6qSFpYiPo2KUscKIr/Kwpo
09QipbjtZUPiu02NH2zjbm4+cQICsUE8hRuMXxs1lyJqvAxIaW1jPE3thILilBfsLqTuYeP9J5vx
pH7A+DC7yLWpL1NbqW10AWg2bR1PvKTFwmjynsAqghum3NGJhXre4Le2P80C4io5wN2AZtqpIAjE
SwlGZ49q/IPqNjQx5zO6dBz2cwHKV9wg72ps5UaAbQWfXD4GGdoJJZCJ1qOOYE86zttRvSk/yF4u
5zQczbjWYODdBczhMs9MJ1w3JmtUenil4MKtCWiEy8zeQm363FY6CFUqnfA84nD2OaXpYuyTXZKr
f7O30ZqtW0iV1CneSrXTCBY/kUHE9oJDl7etuGLffXejX8hdjy9xeZ3e3xgqIKnCq/rHCPM1mHpy
xBA69bxq+XLg6N0KcRIBcH9YF/B7tPtUKC02Swd6e8zJnPJbuUEGyZEgElqqg0ZnXLQW0Fb3HBAu
hyU1ZQBwBSaHMvQiNyIvmLE3mwRGFu4Cm4Wl1jmID+mcIKcmVLVSGNRYE42oIkDuOZXXUuNas/QT
WrBee1NT00CnlpVvykQ1YXy8qca87asuZ4RRHVWICZXv8SDO+AaPJmIXsv3wMLrsnJwGgnPSXiEo
KVK9pXrvIE2pexGLvHrPOXYBgteQkj0CbJqS0C/Md5ke4KZdZD178x9fbkdUcWl3s58nrCqs9qtb
N1vEiAAuTooVnFd1H4KPnadrKgMHQ6dvBJYvWho6d6yhr7LdwgFKLOvpGp/XvKgs7hqZ1x8JEOWk
DQzi/71KmqdO6/idAyjEsx3qOUE+01rkbdIus6+CJdXjEPGPquWedd1sl3bHNe/vjbZL8bnsfvR1
vRtkn1TelUk6s6b8ZW5KhIOS3HFbvd5QtVa4UI14VYz43nsDOTyJfZ2hvmF/MWAE/Hl4VXFbkmdb
QbHFLeyL7/BXP1HiWsTb9OJmCZUldohZspnC8Kga3UtrTfUiQ2ZFi0ulCLO7yfmVwJD8gvhijObx
qJiKBu8OPYprV2yVipE1YL7WNV3ETh/hNWDVioaFlWUOp4loGiDf/vDkCESQwrUF9sQYJko0u7t6
Z+HF/Y2C0zBqVLsIjp+UbBlqZWRUtfkMVYJ2V48pedKprgNC/mzSgwpT92xIIgD/Osb1pmy9T6z4
FAt23NEBo4wAJhDFOKYagrrP+i4jmRkUAIZtkHx11GKZQ4iR0RWttGOtMxMlthvp6MG6huoxi/3d
dmFToK8p0Vc+Dt3Y7TOqoc7BxSy1dMYXsnFpVbOSJSHLT1qv/4/ulhbVrttJuae6Cf2ZfHWfdDOZ
koPNwRzyZP9X6/2A/xutOoPfTf4UlUAtpLk5uJlBdn8bxLtp3WTOrh4GaxKXhwD9RhHn1P9S3k1D
5Ov36+QSjTGQpJ3pCOaLbOV6ynotNSid8iftpRhm8AeRkcZYlSO4loB6Ihb1hTYEOGoRminyjume
RPEoq8wmxanCGqEYyFSSEANV0Y9j8PGxkctKhLRGNd/RT64HbS+fA3g9LSgjlqj07iMZoMx1gEnL
guwR8KR3162BgzbkvMdAfMFIs7tPLA5ZQ1IC4kRhaGXc+9AtJq6D6QEj7jBXOERLdCS1dsIeSIaH
nFfOwtR6Bl/NUH2B3lnAE7Mdw4GfUux8ptLH7xNRfQHZU11RbWG2l6czSLsoV7Yu7Qo2y/U9cp+7
nZ8CLwalZ4s3gp4e1NCHRVJXmpnPaCebOIIKr5ArGD1HzYeNU//8GHCF02S3WgYnuBAbYCxSvHRR
/YYg8jxSViH2WESksFVEz2hqgJ87Y4qTjBLEt7uWq8mJpjaI4I2g8eZEH25BHXqrtXL7W298bp0l
A2l+Kp1qA+bXKPCBPloO8Ib0btCNZl8Hirke/bslYgOBGILCDE4lVUJ2lwMh0cQoB66u/S24R1TY
wxfFRFDfSJBxXWnVL4VkC/QIGtGGZYl1HQvNB9aMkSS6Rk09MiPkAWTTXcC3VF4UnQpIBo0L1bku
GfIUK3inJkJRRmdrt9r20n2/nNeNS6+/GAOSWvUGFSbr/vLDjMydqa1rzndgv696Q7JZpwpwoehx
u89K62vi5WuuTNJlS6mCF5rbvEmjkaSdxnYSVcHxaUcXETYxk322FUw80/GcJwtFC0FkSBtmAnqQ
JO+3JE8g0q4+e3/CyaAVAZR61L3aD05PXvi4HRI4Ul32WFrV9G6SliPctEQA1EOHqU7/CJZsZfRf
gT0clvlYRwhFKtrXzDwHv2sQaCC1IAO1yafxRofXJAK/U1Id/uEMyQqErg0x7VseNFA34ebacTDq
sgXmI9MreSuP8RnyeYu1jIqhlX5CLCqIY783DoHC8htVagJjnIC5hwzoGCLbJCg5MTPLf6FVnP6V
PsEtEarDHp01kFOJF+WoiZGutTlRq/SJGMHYy3rkgHZE8n/WD/FuyQIU0aMcZiQoN2Tpw7qGRKzZ
sd9DX7db16cMLVzmlnC90oAfY8/Shkp9DmV/0c+/Bjw/6ABQmueANSDSQRyEgVgyUGpO9q26ZgsY
FnHPlq2AzEmr9icgQC3TkVRI71B91G1KmYfOdM6HdDhYOrKsvtbypeR54nUQs+3TlKiVmY9QM2Es
PaTxl3LjUuYkBB/KPbVan5eefr0Fdg9X8hxKcE0T0Ni2Qf4AUVdnKHzBjcCBw0/bzl5XPJJuwy45
5Nibu0Ttu26sNTkcY1xmLLDI6w8uhLIYgCRGn4NYuWgdUXC8DhUA0YvzSuHTZv871hrFUP75q0Z7
c9txXsTBGCNz6cwxvUJ5JobBIbgzKouMmvWyk25STpsp0tJYP/V/awm6MFKwmlXuRoy/AzCLZq5E
mk7WLQ4EYwjrDnyTfCkCfcWEt0A7HcCypQ1ektfJHKCPKpXwervSI8rz/f9dftENBQo86LvUwuBK
jyvACfGDpefLCD+42O4YAfzQ/yXUcUua621lmi7h/heEFH4JL9W5g+kPY8nzKQvYIf4aQVyjBKcP
uGDAaQH2GLqh3jfYjceIE/huj8gujyGGTAQmId7adNnl5lon7Q1DuG5XPjIRBgG/wk1dhjyGreTI
/pFdsa/UhKRoGn2Qezz+Dhibna/eTFx0oDcgZzyz5vRLaa26cBKjwBjA+CwVMBdoCQOEmQUBHnhD
sfr/No7bPtjG1/jlCpmiHmRY+YuOAGQsF4zdmkCXFTsByPZLjG0gMhHzPxBFfQGnbSOKBqu7yMqt
zlw4Zt4LLXEBBq78zXvTzpzpTMBvIaE0Fam5Bti72hBNZblwQ/ChwkBmK7Y97UI5AA30fVSnk75M
1nWNs40zGSZdk3vmgEiTNDRQKD6AgYs49zZVDoNHT6LxxZGlKRagnjt7QC2qUYuDAfueeiEjYmKh
GZeuVFCvX7we8VvPyuRHoV+gYbeqp41Wc6qrM6nD0jOdAhL8N2EzB+3z+VhszjA9Cuuf8R+4bYB9
KQGXvqWv/0rXEeRwASxQCyPZ+YeOnsucw89+acaMdZw9NJwNyevVe7yOk1tjhZD1aSE0y5fOMies
MlquDUGNjY66nqg6GjYgWQF3ksXOOCCIqXihdiq2T4FMTbrKqdLis8Ek/0DVDbLV7uW+f4tWeqes
OoUu84xy8ditBrE1k3vhSoLeRPwel7uPWvHwsML1YmK4mpei2yHXP3vUjcSh9fwd4c+MyIl/KHmM
IqBicYmf+S8r6pEJUD2N4MuEAynrK4hf3dmZlcwO/kFie3UUBmlZlFTynoncA6+xv0VBz5fMKcVp
u9w6TuG7g1QnFcNNR0ILhWVCrVy8ZOHiA5cqigNjscAuL6AegT07LKV7wbxE8BMrkRklAFd/EMyJ
ijlrceXRTwqwVUwgFvj6YruGGDk2b7gtrRzgMaUgtbMc/r0qOz1BSoYDoItn0DWy70CzYzEL673l
AlUIKU7X6MrSyrBsCBs30E3hbJKui07pweEHYfg/l0neHZG5vRz+dyF7kosRQ4mTEiMMfQ4F2TPF
QMiEnbn9Or/CmUnQA0BqGorR6C+EAQJILwMff+fcyp7hP5Uh2RjSOp67ro78yyLFxHAhJDK+Bylf
gIOkdh9H+4qEtGpJUDT8Aq9LW7u1an571zx2KYe/bSOxVXKNoT2J+1gHNYwZfAjBfw0gynZX0UZi
qEeJKwIrl43+xW33BQxyuA4Zm4QkaQ/YE45qcYXd9vHfMmrBBkVDbO8cB7jZRMRztzV+J236GOT+
DvtcJKxIerM1qMpln3C7Mz0bxq70NDvLmrRcXiBdXF8HdZGa5TDvwpdZMTEbAEK7Y97Y1DABrKAL
ZYCtgGcFVnisKxE5H61JdBbOB3Z15eemtwgIwT3uvtC2fxAC1zrBUTjLqPqglL+x1sZtd5fS65pi
62JyGpbx/VIuMYf2KzyfIGdr1IG/CGlzcA65+N11MC1Hzccd9PbANCGKzloQuBui4uy5c/Ts3H9c
xURYQMLo7q0PWrqGqc7KBI29hByMIc/PYBHrrKwNK7hYvP/qRvTuho8DHu7UBIeIhok7/CZgWonu
yZQ74yCcVl2r/amFVK8zYslVzbSwUbA2VbQED6jPVO5jZ6YMxkS2SyxS++yu5FFeE9YkMMBVkmRr
9Q5OqLMj9cFWQC/fa5zwcsoZeWynJOogwHAR2F5HX3ds/DKQg15r10DoUCuGO8nltjnIkZvWwaqG
ReON4kZppPDEMu18UH+oMpzMzM6oWfxKP3yUZb+lwCczQiZykx1EgHnRXWB/3RausOFJQNfUfg40
3dxW66gEzinkktDaSYOmiEQQlEObFFqT+kkCy2EAUhH+QnxcGBTWKQnKsxXWF7ozB1WWzPO1CWzd
tHwbXd90EW+0wU/N6SBXsW+XD59BVIe4sLEDpPruzHFtOnmzAYHrYShZEjliectHqAwNmUaJd69u
6QM5y1CVgiU5/RV9AJAzciomqbeokjW9em5A7y8/P39lQVZC0OyF2UhRC5nPaRaJ0yqlvaU6FrNo
FojcDA6iXXX0dCUvC4WRlU9I+18SErxwleQO1tL2BBSX2vYBoJFReV6kMLjhs0UnH/j3J2xe4gYg
EtfDcs5FJVwHpxLfCOBmr0mC9aQ/mKDiGYoblL4nCPQtXRQiT5sc1Lw4+fPqZFueHUMMO/o6ePnF
LNattrPK5i7OGybWNeddh0HInJU1T6xd89By2m6rZaAPUkS7r09lYPhRJ5sY1/twuMBg6cpNbxiM
fZ8NKFsT6yzMxf7h0eWDbs0qmdJ6LGTuCHRj6Ej2KV3hxIBXW80QplMnaH6ZNRyDg+/Mp+A02Eos
wZKip5W8sCFqPBYRDo5AIezYAPhPEHAKHXsSqBhA6Cz7REbK953pDA0u9mZAUUOog6rYjwQRGPN+
fWEXBHVKkY91Y0NmeGF5xPoA9jGPJ8j0DezDw/gIkLUxjp2t5YAcvx1LT5I6CyAw0mbvjufsU894
x7f/6KPmTA5YdD3I83O0OXTqUKfhiLNCfvY08pQhsttPv/1i6G7qSu27+Njr9m492d+SS6RA/xxb
IYRSxoEQhytOsZj/dIT9QJh7yPo9n1fCjoKd3xSm6IqX/oxQKPh7hooh7z3V2JbsPifOC+Zy156x
DSPI7Btx0KqhLD0qohv2JFkd80XHnLLV+YJGfTB3Twe9P6ir0vOremynmJod5yDz02qrd65v08no
VVlRTsVUJKYawy3FWUtqtj/mMGtbY3wj2Ys8vplWQcBCdjqC/3DXktP79iRDICT8eiI8mlQVZKtU
KmDcg1CZVnC3mQtRC7h5lddeeRpGdoRBuzdudtrtrADFidQA5E+s/q4ZkEIoVsk9ULHqbh2SRUkB
vkkyuWQBL5jR8VR590IJ06BBuhCETkrrWpH/KKy0NavT2RwekTqAbW2jTXTJgqiBkeHnrtuTR9QS
ECSQPE/NMmJOtaH/M8GFAJHoKkVKpfkLNNcVANKA8v+H0nYc3zSbc38JIYrL/nsqu//f60Rm0job
b6TYXl3rS49oSomvscYyRTElO4RZ76MLsKTzbkOseCoL5fDrg7z87TTTrcSgZzhxPlTOCmVqcQcE
YKW3aEVIHBUZjlylyldA2BB3lU7ZbsAPNAYgKS5yqDsO2u6Nn5v0RUNF7TqF8kO79MhFYY5Bv7JG
r9cLOT7+1gMg+h59JqkdVw4r9+1aSBALg0sVqAaS2WF7VsRvDNBgsfLNTEHLE9TtdaLoxm7WVArh
ghXyR+oxDI+hkryiobGHk5lyjJ6RnrxLqsAvYa+oYUotYgWqXf/7HYrFZ27k4Y5++rxJmSDmGhgK
nBDymPnY5SIIL79GGV4WE5u++ZsQonFa5rNm6kxA0BA0rdk8U0Nb+iqHWv7Ji5UZbmjxd8LfiQFs
+ki7rj4S053vgsFNKNN5pUBnG4E3f6aeevY4N9qah+ssFAvLX4V+DTBDeYJOpOO/rUnKPEHSUFs2
Mw+aIaCwxMm+2lPGW2P+2SrJIWKNiicOks9vtE7KP2FdFaDaDl+Z2Pjk6JTmApdE2XNNaX/c5Rzk
Uq1MAzemdu8Ukp9uQCbVZNWNTS3N52X8wbBDsMfLWGGRGEcjSb+QvPthXAF655lNsdbkeG/R9UW/
KBlCZy42brTLCRZaDuoosuKnlvj/TDmhBuJ6MkjiStSDqzo3OQfsWU61TNIgEWs7u5SvaiBFLmfv
LUES6U8KsgTVQz44xpb6GgkMEEllj/yRuVTw+VsU6E6gozC3CYZOjvr/ZqNwUj6R9A4UApteiIoE
jkaTA0xK4gYrYEJBIXmhYmorRM6dhtf/PUfAQtCqsrRqsLmSZOuQzxEXUEuddtOSmEOQoDB0Nj8W
ByLCh9CUFbeVsuRak0mgmlufuaX3z2JBXPxYRMRlHAjwVcLQMIn/J0b29w5C/1oJu+uo4G3TdFcw
8eFHb0tNFwS5Zubg2YZaaYPSjISBqVPNBVDeRd9X7UA1FlgWCjzPaJfGwVRm9U9R9ruqLb2L5a0J
drAYfaPtc8miIhL830/07Uk+cfmPZSRD/LaOOx5wgkFRduS7MT+9nB5Kz53BF8ky1Kc852qmzeTY
Pc8jtx0oocN4mnaLI/gVH4QLCw+tYQyLK2AFW46ClP+JWXregKpTXPgErbmqiy4ZqZSvLQ1Rhwr+
mw7+e92e+d6UzCxRtwtbRFA4t5yw6zp7b8AleLWx1OI0xNXZSvk+6M/JWFnK7fkf8M5NA5LMGqP5
qek3OUbsrD/f6Dbg46f4tJS1gJy6t30lT3+G3e4g4pQaKjJMJeWaT3bnS0cnJSFJxG/LBN83sMJ7
kugYtl8KogimtBJMdiP/pyxMoD+C3fJIQP6QbbMfOhR+6UzoLcAZLN7SvrlzJ+FGz7SDL1J2+sWP
8l1EeK/MhHuJmJ5X9OVqk0hNv1GIL6YAEVpWjkZPw3NrogGBCvTypeAU0GWT7hhlRjUd29uSCyrC
cghV1d6kjExxSTUlkFrqgDkUQd+FUrDqVBG3iRAG1CwhrjZvX84vDJzMA0qbNzZmNFFOf0ljfjiA
63VMRsOP2LwEa+pgdqR7AkImwyUCbE1LKKbNFaYumKSn/hZth9ldiCi68Vz6MDe0qGsvvQZ0mRFS
Nydf63QCRtiT6qmfBX993l7gwzVT6wgP2oUrxolDt5KJVQZscltyh2H6+BjWmOk6ZaFAd9G2cb1P
bJjfKycCJQTveiuv94HGA4GcigsV8C5zGcgdpolxESU+8enb+5OMBCU2itRjbCoDqohs+rsm2Fay
xxPqBN2QlxqR8fy6v9ISB18kSkQ/pfoCyU30/tigc4VXZed8TERtpQU8Hmis2hzdYdSGoqIaX4xs
OkYYbXvFwWvkTaG+VIiBv8rOes+DD/9HIRLGhbKpAHJelGgi/jvOmRQP5al1ENiE9IcTg4cCMWBy
ARRS7voNQ2EvBkE41I7q6zibxBiR+zl9XtZoAv/wze436VDKLAEM3ZlONTeyMyMB3NfxUIk56lxH
O1LLmWwIJ3pSjNOxatoZ3GKSsmqIu0GmylUBPMfsIqGh3uVkD2OYiuumLhVhBdXDhFbOfOR/Sjlr
ZXA6P216PtrguCSYEy48I518D72r0aQfzGPBC+NmE9iBN/jiTj3f4cDM1Tl200hmwZKRDIsvo+R6
8T47VeWWzA2KSkF2GnCvLKRgdT/RsqXqVJ3zML7u7E2oZpIjoQXemhvbE/kQXFrmIomHXgw95Z6u
kWlP7nSCEG48/zYZn618XQIRu9BwpMiws3slHL07NjhojAXeUJC9a4IHPIOTaXUBkoi5VjRCOnz0
gmTFGCs4gpBY3fCdJQlxwGsiNpDv4SzHr43r14pKW9g5pDWsnt/K0ahSsqxFGpHJ17d47WtjIMfm
qzfxJwrsEqRh4M0onW6cUSouQI5YkLF4qStQLonKl0MJ7Ffa7TI/p+WQsGva0+8+vVH0disExhRG
ngqyCI7dU7NAhtt4MH9bRhUTT45Q2WhjgaKEx3JNfQKxCB+cPnfQ7G9+E0SRZqlsCTTLx7fvtqjh
sBKtO/ac108/ghzYLyhCVo7l3IltNsOM1vUDUtG7adqyqGiH2cPuENtZLIdZUVxDedOc/nOovDB/
LBSQKoGJF36/GJTWcjGgt+/gZQwpYwTsH7PiucSa4x1XQfR4+gg9AbHWL5ZnBE4XdVgPuykhkoTs
HoBhxtoPs7eFTvFcMRFSPW4IwkeOUQi6tv8Jlel5IYHxQntb6ExJUEkfr+X0mxKYDZU2oyw/Foi3
nVM+QKArKBo8wnYRbs+WjUG81snkbEC5SS1Vy7Q/5ejrPt5fgKdcMcKwraJYHBRM1gE8zRVQsyaN
5V4IVS9XzYMegUvhsVT/9n5Nj6lbnM5ZRIyFf8ZnY/LxEB1oBbanggC4PvpWm57RiJO2UR73sbdm
jA/nim7Rn7snhWWehTsky+u/UAEXWvMCY+54/KzRGf0hWS9XelcO0tmMM+l93K3L5973aQXDl4DZ
0/QCviiV0UewrwphurN70DIltGWaEeEW30hSzzD+0hixqW0+fkDBxNMEihxQBJOarBBUl9GAcq2Z
L4uwzF2T4Eg9Nj/1IvJSjFTq2V9YcLEGX3TUPnGvClwpKQ67PbZAxYrQUgurktiZ2/ISF2XkLj47
BDOhEAQqjjXe+hU86iBDebFTE8r2tR/FStxjMeVdqwwTsLOD4YUoVAM6avnCh52w18BWyDaOao1G
eNvBJUgBCQRXEd55yGkrfrDvdKN+0f+w3TemtO2T5awb7zE9kof4bjayY3Prl4DT1Xlz5ZqkR4rj
MIGjLQco4AfivR3AXS8+p8qak28RUnW6tSjA0vWxEaUwhUFrpUjO6+INrtYiJYOCvDBcQSVDYccH
jttuQgO0eAN31cGcgqyx89HfQZbieDSycyAS/JLEvcVX8lctoRYCL1TZ+o4nzPUPwU/8ipty1iKR
eV2LJk3sjMzSUlyF34h1osPa3vzpr0YUNvi5rJ3+PMUY/YkwreEyUZgYieet58ZHCZj+4MIGe8mL
I2d1FSsQ0D03+oLXWDfxU/oMqnv327cE/5Y9DW+7qp3B9xfwAWGgvC/e9yKcUOABxTmV0nztC9up
rhwV5Tch/nsFfEy9nNSigSj/qaMqmJcYTRZ724H558TxX3JKg/qRwXdsEBl4K3NSYfaT5yKIM4eq
s2z7XAX3gJoroWsK5HkTmwMRtifdBOsJoeOtEbCLH4XaHprVYD2qM2tIvT5N1WCRiL3VXjKZRtKW
8YHufK7VkhGDrf/+oba19pTg5VHAInxsoUGGEk4MPVN8Lpy/neXJUAWVzvXcdw8jfYRCKGSrTb1L
WDYyVwMDfruvr2tMAMn84jHDewIVVC19H/S2AGp1mjofJTVLT2B1FMcxCcSg6JteuOdyGtCS5tM1
JoeNBc506e0aaX0ak7h2Fe0+DUBof8mjCzL27Xwm0ZsV0ur8sJyZKS/LMbJOQ1/KSL/lPKoNhZBZ
4r+YURJSENR2QNcCL/h4ECZoPgXePNJQH+3uSF8LjwlK7kVHfRvtKvYJlOa2Gl1LGbyJDpJobdv1
vPPR+UUYJT8zPgl11dAJiA6GMfLLjK+QecbIkPoJm8hBI6VRAAGYKc3p/Q/Ew31RX0N5elPw36Lq
mlPi9LjI3NuB2jdf18OJcsJHu025gi9RwTV4VcV9eIjY6twkFchwZvma/eGCRE/sq/Vn+BfjdIHD
w9c1ynRJMZah6WfyDp4VTLwn38dp7Y6+lYvhf+Kh7H8GuFMoe7UWoTGvJCQfv+FsBfKe1PNdOels
0PnHWBsOrVaMUbc9eJlESimjWFB0U92mFJ3UWwvdqxX9PK+d8NJIB0A9xMeBTIvFuDjMcXUUxCWy
dZHlcCLy5AXKsk9TM0wa60aACUaRYy4Hz3lIc/WM70CLTKSNHukJ3U8CN5IBI15YYksLPdyLbClq
tzTWueE+3pbta6tJ/W/nI6A5O5nvcSDILkx6AnlAfArLIOW24U4AegfEofiEryV4ndMz+1SFwOv/
Gd6SfecEqPCjGaqW14/UbFP07YX3s7wSLh2PtIQDOEiOHSFxtYiGXuOoSVXexTI2DSuI2TSJr2O9
nxZncDSibUTCKvFsY89FtXHq16OMg7yVz0edxZ5wV8InClVSwWgTJS0Z/Gk4Lfx2CbbChSQ4pa/E
VXM3D9gxSbmDp66qACZVM2rGn5ROn5vmjxEjmRUC87VqQJsqKACEoMHjvDcLSx7eGInMLXTMm30v
srWG2TMK1XJ8/Hu1I6B+5czeRkFShDvKSCKSp9cUBHlyfbAkb3yHNloLwsIv1WvaF8EjJWa4Y+E9
YYXmV0DJ6Mag/mhm3PYp5z+OjryTOB3h3gf9ElHLHtbI8/lVh3xlNchy7Om+BRMH2IlyEnkm0fBs
MCetB7utLWhvaIb+fpMgbpV2yC9C6JIRXBU9+fy7bcBbDLM+FKeOnyFwc02h8416b3+nmf7d8J6F
Tdx1t9w+zBcYMGk+tq+2Zi9ETjdVBIJMp84c+H1WRCZvb05D+LjgSoDb129dtm9ECS09PF77mIRI
bC43s/dXKvM6OmlVlnOliAJk52mgUFic/+J4BlA7+PQf3rr+TllkF/wudYG40cSWCFlg8Z6mxxTd
vgT02snxRoi2DSqin0zr3RYzyq0fmouqi+T8D2AZOK33+KYjihwvbmrPnDPD6QjI39fi2PrOeXqU
GnwCNOskynPgD131A0+2djL934nKRNC+Zz0nZnogJ/wF/w0lyJhxCSbFsH39i5dMeIwEpSJQtgQf
rQWJaWb0+zYi82CVsEhWWb65qEOXbrXuBq7EeWddljpxRHkZyt+vx+TtCzyOn+8llxJEhDwWB0CB
Usikn3UwsJqeUxgx0y+KClsXb3k4toBV2MG0ANNxHNDFep1Cn/bOMHG59u7y1BOQ9i4xg9EOja+n
i6TqB62yjfiX8j1UnjatgQm8U7KtaRlmRWuwGDhzo13TUdMV+9ZvfPr2AeqT2RZ+62odfnOiYG6x
kdVOnKfTmwYBpVA322cMPk4jW9hOgqBYU8L3qo2KhmCPXpmevNsf26Fp0ij2DAUXT2kmfguzC/hZ
gI63+75NWnxR7m9RnfFrPCgw4+QuYEuMFC+Mo77LNm6AdlOVXRHYJoQ/BlxWKZ4ocoAMLKZ9o4Sc
PRdQRls08afezGjcoX8KLEOwYL+27WJSCY8GXEneoSys8/hVeR03P60XmTSzK4gRzkBSyurILDcx
X9Xp6Tki+DdDmYi5OaU+J6aDdmldcRVSfcA+y+v0kGlFPtIAG+xJNkHjFuW1OBo8GnrYTH5iVScm
ISn24JyikFJJokTNCf4sCnrO1i+HngkvhOuNGpyJ1Qsb//AfXvQBkaOxpNO5uRKfLrshVtcxVqK1
ZLEv5HiJM5NxMwVtkzcnL5Dn1YXrO0YSTTZmxicsKhfVGnfKgGgRuu0M6qkDrpeKsKvFlp1En1UP
30wPrP6UBe+0jcEQpQDvIcGdEG2x4XkMAGoxs5fS1HPmMFoXNYswrG8MVGsM/227RhV2dqOk9R7I
KJC9tg6H6jN+pYTp+QQDhj+p8Q7YykeLldHN116i9wUE8FhVImuAPkrbHZUUp7P2YsWzXAI0C4GJ
ko2IALIdlHCTHXcFEEmO4oXg7P4HWMRg/s1EwfL8NKpN7zdFe6rWhMu/JiIdlcR9Bb6mJazNgFah
DvkxkjcyPXjxFuSXRLNH4uyYABb5SiyhA7JXzdCuAx56FxLkwK4DttVNmnTixSOsDU2WawQKvDmB
6buhMMeZgtprx0OV5FZfFjy3CRXADQkWZAJLjrEe6++u0Z7hEjYJ5ZvpIu7EJINUGLa0wKWq08Fj
OvpSjos30cukATW3ivUcmDavwUuNmUfjnpcF6ywesLnA4Yflf8ELcr5o7/iaXpEaKAA5gzWzT9Jb
hsgDj4P+S+Mqjav57fQMt2SUDoPD8XhbsqxohQNe9fAwRD1xJ1zK73p9LEj+UoEOFigygxu4mJ2G
+K6fhbXGlDORaDGvoIaeDV+SzhdCeBLyPxaEXhuiYq21FmETy6BlKUdiM3kzY7P83WeN6gmtkqZ/
q0Yxm+gTy1L+M976ndayHtbwIJwEGkO9feYD8/6vsTR4PJyh3hyO1VOwsvjKICjcyhMNXtXYDfDo
kIa9h6jnuRqfRxMBATS2DFZEqPs42WkTaqZ4ExwGIdAiMUm/+DsUJAoD32NQf5VP/ZShAkL7sbCG
dZ8IYFlXAUbsAUjjrxo2T6/179V1yvHivW5JFR4sdtuahPSb9MZ1mxm+438ELj4Kqwhvc5S4pR5H
KTdoy2XeVIc2xFwS+1vbZocSJmm1oROmBMVxTQibmjt71X07L3h3xIuTgYPt3AfuTY7ClCaoMcps
Gn1fKqyfKE+Ob0DAl+/SnYVLTlyDB/NDapS7+oPN2f+cGYtkdpDCE7mcCdWU+sMnp+v4zHVSszVm
CtAaKfsmlnSpt42OpfV493c/LxGWCiwtn3zunUyox5QwsjBO8/sN8NH3ap2D/LvAufAXlWCcu6gn
IqNQqAokM6Q+BVecddgWDmdL2p12cBGPfi/dSJkiC78XJRX1X1q5ReHnQrdxXy0x+vFQ//C0zQGU
zavnWCkmbYxKLX9JARQ6QMwWDybj7O9C0nYyLs00KKajCE4l5vti4x9Y4Fo194+lbjdzKf+ql+Fm
LmeNrS3B5Fpr6x2sMLGIRnRNP7qtQMhaLvDWoRc8tCx4WDDbPy0x2l1oA8Fie9THCcbPjrfmILY7
BvGQda1TEJVOZ2af9Tg4MtF4s+xqJEVNdQVDtaUgNHV/5fxyhApAhj8W3AFk3vtbKHuMqkE9hnz+
C+rhkfqKe1MQ/lQ2qGScZ7yZMMa4DbzM1ves7fI0m23ZhitZ6fby13qacleT4QTFW2fGF2udDBYw
Z/ctnQlCJg0dnZJcGoWqbK7ECM0N7aewE/lVn05ipq3yo7Pm4KdHympWTBUNr2NnmHVV02r5omZ4
e0Rf5418CIGmAOkOR5lcX0W2T0ouY3VaoGyT0mWwsyEkyzAPY8u1zxJZo45L+ioS83SPRigBxP8x
bugXzGhnUYc16AblXzBpkYCmjvQlkyc/gPAd/0ft7Dofw7IOLt9Y6ZQKto59mZtDBSF+tba0c2AY
KVEAqmyOtFvViIKBTyeXsryJUap4QZHHpM/D86tWPuHOpGSnUvuM+BCbWzA4ndliJGoMQeowLYff
dEkgj9blSS/NMJqqAhT9cVS3/Rs5Y4MnYYkseCdbN2Nzugu86N4KiosfUKjWaN4tVjcB0UeJxFLf
aD2UKKheNn6/dAXvNNfh9W+wgNhMIG6/CcL+RJj365UvjZpMO0lPp7oyaSzD6sUZXy7kV0QiLk2A
1is/z4xcUlBGvLAjOtZf3FCZgICThVFbTrVbm+ji6yALDJSLaCgr+qqyqC12zPkdiLANkkIdj0J0
AS4apMIvBLqiFSQelxsFVIceaO5Xj+cfKHWXyYD+AkDZKANIA7pFPZT+TE2NRbozKkZF/U4tA4Nf
2c0uuyLhvv4jqrybgPWQW8EW9RpuO7XdZwR+1zELfRgjWHGvDHtYTBs3f+IhZ7qbdhrrHz940dwG
1BqnddkCEGFkgrYPvpfUak3b9oCESvRMnhwQWPfg6y7F1bE4n8bVOFP3w06OMb+Li1/fPUQZoaPF
x2BH03OD3StfhppTR3RjgLqkPmh7YHelhIKQmwcxgm1md8SAhaUxNF8/PAzEyVgAufuMKZodFWUD
swDDheoxZgcGM5KQD3cbCPhigkLp5IlD/a9SU1ZzZXhpnr8YN1cqqyn6NmzPrSsGfcXtX9iTPXDY
23qURIUr5IYR6ZFq3DrRQsHw1JtMUcgxe7vIbzBmWNPNeduwtq9UKpdo3WZzMVpS506nGTdHJjYb
2mFvNSiSxqdmZrq+j1HCQkgQk+pUxb3YZ75x7HS9poaWsasOIyq/ODHXbQ1MoSeIQdDmOcAuBjvF
3oeBZfbpyldl9P85wtaaEkcZWhfjv6KAc0kGzI9uMLopFqtDVR5VSUOSg63Sh4nCN8kcbLSYqyqx
UZ00Xm8v9aZ2M/m2CNvfV7F9WfrDC0K7GsBiOoLbIMoXp/c6C30wQv0BqfkxKdXIo8/PUb3DCJNP
VN/HaNJulwSSZuYUGhYc50HO9qLdCMwdY+L6wLCehoq0igVIwaTCVHdsBBnLOTJk8jgEbOBg31Dh
wjsd++sfwgxhGpO6FWXEjFut7Sj+ybu6ikpD6h7hmUVck6CBC3CqALXeru73vgE08qajJuN5p2oU
HUZzndOCRKUsDtyGg4ttlE3zzzjmHXzteD/+rfusyvwnIIEswrdTSLtZoH9PxmKQtHosWT8n1UbB
wZNW5I73zeXHh4zpSUfMCyH2f//a6w4Im3vFXrVlRikHwoea3CjkUd4CIqtKm42LIwG1PNLUtYpH
9SIJqnT+4gRGvMAakjesWRqVo6NlTTtiRQdKWw5k8Md3SfBf7w8Cize0ppn0qhPMOe/D4dbZUkwc
cleSx+nN+0A7J3amBbJDsWTMCTvvdqYpbYzxRp9OPgzmFMTGXZPmrIUOissGbhyvJKAEJ93Z6dGg
JiRbOLZvCjb7G1XBCnMsrMfVMeNwD43Hva2rAKJU+BatSZLUsCvV/RnEUZkSts7/i2H5ZtVyQWBt
sTkhL+wU7/AAX/lRPKZsFcIqPRpUZU7rky8HoY97hb9tG4OfajQcPXK6dGuQ0KryNanAgIi15BAz
EayCatqfkgw/L6qW20bagiH2G8YTLhkxJxTzF9ZIebMxSbHIFduyIJJRxcvqAKVVl/y0e61TDwI1
2FsV4o4xm7Tbk52t6am6mV2bVD+XzRKmrbnbs9yzb8OWDx7Q0sy1kz08NMZ2+cTZ4sOOdoQXliTc
ZBvdpnitT8U9OnZTAI6aGLIu09m//+eGxPT8Yc0a+YnkJZDsp+Rie2CxWHrwnxI7wCFWUH5GsDVI
b4LYrBXyxTnz1fYBautDMjsnS7u0g5cPeri1XM5GCR1LbN8OYUqHpnJeJSjUNWmfc7kCwqCqdmvu
8226ub0UumXQQK9w1oVUJ3iVNuUSW4VMOmaY4K9xncBoTuJzZFoVghw/5cGoP/59NW9Z5TJO6a9p
0bzXwtjfdfTuV0onzPwRrd7phK/OkNC0CgflhXMIErR0CNy1gt5WHqoNZSFIRVVXbDcUPSXTMBTr
craywPQFUtZD+ZefndlM9fx58k+uddPasGWlnsayLRgA8I2uXBtZKMz/dxG8N5+tuqY2R/yRa2OO
avTrX66nZAk0VQr1khTuYOvfjJaJriet0Mejsu9W7LubzjavIfVtG988G6hSnWVXKu5S8wYFTuQM
NRs8wSjxeRVwF7+BvjSu71Y31nxenZ07HnAqDWyseey/Es4SHJgxdSr4TYG6kga1lkzaP6BLefba
L4g0Y7KMYRXTTKMYIzmToNE2+SxCqdXk56gINzJiNs60PLTjitOOHD9/4x/EVRWSpY1DbPc/UjkM
htMaLOoRc6QIFt9XcIRkWkjJ8cOgXQMqno90tBV1eOPhiYUx6K0f7FUyOz+Q9uhAHUCtCxPKI+dc
c6v+JDc+115YJoqxHun23yLJ1AD6VbI27Ea57QwdIptN4vOOZw3gubtDDziKW1i/hc/jE+z/796u
UJpSHRweqI19BwkX58Pgojley8yWy05rZZO//zddGHmbwiABJGF9SmMXP4zAb3m7/BAuS+M+qWdl
dhWfBpt6wn8zGcR0Ntaa+OSkwNwadTSzaImEPk/2PC7GZ5LC3w3JDc1HwApJgka+jTPP0QwMDZCU
xu/W1r+0iKO66XE+smDBsBSYfFqttlbXFXcEkLJ2sSN3jlnivz9PBMCA+U35yiUMcJAPEMlZWRXZ
b3LAlFz5QWoW+bZyWN3hN/yIx2GYyNoCW1JueFRZCT9oCQRxZFDfwSUzQucOu03nOEgJtGSKkuOK
N+OxuwokDX6DACoPtWkZmQUb6ID50oMusoXKVShxzsxbLfzp6LxzgOyJwIqboBiqr84AGC0Hvzq6
8VnyB8ROPH4P3K6SiHXM9B6/jLTJvWIaLI3pxYoU2HdyBTyIeWHsKpp7NGV36ZnxQvFBfIqp+bgQ
mX7wawlP6GhYt+nj8B8DSMapdE6Y1UBcw9vFhKVGJJtT/6yiYCbo72zfMbpUeo5aoMZwW4feGmHp
PnW861Ci7H9dE1/wpvpHUNfczD/SQ3bMGsaFHXI2yKUkCxxd2+RFK5Ni7xFzwwQBa+25X9wLYPe5
jMYNQP3XHPS58k9GuP71iIKud6enaB0xtBspV9NhxfGgOFKTM5UcKusckcv1pou8l/gKEBeDuKaH
IIL8YtJrcHDtKFhhVT1WhCVXJfIo+FGUFAgYr9yPQ3S5iPtcQKD4kODrMXkrBR2jkxHsSzWIPcWP
SqwOd5IKLz+2OJcq2Av1YkCafYeC5PeOAE9KkR6PmhXj8JkN72w26W2NORmanfgPG54oB1ECRhQL
8cFX/xzpYfZ2Qp1xdJ/ErvFhpbDSyTqSpS5KPO+FdyAejgvN2S7jNGUPzQGYUTJ/ykOaWxFixGaE
ZEqrr1c769z3o9cQw2KkmqawYItG5EX0NnG5WECenDTopteZnVNbhTB1kPjjFWgJ14zQl82bmmpa
hh0ojlpSdLUASo9xGhSOrSWO/AwGLo7OkXRRB3F8v+ciAh4dOFk8XY1CGnykuBUrH5McHLmPdldc
WFVsubWzWwgwui0kwIF96zXh9kPhjRDEXs9/OYtGP9Q5ZI4mNHHxhgiPN0JFwPZGI4ITQe1WQ0Qx
14CA2k8m620qLoKwc8vhp1QlxBkTwmasmwSxcDW7xXEgLj9mLdekH6i5frZzHgVOsucNFTosckM/
H3OHiZ1HkYtrz8HPxMt8XtBQG6m8jcxYW5dTYu+u6Pput1L3ImOigF/h/YwEGbQjQt7e1eAWJEAe
/wbaHcTfDL5EcBsUEyhQjA+wGFaD6zCt7WvYbFrXSVsoJ7Up6uRPMVgbKXPTnCr0/y5DngVCpgRR
EaG+ifyX6xA+2I93fy4E0VK5KQm18j1d33WHzG770UJ1Op+pDJglk1wMlS3dBI+BQrppfAuc9Mqg
BGPYRsbgNV4yiWokLUzabcspCYj/4Mzpu5c/WdmUPPmO8Bh+rJB9rSXUKnOcB3w9knEuUcJ7YTbq
0OBrfYvFeToP43ytEzO7jhz0tO3TboGDsGJcXQ6tQ28/Hq7Nr+s4PpKJcZkWtAWYqv/OZH+jc9gR
ld+gmCZ61iepuz2RwQOB32vXBzmNvwaAHohlPA2cbbS7MuDcsBiMYULtCc/DSAGwWBQY+CAebotQ
jYdbZkecZUWtFqV+gyYEOt/IzwmiloMT5d172JRJtSdp2RcMMa/FofGwEb7LhA/N5ftDnMAsLEOJ
XNUNCxd5y8gyeUM3oR3ikTKsPx6krBeYWwsAn7vD0wmMDl5A0xePOCNf3cpdWt2gYiuRx13x7NKb
MUHwtzoJwXyLzBGx0wGTbnyyRAfIomWMjFww+elB5S4p19AGlNYWHAZ5m+2as54ObpT6LtOOr3XX
hAU1espzNr8taQqmlK+2G3y52r9HAbPVEP4haqqQ8QSGtqUV8gYx7DcDTiRQpaQSeaNalC+woDH+
8ai89VEc/dmkYImUxjF2+6xW0sxx6hWTZDs8R9G/OM9mIKUTsn4Bddozv81k04Y1zYXV9F4zb99A
N3ky7G6pJTp6s8E9tYb3AhRplV9rlMHnxe2vBvo+HMeTPqPVyeg6u2VQ26HgWqT9mKelRvLM9S6N
3tqRUxb0BxfwwR6StC0KjkCFTnzKiLAPwEzEoeRV4vEti964EjWX0rg8G0zrs/5ESXiJdkB1yO1Y
YgfS4TZEnAJeanZaNdq3Oc1lpRYtgVnEl9oBVs0Suj+nfC0i11NkeotGOT4Km4vP3ihh50i0lbGh
CYKp3JsTY//T5Mfk8bR0mPzUSV+L84pc8VldtSlr8m+mfUkLVJVo/GZdR/hs2LOPpxMqFgZ/7fWo
G3h3trlONhqaVssElys6XJ7ms3+XI8VUTgD/aK1DtpZTmbt2GrN8PNZzoPW3RXU5AGTQHhVuDcPw
Tt5+SKkTKW88a2gGqvXHhNOw7OyBb2dfCC7+yoP0WDINOgzK0ZFD0cOh6hZzT/NTfIJ0IjQrazQC
iK/6tGL4NWkBVkBw+qpsCXP/iFq07WcZJMFAskFXpnckkrYkwn1gNgxfRkwteAiEmfAWevQhfUBq
8ABBztxT9Gd0sVn+BmxJTfCzUybXaBeYL2dCzugL0VV5KOY5FZq3b0zF1AcuSE7qNoba8gh8OEUE
5D7lVYeGiQC1CNaaDEbOBlxHkSGxGHEXfRqlZ2uWO1iieLrsRH4gFgbQtCk5rUl3Y0nBUeBGQsBR
aIzk8lh9uCyIHBYgJOzEHWgdoEoW0XqGdzBYgQvaGNJ0b11B/qTcF4QD+AYPf37L3AyuIdp43f/0
LOorwWlBg0UnrVxZ+qmAxLDwHRB6FFMOv6ngHfrF+i4q89f1j/OAqeTl6uDwZ0Kb8aW897c6Wu+x
RxnxdePl6bNTO5xYTGetIGF+Go+cZwaT+errJMuK7WYYtenbZCZeSWBa7PBvosYRQ02lef4zagw4
Hn65UOwFHY5qsBeHKna24Ty0k7NJxERQUUeeJbd6nXnFPeSUSVEOjnGQGnHXdKi/laO+6XwGUj6V
fVKAK0yGwFYpszkl+HomxfpP1BvbsJ7zdj4wgrJOZhsbV/blRhRwbBFPf2nVWt0x5j1VG8rT0Aww
Dy3beGnoa4kirQkVRiNawSMtKzVyqPPSyyfKHnl8XV69KG0EYC/sMbF8fuOyC38B+hm8gJZhEvM5
cl4cGYRKyzw72qYfJECKAc3h6b92tzFsIUUsG2jU/C3W6tsB4iHUQ7JV0I1C6B6v3D3dSkaim19P
Et2xv2gjvfsJfTVQaH1LBoZ6JvFI0l/iaxibtSA4WzorXzz4QviWgQ4kBgifjqXOSHdvM2GawRtg
WOAtiPL7M/eHE/dG24kP4GgqfGNBI3aEGoTKwWOpp199dhljsIVCuOKiGe92WeaWQJN0hZLPBczg
Y0xRBBZWR5t/MVK2hJQ1UeCrHX9DQh0RjKcbgUFR0PBSIBlmjqrOGJ7TKFEysWhotefp6S8pE3v5
/C9JtNS/swdirvljW7mLWgJcZA2byLIq+Gauy3eXvp1SkUvsma/MzeUOn5FbYCMlxJcKLBb/3DGj
C1ynB8k3E4EAYXfzOhGSWLl7F8wqtvnKSxalkqpOzd2wRB/Qdea/WTr397RoqxrmsG9ZnA8yNDaR
KbQDGzHx/Hpweb2LA8B08iE3asDzoKcp/EifgNPIjK5XEKkhDZGhNMn+yKa6ft1K3gkrG+Q/z/o+
TIBb2IK0J2tLr6jexJJrVXmuvYohVOxloEM+aBNVJWTFV0EynAoLTWGnIef0rNsNHyI475Ec841v
Fj8VeqcuEnZVM9GZPjaufEaSjFiJ8NyZ7C74VY5ugp7CWILLtbPjoWluFnX469AkcC4hU3em2len
VFT7mEysaJO0d7fkrMtuzWB23f1JZ0xerma3WcslsikekxDJVdTr4dIMTpuWGoNvLBifx5Dp2051
unefy5M2Eq1vRLfvNxOSBta6VXIkms1fwExOw0e8z0ztd5V4gutztxdJf5cdq1YSV1ByhuXNKOTG
naMXadjvmZO613NWLmCaMiECu0FhEVQpmPE1KiSVYoKJio0gwB8YPPEDAXoJcD4RiEcw7urTUwku
gcavYH+ucTOqyP220zVAa85Q6h+979kshgCLIlUnVleFZ9hZMgdB1v5EyFQXe9C1U08FZxLiX4Ti
L9mT5Lcrs3VE04L19VlkfQYJNe/lF6ZaBQyoUgqlqQO7s8gMBAc5gVm9pKUGfs8wsP9mCXWKhb8k
Ni1btMxUPswj+C7GTf2lFVxxIDyL6tiXdxmwDhEgirekaxi1bmMExbdVj7HKwFbU7ex8okGTGbv0
OCwPwYq7ioLoPyzz0KLIgy9LsusXBMb0ko1/1hJ/BHVYWXKuO5Fo+gin8tP48tI1ldJk9BTu7W38
GmZP48IkjFj7yHawKb9VfZ3gC3vYVUoTpnktxT+6SeHhTd/GmGVb8tc78OzEHaGdRsYJuycKzuCX
DdZSeJNLS0mmnXRtnVho2w7KGS4Nv2W1Ryx+yDfh5F50CLkdh9LzVNmAGhZkma3LM8Mgr3z+yxQb
1bkmchpIUT3W2m7qxoHa02QQUgcUYMz3YRRAPx5r32ZO4hLRuaZ4OFNKb4GhnbeKXj4nw/JGpvyb
nwNCeL9GwaE/hRADVV+SPkK8AttnG8TrYIc3K9R1bWZVy0npDJselZJicFAFFYviKhmmUyNDUu0v
2zR3mSqFYNV5qD49ObWZwgrd+XbNuODgiIsjEXUDXpAqmpgtZXEPgrSX2NS0oJ9559776lPkFwpv
3xvt8kbRxmSIRWVqRhTWLQR8HParii4t/lpLHJZYwPJISSebOivGSeT9TQ31nGjCSQpNOPrH8Fkf
Z+ZmZykpvtdb7LOqhtKq1kYrQoKMn1Trg8mCUL2CKTpCsMCTKg8Qpp2KDODcjACjCxY0WKOBld2p
AV1ybhvOVX4bKBzShB+JZLlg4qWZnF6zI9Vr8QOTh2IhRrnfAwy5oi5u3jAbXJq5c+ZmXZdVZtNV
Wc7rHAoDjXekEnjhwVG/aubPI3Eq1TOyVIuopEjsrAxe6u1hQv99fIaT+Li6bIxauUoxUkDUOdng
YpJ80MCN72zKH3M3f/rbNzXFa+TSLw6hSYsnaK/sK4QRbllgchXqQQpaB22Al6S873DlB8Isu+fB
zvIvZn+/4+0a2fGA93zXCu/tC3aWeVvnEon8Pr8QzIfkOKVswQltRenGLz8KUBMpf5jpB8TgNZTl
rG+S0NZb1MfisfBiqanUMUMn2VNmlWEpXacfoUtnHWOAC+yEJSbUkoIAzVKCFhCG2SptvM2gJ//K
f97QPfNT/47Eb2V4rs+HH5jhuGRY7ov+hBtZqe81+ki7KTOD5kPxQUjZKyIkVXXP3YPB9kaunz7b
salvdNc4lxo6QQPsh0K+L8Mz196f5n06OnzrUi+lLa8b0/4MfThxuJY65xP0HlNrsvXcn+CHRby2
UT9sUQnp42azu3VrS5f+jSIBfhBwVZQeK+PBqVWWarMtRI9G82gAki7XeYbbbxOh888bi1CS1Bm1
eUtcHcf5t79/xOgwVNIi9GJdWBnedC9YXANtDSuSqeIWsXOoTsYC11B0BM+gSd2IBnWzA5rQvmZt
G8IS81axm+KgKc1GlpVhJVRnQxE2zyZSQcFMVXiAlGM1pgV56pIYqgsx/iBRPJ1RMXFp7ANB3m12
yzJzQ6k6sMYZvJNZHYQ17e/z9dhjCkPn7gjtjuEOL2FXglxfvaoBkwC3POA6Z8USy/UsDN7KZofT
9aXDAO0R68N0Kg6bIQe4bsDSHs3XK69Cf3QCMv4JdwITeMWEviQpFHMQOoCJF9OhX2KukIdSkLba
grFXXOvLxNOdrb5B8uBudeLmZgozHpvpqkA4/EM8f7ppWRyBQqp/9xdD/e8+ydz5+EvzdBATJyO6
oK6o+44hlZxNJjHO4Fk6ZZlHOj9Egg+XlJ70CaN3MDKf+FAaYq9ChxX+dJqA++250Xl+ggHXElsp
STL1HO17PXPKs03yIA736fpFCe6ZXreeXMJIj360puZWlurzHrTsXF6WM/AP7L54RPsUjFpssU6Q
Z/7hqZF6BgMQ7z75kkVZy4KHwxndpBtVvu8ktUM5AdgTSd2UuBsLlQWYnWRa3bTg1dxzY84QB3jY
M8eIjdPr9iPd1GlX0kG8VFd1vFxbjj65/HU4x2GjhKvHV+heabPf1eaELkARseYJPHyy3oB7iNLV
JQNMZv4TyKGrVSEcYYwIjWYR/IIaGMirrutoFZzHs2vZFMNlZr/PV+N20QNQWFR3fNFnK053lJLN
Qd+MPAiT46yeOuRfiFxnfz4pjnTbdDq0OHhVxxy5YgQZDZZH6dIcqDstvSLzs+M63anSMrCQBPv6
Jg9zIW/l+64KF3R/JRj0t74sDJnLF0efl5hC+TO1dChW7AnE23HfJ6CauqtAET+yav0A4EEg+nKJ
YaAZe7A7vtOPZHoXGkYNS7Uvtzq7yimwobrCQ5kcFdwJggQwgVR6Vs0k+QnWi4OKAqHKhOLBlO5T
kAhJndv16Q1gYlBStjZdUEv/Fq6TugkIMWILr0bCykZ2vK5FKLFeGniHWUyy99COcCGSrVyC8wd6
FCJuK0BVMyJf0Q5WCegzCALvaIK8fmK2G+x6gjah7zhBvPpnFDZbnOa4hGRIzuBVO6d4URpEfc78
oWJ4pUpsicTNOEaAKLy8VjzwbL2036g9FQ/GCWBun0Q6kk3/LsXCS4jPagSAzuLd0/RaxHL8CCuf
LGSYE4+1rhHAiuh/rZMrJILcXvmb9NaHcJl2kViHO1fiN2U9Ihg6/U2guXxens5lR0kX4jy8Y8UC
XDyTUzkeuWuYW0p1ZIbMQvKz7q+e0pX1gZPCed0qca0F1lpyMPFNAkwaA7KWe6RGbPLfkLLWhCzE
nQYiACAHdAI8CC0bqaSq5mNoWCWM7tFxyY7Ns+eqBFM4CBiYMxfY43qbrcsiiwjGbID24Sq+rxGu
amki7/w1ARtlFg9vximw05FgSEcyHPYyBumWphojmUBzOLf8IP+a4JqQKUukGo1grZQw+yMTcE7F
wBo9WzKl2BQ4034yFfch0mljjlrjC/J0SrjlwrS1vYOteM7dkaDn3wPYzoLmog05NxyHMb9+JIyv
qMHQK1UTOgAWht3zOP+S1IwFPGNPzHfdTZtYeAaxQT9ml9BIkdWskSF+00HiDntrWdTIgymv2exT
aQfKjPYqAN/94tkdVWBBybHyAPBGgLl1BUGQWQEI1k9V86+yF0QEZvLuJ+dgqX9tOZgOCqJan7RQ
0Ln47xSp3trdzche7lcbTGrLR5bCHKwp+IsfHxE6Xlws6OssfOsfQSgnNsKkD8+8vzFCvwJc5JWl
Rx7PpSmRMFQWRAe8xEd0fhQy9xwUjO8H8OOFQCs72heh+TMlEhg4uobw/9CxnerYP9gU4vDBndyB
8cvXijdBZbpCaxrGJbAOOi0FvUJqZYLmDbS079I+cn8Q99TJegWG3qPl/+/vt4z6W2rp3S2CztJw
SQ95eJDlwzVT66UXhcwlpfQC3HJTjNyer+RPRnnI4QMsA8U6jlH2EFKlz2wKGnCZqSTZlWdRNGW1
9sY2dGx02sBRLsl4BTg9ITNzY7fPX001va34ypTwl2gvCS6Ij4xPb/95o1Q9TdlcPiTrdwAaDH1f
83iaGLlBnP71xE/ZcbHKLkDUE30U4i9lORDsnsYgJdk5eBF+qcXkbr9phv60kTy3W/qblht9okhn
rfqi1vMXQmUTHYyqfm0AcmzFX6pTWSuzlAEGIhN/GeSFIAxC5MRWdaFJb43GliVhB9Ljl4IdH2jZ
JAQzzvOQvQIQ0T9US7pUJFgkKbVFktxaaJQXHUFFLJ8WMlGFcNT0ZRH2H1fwnjdMUGXs1Fsi+n0K
RYp2ylvOMcrQ8dlKIZtDeaGIVEmeoFNt+0O6l5FzvZYmzboCOWXeSFFnpvaSavAe8lR0saYAlV5j
14gDBuYVp4qez3HCw2lVAzaCSMSMSjBVzEsez/I0z9R7dfZQn2LOGf9oxRigQKewEUK9p1EKQnRB
ugoXSR+7gAzKyxoAKl8bC+lGTiJX0z7yc/v/D7v2RtZm2fl0sgSY76E+3apmFZGVSOcmBzJgEv55
+X9nbR+xp5Qujbs18yJmFFY5xmNeIqpHr5qVo4tTNLIW/emUo2oy1XWMKzXscgv6ALufCXUrDwn+
TUh1naMlUyNoYfH/jSZ8csJpk9C023MS1lCSL98ZjNr6QVFWD3X4nL7pSD/HtzYUx8nvcZA93Tbp
zpHGUoxxoFoXDw+Gyj3SMyr1X9htsYbtpHDQrDqxSq0kkU93dyJmZGOM1Zaez1B67nXA0v3vm2Cm
mHpIRlBx0DJLq64Rt02IHTZL7wVU1/wA9Lnaxo+vuKGEtXhbN6+FaQC4tvY3cQZfSsXP5QhAOZLA
bqspGMZLfKYfs+1O8F1QzF/wiIcIxX6JoB9tuy5A8OHGRGan4QgdrK74Wu/1onlg/0qMWzTpzORD
ahMk8ORGOJx+3pPZNa+LazryB10iYt9lkZv311t5BO2OFIAZ+0WfuTbs+IQORcVJMC5EGIQkfN8Q
P3J4yQJUhJZDG4bkIcMvCInSGCoZ7YTn9f9BsFBZoHt8WZBPcfDUn9R5texcdh9Vwp7KCZV4N+/F
qkik2EQyHHhYiFPRuFuVREEaoFvdcbK3Xf0eKbCz/90/kPVE7QeG6/UBR8Y8FFhMDoj5badp5ia/
VVXDRLaX6AVIxG6/kd/BG+wi0jhi4ZntXYdHu+Rl20pxb8YV+UHhGzRRnZXFon9atOsOECnCqtmd
KxYquZApOw+mEtf2VUlnI5D73PBeO2CHpn4zt8wJ7ScD/EeOWrVOszHx01dLiEINjF9GLTgDTjZ4
mwR4Qmm4pre3MyO6Jyi1aQSlEvVQTMBtBhD816G0lCL5AGL8kRSAtzZZTOC0u/SOChbZi+a1WQ4K
400F0JucYE5geLjAd+ZkmFkwY1wgb/iAoSqQFad0k67C0E80LSw8cYtKj9DyMAi+OEKYzuWabFka
jmCuyPgHaxkuRvyJXgIvfQTDhRsVxihaJDup8rhhjcnCrdsIEdUYt0FALt8vgmIj03GEyN9R2uR4
iT8zKfRdgZeKkJ5IaI4/1/j9pCaLgbGszy+qb1XR3w1n4JD97vLeaqyuV0s5tnpYB9JXFRYg9xRZ
z0jmPPBJzXrkqdrc31OajrAhJITQeLxQNba536oYNflxEEq2JzXlfQrmUzTR/suMj4SmJcnyR3lX
VA/5RKAoHh32VRCGRe23UdlG3A1DXGV+Q+w+p8aEtx42ZDspLPwUaSdBZaz6A0Tkgszv1RmybpmZ
zW8zZjRqtsBiHhCsnAv6Spm2ZyG0VYqWLsF4zeSJLlWLctCN+YJMxqFGS//PfXjsMqrmzMaWFO52
zDBKXChUVw2B497X1iStqT0bg8hDnshr1j7x3JzAbxgp2Mjc6BVPKaggCuwDVxTvFX6KwBQetfWM
5bJg0jou9CtcFcVRSvG1EG2akE5E+6PaW2cwPdednhkFU73KGoOA1litAMi5aAZMF/hzk4QYlgsw
cCOwliRDmy96jLEyUyoKMfvBwcjVUaBLRESr0RfS4SWttmDDVBvh8WDTT3aZMzmBD6/N3ZOh4n89
/s+4GTDood7c0dh2xoh6ymwSmSgU2O2e8A7iTkWPWWhD/7CXMylpbHZe7tKXRm8/QeBmyzK3fHUB
VfSutA4bSRuCYMrNfJOicTS128G0XX4WwU68pxXy6Q3iGvopbI5BeUCfIIiz7EO7eTrRog8f3mfd
jFx+bNTS6gCsnx0n2bqAmy1AuFQEVXSVNARTO0TwrVA8y281LY0TAluyTf1AH4bpw6ehUlGeqsKp
EGV0Fx6744mqJziit7KdcgtDC5qNzWwXzw4gYa916pdROjWu2kSlRdNxouHHGfj4E+agc/kY3uNW
uT67NmmXBnTF7J9VT/EzZZk2LCdJKewAzp2GF/QAL71ma+aiO8+FRr2D0VG6IDqMlFDmvu2Mx5Zq
vhi+dp/+kYNptqvHRP2DJfcnHT2iNmh2eDfA04BrHiSG+eNLGaiUy0z1xjGFbxZswtwyVK4UTDUt
jxhzjfB0G7Rul6yTW51drGyCVYLP0qoO7vyXXM9lE6uaoFZ0OQjMs6c3P9rssoecZO5y4/73yMrI
G9AF0ai1qNOd+wuxLFcGn7+HcGoV37wjPYhejV/ZDMJ4Ptw+mJIj4T9gXD8CO0ZDys7jmPQaqzMp
yD3RHpUB1whU4LHv8DZoy8XlU50F1WZBmasK0KR0Pnks35e/tooh5EeV6OWmzykI1xtazTtSpeHa
pVdXlQdMP0W9Cghv9Pcu2KnuqqQw4qocXj25/QW/uMBwACzGYeeDUtqOHpkNNTpxj4/zn5MVDAve
AhZNdXww69Q3IdEHrkhx9ry1v0TO3nZkjvTT7MAsjh2ZrxSyDf9q/23dLB2icymgLz0KoE39XABB
Tkmo3DNflfyVJMs1HDM3X7/PxFE+SOjGCdH7MfZ0Bm9nLlQJzhpn54i+2pSuj8Dq50F6YfeS8vPT
2UIgBWPpyflZTrGN/vNbAaE0p51l3ojwdE+BjELrWFzZgyrA/DM3hU3jpqSq/IiD/L4DaBbztYxi
iBupYL7+NmILMA7TTA3LPC3NP/y+F+Vbl90+mWRpvb4b3iqtoqIyz2vNoS9zzUHBJCaVgwxuM9KR
uCiwmDrkZfMVG/IFyeuLeaeYOXFbrunHrpRdo8LMz5yS+Fk+++sr7ymL7MweN3eHRWCeJ4PJ399x
Eo0Q7Mau36VcuhlrHqLWTAp9wWrv3LhVb6eXKEt08tCEvoqppf0rpc7oxy+6akujJFE42TYjeCkM
K2az5f7/H81YKt6k0Mm3u/t9lqU+ePdTIZuceLba0tZHlklfETDwop3yEfOYms+s9v/OkCpY1pK2
vn85I4dhsoULexneIIC04d1L5ZAkIJ9MZl/xjSN3SfUx+8K6JtcTbQOJ37YAVGcb7nLAgv1COomP
oEnyijc9EnORhQGGgRetNm9jM9oppYIShjwJR5phg/IXco+3k9Lw+NoVQ9A1mV31d0mcowEd2v+0
RskTz9rKBfD4e59kQRtd+phrkiXdC9oNEWl4Mbg1i9DIgfprbOKdgF3t2KQesIWUT+hidjDWGC5Q
uZjIg84Ls+Q8zV3FfNZc/8cXA5sFyueT8vwSWYEgtWxhlRNL5N77laEmx/e1hLynqxQO1cLbgQBk
fEZ44tJSV9iJ3bAJsg3vBddU83S8UMRhHDCCi1DrZ5SXOw4iW7v8H5ERU+XcGq0VfoYKm8OPD5Kx
0O6BMJxHcE1vHtC/nNYXWcw3+SLdU7snndtlSn57yz6BJJk/+RbQxMcQFP6zEsXFnf7Tmbpr79zj
X/Oj7mbGiuhIAp4aQmoTm7/xwPTHvSPWqW/8I37iIG1Uav5ll7rrUQLjcIkY2Z7YjgguOYTM6QTt
eQYqOCR8IoYZoYBrP5ApvuEPd62/Be8L7YodX/QoxX7URGB9j/CNeMGseigYxRe72sldvpDgBp05
CiILcXOf6DCIwy8J0voQN58SP/HFU4HIVM7Tzeb1y7GtBK6h1c1db7iAAJv3CRN2Mwe96roQHjLh
upYYjmpeinJnSqbFXTb7GSA9YyMZNz3AxHxS4wL/HixJv6lfBDnmQ7zVwjdm8OV72I8Hwb4CXsHs
yJPwGwk/iIzfzXkz9RrCbgnanB719PeehIWErSYC9EaT8Y/8p570mJbhzoFn/tYp6mYE9UdTZkY/
qD5Oc5urnpWjyKj0BF9t9tLz3rahwl5fGEQhVBW8wBq9UyIKwOez6Xfmcu2uj5udoqjYr6ZnxZeq
xoqg81SRB13xttLKY9+q2ZP091fy6syExzZUGfdGQpGBrjnaQ7hStJWAwGQdMI77+KubSNIyZUjs
Aa9RdHLC6ir9KimTXFviD0zW0BtGW3wii1YbftKO+mMSTZZypnHUYAFGaTZ9FjVPiM9D2MlXW235
OJkwCS/fdH6vGQ1+ty7QClk4Ly2FstqKJXV7mJ/UiF8Gh4cN2he8OP5MU/b5HugWdaTf6bisChPO
d6lQXAJQAgCE8EEDycpyl/IfHSVB4fHckVQ+yse1b1wfaLrbUWmkFsjJBaoAEBR9cHdRgCjgJQXS
wt0ET5B8ac5Sjoez5yqDBmcGdcxdIdY9f59dUxMhdQPR7NrFHo+btrMQYoZa4RP6kzI+bMW3lT38
ykC5nec7KMgBNQF43XmjOGfZVUpcUH1Tl7Ho+ehGgBTZ5LalbEkuy3WyTbZ9KTd00lX5PkaPcuaJ
VDMdP22bDo7UEMlrzx1h9et+zIG7WvY6FZUwiTwZfhRGvXd1DkvpBaGjX9N37WlEmXvG7dcBFoa2
3WpDuqpTtkGKqk7MBW8IHS5uX7G5eEiz5HSiKNwB/3/ILprbPEyWAfyvQmkVh8u1uXbXgNuZ2+YE
u9BcRX78Si82W93s8QqsmjDyxG20WNH5g931vZbANwR6ncmpL/Wo0rldNKELYxw/3Xc7adB/UDCs
p6dXxLC0HhouGu9IFnO5/1jYT3C1W2RZitU5XEbzZ1tBHK40eucJ26BmeHCTnkB22JFQ+NdLDh8X
1sNAsOYXBhs2aEmtFLPnzW8F6EXpvyDOFi+xVjrnR8eMGG1zRuKPpefcp0mOOHePvXBy9v0EWnp7
J/QBPqx26IUOR4uGiFdTtYDkC/41dxWY+2GqxeltlumseMAg+apqHEc4jrIagF7ArQBLiYtECCEf
9O2PQwDEmKVRiY5EC2E7gBQ5h3G5akxAH3SY/D8PkjLWQNrTqQkkEnYF/+BL6Ujke0WCeU4l9QQu
oCK5sqIaw24dDKbW68Hp9WWciN/+t1xHjQCC6trCJQquaH+v9d0y3xL19RGtHKf7eoepL+5H64UH
XzZzteNzZAoWk6BNn03MG8NENBmr9rb8Sh1QPwfQDPL9kiEGR5kD+ENpKDYDF7M2IUYKKly947JQ
DWraEwywZJt9n/tu1QJC4ZOvA9enKd2eJ968fOMZEZA0NrEvE1LCGlwGnWg1di+qLq0YWeyP6yDO
PYMjqb8Yi9Zlc4qMaLIb15NAqpNZ1IykTCM5OjbUuRIqGrx69uuIq5wW1BDP0M0DxAOEAnvdt0ch
Mpoo1OoFOvpGcTp8Mrq0aWNBdfZDmB8JfP9ggQV5by1lHEbsk0nCc8DYOtDWaSvCmd4JsHOPz2IN
5Z5c4JyvEZO5tPu6/vxdSaGN0vW0hIhzB1o0iTvYqUk2etYYCybfILHrA9ReJu9MtIf2AHO67seF
849JufCou+mN0D4fvaVmiztROrGWbEOj7KdICtu6wKC9bfPE92d9br9kJb+O16IZvDrDLytt0XfB
rZtoV0+PIWGOAdni+/8CQ/mwLhVr3TlxoXEuft0rQFlAekXO9WIhMbD3d4UTC6i86XO4TUpkDjcn
RarceQ+OF9IQGc9f2x0cm+Y/5toTzGjwK/aZ1VBqhx1AZHoDbfn7cf0+YJx4vW31LZcOZg0Vw9pm
/k1GTSn4PG2m7AAUNx7YGekn0jzkeJfU+hbscNKSVbdhvRJKwmzCvDLpCx68jHpPM84zOI5eEfSd
d9zAR5+yLoL+Hii+kHuwpkFX9RyOx9cKhwTjeKukJhRg2roXYUOU94kAoZs7l/Pv1ZjIv2+vxcXG
ps6cHuHqaZotRReWPvYkNmu0481ktfGCfFRy84TNAOq8AIw2o1jZys8voAzrbGyccZmEa6LV4gNB
an276qNnLYkGroOU10k4S6u6T+DRq2MYFBrVSDWRxReyUKO2t5BV1LX/hJPdDtxXTPQrPoPoSVHF
22AxeskIWS+WWCsYSaS7fOYnfhN82CECx2rGm3jWRWgBN2zVnhhDLfbdUk/iLZ752rgMrO5Idvpb
3YAOWEj3TpCY6uTKG/Qw15Ib+IcuD4BZYZEpVoUnAvnkwjk+AlYe6/Gea+EnD1sRiwnrbY30xqi8
PxTz/3pa10xRlESpiunP0ain0Be3xnVhpCn+B/AtUybCgk9dVtNwrXsqYFMmg+GmrtcBpFq6kj7d
uo7IY5agHfvQd9sqqls9LXDwQeP/thCyQQbUglWjZR7UTPk/mG3ik7izpnaD7WODYTOCG1hcyuCg
nOnDG9Dn0gf9gQS1OQEjSQclwbrQuptRPJD7uvqANtiNXTad3q6ahrGyRDssPZqp6z29CJsIcLge
2I4Cn+luAFPbBFVqLe052BA1dft+nicJTWeF22LASrMvEZkfnf5+TqDQ7aC+1VM15RCh4wVAAkWT
VoZWfoDmRcRPm0sT2mkbtkqDRlO1qfKhRqjfQh2vZNA/JOc93J9GA5PiasJOx96MD1b2zG12W8PE
D3DkT36Jskwk+bVaiuR4bLMkyQSqbiO59KL9R5002wwNgrTL0UVBSZQMNCESF7jbg6f8OSNI4nkJ
41f6vc+bZU7EiDjIxK+cRky/uPnOMYYNS2CVDeTGOPfnxRCJ05SVTk3n5pejDkpSQLpKjRNm9jWN
ry1rLmJpc1U9/t6e7/TBuIpzeSLf7RB6hh62hrQYecb05eOywcmMSEuuo2Ty6EbASqogprGtRsap
7RFNpDqqRUFSTK8OqCDmawFpBsn4yjh9CKOumepy2NG4qTLup14nxRqXWgp9IekeMV1H3ii6UmfN
uHbKT2mAxH0N5jd/mih2MTka7IyptqM8Yn44OFPB0Fsgfmbg2M6dOdX+/zqEVW+9/ZklOo6IadOI
t+UUDYKCERu+mr1zeliOlOWJ5OuaM4m1m4z/f/QgU23vXJTTclByRjfu+vRlUVdQ8yHCLkFp9vVC
euWphviX/GuqmynFoWOUgcjweTQq+/v9EdW0iiNqXTo6zmafJVUMcaSxj1VHf/Ov8xYVdoDsbi22
1PFLB3CWYNZHWR+rFIYuaeL5eT8xXMFP7hXdTtNnRI+nk7LMVNl2J7oAHIo1WfRrbXb88yah/2OP
u0mlwsod+blEFigjAgNs+/74ZSDruoplRZQpulGrFNVsDPGzitOBFOh2mrFLBEugfHv30EI1qZHv
hh9F9DTZBxsAKB9XhEjBDhugVnyDIwpCSHpRH4dAG5R4Uw7x1J/dzkZiXoGqUjBSgz4V1mG95hC8
vRimfHDVZIpNb4LWL2WdS9c7/twjwLPOHLwRZv8mKfU4rSwPRl2wSR1DmdmP3PoXEtYPisPqu+Fo
Yn9DiACo6cfQoMW3v1/O9+Nq01UnNVXW2JyNS3xZfXk3+Q1mSqxkBGYGluK0IpFcDFSkmoZDPRPR
AJVmKw83oWrs7djirjiNvTgfTRoe9uNq/JBkPPvuImROZclNlWDCZjn65iasav8Hidp/xniyqA3o
AcYXKqYVhqEQ5x43HfDLMZ7LauxbC9MyGrOGoOCrT5b0Hp2yZmdrPHyRTQHuyKUC29UfAPrFimU1
lQN7+OBg47wNLWCtXaVoCAufSY+wzo004mTmBgjBZB05wwW4DXF6eLynmndV1wVvxea+2MTVRstR
rsmB0MJw38YQxS5uJUe68rtaw+aNE+6hgOOMTw2mobuX6/3c5wIoLZQcxGKcT0sQjCskNWXQL+5d
BZRA3D0My+N/XoDp62FIV0p1YB+TpiHJ2/ikEh9x91VglXJai8hnJqGIQPNaSEf+RunXYxn2QMCG
bvLjW3e+wNED5C6pGVt/QNDR08wKqhkl44cVHaOTAESnJRWs8p805sPJlPyPgCoGwHAFLs1tYCpI
DCCu3WMcs+cHVPzYOwB/CBiV6YNjz1zgcPTPe1JkS5IV/Fp1dzsypRxNfI/UZIsWjikaaJVTVIYT
qa+VKIBh06OpPBnRekxobEnXwWMyDIX9XK+7a+wMQRaeHSe2JxJRueyMsz6CCMHlE3KrdGE/jTTo
9BC4P5O5hdBF5RdQ4utFAqVqYrZDWYQMLt1nZkJ3rgyk/NqS/s4qkAP7e9TrvlHhTDAE2d6JiSIu
gPg3HQsNYcobV5gULys3lHsIBzV9NxeUzr5gMGLNU42hmRESoKIy0tOJeB2XsKuYtM1QND4ZnI8U
U+P5ilojW/kcheQqmJxm17Kb9zFR4I8Dh0E97Jknrk9Vh7/SAxSR3PuJ+5bBzPnynP4f/fOWGQFT
OI92OG9UHg5ZUoFpbLUtbaadut9eBH6sraK1txjAAXB4Cq1y/GMwZm27a9TBp0sMEc454ImCsIkX
osDI+EtT0/OVRN0WuilbSEUHYEmKdUNbLGn/OUhCCgDSM9pT6C8H53NFOcSmd1I0L+9B4Os4GIOW
ESYyKpCl11IGPw1jaI0t+PUchnueVFEbrlDjeJI2VkqgE16KmqF2SMi02Shk3uWgE6GIfvccHFcq
kDuWsCSMJi+117WRuqUaqN5KRz+pL3EPrqdz53utJLIbtn0YQM8YNzbBNG4FdEJXcpeZNsUuAzft
zcIvYlN38ldWmAH25U1b1q+4bCACzcNMJNFV7aH5dfvLS4QvcB5ki+7w9yirVKvzuvtoCHoXqhwW
Oj3j0eIdE3NN21TAAcOsrjI+ob1F7sNXXrPsGyixbY21hJkPovSCcP/t5VzeyX2jr2YciwJ7dJF9
I5rcVU1lVHVGHGbOEfQNnIZslovCUDBoEU8Hnfwqj2pubyBKbK9Q9x+l1fomWoTG5vc3L+fBDm0X
r9yr6fO56mrTW8/x1I9obFtcd8PIy3ICTwKHieXXgtT2IvjrHrQPr/mhIENFYwld5N8r+CgQbE3J
1ODrFtMuzNhzEsjWnYeupH2+69ZIFEAa/Jzwg3ANiMRnLMuBwh1jvRjiC3rddprDyMKhv1PeCBzr
uyBw39It3LmACWf+cv/L8rqqsy+GFKPqaCgSgvfYV6TkmEGMtP70x9gba+qOJoqJocmUwmTJaaMd
ayw3Zfv0z+Au+mRcuqgXkI18vAL7doVHA9vfBN2pXpwmsX1dKeVI7AtYsgZ+kDXZEJVDzWFSNbxf
tzH3j3nQ2mu5vOsFAxvrlRGsxPixxqW/WfNFE/JCe9YV81H0V6nDbKuYZxHgiGsaxSuhw653nbDf
/GQuhdJeLHk4ZzChOHrkLJmzAgQ/EA2Qqq4Q4HlgO9oM/tUZCMRQVeIh41cOcWNWAxSJ7XG89L1c
1GORSAbEhRQ42nOkiao6DD5eAuScbOvKjZbmnQFdT3fLOxY2ip8qmDfCGifQZBAL1YBzJWajrlKP
ca8LMe4RBAZT3C5/WQwwQI0L0R9mFf4C3o0/8kjxjgIdGGbq+L28PvykIeNpwZLHca0l+/11HRVn
R7lwWSwna+8EAlYz9veJRogTZ8eFDk2bLqaRoY+eyGX4oy+EEtbeQooR4eJZ8gvp6uSp16exY0Z+
RXhANOVRuaI6vWOykYQz/3t/mTx0VvP4zUycXNdwrDGufRRFaSpeM9xcUlJ7AX3WN7CVHfI3MyTR
a33grTRe0IupAGWG7Fg2CVUmqLxTKixT4/fmjXTb0nJkDkG/5aoJwvR2UErjm2OL86/1o8gBD99T
bO89m0ThZl/Yoz0E7flcJeDFYgwNM2l2ypP98geIGLnF4RMPEpuJn+uTu9eg6GIynUwP8Mm7Cit8
7WuJiVTwLyk+ke8jXI9Spr6ojW86KruCglm4/scaZzIgpljn+APmPD6ACyT7/6CbGXT13Ql+TM72
nZkO4I/SPLUyVZLfgDm6TyYSkbe9dW2BPvKRewDloFWPWXRYSu8FqPTfK0IjfYLJagwMXGX8RDPC
f0ZCPY+yqTPO+JaVEWkjljEVbCbQhalgk5XmVMAFfkLnHjJQm2aAGts6q9wZ8IvTwg3/0BWVD5SV
Tl/dYOU4PLDnPi+dVE4gCrHDjLoBDfirQYaNkfBOFJCjtPTjFAXnQYeVqn95jkunEwOmRDA62Sv7
ssADPVi7lHYZtZ4m6V/X3imiiptd5AMgdypHAbWePt3BCWHJNhFRwU80DjF7tQWv45eXCEQoLN0h
0DHj9g9PLjCf4GU41gj/hPJq2zJQh374n8+uKhN/scK5tK8xp/KZLgtNJagqK6XcMY6GXiIDLFK8
MVHM5x9PfN7sAyQ7SJkeoFyHI0U2XUvxm5PS9QM40BS0dw+K43O/l00El7uy8peFTNTEYGTX42z+
U9c41AL9jy5jPAd486WDJXb0HDJJtD3tcKADVvIue+s0D1g+782Zb3tO4R511vfCGf+37hODs2r0
nbOxSVFYmtuMYkT19fdOwf172aY/u6p91iqMK9pc5ClIytXNxKuq9S43hhh3MOVa11w3EKcNUl1X
XQxEu8po21dQ+GmYEv8iouVSWSBQlhUAI1GUYZEYeHzEiYOGz4d9zy9TVoWRVs9r8Ouia1+Z6K9u
pmxu6OlowPNVbCjrowstjSzg55Pz31wrQ6I2jylX1pkQZmuMjtyLKHPU+Uu+V1hReI9Cc2lIC5iQ
p1a9078F24zML1ICse6KyXBq2kGSyysnP6nYq205i/nAyruAJWAZAr7nuGhsU27knNZTWdgoAQTM
+g8kZVREYaBw6fhOVVduct4cYV16JBxi05jhEwFUzCMJz4RN2zHjjSOnfTn8ujtRAWKNoSrc7T4C
ZlPygdu+zZNLfqtfB201LGC0AgDxc24iLKUeMk60ojloitfEtrseBWOr10yUN+g3qQLz4sHkoIpe
e96LtnVHzXHfScdeF6OHkWxbqFXG5gmNW9XIytOoTXFlwfBYriFKry2s3YJmLe7wUoNmlLSoPZLm
HQX8zFu6z97Q2VprYzp+DkylRdBEWCNVgp6GWM1oln5gYcUPVUmeK6sattSmyH4N/jdbSyfFPqru
95kzzCO8nxbfzw4rgeR9GRZbvelz8z33hBCKkyWUkD3bgso20niOWSD00iMYo2YxRlB3ZxMcZPdC
hj0FO8GNzy7KG7AGUyLqwxV7X6sl9L8GKB9cmghuLfJEIqGPdr5pSrn9r8CVMDhhx3rYSiU4wjyO
wuh7L4XKBxngIbFcuJBu14NiX1x/lswV7owumh4u6hIyFCFAb5ztnCmzsKGRJ8ReM8+2HJwxYUra
GglFVxzNzGTI6iw1Xt0ukL5o3gF8xbjQesc0fVdVGc7u+KtAyfvJwtz962ME85Vg7+koNdxEErDZ
odEGMHaJPnkq9ehf4D8o77HhqJ06da/t/q4wSbdB3fVRcFjmZLApJC2/rKw/Oppu40qjlMw5DYHZ
/mP3Rc0SKviVu+LqYLXDwx/EZw8zZEMGkLFf311h+w+CwU+H3hPgcP3C3O4kHxJyb9WOCt1wRyiE
CigIFULQTnBvyhUXTLvnZ9tKt42MQ6XUO8saM/ODnu8SWJCJmtDKiMARKIOIdspgTvToqVNFElUN
ng3RTTggCMP3D0G1Fk1c8yl80KqMcfr/yN2T+LhvUGJU9jmw/NWkC0Kjuo8lHziXWq9MH5+lb4nE
rULBGwzelKFDx5Um5I8lo9kZ7wjANL1t+foVpD8tRDB62VRYUP5xhbDpnqyu4k+W+5VA7osbKwvr
Z+94tRUygbjbjDBlY78GpU5AzhV9LTxZzjdVKL0kShLtPCB+38IzjBawn6iSK4bG+vPgOKQhRoN2
lsDALPJ/UZMTJwvezplKcPZ0aNWW1kV9IP/2c28T1679Kje7u7EJTSS3+sp9NVp8FmQ1ltARa3Vr
iQ1fs9S+i2S2H971LUCU0ITwOMT7NCzQCXHilOtik3Vekt/zmy0opp6Qwzn7UFSOBqclW4faUt4l
54h7Fqw/mIWGTs9cEfdGl8GnpttQ82vHRWSFSL0r9XvRxub+Z83XIn15fqH6cpCnTtpuE8Ke6E37
UJqH3/fZizkIJBpcYnBiCAmeiaA6A36hlZ3Jbma4686ri25B0SOXMS9eeBlcGKf+T4ER85SO7h9h
fe2dYfdUwn59wROONNtMyYHjsD3zwvpytj+KCFqDILet0KBFVv+bb0xcFTrb7oa6ZNxGUxGfFhAc
zjxMaqYXDaWWIJmbKKTO313sNpkG5XinLJFGwTABNkNtusrpRXc0Q6lB9+mnqBneG8xjS27537In
JBjjwH+lOtJ1+SBznzY/5gL/JGWv3HbsbB+xSBRK5YznSOLcj0v/RbJKQ8maLQ38nQ22npI6XHsD
oUVkz4S9rgD1H9gVjGaKn24fenPK+C4MGDfe14n6ZJJSEDRiva6gjCBqezLrBwUgw76dVd6mnS0W
Rf5QRYUJg4XA3B4v1tNDuZHJYNenvGI0fnba7y1XNWu4o6CDrIMij6gfZjqUnDaCH+/94BWJQT6b
m4y/oglUrB03oiZ04oDiHek0UAfbEXqnT0VclaGm9dDba+kRlBJiePuFk9s1dZptfHeFz5uvaxpZ
aRFn11iStXH5khsBJOTtVkiVPQgb0ifC3ykUDTx+NPM4OdtytedgMb+/EwXCDYozvvlttvvls4PY
TZYzkUBYOf4FTNrM4h2Rt8Fi+GX+JlNntlvjBxjEyHaHUN9HRPJMyZUrXm1Ftrv/GR5e9ZFQonpW
eEllDezqYAsopdCa7zPgHzlJriie1OEBA1b6QCGYW+MWmW73SAo4TnYUjSeVfsAT2+5P7Up5EZnv
y0bKCCu/D7evAiIZGl8QrDs5Av+TWYbnkMK8l+KZwSK1ydCSrrH07ZOIonpKoXsmRCGms/i81o+p
nelVOGzEL3AUcSnxqlr3zQwC7DElp92+dl7BZHHLLhyrWHijbgCZlft1oklVt81oV5PJyjdOM+ym
/W+MpHTjaoJUudJepwjadAD3/ZwKwiMupsrggpt+YRBifunsQP+BzzcZWmma0k/BQt4I507pbHvi
Bw57nBBKIsvkaQ97Ofar92tTP/51jeBRvyDvpWAnYKHiKorpBiJjk/xGdbbWsFxS1aqCZKClipXQ
ZxHqDFGKvtlBOBTux1mQhWgovQ+W6PI8Y56cumrknFOIZn6qU6BFqKDxrKEqCoLo3LH1xoP7qscA
Ytz+r6Hy97PPcgaSsO7JdPXd7/so4YNM6tp/eOzf38bNWb3b1YtXKrpMQnrP0fxG1hvf9kwGhTCq
AiSY3riKWVlCru2hsdkG+SsQuO7UGtWL+3UVTu0qXmWZ/GbzuudZLkjUaJhTbto1uuZrwzrsS/K4
FSurHndXaxN+Mo+k4kXRJ9T+ML5S3sl56YCsAL2TpMiEG1p4Pydh8gGNrDvTYn0AIt/PUWf+6HRd
oFcfS3KA3uuYylT8QGNHiTb0kP1gnWWAOC4yj8V+Z5yxJDAWTEjJmoOadx0U66tHK1g6HqqPe/v0
tmomGWGT6w2wueKQsDjoPKwlp14IbVGFJU6RWSs1MGylx7yrKaUMT6Myzzi3cKiB7HnT1KEEwIUQ
Ut5cL2ogPK4YSf4vgnYKV+Ne7Zx3yaFWefC0+SncJ/5RPsYaW+n0gC25eGvglyiLjWI2ClZ3yfSZ
0ygvbSRzGc9BNnxyKqOgII8xXrW57ux/5skNxre4hMKzA1u/JDoi3PWKmYGteNhrokPDr6rqyFEK
jpdoK+PMhvF21q3Iquobp+bhgx03eqqez/nfbx5/WmfFnb9qmC/mGcQMsctgry8egj+aUIvNlyyF
RjuVbtSNen3Rhk99NUE6Lcwjnn9Upzm8TFHRLgN5nKEyCrSKgbeqP2A71znsYw8skp/hUyIUqkP6
RT5qEGjo5iUM0ITpYbilJ40N3aJ+/oc6S8OXdYwGykmJp9XunPC9TdiCfyt4N+W3Bze9+cggwoYu
Ofya4qYGg1MPNPQKFht/HKI+1QaMDedy1XWvsLnO2Nmhw/evmj3Pe9Ws/edx0mFCKlO/1KQJ3L0y
Z81/zW26GlMP4k+y4heWguRtIPYgKFbt7kR9dE12RITiuNVZiIHClQsYUzaF6zbz3Yhj1VadDjPx
QopNYYiczKKoS8sQf63Vqv+n6KFauKA62UK/oOJo9RDbgQiT28bDA81af/p0XE7zGOdzVIwbnqo5
tU6uhxIyk2stuRc6pkv3l3k56y+wo80gC1sus1R/JhJc/AAbj32cilTUcA8cbTdeMtuYj/e602n8
xH0F5YJ99nPcWhFzvZ95p7iXKYgNHTHHm+rkAeFCucAQfvcSlESlpvhkjcUJAPA4I7KC7mk8Toju
kEKj8/wA8saNjZYpdscjrqciq/iUD55S5KWX9yvhSreMS8oyKsFNInJMaQ4bfvJt6FaQR57uljnS
LBr1AYv9JCdyJyY/KkrT1+sGI57I2+qHG96oqjnIC5ZXrltPRQi76rT0QZn9rw7isgHTR6t9onHa
8Kdp/+pkCaPh+UOHRIkIeEohYm4PXfPXqBz3Acxe3ODH+IOXInyZX9jImqeTIehT3bJNBiD/Qj/T
VcVNx0qoTwIlc07FX+tYwOLZyxuSbmbi3Jo2mrbnbP3pP2PBnflX/Sg+l1QOUVRd8pjhY3P+mjTa
EFALFjlEPly4CFT0j1wcyiPgwdWptzwF07QCjrMTVEC06OStrt/zDTcdx+pzkB4Cg8nVxENsgKvZ
dqSpvL9SL0NsbTf5ynZ64yJW48TOuFq4NXAqmFEpfVuKXWYEZxB4wNgBlWNY14aCzd2B/zV9a7yE
atu5utUDUhdNFzDetT/FBXdqOjoiSJigyJSuf6itxv0ZTLhfrBdQpcGO2dzmVJt4aeFm7KCmcqyo
Osnld/Pe5KFaxcN/U9i3Y2lH2dlR7KIJYORnaq2q7HhfQVc6sbkuVqQCNHqZErOICfQfWew/W9FA
dz9KVa0KyUMlb/Cd551sSdg9qrIqxLzi50tstHOKooJdx6QTGdaxlMvT5ZmGzTsibCjG2jH96IeC
j1+pw8h+SguthxgIfFRXXL4Z69OBWVH1281gzApqfAG1+nBZGh+Q1Vf+j+XzFVsnAr/tuReGY8IQ
zA1oXck/+T1AmEfZqpRK8HUvaK2h8vKCqo3IPcIKW0YgYZ1QsZpbjdVwReNz1go/gOGl6g4j+q70
2kv7iChIuV76SdMqEKWx0v6IdLztZpGpLQUkClaD2e5mk+Rv/s/wcgbD3y6Kdu0+5BVK/NYLwjVa
HLYp8s4zTupJnTa7PtKyrWetAwVwn1YyV+CZEFe7ogruzaE2R/NwVthqjoznTejr5xArG3wlL9kT
PhW2bgFX9XmfRFY41+oynXAjn7iPFWpE68kVun0RQsnx906FR7i3t3JEtIUwHNvHFSaK1Sv8qRCg
I7g6B4XhK/b8r+dLa9tAkJOKz5UED7n9LZ3+Y8ZbCLVMZslFPpdWwuQAWdiIJdIr3gC0wHWbOejp
H/PCwBKOuA/O+WksDFvA4LLwzBj1meFC6NJplgq7UeVvqqjysUn0GK+BXrSEeRPyZSVqlHSHtBiC
rq/gY6SESqlcqio8BFvxcx2zIXbZ6TrjXoLos8zx7Sxd8TnGApA4wNVXaQ7qOgXB+2G1mOp+DAa1
BPhq1dlMtJ9mDWxEDtlFJ35EI4hk3XFy/Hm4UVr3XlitDg2xmVmSd3n9YjUrOnxQYw8b+fkSLidy
hpSxuT03B+gH1DiEl3A6QCaFdQ7KsmseH6oEC2kstN23XvUH1YIIp8tEfd6UqPojeDOfGGFlO1A7
CJSqk9Au6E4hHkVj0doRKXBSTt+LUHozigBMwL7mzJuVHKw+DegzfUvaJ4hOxjELiGSoDcqARZUB
F8ujfQ59+V/UbvQFjZhBBXzc552cFXfYID6QOUlsPCAJCPodSKVJWhOOlKOa08rM3DShWMubuQ/u
a1ithfh5OH1Nal885JBAJHcy4Ncl5W4kg2OIUz4yslM+6MxcIIelceRhUgm2ecid35sseTLh9gbO
5yJMUmrJ0gZmAksR93YUby8+zgIrV6vMWy3AgYLkUKeLayKUZ9d/Rw6meuJOe0EED91BTpcebEiU
BJ8TTuxGYRiTv/6v0xN5MAx8HodLc8yif/Y2cBk4Lx4cdi+KwIAxEa5yqYWEvhuxZ0rHNsX6JEZq
XqmDD3dX7CXgD4kLrgqIoJT/uXiaIyYHvmzjieVoctD3G9oFBMm4baASXe7lBf8KXNlbR6uzisNX
LEsqHC865Osgf2pQrFgl1kNTGetXSBzj+laTAnxOOiBtzn+TJCCSuIqCz1fkIvwZppYkQep2uvII
dKYRJ+GAvgSK1n55vcI7/zqsKLrYHq79L4dhPwu/ndWHfz4nenDJ408VMs47caoEi1ElhQTOcY3p
ci2+3C0QOYF3UNGoY94v3tdLl6FG9Wmnc9+/Iysl54WXe+Z6O3/w0NaemgetOgDStE/4ogwkVZAU
KEZY9UCabE2SqzRT82L3SsHcY0GQO847c5/azbd+Tdkw8k/FKr7YRyZIBtDFFIG6CJeRxVR23ipc
EfPmFEMiSt1U5/RqD+xdQ3xrA3RO4Ka8kTHBi7pJFbaGL8TAMviiC2scfGlWlExkYCrS86zXZXs+
LNfhg6nq44y1cioSFS3VKmQ4st1mQwJSKQ7IdF8mamCYgoDq8vScxjXrfoDK5eMujevgrUV8HDz3
Py26gjWak96lHoPvYjQEgjfraYQgee6zdA05Pu+b6+KouhvrBFP/ArcZ6imab5KrmFoJRKZYkTng
o/Fjj90GdYvTp/abxp0H0FgCqH9nVWpIXXmIVqF+kHw75Ix3Xv5FtXuwHYRF800TpzTvs46IRjpF
8df6KPbg7C1MREzIaa4wEaYBJH1io2hu5y1oacVeeHRlyeEh9obS6D42Sl1iNIms8LDJ1OHxYBdK
UaLElN6Tpr1ZMXFAzVInRSdpxgaOnAkS9Tv+mgaqduc3L0mwRejg0BM3u7C2xhciUdFNMwlboBWY
dVkLvfKCh6MHWoQJQFli+GONI/P2oi4oFDvrTFvGeQHXM1kmp1bYhs1kc0PdTNnlkiGSlmftqc2Z
MLWsrWGbHivexZ474MbIg8TnDTtIHHueR7oewg7FRk6XpOoEJqOnKbGYy5daN9Jv31V3NYzjCOfd
d9N3AMgdiF4uMBKSaf/+z0tvzn0L0DE/OYRzeux7AtbFTN3fsbTsrbJFkTcg8LyNjiV5EQ7AYPnH
fV74I+2PUlCv/57eSiFXsD/g2lYSOP00BCSvSq7kYQnIqtPWnnHRvauRgY2XX/GRQfi7NqkAIbfk
1PtYTFYZitv6TXT7sCamNjTp216IU/yvnKZXGV/DaVHornY30eIw/+E5B8NtEUC7lUbsdOsWQ/HY
1PdJoDPG65cE0DKfeLB2Cds214TmAqOS0nbLicBdEP4qP3uoOGlnfYkoN2M3BB8v6maSjP/bqBzY
P6iJlTO8xMClBYnI/nZ28b3PwujODL2qF6hi23wtadYImF/d8mGwDj8v9uMUAVmM2MU4k3k/DFvt
ubZTFlCWImHoJYlTwQo7Rboh/FsMFh4CwmVyXy1/Fz+qo4fEfbEmm7ruAQtzYtKmaD2QehEOeyKI
Jv2zHRrYCHDkN66pmALprDIM0na8mk8mDUEMpscEixKaBZe6jwMZk794yO7xBrZkJVCCNxbNTV5Z
F8t38zIt73/yZlfZ6keUnkpW97A78omr2UfN8rivgzL5npSOccKZ/QVgKuAeplhH64RP2IR1pTJ7
ZMn5AuA+Fn46P4x9y3KwDfJkNdvIxnbLWaXDpSc4phw7gZ2+/q2Ws8nJ3PX8lp5+yytiq/E1npdW
QEXQpJk00lUuTeCisJPvQlZnDtkwxHY505Ezg7eFnw8P+RjTe15sDjs9JszFaks7bQS74i3h14xz
f11PR2EV19sfRNJXLNV7lAnLYBt2Kf9qu8I+DHBa7vGJ54cbGab93BIixjouiw1F9eWzZ9ZOtm5S
eEHV47hF2YaXiI7h5TMnZr11x/ygSayEMTFngTsWc1ZHMzDJa0oMnhDu0JWuu0zLeiklbLVVkM7W
R5JT/GkXflVfm4S0dN6rOyoepJcRU41cpOknEJQzuxG3vb0sxwWvM2vrmF8J8AE2DbfyaUuESv0G
Rq7Krh8v1CKep2Z0xde3q76Xqru+Tww0xYghsHHzNvQmyxx9aOBAVbbLv6l9GHp1NV+MK9deWCJ2
kCk/25CHVLZVnlTj43AQrrVhmwY0wFsfGiLL/v4Xxv53f8XYkuazv3k+qbc4+VA7EASI/AtTXCsw
Pc2hnO7X66+9nPe3Rh5Gi707H8Aaqax/NM/QtMf5jw2Vp2+qY2U2okF+F8ul6OhG9t026D7+Lmuh
omLp3qMzdG7h9MIrCpOG1jg1bRn6lkdSM/FYSlTPmpikPoZIbFW2xoPYcYFm36OiqDkFVgB34gqx
ClcsPQ7aPIlzsI0NeB/LNbIYZ+/njpIejjswLYh/pKhZDlbhR9OUPX8QEB9iStRL3DWX+SYuosRe
qUgXqWKBvRpMA2jt1jcyXWw4/VobzwOdZ/XkPHRJHkTfYKSYI4+KD9dVzLjDdDLtnA9P0417UGzY
h7Ft6iLaPHekRTQBuV/O0yhtNZWBw09Yn1KLlExT17DdM9a8Qif264H3tUSj1TfU7t8p8JrCWH8r
NBQzGBw3MKjxqaf/WK+oTCxnUcoyLOVJzs0TQLZ7/3Dsn3HeBlTcqRFeZ7qQ3zZFXjjSVKegdCVb
Zc9f6cu0W3I6XeATAP4Ccy3Re0YHpQNxt1BW19BIKDGk7syoTHbT7qccT1o7X/zkDix/bWmurf0D
KTtsFN93VnPO8zJYcNxW1GZZkLJG3NcQWgdvItaffmSExwm2ll6lJM34Wv/NSmgs33YW4uGe31gI
pOnKEIQ/nULnlVwP0oGK5qjhzI7HtH/AkWqsnujUHDqcsEbwYI1TcteZfDY7+x+EFhKKzjosGLNr
a3LevnPnhU4RB+uxsr/9rMoAakreMCX/9bh3GGTf7uSo4XJ+A8EeOildP36uePnnqrj2pNcV7vJJ
Q/IhnvtDTZL4s4Cap+9ZN+2cSI9ccHjR//Q9fj9ZSmMYUbTpSpXKw55VsDw64ZATYqhl5HoUMJla
erMtgMYAUsTHtyfCKkNUPnp+fTLFbsfhFzudT785JMFBhQ84YmDFH6y2gchelri4UZdHgsRfoNEC
sK+aKwYyZ8Q9TnsJ69lRjWD400OXidcNL5xA+evT0rKJT5tvhpfJPrZBcr8W92PhWhIeocUiV6r7
1GvRJiTTEfar26h9C4GMiGKup7h1A+p/CRGm+Ly+oHmeZl+UOClD9Z9RnJ6lyDs0MTPFtjCBJKzv
Zq4ULH5occ8LTIkJWAns7D+NA+3YkaH1URI4st810ke9N5nSe4QtmPfrRs9h6IB5F3DHeHpAcAdg
ymDCq/Ky4r+yyhTJJBQ6wc+hCHo2HF8S4EsUcbLXql8xNXlFJPxQdzorRKcuBLu6R6TeM7gdDLBo
oWK3r4L5kOLh3YApAUpq8r9QnpAkUXQ7Tdu8MT5pvHsMBTI/oGAvCc+3ZDKgR9tlEgKVBYGuSdkR
vvVOOSBE4ht8SrWph3DajFaCvgEFC1Nhs2f4IuqS1WiNNe1FKEsYBQ5Lx8/BOjONXAQL7ea+rsDD
SGXo7fcsAkmrMLoFBianj8+3YRMDY4PouGOsH9PxMiAlKOmHZiz9mAHQ3rJ3lL3GkgNtwllk9V+b
7H1U1NXxrotvEtMDJzVX8GWUlbECdnIkuG3hAp2A/hXE0fd8z+JqO2ZJ1a7F1rtvnyWd4fX/QVSi
CC6crwd7h+6h6XFnXarLVb59sbhnZ+7X9ol90Yml/N3ndVrv+K3I+qTU0tGIiRrBPNYVZtyPUiKJ
q4VMlqAze/oe86WtdawEcgz+mQ7SRZXOwYyg+0fov6DUBFyFi4ghYqqDCGc+q0Ga5+Tb4vGq99ma
xopHLngICqTwTOQ8LryTOccGiU+GWixJsTzqrxflQglqCUbuge8qL/7NoCrb9YkzuO6bVE2fpw7u
WCIi5HNveIuu3+IgX5oHYYrZb13N/tz9sD5jWSSop72j5TCdqX9FqndzkYxbJSur/81asFYsRHO0
guCxXEzf305hcuGMEkX6UjvLTPnaq/jQGLKrTRvzPReQLiODTRqjRgh8H3xxjTC1SWMq3gr1ki02
22ZMlNuJiJ6gmN9dRMwCF0y5jo5g1X6zPyP2FBJJasosQN7eMfhuTiAucuFeAvnEkuaEQ2BkkIwC
aaIg9gTb5ERG+XzO7K2s6TSiSz2ZUBhmy8BEebk2cf9/i1H56UySJmOllUYl16NU9D0rDjLhGmIs
nkxmurspkuvraI6Lgphp6z56InejP2e8mQXGGShp2IIADm/bFTlx34zwpy9dF/9y+tlE1cgo5ghd
6ZA+70UtyLfkPLdu/mHKf2OkdBbm/xk6Ed/l4TgnVFq8sBML86HCecS2XZGEiHzoJ8KxcuQ9IwN/
I/cwT5IvGXS7r6pYjCYXcRsd3nmmqdAxcZzwk/KTmseIf2ZzmKaDVv/TkvtXn26XbxJD4IcdLwhD
5Yk1S5ztVD2iUv64qTz/NyrH9a8+k3+D1SLouLuuPiyWVzgLf2nVyBcy/K7mZYr+jGlLeSATuyro
Rl4mj5K3/Yu+RHrwSg/1OG9pvdhNhYwYqw0u5RpDR8bVCoHUG71uwkLi1fyjKm6jKTHNzFgWUrcc
xMZOv5il5tDRvY6FpKclrizBrR1lUbeKJfX/Qd90AfwR3i8Z/fI3y+VguCga1xqbTYBG7WmXo2DC
UNzGpNNc6DKeT51oAltdBXw0E1bs8fCGXA/2XV0znLB81h/dtdxB68cZAbxo4i3Zudf7m5kLwKwy
ccamqPvoAGbdxZNqenQDslrLdVIB8T8WAryRRBIMwCHQWcYflGBBJTVlzVekI0Ft25B/iRW4Hr7q
FoRvOsOEtMLpaALRjLQQoGavQzKPlFkUtJTa8esBj+8L5h54wtsI93rjsnYtDx0Icw4P8WUn9d7Q
ZHkljrxdlJbbh2+bWB7uzJKp5jIJ/chQmfK0Qb5K9UB+1KhV6oX6dtrKMyadMpsjMdz1ccX2KMLC
i9KYZ8kEomJU0vRnD1MYZpvkDxtoEW1rt7zD9o6A1OcGtXPrlxFhojfhfamfU15OPzVik7dukK4+
z7AGskcCnlWn1VIU07CfSwP3a7qxV/cVksq7+pWcIX1sgFpzF7e3er53/PwBhayK1cFJXd/DRtXi
0HzK2zLzKQIln0yU0r918n04mS0DpvojzkiSsAwe5dYVEbsrzbXZMB9cWXJNtsCv4SxA9u9kn6Nz
+SSR+fNtFdEPd0Tnb4tyt2SXXVR2gzKlTZ7/qxeqmf6wVzTUPcz6VGgIGHjYICtqGBshYeqs/HxX
YAumgHdt3qw0TPWT6L97gQ7xG+DPB/PGfRZNkl31OJ3UujvtEVBcskHcc7jkkBdU78XdOmx31prB
OCCbRM+sqjlKeATEXZI4XiKtopcWCSHQ/z9aHpFC/96Z79UgltMrR8NugMm2IfHMNY6Xm7m4zKFz
OpmoTU+A7fDGCGMyHLBP21+dOPHkjO1c8iPLCAtQKiyP8tKS5x54Vf/L1ixmxxukGHiTd3WsmsjH
6JBNrQLcEH7QvPe0ea8XWYgvIKvh5B598pntkk/Qep+PYwZ1rAvQpn+q3j89QHgJdiYyTvjfL2rC
T2fY2hWRxxoXo/tpsSFuKdWV1+/eoPtWDo6T55DdqswPtR5ptH495wFVP+Aib3LKVHfMLHmrArhd
MW9/DOQL0hLMd7Wl+M6mZ2RLyB/AlvcrDZkTSwKBsyKQ1YGdaJOOOWL1k2vLsqGqejbDXR98Weoe
IrQ+Qt/tBlvV5lsh14OInVzLEekFPGxm0+yoREI3Pe9TZcmo6yF2T9K9ifDPiN5RRMxOFTrDqTVd
PwoFl1tUTAnUGVAR1QZ8O0ilZ+05dGX9Y1QnCBuDBtVKUSRR5yFzh/V6xPlGOXF/EOxb8tWHWK3O
HyuAXAJwRam6kP5viDixnx+8DAF8DKVs3mhOGvnUYNJgmt2k5/80oqqvfHzGg50NNv1ZX6k86o3A
qLmVDl0sJqV+oHgNT6W6git+wlP6zNGnBsVRIrCFB6tARcf4eY/wq/xVF0wDGZrN6f1SqlXF7h7s
qNAeVaudw1hmYgwwovUPWjNy3sL2u8irj1cJWenmCxNUTzhvW4JHeRULwh71qxBZjYDdJPHEXYb+
AZ70BljCUbYhVopPmm9rlZB8OBXkycfBh6/Fiv+GKbecnWci2ecOwAlBmIK+j7kvn7qHM2aQ+buh
nQ+TJXAWM/LiqRxNLL8cvkHGm5lBPfRSQwsV3Be7mxhTgq5+GGs6TJ485probxbNCBR+pKuitMYn
LLEufw49HUR7j0fXyTyPgz3Ei+5LP2gqZBZ8oyew8JZCbhAhjsJf0PpuD+QFHX+0UmZeHIRV/fS+
akyKO2XC8azhk77hKd+uSjgyAyjDr+ifyRua73Y4FMVhIodXcKNWFwbZUr+OoVD1RU+ut2I9m11b
Mwa82EgEHZ/p51/XlJqlgdU3JVeyRFYkfrRpY9x2fKyiA1cWomW03RIaVWCvUtSPq7QyHpXtNYbB
uzv3pldhcHxdAm2FPIZLkc6KwVhA2Xbp683/C3Lnmdbk2Ec1jnMPNTN5QZ9JhXHATZ9VOnE0efCr
63/lkF2kQ0M7kifxyG8qexI0R+Uzets3qJ0aVmFTpUJ3vtaHGpcTbVQTxetOUc9eU/YRUTmPSBgq
ft8u2H0ctTyZohJNS19lSulQMh886aKAv+q/TkED//Tv9RN15F6HjE619sl1Mro/Uh7XsVJ/LpMX
zGzjJHDTyNmq3vtIKwT+ach/pykO9VgN7RgpqR3ruxfAgKEz5XBqwTU5eFEs3D2bJ6KE/xKoROrU
QFdj9ypJ7/138RQuA2EQXmikvup+2aIfZuDACKOgFARQ6qf165lum1wF9ur0L0xzxCUX42G2Hite
6vGUTj08lN9W2HI5Gq5gv+fwLBVhToyWt5253U5xW4PLHKSzLpaCaU3uGQImnk9lzsPZIBC3c9XX
W9+Cuk3ZMWS8yey0iMTWtjd1dPMgClL6zKr+CqMgvapMCuu1DT004KnkbX6PoykBDp2mW7baj8sp
6DLu+ZvRyjivGftLeHyr7IYGQhcABCi2l0yemYeuPYeSJpbXkmN1U6Gob5kj62ZA0/MXKd1QW493
C3xgZ68rfZJTsvfOty3cGQG+wWCDqggfYNVNVdA8m/p63wzTtmmn7LmF+JVTbsXjywBoGhpna+Oh
FANQR0sgtgzucKFQJHFCSBI7KdRYGufXjYkEVmIaxSH1JGxWT003If33m6gkr7pxM/pkb20tUOpk
Ct1XKkcJhCWxlaMKqMAOfUCI7aM/XIYdNmBydPhEwv7kCjuVWKWzla41x3RC3CHOShnUszDC7Peg
ul/fss/370t/lhzZgRdahjnCWJTiqwPC3Q6mSpofIMEIrY8VPdAGhh2OifPNq7+hqalzq9MvRWaa
Jlerhc5NDsZUXno83i1grpHPHaQHm2b8wPEyollM+9nvUXrHHl9f75pvTQMhfqQLpzZvMDPJWkVV
sttrqDM/CBHnHcOSBmIJ/3xNcOXI9kBAXu2AU0jdDNOnK8ak1d8FhuzG3tZL4Wg7Mqkut1Idb/22
xANwBgp7LRm5qbX6sgrGbIHRoym1K17qstsBXTMQmqP7ZMwYA7JZnuLeRRrQIM/fil33X5ekstHf
SKV96I/1XzrfRrPMnKJGwBEYklLbySCwK5qYh1z9r7F2BUjQgQ45NogR3CIkXIO5R4TN02gXDWef
40osEiEXOWRVnztSPjqb857aE+45Cht3dDpZd8yqVHbG6DI4B5I75bp9BeaLU8uRRcwiDEdiPDVy
fivSXI47PmRpEP6+rdSHDyuSgGM/zxssGtUJX54S8NT8MdXU3i2SpAlG9la5/eRz5Moz+hxo1Ci2
FWqa5hB11GNg4uTCf4tspBjak30KXXeT/ZVKduWtx3O2QPPczM36PSAxfXHSdJsmJgOVUftIyuTt
hbVyYS9tXyZ1wb5lttmcOY2Ev/JjgOd/ZZiKyJb9oNoVpH82F5aZ4NfOtQjpN9OLEy9ieVwksw1i
f3vAyBWgHLuq5lD4hlM6IYaSu5qMyp+bNwLw9ySXmeYyKjiT2+xGJBlMFZo7jxcUb/v0AB+VfJvp
pBdPRGHPN0M0YfZiDhX/m0yGvBa6sK9phsmeQZPWUunlzLRif2emUvS89dsw4/Fmu7n6X4FEhHQt
gPh/bd49boMhSTnozDxNRIaQz/Xku0U4dYrAByzXflDFk+Cnb9rScl0SLqFiwiFzOS6iuNpMj6n0
i0ZsjZhgU+OpK2aCy+RHLt5wADmQDdiCY6YerRiX0D6+MOE1DeX527xwOA7iDo6RGLBwcGDcNnqX
la+EnHzyB32+KtzKJR0ftLxawAWHC6sb/5QL2QsMmWmsu+J0tRInahaccHzy9r/v0GmO5EXgt/vy
o2OfGnMV3yAytAFZRnpTPlkIARRuvz0WaeOzGjqAEl0AlwKwjC6kmzgCtWlxwRb6YhLL/JJSv2Z/
i+bmBkXPiRNRwWpH6zqS63+JAfPTaJ5XJkWc/Oo/PsxTAU+4apv/V1yItUrGwPh3+IVlRD1792/L
Ou/qWITm1VCGsdf3XXM9rqEJ7TIwIK0Yp5mPhRzpOVBLHqlpIYx9pqEB2e1B83vb3gmMhw0QTb8Y
vXqGRAxXWD3gTeSIZQMcBiGVVKKIeq+1uMUNvPU698oPsQt+Hlt4IBIxJj/DiosnqxegToKUdzmD
D49v2swjZ9kSkM2u2jbSHl1Ing5rBHnBXZKSVgl5Ec6zod9so+vacA6bzzW7sQnaZWavTZX5lEyU
O+pQD8KE/9prTHl/LNxPbmBBoTViEn7XNfj6kiznY7Nyq2Tej9gb4yUWAaK78Jo2v97iHgi+0vDd
5jNMYXKnw8k4k2NUT0m248eHc0tDi4bUXQESTTRkTqDSUAqkaeH2WOX5ourfhWEFrLkCtnOY/5Ah
CDbHjB5xA5vhhOwIZW8TViINzWlZ3LPqraNkOkM2y9bDCe8XYTZ4je7huFDxf5InNOye9JseDP+M
88IYTINZ1ocUG0thy5uEeAzS5uVcklZe1LGrxuHG1+Egcngy4zCTRcYdV5WD9jkGpGvPE/T6DLU9
pJkIEjgUh5XnBh42zCl8Vj5qn/Ab+6V5kizYyoVOCUQ88hYhZUZuqAm53McxN9RLHxXG+VWiXCf4
BnHjjPXPcWlhdX7JKAnH4fK5Te+NDDoQ6Ebmz7yEOjsJPRX3whvnAqluxKyhVmHXQCzDzN/4gHzv
zs+O0obm3ibS0QOqtOnw+O5aJ10Jrv2fY12nSsw35rFJVXahFXaU+QcCEdtJ70UpfFHMCFQeJ5ny
M6/o7k6G/crsOUEU5E8wHL+Ztj8GC7N5ST7MzqlsvNjKFQpstLZ7xtnT4uT5YwkfW+JK8xbG6VGu
neYlpmkRfpzfcLX5PKnBP5Lj+mY6mB675HCcLtUfOxTvOQabGNIzEEMSHlNFm3QznEzIN3zBNkfS
JrVKSGp28YFqbD4MAKTiRoXIGxc5ZHoGg0/9rOxFKLscoq3y8bbGFp+KWTttMCBtnfmrpfEYUbni
ES2L7ghKxf/MEtOgok7ODuGMi7rEU2uECD/7Kby+nDgZCTwLLcni1jcv+xApliXRYvzMR7jOPnQn
7YpEMGdfsnhJnYc6/AZyHXiXmnTDP5ozHs2uvokmkg7aCGy3Iyef+AYv2e0PsxdlIJ5v1n8zXNXv
bz51A0nRxNWMwkVNn89mv0hWTlev95XSH9Xk4x2Kmg6YaA/rml2mMsty2nbZExiXkSCN9z0OnIp6
fZOBIm3gXmaLUqlXIYxlreg/h6vHsMB0dvZBxqv8cIGWgoxNdHTrYi1yKMM7s6djwo402k14K2e5
NjLR+Tj6FhJQ76/+dENQ4eiJoeIRhHUfQvlu8+wX/+OLNVIDTO9sHjRU4YH71ig5iu4DMTH/w6lV
zahBZNk/TxXq1bSYgYZume8hMaey/vJbnOdv0E8ncfvprvoIvx6xNyTu0bUkW2QHuAUp1m90+Z4r
P4h0A5KNYeTBkDIvJk6XZYVKTj4QrMYDm4lg5yhbTlgDoNX4dKY7sL9SLht82L3mWMHYpJMzhtPl
O3NtpVaDHItl4AgdFEDQ850niQ2S2F3WpS8X0NSNubKnFoAlCq62w/xAJhkqR1e2Apg6JiTSaKbN
CBH0P4abB7q4chho+gsNSqonRWKalJUNEJZ71WbZIqG0GOmJD8bVBZ4p+JZhemWsO1DrommPYKK7
AvGnwhDQQJ7fCm0NYE29xXJkEVmb6x6AjjgyUlAY0pBpvhq/tY+2xj+K3+zlSbnOJTz7vXh7syZr
iB+UESRhrKiTHVLA8ktca8f60beJFVlmTWf0Nij0DQEEPGwkrJB1aHzuQdn4LE/KDEBF81fjSz4b
sDW5EbqYSuDE7Byra8t6Jfgk9EDSwvMPhtBm6lwAgkOfOi9/WdE/YdgEP+cKhMIvoo1QEy4FXrMG
QBEa4DBwh9rdTA5pxC5wRRQihf3hxITLvKgJw5bf5L2qe86eMZOY6KlykCPYbPotHqQ/ZyX2e21H
tYuo+WY6Tb7n97/LVaE6zMYeSVzS5Wo6Eo1jI5shIQJEl0D0fYegDkikEkum14Jp77PWGI0Mia3o
1U3fvDF2pHEgeofJsRKdufBACssuxm9fVwjazFB/j8NIrb//38I4SQnVVgVUNLee4qW7cvpv1WJD
OBk/nis8/C+d8z420jWPSgXfPfRqLR1adF4yDICb6BD09yF1Sxk95RzAm1gEKjcMJPuXBeivmtwj
xGyl/jMLofNcLXCWU2OymVAJyhZ2kNp5m/73fcOZS+mkFJU+O4mARXcAklRB1WbNYbTClGU1a+xH
4QaSMnRaKrVc0VDGhHI88IrsOuunDjsEOXPGpoYwqF7iaInBV35/gDSwAEZ1+2og0qzzyn1B6gAk
aek1eqnAtyaQcUwkBtkZ9F6cp/CAeHi27TqbnC+BcyCF26y9YP8Cwpd7/WmSqLCU8RsXRXRwxQff
lw4VvrQd64RNzz2PFSrB9Y47Vn1O8gFr7fvmpACIXYFWFmvz5pn5W8uLPLP882IFjI0Y2sy3a0SS
cg3ZFalyo3VPLacGw5bRIGUNrGybmsqdSNMn+lh0NP0qU97BCieWC4DTEROn+nKtLoflMUwWmYwn
knpTYzQp4PvaUr8B4tC1S3WAFpwmINx+PoSHppL5S1+YAAabne+wn+h3cIlDIRebgN+cCivak7V8
m8r2MJuSD3gXlze0pp3R3Nbezx2sq6b2moeusNfZXH3Y7D7anEHYG2h5sYWT9m9ULovcw1vefLny
69y77e/pilCZuphSi8IaWUnGwWss0J4yE+bbpoXEB5TYFyHS/601qLpUVlONxVRGT0KZVfX11Blm
vpLBKU2mSWcZ3LLGC/n3FTXA6SLKEfGCZLy0pRHU2vSi2tguV4j4dwY+AiaWeXvHy7RJMFri1eWD
OtD+ejw8kyW4HvYN6xbwgFayYjCDD7VLy223agsXis+N4f8+R7BE8dJ34Xe0ya/oj8fTFS8JwrJE
OmcGbXRJ+0DQcVEVfkGAcgxpY4Sdrd3Ji05/NLgbqXYb6q7PEVXhhAn90XWx7T6zYIqYp5r/ywRV
WVOuRuP3cHkPCmuANSNRjwAy07jT0U/lh4TyMDlXZk+6Zj5cxj1k7KyWVik7R9JBr9PlfRMwK9ao
k3wRmZ9hLMCVUw0PWg07W7cUPDRXILL4SbHuMyekRCi2p/KEELqGCISmdenifwwv1wfzIH44CGsR
Ae4X2JuWFCJQ+B1D3FIz/ZtiFsSSFJ5ottUfn/xYEDF6J1C7g523qeH84b2oV091mFIHAOE1TMJL
xJ5SCFim8v6mZqeAJzl6QNN//jBRhPQlrexiUdDVC3SuFJ2lep6RPC4pcNvPLzJoS4toVLAduyX8
/t0MSXZ9cZlqcZI39s6o9qd4O0ggXeBjys2oLjYltrdJzbN3pZFyVXqF8x5CuEwfqsj3bPSzFJ7V
q1nV0pUOw7/LDp+AeN9av1AWqfC38Q+Kzy1rlgp02PUQxupagyfMd8jOhogXEUdVD3ZIZcrNyD33
RIelNscWq6QmXo0zj/Sv5K8r9lpcjp6kcNea6/CXGwwCtLs5tgpCLCtLl87DwC/zFHM1f2grrh8j
9I/JkbvzUBORcyJ0PrTPBV1KZ+PkRE8kz9M2r25xn2voQ7WuJk7SGCvqMnTjWhESYPQ7db3syoLw
5tSsLnCgMOiesn0IpdNdahBERwSqrVcqHMF5EwHAlH+0waM9JhGBh2M7/GR3AapglYJoBKowf3ie
qoE8aCnVZNYWkq+Novyy84FKrn0XBfdyBV2VQJR5nguXK3gnia4Q30mcnHAFqmmeIqFRkVPIzHJZ
ONRT/ZZQOqg4Nx8vmTdT8TnvhVWoU7bEPsx5nVCYb5YbNiqZHIOFHVcuijvuhEogUZg63wvtHxKJ
X8EL9D4CxQ4onRSM9mfi8QIK+hL2mSQsON85Nv7UMx1vz70S62OnP+DGfoCweUaBx41fjsRlSbyQ
2fpBN6YOf/lwc6BBARXNgAR8Qr0N4BGkqL1prgArUlpfmrSFqqBM/LcMcCHH2t3Qn5M5D+kvpEHI
MmUCkzFudYVDKM8FA5xTyV6EZQRm4tNLBizPjVoZsr08T8BwpS3aqGKfgSb8EPxUL2SiLTdGYOCd
7+muQB4BHwuZiQwcuU9q8juBPAHeJIsWnOGROIXEN3ljvl1i72Es2lEgGUTS9frpHFF/0LRyRYox
HQ2wW4W+ZzbgzGnvvMBdZPypRh6MlLjbbq1xpYzXMxQKRslA0gdOehaDZO5Mvyp+3+/YWlvZOu11
Qrx0W0tLCFN1juRd+exJ6dBHrnwrgmhbLFsVTQg5ZOhAXUloubqveb3qWbQMaqyx9vcvX2CEf0VP
ml8UG7t6QDfF9ZROUDRgpprJlqzLxRnmHflVQ2szRPZmxfmAgcO/QcupX9bvDxXTgmxbyei3kvr6
ybAfM2IAFAHkCEGqSRlUlYz0c1GJACukAj7bhOCUiDt1gyLk2DhljTNBUwkTdgzW5cYciwZ2dKSe
CY+LQV8TaH95fpPLAWuMLg4/ioyqCZXSOjqftsFnvQqjw1KtEbJwfOcorRvZ6o+9el2GZTEkISH8
m6R4/09B99uklbZDPb8QCrqk/RyXML6m3am+rMSbkFHciuII10g3/y/RSoDuHEkC1JJDXeEv8Qwa
YPvmCfw7t2C6Bu1pnGDSrUCBS36tY5vPiDEpkiFCMAmwpdJYAdO+qvbdNHbU6V1T0T1BzzGnkMcX
jS2fvVBComPmpxFb/UCcu4bHlNd+H9/unSVZHwpduYtA5R2IziJmWcFAzKQq6qlT0xdfe77QQ92X
wodiehoDHc8a73dP9gf84SkkrBMn5Yt+fsv87BoxjGqLArX7QMseT7lzWyNBnhzWWC8qTJw79ScI
O1StpdOgGu0xuK6z/9SISXymOGrla2W0WAesmOMEmdhyD4w4c2e9+c4W5El2QvQkPIhZn5+1KFzl
e2eHlcjx7E5CVJ39YyUpc/MemDlTc/Slq90HxB6dh6rUA4lQBPDUTG2b42tTFvU/Bl+TQG6/CdbG
y8S20PFZYUPIB0MQaSKtXQNoaS44CPWbPU0DIKbF36Y2LxqCi2gc5Btd3cUgz8lJrZpCzI0Tim1C
359bu1GpXNfl4ruAw0dGdFSxctQ42FtlNqI6iY3H4PXz5uL5jfzDKvUqPEwwMBCOhPm8vL8XkGjF
EjmgaYIeRuYBUlgMB38wdsYxUhHOQPJRgiVV/1dQjbPO9Fu82nu89hHEjEzKppBgMFKIofeOXLSF
Iy3LWF/Eyil5hFlqyYyLGraP7oeo9zG+N9fTNsgXicWkr835HyTYuoNxXvdLvxeyxuvWM4wMD+MZ
91ZBh6IVjqHTC2gtuB4fZqAYUhye2WpI2MWaY3RpSSHqA5z3Slri3MqVyoM209Gw+A0KqjOaoLEE
xkS0Emjb2LA23szOKFsaazzakwuvPvcyvAcAwvBiRiI8nSVEKA7rHWD27nE3T5bpZ0sHDW2hMPyP
c8Z3uTp2d7YXt3xD9+mF1oSwtyME/cPoago34w8HAdMZ3TrWIaWnn1eyvz63EdZykhvklHvRpwv6
GuEXrZK/fxwofuz6jsQww7HEGAYtf2BHpJAj+XqvjwOx9E+L9fK+i6Ze/fb6rYnOSTiTWAZnDkq6
ANJKZnUlszSKtkiAdJYW8faqVSs6CvOuV0bG0x9OY7BxCtuyEePvb04r5I52dWV0I6baoIKCWXZd
QmJC+0p69Pxwe2prJ23LPZBK2vUqoDC9SudYU3M6gCvd/9L0ox6LVpElgm+aHt4YxQGp9U2pEjUy
y0YSeiDjzCrJyBxddIfYNvEBlo/mLTA5lZZspuPkoWgeEiYVz4Ebzekkb+liBPPgpa5CG5G+vHDW
qeK7FgntYCLdj+TFQ/QBd0oJDEpg8LkgZNIJJ4TKeLSv5ksKbVPFwHlk0HA63H+b9pxYZlMQ/oMj
cEGJfUgcIe+MNCBYBM6melELtNmh/9fxlmDspBUa/e5CqwoSgK5oIOMYYmayvISxva8NCIw1x8Ae
6iyRlJ7sGRSuC6D0cfYFTQX1G+9sat5BQvB4/1OG3zngdr9fhZ+EBOA3hZso1L+1LucDSSFYQGtn
Q6m8ftGiHupLLBtwZCbabE6Wm5QXbXM7XxDIhGXNb1xs6mEb+61W8xTdsUXoN8lixBejYBYfIeBw
nj45tPkZvYpRgJO138LjNBGpfdYB39C7sggq8w+SrKleXuFzxJPOKBrZ88Cy65ZDkyVWSYSk5Z4g
jiSBv/3I3GukZenXfyzyWksDqk+RWmRDDg/p7TiIkC6BcpLdNtDpJlJnvOVQB06C0bJcSCLyYtHt
1W2wZkt5MfdNjU69KAjDA+ucUCJzCquyV7SuE9Ab+KcyGaAolquPyWXvpZyztBf0SE0+DN8LFMcE
0D8/KgAtbAALWP9eyfwydYh3js32bSEVZGrc2PmpCO46nwyIGRcAO24XCQrN8bHjv3KBovL5RLhL
RLar7JqY4Im2d/NaI2dzlhMZ4BvnOS5nnrG79R9Ol6Ib6XlfhjRRbDiWQTuxisJdgiBZNX5WeFqG
I2NUNtvzWAfFgruh/rNPLcEOj8lZlePsoKStVW1p4W2bGEKrIvquVdhuqxyEYQmYaoaBJO6cdor5
YYfS9ioRMkdRPM1b+j4efIGujJKwMZf2tgt++ckUFPH1+UgkR31Wpd47Utzw5s00gF+MMNLFpl+w
ujIerSdoY+3ymXSkB3A6IsnYq5A7FSbXSdWAo+hgJ7nPwzrF3WaAzGSywrROcqr9yCEJeNqiV32q
OtpCtP9ZBQZrqCfXesYcEPIiJHJMsiBGU8Lbi64V8i9+z1JGai0QqBRycTdQejGnP3wq2hyxzMbP
nsMkYJ4cx+cpUxIUvqhwmsKhNZ5IJJ14x/mOMlOVi5JyBQ7gsZM+r3XyuhTpRFFvXJc0yEXr/qay
oEIxBhJ81GVHuA1ukYnatoJhpsfiiThoih9jhJURNFHDKr1mOPH8K+VvT0kBpEURdnjrzjy6CqjQ
7qnJFQGuZvuKWf8d0PKTwjZBdc8M/jGRWM1sFf0qZEXC6mdrnV/o4nyfKzVU+ADUsQ4K0MwR3ifq
WPbwxQMzbdthpHpnDS/7OlLZDl3cy/GYoJ2+BhrNd9D0fZSQ0SZBMNS9lDR6djzaTD78+23bPlDG
mvkXQHpMcFbq1zsWpDBaZ3tbSMYyyudC+vd/WpCi6zRwLQR9tWGMsDMxV5lvoFIRwzQSenfgFwIA
e1JZw2PRd99ZuB2g8guZgFzDrcFjiMKnfqI+TuEF+9X68SNGy3FhuOWmQUGpyRdanG40zdZ6NjTp
B1J+H6Y4CaY5qjewYAIV76xGv9JRHTV02AmKQPIiqcMytY00Vjviwt1gbSs7OqctekRYLgDIE5Oh
032WNb38M95jrhl619JweQv7JsPtQ2BdGe+vAsk7iazx0PIjrSPdtH8p+PPlZCF2eEfLIGSR5OZB
baq9jwvzU9ppfSGtTHXKGCHlmzl8QAq+fcKLa/+LKbGez14Ur2cfM1xKFWQBtsYn1xe30mwHdhhm
UaMa3jnFY39YE/zFQjqFJh/AwrU+RiuyaqOwx2ZX6tv5LT4AgP4+1ELlwQbHg6Z/xEukgl5OAGyt
H3q+ZFi0ILCOy0amewGSTS64ZLaf1WaDSmXDFGyWYiPm9x3EbD/HgPWNZ0WeuBiw9h5I1VMyqjPv
wcXSiMwBudxOA/DX8QkOxwW5690muFXwbBM1uggjqAQldYfgIfA+moDbPoXBOwNZEFCgbDECcZbo
JiG90i+ITGVikvgpc7KTPWHV19RNse4dAykZgMf1o/eJWQMYI7sPjRX+ppvwYw/a+avzXl8x3c1J
pppMqSi7mzMLyLl6h+sCpKESLR42wpxUBnCH66o39ZIotjnvLDMPMFMGiTZJFKR2qjshr3X/DbTc
HAAJOQCRfY5vVpB+EutumNu8nz9J9KBPsJ8t0E5136lA0h+LYiNr75+zojPPYUcDPVW2AYNeBBUi
cI8mp1mWg6MBevYi4hxRPXU55frf8BXzKVRTWHS8i37K6FGcDmEOYwKRjevbWQJL5zubBFS6iC09
HDgPQ/L5ZEL02IgwPXuZuiYplRgqCcbUwBE/Qgb0h4+kF5suQMo9izBWGls6jGZm5+KdxeDkCXkS
M5aA87QGQCNofpR0mxmB11S4SHafcXRlY+Hq+sUwNX0EWldSzFiG//TtS1JXwH61BMpGakCecV1p
PGyMxOdsZ36hn4n9oJwrjz5Fyj2TWUxl0onK4Q6TiHexf2EDd4AQ5HxXwUqZp8QokF1wHLarehZL
RccvdxwoP0muAQjIjL64obkAByUuNHFmGO5laHeRlT+SmXBR8E0/I5viFSUJQ7N0Q4h7Pas7+pVJ
7CG9V/cQ2WpiHuwdEjCga0jEAPkNYKJQ0tZn1iWm7GSnr7JRaMApTCBoWOKQ+ty7l+hlxmgW5SZ6
n0296dNdeVspFBE0Es3FyOlaFYR5H8wb5Ff3+gGDWI9UUsVIkmZdT9F74CcbU4D/3WR+71+HhR3D
/FQhJM9DZj/ofnyt5aZqvbzWwvdJr+BEplAM/opBzbreN41richgG8wp7sM9cV/T00tnD+wzhPKJ
+7YIFnOFDBGbWVp3H/itd5m6uIoSgHEwjuU4+G5XpwxdsQi3+2P/K/aJ0F4atl8bGWoMBcKXR9Zu
jfjYsSq3kgTOIah5t26Bi5l617J6/sn7PWbf1wapUW/l1N1w8oFSdiIVX6QRENF/OpbUGEEJwzO6
JG/mI8M3WtdA1MKgFep+RBID04GEBJK8t7XJxabhVGqf7PAAJDZqfZJePyX5r5WxAA86W1ss7n20
rqPDpw7/KRxt/dl1mUNUrj/Vfv/xqlRIlxnAaEG/uN93DSF7sIW5sRnmJZ5xAUSQ65fFhu0H9Ae7
HOTMb9356RMOQNI2oqkmnmZ1I3lJFgXdbr2p6UmuWCAfzDSe630qTx5ZkcraMvY1Nlm8BOs3QLi2
1CnBv3HEPNThWVjf+LMecLdXXvtkOGxyQ1Msl8ATOCoiWoP4L9C1dmDWx7/gtrCtFMNR4AlE6b9g
UU1yb+5co2S7xuNyZVmXuD3SaTOkhX/rJ4Vtf78cFzOQAIM54ZQbXG3JbQryHVap7rBiWMAwdPCh
LtfiVGCd7459t5u1IO7f4plM62fuFHAOs1EDUxSQ0bmAtrWllEk6pdaalFrtxwLEmM/ClVtlMkeE
T3zgAx6LABcVS2BQLz6YsrtneBtq9Sz+M9X5T478NY1kSERMtsJkrXbcL0UD0r0JM/bMfeTp7d0a
+4RHjV1Zyy1w96iZ2YF+AUrbxihTrFCVpmkPQGLJg2Xbwux0eJWCNr2/6ljiB/CQgkU17up7odnX
FOmENbPZ9gLk1TIpIVeQBtAepgk+vZ4tgreuTXYtregpeZQcYu8iduU48mkk1B84bAI63YYc8qbN
tGtZcNEYaKypmxSLZPb3kkzCjkmfmmvt8ql0+zDp0qbRKXyxzN+WX0idRk0Og/yjPqz+VX6wRerG
4IaWUe1UT4CJZimFazcNP/jdHr24aA74ScQFJSytLvp2UuNp69wIt8U9zoecSiqNd5zQEPzlhGWo
nvQmFYCeUel4W2cuQNCL9b+PBj1a1AjXhNb8VwaLhCOH4jph99NUi2OPo3Z0K+jP7bxz3nHWDsG9
aqND2HrvnH+h5816nsOlaSFbEoDtH61lYXl69P9k9zdM75cgSaU2Cpye2vWQ28UK/mpA+MuHf06s
Zy+iQ2gpjx6gidWjViFahoJIqktxobp61nZKtVqz6CLWOyhwHJQm2BNF+S/Q0wnPpG6pMW+bP/P1
s40f+X9kNze7+xYrsaZ2OC2HJo9FV6FQX0C0m0/mzkKoXOiR1wzZh5soJxc5y2PIwuUCcioMowZV
v/400R3oVleXJJtwgPU+dKfMkmdruq0g5p3Ip4AiTX9PGvJr1Y1uT5jdOQUCxC5xyhSiWPbh5r4F
lD09NERWdB74ECngbTFJa3UibjITRmM5rDKTNkE9SP+cXLVjwbwXkqp5FmiA1mN20pz7v1pEs2zs
EwM5MhY0UE+HtEJhK3tIoEdAvnVYkzP+O4l5kHk8BuyLGSAwdBYe1VmuoI87MGeB1SZZobgwEOVR
0YDuWF9UwbT+Np2wsL8q3DFmduhZx6LoF3qRIi2gQLZpio8/MloHV4F/mkxzu7YXfCp6FUSIUzqT
ZrozQXKB8fa6OYAuHqkgtZbNNWIscJuJBrukE6XZhobb5tXQ9MFZdTU+ffPP9uBXKxJ/KNdXv5qz
Rup/WNNjhgGsXwubXAzE1q+XBHkBUQuVZwtsELDsFuMfFo1hiaUioyP87K4uGRyrP0dcXueioNEm
ZrOh4mX5EjUJTpUqok38YV0gBeID3Kg7HqmytiGJvTxoKApggJgk20XW/FdIOnMIweM69Tq+k5EZ
a977epax5qoDY38n3ntqorgyPlNpc6uHnfIqHNiQFjql6qLw6b+ArzVaP+DlfeF9rs4ywTR3KTSK
dLRkQ6kqvVv45FoHURtJNY/NLmNJIVF9tDtvNDn6vFEs/WCMcv3oz1FvPgpF4ejViz/d4gXVHyvQ
8b1s+4QEAkVkrwCC6SpgPKluIN1iYRrAxASRrwf5iOxT2nh7GUAT5tLvkCWft3lG9h0ou2GvYrkE
QFhZBQZ1GqHZjVxQ1dkdbFDr2edh+92IfhAAWNU1YnNBbcI1WP56CzeijuZkpGUha/w0bi6X4ed5
dopC9bhl2co8/oCs59xqX5ofy0PD4/iFJ89B2VoXFX6MLkdXr5ELfQjTRd70maj+VGOdcVU6gm8Y
x9mmF/0ymy9bmlsMDuspqD11wdonRykHuZpxzp0xSEuTOvlqJ7SqiGoCRH90HrusAr2BJA2qLZRq
BO+3Hatdck7T7x63LpylCFfpSXuMueJOzQbmIHYs8Ej8UOeaT6NQXNV/FHS28E/0gguBMZExPSvT
DsHd11oXROnT7v5wtIdjda6u8jLQnWtR8on63rWK3Pe8tIQTHNv8RGwiTjSe/YCseaA2j2MY51k9
omtUWBm7M8qLWrzTnz2DsxjaTrQFp4YR0it4g2pZSaGBU6YBeW+JLk76DE8Ou+agUP5C9fdMDf3x
wL/H026RbzykujGWGjk8X21wbugZNz38nX/Erlbiap1hW5ezRcUXazV283+KSSD/7rgaoXZxfe07
kl2UoMy6Jmt2lYskw1igX+BZs2ElVpmIHpxcSZ2KTUdQO52vEbOF1A1v8TopVGwzMBi9z8hQDq+Q
jTBJp1jofmdctmjvHkCV0MhzAL1qBm8SSAch/Lhtzr50PYUGXY2XkpR2SEcTRsrDLwu4hmvV9cik
dVpj1XwVLM6zFSrmylYHbXpz7WyEOK4cSt3H6xIdm46w3O21lQ+x3M0h3yrQ+Bzdx55VjamOqvBG
Hzms6s1yawvzl+eVvR0eX0zQQXYI/cgLohYqWK8g0CPmbuUsBa4zAW547kM+zIgF87JNaG7y5p/z
4RKWaUB7/yQJAOXNPXxU2b7uUWsK0GEzPcS1+guJziqyq6N6jFKCuE9r19cpy98FgYEvYo9ECCQ5
grPrLo8gG8teiD6YbEMdFOULPpHVafYS2HW75lmA/cKy1SwcVJ560f2UIy7eXcit6aRHsbcjNjaO
wSVnD1cd0ewB6QrKxeKich/bNnAbodckuwcce0+3LeRXM3GZTmqQv4Wg1KSRopL0rxcKWwENENK4
+N8ZxWYZmTxNAmT9yXPgE3M+xjnKy5WzJ460Hq8DR4OunUrax4e82MWlf/Wq0vjML6Iysx4cl7rA
qdBjFXf43OIViX8KKddfG8o1o3e2hqzwRry232XqFWJembXgE9C/mdtKgvl70vSfM2lSIu3C7LJU
qmUgDozym1xQN/Vfs36dqhkmhmSGM5VdApq9HaoJQ9ZEaIxhA5TYDVa+D6wk1p2OzW1tQwrNzInX
qCcfGXCy86RiTgnMEhkfeAv9W55q5/8swo0uKWEr28DATFkO+/7E64qhnYxmv1F4qlcNldtpmSYj
QYQYoknQYqGpReMFon+NxfEIFSeaKx6JjKsJFyM395dwjfkqqwWxUN4MsmOOf4RXDyelnoC8Fs3B
S9ndAbV2/7uL+CL8Wv1Gz3uACk+d7XSmy+VoILsvLIs1xucSbDtam5ywjcscKWQMz2baMiwogyS4
TIlGiFwERxkEMSFt/OIScUx87tMLhCCaxfutJ3Lw/SE/YjVBwx4yDaP/ZYxShfDHumil7rJUBMaP
UEuxQ2du3qxN9PZStUgG3wOovQPSJCFyjQz/1A95gR8uY3peZJiJdxh9VTE6hyUI4Kb1lr15QxRl
n3ATyMrOEvoJKMZjBnmvT9CzFV8OwVvKs6aF8yF6JoksooPom8hGNvYT8+OCP1mKnzSvmIO/0pVm
bTaVw9zOHv+kQpOGxXjjqCnpWGeP6TQSZdMGwuYSI9U+470kzNgknrJfGwQvT6IWDXlgtJxEts3y
gi99m74aUO33ZT7oZcC8EwM658R1W+DTdp5I0AgV76t706OnqbTSL7c/ps1JidM7exclZbPKDRj9
EtFl6wk131KvvYdJWvmjyuxwE3C8KbAwxuMPK3AEMz0sdEfwVOqhVc5A04nXXbzeK4kJlTcLOWj4
WaQw8LiaLcuHQbOz2kokXJd2TqBzWXmlf5Nq95UJHQACzem3+pE77XAQl9AqajQwCSsdipQ5yNi/
mLYVyAwnMj0+eYzJNABfhEmU4/abckturV3qZQEuTHPRUFVmk558Wm/0bsoG69D9F9FWpGu587Sk
1uC+/e4f02gHYTSANQaV1XKspFSCzkw/i3N14og1mEhtEa5pOH/5GFKIlDoplySsesSeoKFjhUiJ
W6l1ozin+S1keoLG81KWJtThPocjDCosm70OPf9ZyJ2dnTXm+PASzomQzmSX+9qlxVRKpKZT8+AZ
qSR4LUyIe7V2UPLLCV3DltD6K77YkV+AKughjtK/jEtV6s3lX1zR2fjtBCv+YyhmdIskEUkUZNWi
ywgdnZtS3RmJgJYhhSDYjg78On6c9UTQwVKnUCbBP9Buy6KrsFO3/62P2vrvhBsnp5GVTEWZOxpv
UfBInEBwLnSksu3Q0QYULXaEuhPYoVI92GmE2RFAYuj1xqbz8qKsh3nVQzXUNMn9ZjqZERensoCN
zpQou2oUa/qo+DM8a4osuZsYFTnwxT4m6ogWKWWvu64AfVs68xSLVi11LPoIZmwTcRdkcown9GYv
cHlHyco/lmMpJaKVqpsLjpP+m+2HAhXHSA2qlLRcRs2v8SjzqhDNszByN2CE1IpeAs7lCMHvkeM3
NhOgkZY4R+KnksSrhBQPoABhhv9iZKs2GKBW0t4sXpcZcyeHMznxroyyGCbkUhQkuWpWzmDXAIHT
zVMhm9/+B42oafLD5AMzOfzYdvyBQ2ZDvf1Vn3UEDUJeZkCHBYkPh+XLtONv/Lpzq0fc4l9rWcar
WmYuXoe68R2zhjTrEFiL/8M/HiwhxJ+tOUR8Z7hxRx5A8QOXyMfTa+a5Xs/lG1Duce8SGzFVZRNe
Lw53aNpf9ZgVdPAqSPNEfIQGDNU32USRCBI8UbzNd3ULhavLy9dM81J1uNqW6Gc5JyuMsbaV+oYj
ZqyH+CGurADT1WNhsBKHX9bi6LgusiUC2JLC2gnJW1F7Lnao9K1XYq0d7esoEAD0NiZoSFJXU4VN
TQ5EhB6RaGjtU+n7yMzjZA5zMbjquuHKUCibl2G22vdEjBwzzzkstc6K6ah75uajPVj7GCWE8Q3D
A5QqVRd25udZIKaMMAVjXK9vTJNgP6+zaHIbxKPsyFBw4Id45aD2kIBjRsG4Da8uq+UuSOQjLyCN
EpTbBL75XzTO4M4/S7k1fVuHaZhyY9H4RzB5T6xEZpjWAHeEvac7bLziv+mG/zlRtOvImlMo6C//
gMSzbFnKYFx2quuLOYb1aH3d15PuFLHXf70DEE+vpTkiE+cokHwKxUU0VAiDfKM0xLwmeFPMrN3P
oEzPn5EBuxSGQelK1gkyqt/cj8U/HMr4p6a9qswKHZ5MvSQn80psgc2iBOx/D4bRTaZDUrt9h7yo
5qBmdYCEPDk4ntjkXwhRPKfq6OMZljd46l7t4g/SOxpvbv5Ap1gRqoG3Zm3hTf7o/SmrD2e0WuhR
vvXeT9zXX3oHxsBjnxQznsC+PyPcG8QeAyl5mhxZqw2OTC6H4SypkTheJQ+NV7Ploai7OCQG6hoF
MlFEI2KY9hYTNxLV4XJvcCuEToT4oEME8UM0irPkAKbQ0NM39Y6GpcR/AxoB7BDgxA2yE62lxeib
Cw+N3SGkB2EzOP1jAz+MLnRxBBN96YrT2Xnmk886O21s9K8hil+xbAkjy1GkddCqrZp5Va+MhLvt
rsL6ZNnVE3TEz61lezpF6s6iLqkJApXSGam02NBDMupYDSZWWd5UXEr6pKblVk9Nvrpq7sgVBQCm
Gd/O+RoMlLNCZAeQeQuV1aZotR8Kc8R/NVKl6XL1Nhk1HoFsq9cP6ZaFeSSUZgsXTAY9iRwr0e2U
8+przCe28snhYqf2apn7oljEaR7d7tlJ9ZU/rCD3d9mjdIT3HBCBVAIaCI3fkOZ8Wp60ipQWR9ez
IufxwrzqwDzvT1q1hEsT7pwpM+BDYadil6msOPHVQ9crUaBUT3ZLNRwnw0GpvShZAEuNuTI9IW+r
2fL11M03njrh7hYxSUWEXeQAHafrz6ko3++OopqGoRxF+WMTE1SfIsr7Vd0spr7/ideBlq/kTw5+
/9UTfSKD1wP2VZguzeA94kvK4iiV2AlX1Tt0iZV+m5YLc0Wq054yeogeVb0oQDa5FjIEnL7HtGpk
nSkjhT5rnSwEYwGJ1gNGo8dTDICcN8pgH1rSwW1NXYXT9VwJcnbrFPOvJAGD7YFhpOdA8MPAzK27
wGuxHzqKRLjJClexRvuqAwjHOEV3sLUp1cW85SKNpdo1LUpYRO6vWLXAA+4YnZoWjyXWZNivzSBK
DwktqOjFmNaaihsS/HtFuwFQLMsHzxxuyEkCDL3Kh9jZoWZlMAm46cRoPsx/kCHd+9UC0zEVweIn
JyG5CLuh/sQXo5UreqfKJDA6AmKMRYisu4gqviOa/55/X/3Rye3lQCwWDwvozNKVcbVz/+jZ1ndo
2/0vGN6n8HwhKAkuPmpDE6E5YSR/noAln13UDfKTorUQPmcOLSkNvifbVLMLiWs1LkQpnpVpsowk
D8NfV1cYG5Ob/lj8o6g69IoTpwloUrLvk3Zg74V918WihvAQCiRPmx06JUaz1iOC9BhR7y4ESumF
1zsPt4IwxEZl7OD38Xn0lWvsKmWCRd9G9ufh+2l1fohJAY5VsgdqVEtMylPPMbrkvYF7KkT9GMi1
7W/T90fYhTuswJnIBTJi386y1rW3OcxR6jAVA9GYN25NMO1rP/zAhPC9VXibkPiw/MaraART7jIx
me4OhnGFloLl78Pk0/ht/vwMaFZTuSJEDUhRoogAKMamjbUcM0tM25If9ohvIndb3L4ok/MC/dGQ
eX9kPo3/L1kDFYKYt9Zok79rcykAzembwU6yk+qrfu99kCuLNuGt0NlWY25o8zmlj4hk18IFsTiV
gRUTqMVd8Rc18vELdZayoq9SUwRKR3EHdquH/HK72AThfLJm1JAx8X9VOW1DUC9NQ2Sku/A9RxO1
uC2NY5LFtAGeOdYU3RhG3hQq2PRuMTlqVtvUMzBLAieeQph7ESDiUVwEsVGgpBQiA/zH6Vf4UZf9
nf+wPU/4/06NVKNYsoxHWQau/FGnPO+FkVDnXdvNyDKBxa97gPQOFeIJjxnS8nao8fw2VwAd/a2D
hjBBERmyyAlx3sbJUcx3I1IAEYRiNaf7KMbSP/2f1vVqz5XNCSmHLlz6NUMtK2OYcOD+GkZF5toi
Khc0wx8YnKNCztc5WmrSeHHjHfu22LDYpvs5++HroQ7FH2XYADgehaZ25QFqFMQl1NyO/fyUhW08
6Yrwk7i+oNFERX7n8je0Lw6Q3C+RdoIHp+NHPTHmR/sOJPMw4VG3jXRb45VV9EFOB44Ixk2O196T
AFjA4s2e7kAf6t6jZNgm+exJETJDyOP32kI5s3HW9KxyYSnj+HFTMFV7nVX0m+ec92oNKRwELRgx
FW+e5FGkvWG8I4BzKKrF3mP6BzJyv2LM092YALm/oR2q8eaop97t6tIfD5tiAqPRBEEuRRZB5Znp
giqr/cGEjmf3o+HbdbOG6O0KWD5VA9xtz2XR8E+YZQixAiAAtzSZt8ixXoUCpwOAleXVzPYGZYOd
IypQ+lUdESSO8srUDjC3SfFIfGkPMUY55sJ4GhFv69C8dFD803ojreFmVzyOT6isDIDiBlXCBXSm
gH585h33AXLVw2RthO3uB21Y4C24nwXh07Y/qdHSGdziN1gqVp2pkVmr8aGbMH/WQb56XCf0ALIF
i2bp59ADwCyVRSqLR3I5g4WfHkiE8iHRA0b5VJs/1Zxug5CB9evVM66DvnrnDXrs2tmxsZiMZDaA
ouTnPWdNwmcITRrUOcQYiLuUmvcdi5tQmlbYaX6TN2iXMpYHnOrkdDyvP7SIuCj2u9/+2vIFh76z
Yy2moE3PhBdSCH67ic3+GC5+xyTTkDtU6JpOJXglEcC2EW2SaGqH099zRSb5Cp18OHSYCXf5WtHH
S4j0rzHCDhHF53CDBpNIANxdQI+jw8Lv5uPRanP6Hgo/vlNpOeLGzc/HSQh0IcxEuLZkOXX/oJ98
Z4JVtZWPR9aaOx54kb75bXUTWf6I0gzjq7uhyjw20erkKAnCa6Dz6pzBoPaTCKdwDRDEbak8Juea
uXYX3R4MCk+MMwfih8KYPdQXMxQlTWZXlatFr4dEMNkNM8pYy0L4OfCUeI4rWMOld8HTX8UBcZHj
9LC9v7dR4bPQaAqX6sKY+q6sKXRYQZtK+UPl3j5VeSw2krdC7M6SrXRr5+OT8S3EeYk3ubtOPfCP
K/G0s1LuwFRswNzLo5gtFn+3Ag0GrlfLW8RG9pVfxY27FGQ1uqe0RCMZZTe52y7SzUjSlBWG/gyB
YiHRFZvLNUo1ji1LEG4CBtg8e2JlUgtNTROUbbdzqTArPSvhRQTZXdtkE0IQox7Y0TxEToA8XiQ9
sawOXBMEWNdiYffV9Eh/4JZ6/WWGJISbF9jViY7RIut+ZFD/zDZBORHLe+rz3ktzN2PaVNqbWMnH
Hx0kzug2o0HgPk2P1ZwtWjLdgW/2T7+r9//PB61mIFCWHwY5m9mp+R4sCl44c0wHTQx0xT6BZkhw
qQ9iZhFRTYN06pQR1mt2oFWKSDz7upLc5BaSgBL6miVhu782NXNKK0EyKSyGSv63TbEDUs0s8DWk
ZrCpJeaSyv6DtqQcxE0+TK2AUnltTToSV9391+QBYDwxDkx8lgZsYiodudYe6CUzJwwmXFvWh1iz
/yA1vobcot+bXG+Qn+/BCzd3CIHxfdPeGRytLZFympPP4B0zVznQkizeJ8YJ1v397ykxEMnl5axx
PXPePNKVtuyQboZSOcm3/MenhP/g0WvQLhnfuqTcDiNxHe0XRAb5WhTQdpAsDeukMD4+E25nh5U9
dCG6Smk/2s//pYqexfdxzBcIxB0BNM5XtNCDS4GbTych8p6lyRUASm7E0X3usndJ3yhPrz9vzZml
J0pGqYPWSz2rCfuoRe8mB7O3UDxbFvQJhVEUTpHEm7ePQfugV8W0XatksYAOKoyPajMPHXncXQQ5
4mWw/KXFy/4WmgYRMtzlGmLAssaeYH6xzZdH+wZt7jpljE4JgxPnEmgudFfVF7VPgpfYFHvSljTo
FEjoA0qknpokd/K1+lnx1gi3AsBmuQaevHQv4ayy7gLM0xvXwXKU4gnKJjGljnENBPQVEY0GuGrU
mgFDrVvf6IuNYYSPfs0UHkA3KCwRNa3iJJu+zEp9YVgVWdpwmtDLFdq9m8Z+g4Xl0V3vAGsBIU4n
9HspGP+++0N9Pv1l8dV6W8dRvg5uljThm48DS+owvtZCAcrFLJSkCNvyz/HxMOTwQcH8yKhZKEvs
GGn/YnpNWfpkgQBLNFiFSzXYnKVm/vz71HLSkNz0bqoc/hiWFnggAjZMetFRAif14F/Io8GEPKmx
31bJ9S+ZDhQG4oyWPS+ohmywDHPBG+lFhTZoP1rknN7KN2k/nNdzyr/W53Vh+WnbnqxAWjLdSxBp
SvO71UPMF7J237pqNrgUYaVnq/2H9Yn+PzSd9A83UIkY+zH0Rv1Gw7DNZo0wBXG+5Jr9OEfBKLW+
a5SV7WFepTtHjMnaT2Jh5cNW75Uh/s2PTcR5U98b8+VIezj17KlYavoUfNeKXmP7fGyC5r0xY7by
8UjwsNWjk9ys1HJocuycEcFvy9+s9w3FhKN5NwqdRlvrwuveRJiCZEahpjuBb/gPuaLjywKTbUex
B2nKFDyGZeZhqbE7Zf2m9bcfRx/1KYg4jnBgRYHyT032OdboQ+3pbxXVHy4ivC0a4wYp0ax2tMsu
+9l4RCxfrljYYbMi3D7ERxFHaMgRsllezivsib50V4xTQZ91ArF+ddqpSIJ1A7EaB5AKbIcNBwi8
hIhQ8p6d90GRBd4RoyfAOiPiSp+/lDSo008UiIpoGwFNTLCcXoyqR354n/b7bS2afGgpRgltlzdB
eE3VaQGwm7dfPNMbm0Fo/dJw9TtIRehAfViMeoA62iSsNMixU7MYogKd21fPJ1LqSoMm5LUdLURq
LhcTl+s9N/SD1IZhGJ5hcNUw0L5oVSrRMBVGdCiz0noT4PK/gbp6n2kQDCwRRBgU6BF7XreItnTn
jMB4c5h/+ZM2RjjHrvkWJBJ1apIMKRLGXjeMgzoEQuvnUPf3X2WxrZPGxYorJP9BTYQ9Fq77EZZR
9vN3WljGL30+LqbQjp+NKpvl/HsUnvmxHOmijI8Z85M5ZnsFbpvGGyijKheitxlf00ZpVMEBjoVV
nNRgA+t/+otY26PQcUnlWGGO6XJ4IVZYRWzJAqmskZ8cJs2js/rv7bZzfoQszWsGuRqlhCto5Sr3
E5SNY59s3Aa0F/eSdhIwS4x91XX4Db/cuNrcqcjtq56tv33dBUU9T2ZkFFFQgelNZZlNOs0hpDtw
f/etwI4Z+QaTMiwJ2XauciWeuAbSEavx8LsKkZ9GnjNKOLeeoE43uOci9wlfH8H5cHOkhZD5iDEs
4ie7A5z03J7utA3x7sDa8bcTztPAel5nbLnMSDemNuPA/F5j19cXiwcq9TrkXmj3llfUMaYVoZi3
29RUN+NnfQCabGi8e4J7PdQGPQrv+faJ/QUnsQz+MDzSfyiaSh4UoLP6xOVPGOjtuRNyyzt9HBpV
dY6XeNPOTg3VwMte9zUvaHRD3X8XIHC9xvM66/K1HA0fuHjAPE+YiOVtMLptwlAW82v8aRptJa4W
FV+KjF6ZqrSsaI4lK1r83Ix7wFpUoz7oRnnou7MsDXzyd60YmnqTMWIvVL/gdMBqIgZvGZhhf9OH
En8pjgrdxBEb7DFIKEn8oZuXd669wHzKJ1XDQ/xbHYQHo3GUb3hMbzaNY0B2k6Kr06nijY8LphWR
hm8WuINdBfnkHUS8Djk1nZdgpsFJ52ksQgHpFyz7f6gAB8zmdAjiJDblYCTrN1eai1nL04i9vMqS
Xcm8+4PY11bN9T6JMLfQ/zQM/jay9JteSsMN8VQCMAGikK7fX4CGUqFqWCAfqzGdsfYDxfQJEB4D
S3ijMu1OOwZxpSmiRGqlRtwlfeyhYWnGr0MhTlo/pZotLUTCNqnuaAI5HFqBkBYTfR9JIYr2c0wG
RdXo3H9zmT9gGNpUvj3mbqYtl2lQqHJRP0y8NayWXAQCdfppZDX3kDIMvrzJlzeT29k9I+2thRjO
0g7teW4uqXoElYS8IbUPOjQ/TXK/YVHxAs7/akKe4oXP17ACHZz0EQB+8aRBqRAp9nzoAA5L7CAa
aX3Av0Oxjo84o9AOavPgLaglXaWhck3I/b0fLWQ5RsSZwKJ8M3uDKcDXYOU1lYsWjGDYk/+4y9vt
UZgBcM/o5h58EHKTNtgNw3tL957aqphfoagSrPx4XpBHhGXOrA0UbNSK4+L7nUl25vHi+U3rRQGo
5HebWxOgEKxNLV6RyUP0STrNip+9Qycn7QHC9pJVH2E2NpJiRRFtWiPtnOKlC0PzZregTt6lAC/O
282BX4LL1Kj77QRn7Kw8XcJaCwuQ0IIlyLBAi4qfP1FOHd1/9UOUyk/Ne2OW1z2uVDUMLOv/GEwA
HDscft1vZqDyATcSiCOGnzrzlhxEaAdJmU/R3wt7IffRCPZV2/W1/N1Ap6zjar2DzcJ/joGtK7XK
kt2gUGRxi/rRoYdOlfXT0+yeTDvj/h0UPFonhpJSkRkL/1s+UXaxxrHGU6in02RQ8dgqMOW8UpvD
Q11mU8ZskobrmbzxXngCVvmAcFq7aXeE4vHfqPVndUxCeTLnerIdqq97z21/Rk5mQ69I/eyODBPj
2cHFc+/Xs/ZlDWnpEyQAx6f++LqOxKNlbWEEc7r2988O8FZ2bA7ncGgePZI0y9R+/TJcqIURJ7Qs
Hfsnn2pbMWrc8uEV44CqGZCX0GkuRmdCwPqkyjKnnxwjrBMwqcup3KhEbLw41ivise7nwxYBF+ow
BrWRidpN+Kr++EOgSfLKx604PtcGfCUMGu7Ea7kcntowqSLk3lBCTJc5oMcy+KJTirnP4HqLM+Ce
ZRJaRGYCX3ubM8sxhWkYSjUumBKjc8t2NnczFgrKH3FekAKPCOnVN12VXq45T4ohZ/E5g4Ao16ek
D/Kk425CN1+tCBEOzYnNiRk7+lcN7/7/fghYAufdz0O5Z79MKowbRaW4rXkXdEfjSW1xQsUgjvuV
Erke9bNokVSvx+f/lbHY5EDNIuvJoGslt+bW/qLx1knmNvEXD8EIhuo5S1DGtD7tpI/cC5M5iItz
Bz/beh/m/Vjh5SnE/NZNvQY9XjO0KPnMxYmmF9G7uUR37k69fx1rqIRWg8kZdeAWcDqtmkZDERvd
oYhXL56owfEkOpv5fLP93HYg9xQ5Zay5nWoSEg+Datu5+OAQoXH3pLFJ9CfuIDrc10BnsWCAOzYI
QYE3r0WGgdl7CDFLs5E7nCmlKtO7FS2nhjHfJuPEVBdLc2kYW+UBW3OdMDGI/OWiv3FtQfaOJrq4
VHatZ6oNFxxd18OvtiCAuyh1fKJVmKIKCCJZ6o0twWfpvKgAxgw5GqoA70JvWk1+FGuaxs3Lz9fw
QTjNsMHauC+jhtw+q7jniVSLbQyURIXDcg+aGbBmqAxVulJ4clh7rsgqPQC4uWAV6pwlqNY2ecsw
QsU1BEMXD4gon+YXUp7I95lDOs1GHwQyvnWoLFQMDlvavND6POqq4u2Hnn3t/dzBvSjcuEral+Nq
TtSvlau2KCpLDYu4SXY6EHyFYp25XpG1zPQQfTbGJ0DV12Js8J/ivP/MeD007kQqhxQhc3WmMouL
irUQlR9zD6msMp7/Q1iZW2pU878DfjlyGBARHw3MVp5cgkL9t3sXLaFYKBvlECGtdBTcKG7eVbaW
jgGd46mBzRadzcDTmzmgglHVKYnxnklFIfmyJsYhPaDZZj2e1M6sPfq4xxfiV1PYv9ju7S10vzul
gqdD9D5S9Bh92UBgAi6V7sBhBmAcDoJTUkxWdxPoeeDGzqOca7FWwTLAEpuoawA7ipv5I1HWbfDU
HY6z/4TJYYqZUfxvGn80fWQ5BvjMsi7pmzcdF+n/+kCtPB19AHhQmA1kAIntmsW//uuWXDPEGWWg
haZCkIlDjHLkaShYsThRCga2mHCIqASRyQdguMf+LFISs6k9WRqd0rH6zPUwYv75j7wIQmZuvU9e
X8c13GlpfUdz8iYCe1+MZPLaflUedWJorX5WynXAoXAbtxF7dKL1USWfgEdcLaZRf1l6QDH0tZha
SY5wYn4FPrNChtTIwdYV+x8cpJ0CW0YV1I57FyBNWPq7yx91ecwV+Do4tgnP0BODK4myFd5E5k6v
VD9F97MxIKyeVyni2DYXXUrj2ReGa9OMmcFgIa5VRNPPZ4lKQ+bKztJ4/JGjlNNdWF45WxxALgAw
k3xPORVuX4mCIsPgCEW+gypv0J+M7fEPk1MeLFsyxRLaK2rsOzt3NwP8Swoi2/uVAlTksuCUIXT8
Ihwq6cS+vG78qWLeEqvESV0a1w1kdb8eVH/VNxD+05ojmddbNzrVo4kH+u1QQg/VNmxUOWNOZviJ
19frjoRD4K3RndtGttfytg6wbfraeDwYu9RLv9whEhn2jhdW4qUEROHx0WxeQT5hnucUP4bokPJG
6Lvyibs1sEMApiJNGdUb4EXZ1wehKq2mjvuWahRpyjQcmfi9HjTo/Y89M2mtzKxaqkcIr6wZYzwC
CzTUxq+hHpPDwEtznbEHkP7GhdOxKkwoZ6+TE7MVVC9dMowNcAGVh4PIdYPNXJs78739mcwdG60C
+GhNP3EAlTarJ69Wk9CJvZb0AFj1Gbrs59A+J9ac0qkLFtxv2tz2P8R/78xxO5WykDBXEHg8HhBs
vBH5ZhvNSh3LM446XjR+qtf6mlAkGxrxQF9AQ7g8o56CbUSdYtwSDx9DWayEeLVeCUoPiTGQxNZT
RXaCAWOxcPBSGnUXZ3zS+/626uEZjBlhnALJg7SD276aN5j8FdtIiAtGFJPEfVChdOYVwMgxOiNQ
qjLeyP1FYZLoxHi2L5We9HtDJcLWcH0seRJq81SfZQ4qOdysZgvlIZXnEbrbw9319RB68Fe472cO
1orPv+bLYf+nPxm0SpDaVgBGMIpdNbp4IzZzo0sv4ALEb4/1Lr69IP7y8IjVJiUongPTowS4bbcv
nAZBAJwR3TJ/TqmWoIFve6O8TvBbNcolGot6AjzLdXM6wxwPXNBAiflIp+PtSe+zbqxkggBjNpAz
GLj9gKhD6AoKy+tnlUzcafmFBZupkgI8xFgguEiOXexwctxhi3VyVKs+SwssiIx7x4FxaOI+HQMk
gle5wn3dxh6HZL7270INvECkk4tpGhR4Vb0m7HISRAUQH6owHEURLZkJB5ZCrmCuRMQwkEUu6zyB
8YMf2wU03wmv1AnCSVz0+BdGegQykOW4lzmxw+Kpc7Xma6HD28f/HK6aP/7CGggGSKUpCGBrPosB
3g1hUQB9YFpFAMcG0IQ0pj4CP4PuvgnY0rCxiw/YmcC6tmvRpfTBol4vWUo6letPoVkxFmnmjBAF
SAN9mMd0ldABnxlYbnJ/nTuYARCEIM6zCsZkGM2QAFaLJfp8aGMwuov3zZM4/jYxE0zkj5DNbKZF
ykkxCqJsOVhj0IPHYIRDe+YaQ3jUmWr7Ms7eMf/bOqJlv+bjKjODhnK9XHvzMju4X2DK4RWqwjLO
YPe6SdE4Ki8Fbmee+s8jIUeqRGUbwturUW+3aI4A3YwkQt1KYhHkdZb0AaZ1I2X3njiPlgCM8CEx
pXD16cz2q4geM3HA74s6uQlZw+SI9jXYRw8j5kGcG3zdUf7xYiYJBh1DOml7R3Dg+iF7ySrAAQe4
TDfkdcOy/Y/7SESreEm030HykOXRQtuizciXl4ov8rFnxqd00tYIF0958J7/pRglkKyxnXa6RuFf
QzpsxEWUwF9Jhjm9Z2TkyWQAMlnjmVliNtVAHqHpeR68GAvHfdPPS6BvlZEV1Ns/woWCSfjfhEiu
MQukklAuNfqYiMRgUcJpob6Qfxeudy4JN9NQvkaGny+6TZ5epWNOI+0YFM2qI9am25fFz9kc+hnx
awwTZftJ1QAkVf85cm5wTOcV6LE2WwKNHBIqh8vuKKpJJf+qadCP/CNv9YezrX9BrZXnJpNmFTzC
C5L68pTgmRCln+8uV3ZFU5C+xkdMGbLLn1NdKRtymNuaPyrR9r0MK//wQ9ABUATljpNsi6ErL1u3
mT8IekWOAmQsx0mnXOC29BBWQn1U5i7LARVtLNgAtVgm0++cmU0xADPGrxDXoLj5ja8I2jGkOWoT
12bQvwgKG/tMIiBzw5AcdaNSfmCw+7M8x/LrBeU/H2btmylDo/2tA2KjzWwkE6enp4P2WrL9+451
kS8fMwDZRWSlsmcKoBNuUWyosSEAAhD93CGBgaKF7IvuGQqaanpLV1EYfAWFi3LgdIoDUP3MCDUv
UKwpx64pqz77sqYTcuip4UpAA4N7r+8B33PqZLGHEWCPSyy/vXGC1N5HPdMwFy6y8o4VRRtf7zG3
oPHRQAL2QV3lhsNAxqZQoRiG45URQJSJXWtRDAZcgu44XOxEx1WMBZ7DxQRJ7UEwI3uUe/MlcI20
ABhDuD9suYmHdx/cZ5L3NDrOWWl/Y8JotdiI1oreyjjLhwS5QYHjNvLclQ2W8nQMDsDdLm2n04nY
bYZGqi+TdBUCNDOpsQ2hjoY5SwY8ca23lmXDbcaSIbU/mcAY5jUX3WpHy4QQbiKCB2950gBz6Xw/
NdwxpYNU5ZfuW3+yvzli0hPuvrK51wWdx80Gm0gYMUpHzHhW2OPLIGgbtYCHZNFHXjegYY0PmM/7
4GDQ1USEOwKJsPK7mte5UVnaJcqdfAXOgxwmDqAByFqus4dfyzLvLZKK/CwW+vBaa46KZJU7wJTH
mXFmsJT/TmI1oG9gkbZ68J0zQ+FmLQwZJo6TX9HlG4Hu0zK46S1zq7ySnAb2xrVEdUunEkAl6EBj
s+fSuGsdboIPB5ndWRtIfjiI7QYeyW7iDIWDkKmLVxyJTCGKh6uzBkddcHeyuvbdKCeR+h9/gWtJ
BdQOau611axiBURHxB7rjV78l7W0dsHZagU0n3O5F6VfKewNf5ndZB1M6pmp4wPHHPE/Cxu1hwEi
3fCz/xIz0PdO/LbGr2lcxFG0Ed5sMC+gTENedjVQ1dTVn/KFBR/UiF6WBCpwUGlt48lxQHYJDZVq
m6qlUJFmTRsNYRPg246bWAZbkzU9EdbaaS742LaVBVn5EW2ZruKrOqzPbZiJpsGji4qp84A2a21t
p15m/ggRI+invQn6gLhxv6dE2blcpHsjDw58Clsao4U6g9/h/CGynwEuiyPTASi/kYbwPrXBikit
MzEHtyo0L/H33tVd0Laxz0XKLx7159w2y69gvo+Dooz/P+eFmvC2arZUvBMLyhSp01bdi09j6KSw
jMCsPGmRjgmbyCpxwyKGxi7ywlES3rK91x0DWINYUfhx7+MtCkmR3cx+vUN6LNuqPCP3tob0KijN
KBYV2IkoiR0MSf9zNq5qOgazLYWEmxw2yqIr0vYg7YMC/FoBLsxZcn7hRaAtKhutzRo+DZh1FqKk
qGuD3ir514AH873XZ807L0uvrostlIFlTTSNva1/xopMmZVAqjNoXXSJentGVyzQTvNAu+Q5/0j3
6idxy/Rzm/+0Z8Je+RZcYMMQjSr9WJfG6GUJjtNaxv6FGpYQ/tgfgZdyBY5qMDd0qI9y79dVJSYr
qrIKq0DV1e3544ttVGWS15P0r/Jl/zJQer8dzERC3ubSsgkwzkiCnaoC0XXhdU/g2ZQtsAW56APw
Xa2xjMui1KHV4HuBkI8tHplvIE7GU5eGebMhbYofe7Iyqr+3N7pCvMRBgX/sSzHxC8JGPs+4iY9A
tzl29eHzzdJKlQjDO60Ya8WE1LwpTsnMUCSQIIxDWblGTyapYoSw1QXkZ2cvfZ7HeUwDLf5zEO57
5A4dEqeqkK0Xs5WZXJ7VSiwzY7n+A+Q0sdp+hjzLAjFpNmlCeaqR9pzrvJbVtR0ZgkZEox6WrwvI
1SctUknvaEZ1SShipfkqJhI7ehPXNZDOzZAq8x7gj4yJfEr6hFkUUYrTzOpFJZ2iEOt+biNeUFbC
2rXySjEOYpvuQqj7iv3uMVs5k8HW/M8XvqdyrZpgKTH/yBv3azJNdjsbVjIxZ+l54WNNz3RIGUMD
oej4BQpEcrG7cH7NSL8cJwXIIjzSomv/xFSc+//17LTXh+3XFmK+CQ2sRfA4LA9cD/2DXxQ1KMVy
rEqEcX8BC+7qkZO/ZtKP/ZklVK0se7dfRAUqF+8P8vq9N4+Z7B2rbIMwVN0qlvx0gVHMUHHT+ED7
Ppr95qGsbZWscfU3jj9vskg+JeHibl0K5MVxwpTCqr02ptFD9cCJU0XjcmC5nf+VyYfn7DFLmKC3
G+L19M99w7vf6K4cGIhSqcVos79PodnSUpSpCWI1Wogu8ChyoJ4HoaP5P9MI3UpFq3p4jBbRiM70
Wg0P/sxa4TrIbWdYt1wlX+MI+XHXEW9pnJzw1lflHUNeup6PvfIjsohJnrP89FP8FDbbwWsqs24l
6CcjZM+He6Xd3UiXhrXlhSVGnBOl07DhALlYEq1GuUn2vEOijpTSwhC7Cv2p5gIk3f1FxjbJR2s9
+zof9j+uhOfGQWYPsDPAnjpKjsTY74ThDgy3KAfWsczH58o8nCIGU3ZbZ2vYKnrNJajMP/fCri8M
aqicQe9Obp0sDzvtq1+GjOFa6pEl8ftFYHTDjbn+2HEdKW5P2bhRn6lfN8fS+ONX9qTVp2J9DZBk
j0kxesBOJ57ko4kL4GHJ+Yo/z/OrRbMz2GJPNXmJIpoEffQSMTzSv3qWQCWTv7oFvsh+MnJ0RPE0
7nN2Z9r02QP4fQ+N2zfSwRzD2xLSmuu7YgNpLkPc1uhBIHaWxv16+2neUAekRt+ozbzxWxDTn8Fd
uJ/o1m6ulGJQSZqHEcq3Gmkm9oiH66LHYWGoJTkB4emX1ZIknHoF0eWNUncbXfmLkvRAtqjeYaeT
GhSw5FPQVGMXlqxnUcOMy4L91b3NmNpE2qF0LXyAVvjP1ZotzFxMTMKFh9knib3oy3Isi5fp64DJ
OFxEWBJTrKsPLHI7/ZRgHdp6fgNZoi5YWhM72VDYJZcObyGe9lByUcJQMACxoMHJYhpLRYySrC2t
YNXD8ZrFbWRVCQEhfJ7UtXL24S3SK08rlGlW52I+dV9sypIzp46UV5pkgepaR9PdqH3ioo0jANkB
2F5Xkw16WKpu7XUN2sqoWYGS4P+EyyYGSty8aDY8bApSO4yCXXbvHGeaQ651OIU6ZiezChYJtJ9Z
Fc0OCmDHx27yEDi9la9OLi1I2mbmecQEE+R4BXCP6hWFpibBQ1hLu31VmrYDQka18BPl9by1EDB0
5Q2rEJf1UxD6Bzp6Z/b5GACkJ+6rS5CEDSQu1RJt6/56eBFpwXAU7CZ4TxHx8KoG7n+Skm+nj1Nd
frh4LRkqdBS2g0Ym6SU51AC6k1XxrJ20iH3oVCdG0isB1BgKimHonctv/23TBZClh89u5NKm33U7
2IMAuNcxwgXww8/utMimDFnajRUgLCza6LZRv+/4KzTduACN69VRQY4dpnA2/r63PJnrsTJKPEpB
UcqFYklHYD958O0PI5FqBT5i9leqg/5yndAtNMvaaKCA3ob+hTN1s8yEp+HIAbnmugrcGtx7VP08
/rPadiLXN90RhXuqb4cq3+ms9I1GEKhf9yxt5d23YEGMW5Cu71tOW03cgECSUrF2O1cnV1mM5S0z
M3i56SMQ1lXHTuiaiIAgDWxpSOQvlW4L4hiKmrGNU1LFjCKG4YbIL1HGAvWU5KlGQR0QAcuWQ27R
/0Om7Jevpan+DFjEGvZE0p61NCIvqPKc5OxcmMkx33OTRf1PrHhdntSYdbfbNL06ThY+f9E1Xtho
faRTk0ukMsBXrZtM2pJvPYjUwLOtRZ5LaOOkn7YudCsGUTHipLUFtz9CVqrEXn8dVQvw5aGP3SdF
1hZ+DIljJuLyWSWi68v6egM5S30Q82vZKi+dRDwliHRlnxEK40ajUo3vcU5dxK9fa2ULnJgH5y76
FtuZLZgEHfEBjcULD7ySJno4HKcRUrUutdO8xZFo4FH5dh3CPBs1GmYgrDO9ahlutCHQXEqt0dTj
WQi8frWUe6EAE+3DzEa281IGVrTFDayu9qt83Yg1xQok8sirGvhKQYS3sWz60Q0mDby/Ero0beeY
GjN6BSEYU5i+QwqBFepHzn1ifH+sZikzKpNbvSjvQROXEYEO4iDfUWBKsCvwNYU+XHel5wtXAMIh
RRHvZHc3qyZSQWVANQjec9y84M/neYkTosD1Dnz1LuF/WuH0FLdx8i5OfKG+bbMGNOh0oBnhYW/b
vJxnl8QHt/7Deyb9RgRYMbp6ILBTlaOuHgkgj9f+mA9a8Fb8OrY/m801e2r5Ku/JMIRzvsKeIUgt
V6hWxmby2WH45XxKsl/c6VNGI74zaHeQuSD7Z0+IYKtVtcTT1Dix6ZPF7u+VhMh7FJfkh92IoIdF
aVpNaPoRsF08jr+Ss+LVXpLWWcBAAhR2MHpj6dlbeW5wMu1Cz9xBZE91ykh+IvX9axycLvUhMR7l
SBSQvuC1+LT9kJnGo67+CzskO6w93Kc5+hpKcPmakUhW5J8wenfus07jka2I1/S3z//yPYWWvHYD
10DH/KvOMsWmILskDNyGCm6nKWD6bR6k+w2f923T/RgNbxkB8cWzJszfz8rZU8m7zSJLDH0kDyY+
VsJNL+RwRgqGtsEAehdwtTITlUrgi2u/BCsMYm8Yt0UaArbu/K4Bt3aHx8jAlX+7p2bstfHnQvCe
lOqCbF6FgBZ1++88Etsq1BZgMlQe2m/1NghGA0R8w8q5iiTk+vcULbh8/PyVbuuobFYY+6iqLS/y
ISsKiLGZzKcuFgxWouaZrf9ieirBF/N2jfdC09anLpz9cAv79UmiRHZHIrh+WZBvIc7O6j6YN6pg
+pT6MwUeNoIwXBZYJcYtrYNU9HnW3AefMVCyf4MhgbHwNdpbM7uitr2/BFpbTkfE+ueINH0+SZxw
771zd1kBM/VAHb72OcPnFLYkbisC57wAB4PwCw4Sz85zGfB7pYayEpAavL/t00mftWbgJd0CfALa
Bt8fOODrDxVHuWvYD6hjV5CoZiT0Y2iSXAQie1MyXtrj6c4qWdJxzaamXJVbMCIiR1cC035ukkOF
HeJFq02hZTJYf8j3DgtIoePERv+anqQqOX5+ujl6LxqzhWYHFtXYFWIlFGhazwLOak5AGTF7TX3Y
RGC9yJiNE3lm4rKHXePuNJbZCPl18J0S62pXs2ERE7BPZ5kfCFnpHRNN8XImgjgW6TqnugY6No5F
LTZHnnQ6ohqEHW5GHn/zYdCkddsAztFCDmcb0x192BQYCAeB374iUeGOtv7sLkjDfGURiC/h2fd0
/Dj8vFkHxMcpP4cN4xnOzxYGj4IqJjo7lFTNCxfo+XZWIQ1PymcLTZqjY2YsK8scFfLh1RzJi9+I
XKRyZB1GFhjZd3N5m67E1Z096PtF5s6j/sFjnu/lUCqoJ19iiKmcQw0rhob1r9C0LyvCOGwj2siT
UlQp0is4q/Zlr10PoiwlgU3/CFg42IwXeReUCTPAx4RNhEke0BvAI21r36hSWEMJFDD3N+iLeqon
Rg5qBNUdsCyxugdMSZNsxiV8Ct3XiqPdUZfUNXa1cwn1ksaqHsW5pXTm94BCtQW+mlLSJL5EQHjs
WyyeY3HQA475yBbse0RwiRrDO4M8QgAmigoPfuaf87PHwwRNqCEcrfgl8MqgwnlrRIWMAs6VDRgP
9Kr+JOJCRwbI3ozDuvH1i9RIakddsrZX+K1ttQevR4uqexPcRlxvz6cj5N9j8l+Sj541muWNFNDO
hNIwOBVJaN2WeT5VhAIN4pD6rkooiBfVxFsqrG6iQKnVReF8w3dUjq9F3J/YvtNPvsLs5O9sBz/x
LUTBg2ISUm07bcaMAB8nf3VRyAY1YygscJVzpdmJKHHfZ3pYHhYpsBZfpAVsLCi7ggj99Gt+qSm3
ihe8Kby8J12VJu8l35zWUFbSR/l3nlbLQuC4oykoZL1aMbz3UdRTjJM/TV1CyQs+5kdTeibmtaNA
ghXK8VV9r9Un5CbpTjEnV+dP9pYtvXkxLjypBgEOgUUDP01NcA+yYm0sTFhRHG/zzA5dKZWGQf4Y
vc0h2AXSHwm3lOzfceAPh8/tYBY0+MsSZ0/HK3xrRnhNzERWmJAWMYB/ULsFml9L5rKskpebURn8
yGw2HSE/JUdQuYr2vQ/WaJZA0DZ4s2G0XJzHCv4f0qdy86Dc4ECwj8M805Ol6G8tI1qrvOny1AJS
cmha4lkLW0uj0nbPIIg26T0Kxhv3hcd4DRKJI5HzjE2rt8dNV7DiyAlm0WHHLZkVaXXmQZQJipGC
575SrUCnW71KaBYQqoOSBLyfW81K5UIdWLxDrZUtQDfOG5XLJvTHi3oSDzvwTkkkAPTmKVG82Unf
LnVomA8V86vlqTPqKSSUQnSFBlTDe9ID3Vx0l4TGo0MyKP8otVIU1dqupGrXJl+tFFN8UxEG0JKf
WjRbdEXv51YlKPF2yNa1AYM5wc+1gZizv9M9WQxjVDpbQlUUbB2zg1qWM2nvsEgMRqrM4eY5jI5I
YN1EZyGllOrI4Ilsxou8rEauY+7xnQ7TC/5ITwyjE3BOEHEygWfw5K7o7hDC3/1dDZVnNlnmMsyG
MVptPVDHnDBHry5T3EA9UzUbfLex/1KxcUFR/UPh+Zd8u2vu0g/CHLMXNPJMKSW/HR+3MfL+jRLx
HP9Wt14wkyG7BmiY8YfjStrVItgU/vzxz2BcqBWRqPcLVvTZ3mERi3EqJpZfihUoWIfeS7+n08Rf
BIdTV3q2+wGJRFwB2h5Ph4Jt38bvL2JQnll5HjtnWMmmLrvJv8hU4RIqbSBLfk+VOPR/s1GiMNQn
ZFIInKNL8W9gNYbdRKUOZwYaZI81tJzy+sA+8/+HdITFFBF2N8wC5bzum6y8AkU2vgmW+LlK8p1l
z8ebxaEMQ8r8voripLrqlUjuCHA3Gw0JyI/cl/6lxWzERQdsWW87VxTMLwU8B5atbmBJEDo4Dp+j
NYuUKrV4pgfBPcY98niVBlCGBKnh9q2p9+VEQU3cBX+NRXXXnr6QoM9+yjQcqokxskWyXUENS/88
Zk0KMTk0zM479GfB7Txs8HO+u+jtfVLEjkmq36fVvnd8OaByVniLPtKuUZe5ZYG5zyw8Rcler4Sk
zFv0dCOxGal0CnPh2u+Wog7v0BapW5g4s1Ns2wv4Zkq5pH9+9QRcyOCNjgdQmpQW8IS3DjoG+keR
QU5PxnyZBZXl2G97Rh2BxU25WcJfXfOR3RbgXFsiXouqzqC7CBPbHsMLNcF/NlCtB83M/98lbkMw
6VSIA6U4ZxMKg7FxeyI0+uSo5YCsJKL+Z665z++e1SR1gcU0S/Ajg00u9uDIVR/EXXpYY8NNmfCV
udzssaWhKrwTFu6dMS5LwqKAWXEKe05jZU/WTA9nzPNp/HQqRuDk9HIcwije1vGj9AWt8sBKRZSw
nENVWmSJuBrBzigTZCiKAFpIa6Q/0aAXDh8uMoiYFSqvROVhmWiCtkwrFCrNW2geseTR0QxTeoVR
m0aEAStk2LGiNlat3MlrS0eekHChiW/r7kKFGoI1s/hqbitZWJAnPz31VEAx7KHlbsx6+lu1TzLY
nj+Ym7m7YM/oJhyj3//Wg9U7+oM+nPLquayghOeSPel3dglPolzIKVrkrwgllgziw9B2pzh2EAw4
YE8HJ/vvyK6N18pM/d4nEKgr1ywsprAFEWkstCJyLKbfANHH6vzJNg9191aNtfjOV7MEDT2wRiOj
VSyMPeFU7i4oT9qA0q++9LZg2X7GFxBYFeQH+N0RRQPPn855/Um1NRvE57AvKm1Y6Imh24h3k2cB
DMp+vINgBhEFwv6i6Ri1RXOT63NzNbM59SQUy7aix8Xva0cmv5+WRAxnbCxUk/mc2G3JQQGv4fyS
wgbF3cBAdtEhiwRimuMRjMn2P5Y11He4fSZeVgSYPFvQjUGT7/mspr9/WiFOCBJgbqg+O3VeGfZn
IIHwbJMba8pMOfzutIiDKm/F9r09MeP+jbaCn/yEszc8yPdu4p9Z8se8hFCt4aHDT6B+DAS5X3Pw
Q4pngwcyfq1dE2we9ydJOaF0W7dbGt5ztCCOV3cPiZI1pgnIm7k+u31QGmaMjvS2wJtdUwv13qEu
/RRrEwGJ11t44+n5YiIvmDhbVqZCxv5i5mJjGGWSMtzRwulxh1KR/4T58EuHZkAFb6J5oczAy2QV
nmEuX2Fwx2ID+iIhKMFl2Lg+T+PU24ly2W1ZnUN8i77oNfljAp7uNSSX5FddzxZtQ5U5xG5AXMct
UwgX9e/5qBlYAg142Pc4dRPjndrniDjM7CX0XCBPh+3Nu5AvPkqqC309CQ++h/DXlJE7PTEUqHFS
72KkyHuSe3nN43prRhqcMWZ35AFg398YUUxBTosmuylwItsr3ksECaXpQs2Er8aIOTCKiPPV1rBh
fDFCK8ZpkPZPrk/n7tNSRGkUbH+NWESgBv0S+LbOCq6w+hmX5qFhLd3XlI1poFQzCVdg0KkvNi90
pOOuFadsum06UFwi315TUuArU5TYiWlW5yyZKe1bwL/0frD2p22ff/US7tQACWP7NKRt7tTxlOT7
A2FJ7hvNFtLfslrYYmt1r+9/ombbiThSSPZPxnQyt/oLp8kM8tXvg8QHcBNJmbHULueHdGi5tYsg
KvG6VAra5nF6hbgR+a4iRxm8ud2je0Cts9fZ2KBaoSTdoMIDwIOj45J0U7+e0RBgLGw+Fy2OlQBD
6YqTa8KdmN4VFwH3CeoPAuNA9uRAEzwev60LL0I9JX4V85VnTQqt+h0Hdi8pNqK4KuHo/PRHGNwN
EA6cewLSAdauHKUKglTlMfIUf2eDI4Zg8Gh617Ou12cnNXl0+oEXezu7HOJCAA1QKjsWHcL8Urwd
kzUqRHMr0F3zI2+u8RxSNd9ee2oRlFwGmMy0a978kU+eW5eceMNhG1+hZWBVK/EVNj94MCxeIOmD
q87F9pYBlTDCxRsYQvzuAiVUqPcKK2WKAA2fMJZhyd5xFPinb9JvYm+akXGCxzxRxZpSC4VPY/Tx
itro4P45LCwyHFVAMREXDXK8WwSGZICNLBl+IfCC0y18wi2tpPCwk+lgglK4m45n7uaepE0E6eRf
m2sDCDj+26aU44xJG3eORT47ovmuTizbwyTLKu2S+9O0JcWgaKq90YT/V+kR8CN3AQmue7Nll1An
kYAbvDYfWRJ1Gbh0IvAvBVW0Ov5D6681/B62g/TF6GnQl0CbeGn1ZDitxOv6ty0NkucEBCwvcBMi
ynXytB6nb6cJmDJz2nKGk9CFiCBPW6gqI2IQG1jFWo4jr4MZcyoRq+bGMVKSsm6jSp1W1UldQDf+
xCOVAa6kR9oOik/FlcbLktKyW6wfNLgNdzks/57OnmihGL2zBp3dcDrAHSlW8mcpA9T5Wq5ykfh0
Epn03QiVA2OGl7CQoXpQM0NtzwQiWrJtKdc0NeZ4TclQIMyfdMYqxRnERiJMIYeSJ9JV9nxm0RFm
UpExdmhK2K5NB+8n6I/nfSfdhiv4/5rI/FWsAJZx2ZlBTmDTfYo2XHacQa8y7wYdMDbOMF1xZWJb
4XbJ6cAgobkxdmAXt8f5jU+VY8ILf/6MQsPbVQLxlkcoWcaFrcZdnkAEyMAdshl+KxM/q4CIG2y8
2CTe4jp1QL6d7TcKrFPz9d1XqwYH1S92Xu9q9pYHQJnG7KdNd0BCjBbj3Qh4npl3W3NNRtZntYjV
9JGGp9zIaRPaWMVqlwfQMGjHY822LK02UuLHIBIerBgi8jxoOEtAdebrJKGzQEJdGKda2ukDAUin
4GmdnXN6bofHHGIUxqbQKsBmSv+sXV34hMT/dpyLHUKpLOjVqtVNfwQhqoBQ0V9PPuusV7ofBpGo
noskQSaXTV7sRpawZPmkOQogH0hzHCqBjyPnKI1VlXVEpfj8c/0qUQ2L8BL4bEMpmaMi+w6+NZAL
5PC4K87i1pqAvvH7VJffHK/25pn8xysclRaDH9u/VGey4mR8eYARlc+icpqm6CoL48UlTFQSLG5d
3Fz5kZKr5fJlPskOl39bHrwW52hnrS1YB6pZYeC/nqRKG/TBQfoKZTFy23SDt1JJKOI8RdIv6dWV
3duaPehTd+42DP9CcofsDpO6GJMAy46VQV5vjgkZfIJ4A0+ruHpPKuZsS6t3zckXN679s7D/6g9V
ybTm6Yr7povHd5iAK1SLt1e9uNZkecENyvpVzlHtDzU4TJNJsKqOaAkG9nY74vqv52gU7gxCtCsQ
S137wKl13urDh43ObLAUQuIw9T6yN+Kzz69DokFmPkWQeuJNYb8VVI77vH9auvHTmMa7xeD9UCxJ
k/3u8dJgr9SovyNsqPHeWo4RtJLxYivk4GBxO60qhbBTuVHZ5NBpfyYBvFe97yn0J0C3OrL70dni
FZjIRv9JYZLdO483Kmjj8yPCdw2S7MhaJoP8vynhwVYMX2VCFZ5l83ruT+e5lg4WK/cduQGexijA
JdQh1/f/YKi9sZVQdH+Va3fixP9JVsmWOwGDjZMuz+y+EpFxMZwfvI7yI34mwjGa9jMziOLiuvrX
EG2edjxbCd//o1WrPda/eArEjj0jbncBSgzvhTXR6agiQCu89zH2JlvfOtP0TkK8mEeirwpHz4WL
1yGXpKVHKb9UcBC8M2Zexi3gI15S0AEG7AVOLFep8xD2MKfW8D6j7IaAOdjoFBE1GD9Vuj28W2UA
sAYFbwPBrrOd48gHXxpLSGUiKCa0YVXR/wmU5SdH1wSRsSXwi34TNqE0Go0LEDc4NxiWTJK5lwSE
E5oXNPm8IbPaZ1CZwPm97Ipm0KpvzTAqd7HMMPytf2UlSMwNw3NRoRDIPo9ikU+406ICmX571aPZ
SvRpwZaVdUAIGnhZMS7Q/sVX4XZOnznoVgBJJyXJ2HnFKAxYZ2RSKn/+J3mC15l2v189Qe3GVFyd
vvpKmO8bsf1r4P3zpw4kvK6dw3zD49KxSBZm3ZJ+9UW9xHGKNORaWHGPpvhv50P2UA17vbOWNuci
zTyiDC1sD2SAa4ilwUN3tLmrV/EUIxZ0q0LapMUxbV7vnl12LOunUzAxnjrQi9aTB9/TTXdxrQwK
1Jme2mF4zvWlE0II+bje6wtyn6V+S/XToKTQNrusqOjhRtEnXxjyy05IH1+7gipEvlr4Q99GTF06
L+vvlkxR96eLN4NBstL7MpZ4Uqhma4JXVKe3vlRkAgN2DezoYz5pPXURpE9wJScHuNdwPcbPjhm/
PDoXR8P6PY6bFfI+iYmC3elZz094Iu67Thfbj7H+BXP7/Dv1p1olYbVxezoEwSkNTAXhDbHdFEpV
nCOkIDgWuoEQM7sIY0ZRjHUHFRaBh6LJ2QeICijYAPKZZIMmJBF4TKf56dX/dnKKd6E8QUFQ5zKG
YjucouJtMoPLUFKxBFVAhYgHILbcdbukbAcWDs5AjDvw9adauRjBelAHqIzGXFOOI523WHTKSw47
dYTMn6EkOEaflehBdo/+HTClBD7sBXkZN43ab0yrS0QEdTwgB+cC66ClnZcURFnJrhMZf53iiI1M
g0rJLgsdJvg9PZnOuMIWdfwbFWxh7WXsKOoEyLK5j3betHStfXN9aM9eKTI39NfvvNzuUe9XxyER
qVMqqWuX775YHH25JoxkKcnKpPEUW++3EbF5FHnRKIXvaWL0+FDjSdl5Xz0SeDELKFqAJhwMvLLu
Z84X0/Xq3Lf5kaa78H77x0yqJ7OurIQmXaVuuYW3f7HBxrgEifrRsdieGTZDvqsu6/3GdhCi/20d
z/m7bVR/uRsfFi0cqkZ5rxDSdS0kScMUBL52m1IzmRkxiZUkQrVXXAeJwxFAO6epGyS5LYaTMNUi
QMfwyhF1Gv5poaTIibt5wOr82SOrfmr8zphMnuLQQvJR8r8j0ypoR3WX5MKaBRRwj3dQvR1Pz1yn
u9xdK8UPaZhDq6B7D147yhtQhNROha1sHZypZSyP9osfXGuRp31cLx//KlY+ItYMEKMLgqXNMf4b
NHnOB6wH5YjJWIOkaLk9citFkC0LmMFygr7GcLUqjGp6S5nXQm2k6yUckrcs6OoAcJZUFfMKVHRu
iAmyB63r026eHoo5/l5VylpUSuItUWdLL8fKOwPPwgNOTrhQ1mChsUab1FN9oK43OpqXffvesTl+
v+4jeVx3R0436mO7faEa45/k+H6xj6VE8Nf65zXSLlwqadRkt/KF9k6/n8SSYOvEr08DUT5GDfTi
UwmD9rbb9YNcH/kkR7ABebapLKWQgqZpyMDGDtVY0AaqZTVFIqyqP6+Vvhzaza+TjmkJupvKQVPV
nlTdidq7fBdsGc0U+C1oJ3C7eGBEC0gb7vGVQgC1BGdiN1+OAwn6TlOWyI5O0rDAmZF7erMHkD1w
fZJq6KMdZ0q9AyJ2Jf0UWdaGYwmCeD/w+3T3LlFgOYVIRl3spLlyQVpfYrXw2LK4rUuYx1iFla2D
t85N9oq6x+9wlO05cFdoTU7yal62nydubSPsSaOf6ZWdWp9hsRoaoj93MqMIGs/k1w5A49W9DXKs
aI0kt+DKREqk/mQ0Y59LYP7HH3ZXvHEiR8p3EPFJmaJ1uUaq+vIktskaZ1E0D9K9D3okaGXiGmI2
ciB8+M6HVLYAC+J4RHLd0KxcZLQzD2ANkczYmzLk3gtAutLJjgF3FktZ8mGK8o/78evIJGXUGIkq
j36Nwv3P2lQDLHGczo3iqQ7/KBAdDgK4tkiybgCDlB/ZBSTUlIy4wV0uBkeBGwo8Ydem9nEKYlhY
qkDZZ1PWfzgevpNRR24x/Y077SiFpRgAsNCMYmO0HPt4iHyX6MV9ke+B2fJYKIdOuVUnIFbyylSK
Wzo3aXWqhjHFMy37qcEL8v9+PogSL5T3vF2Zf3uSxKKd2RqAKuX3TKNo1kMHiTnyQ+eu52Vz+5Oc
d0zNfRXE+BfnJHfmO4VDi+1kfJp6XLuEPc4UD8D9HNEXuyOH3Kwuhk+4FMJjt2lUJOiGKr2Ea8l9
4qHCESOZVMRNA/TJN6EmQ6npiHNetF3e+X7502amCFa0AMMjKyNT84E1lIu9y3/mdkdjWfcaWjcM
uHz9Iq91SD+hIokKqcpIVDgMelaMuKrERhsGHhyMeO/RjYPZlNcwD/7CWtzIFenNEhlYoZ4BZ4gG
nkq6UZCIqt/apyYdFXaEPV4pxtQT2eQE9yXleXeeK5WKoY73x3cgP10ncgW+czUKKZEQGufzu9td
Cw9NrBRcJ1ClIyKJTL9sxSiwOx8mWvXAfwB3X8n88bbR9tizXl3NSi2ouvng0R4HhWZCpe0CFrBk
x3+tdIAugz3eVJfKvNF+gbIZYVeLvsQXelKvSifdikiL9DYTXwXU+HngsiE6H4QB3t9gK2RhgFwH
21m1kbrtXDgHj+wE7tHgQDYExmnBASVIGK0pjrCOPcZ+Ii01Aewhac6QBMQTBbGg4FWPdKv+Xd/f
YD2arnVzGAHDa675mMsAJwO9zp0UnjGPch2kP7jO28GwecrxkEudRZIz4PvtcHcNMWqMBn1NNT23
hXy9cV9ozdSiXr7d+eJUaJ2z8D1Q1+ygSzFc/v/NgT2aO/E1FU5VZtm5rT1UwUjQxldIMNnizQik
rKQ1k96ycm0v/5CRD8Jk7IXOUwrsMsRhcPAmn2le+pc7xvCieLNIQjJpBOy9kcrehd813pSTxT51
ZkWoOTKX4NVFqRWzScEEQyoDIYe/5VtCBCCLRn6Zkw3a7NnMYzl/WJetv877wu2NaaiGaD160PZf
sjHviIhGHyLkNIjkRM//3RpoS2Kci23bkzwehVDlo1uMe+MKSpczjRuDsF5pY5hx+EllVQQkujnB
MCyRl1hnbNGmoFTmQZHf65tArxuUa14I6qO8bCfvek37rdZm5ryUYeAbrtzAC8sANIHnJmNZRUWa
0+KSab8H7++/prt0DIcIhsikRlb3MvlnFGGH7KnsMgEeQjs06Ijy5FhG0jCyMp6SBEGZy1TQRW/T
xALd31PeyWN5GwEw2A9z1qFiCyQOFcwm5Ybf5WprHYok4FK12QXlDgnHod4Huwn1FUUdIuQAoUq7
6QIcT4QbPPhTbpYJsFkC8J1PgvLXdiz8z15RCGQOijaQZpz0C1cdmlLpnnsNf52KD13b+grE4Yxb
Cn346KbdIIyEw4SMo6fy5EUFYblScb7W3jQs+VpSWJXueZ9WnnsXLP6sm8vFhvJgdJBJBS92Bp+c
56HAxLox7i7VXv2T/xqF/izcmBI93xLHeaU7P6NJ2tTALSgnF7DKJYhJVWOVOtvZP/j2YGRd2FLs
+8QJLWfnAv9uX3sLmU5FHqkyAr8kzVMBSizcqQtRGfjy8hnnJIij0G9q2s2K5ihNVVv4oyWyAiwi
jC3d+txHEUHmpW4/8JAgo7C0941RotcqmLA8RsF+FtVtq3fyChxDSp/6trC13QCWGMjApPY8zhCZ
6TFilzxDZWZoSBl7/kkaXuayd3jaPTlsSrz6v53SzqZ3PWr1lDdvnfmsWsyFk2LW7+Z1Pr+zQNlA
ivPlFMrvpL/hUohcqDiLWKHircvPwoYntF+KeXzXmiBN5D5joe1Ob5bO8JxyrC3TPl1kMnOAVCp7
L+vOGHfLcsb1InnLZBKEv0yUm5kGCVvPpewFKhvuFLj2tWt+TeGQtCMk/VPWvV+Dm+v99KG76+/f
0kGt48a3/DeZqTOl8hLqHWtqHPfaK1HlnqUKNBgsF6wKTs0zmpeu2vGaAVOpB1XefqEsinv1cAdt
IZOOMN7IRPWxrqFzJJhibyuW77SfQtTETxyx5TEJjGkj7Bu1+b4C5UewOr8ZBvv0XPg33cEUfyMk
sMgGXb76iksqIMnZxEgj/C+a8CinVbgk6QnVbZuqYxWkM+Ix+zoew3AvH/TGdTFHsw9h1BT7dCix
1dy/eaJq6H6pt3MW7Ahv/iU6JGTYpXJ8auhwtfN2awV4jsT2+ngLVg+RJNugbXTUTowA9drVP3mG
lESpPNjLgOrGES0Yl7OCZk1N7QRS5DxNg9thyXI3DDHPanTusTb2DCP/+4jRq9B+SDaEGXY6HBW1
9gqcPSAQJkmfMIDbO3H9dDWY8A9zUTi1ezsgtJQDBDhY/msk3pQjwjyCKYxyvSBzdVnXtOtjEio6
Q7QFoquF91l4PCs6UfOOkj2pduNdIw0gKXibaz3kq3mz5xCt1LVmifNeWEJsTaTfS4T4x2lMrPXO
dLoFaTc4n1MfHqXZG8jiFvnirc8Qzx5s8eEu+58sF8sKBuwdHvrVpEuqj+3qCF230bmzXV4J/MhC
lqDIRnE2C6z1AshERsaALLYOoBRPfYIx8icjj/9D66fLSNRtU0nJRmhlcSfCn2imTPdCp6cGhNId
crJb5ZTZtxwjWMUgC3edY7HDVJ+1DqoQNi8ACT7iOZDitAnc6hw2C8SkM6cxJdbIxWyhSierfTc/
SKjjNYzBHOAJic+h7kaKiNkBXAME7bmrRypixsBI4SEf4Y9yyP0exnPemyEc8QlOwsiWdwomWx9Q
/XnCIzL4/W4ksSGrOOcjTCwX/skcieR8L7o1FCYGTY3fa8D/kr4yd1Tujw1eoOQbC3MVGXyqi9CG
NFJ7Q7izDGfApaDRDLlTwLrkzJB7ub/Pmq9uZ5RXCWuEKJH9xxPR2qpyyutSMPjtq99Vj9s0W/eW
XEMtnd6x+DdxyiqAzmWA7xi1uIoe8blqtDuTSzY6NsRaOfpPLnLISvrlX9mWCNGIOTJ+ZvOwgVNA
nFQtjk4n4c6vR46swVe9saB2DdcSgDA6ELWq4yjZVeDVD41YEisXQh1zOPJeALrRHRtskljXlLET
BrxxNUyrLGlx+9BgUaePKlCMYksZvSLji/pH13D/JLdSzhWM9QfMuuBhvueP7eBQppHklCgejwdU
NZkuxuQ8rBkRuGOCrysTx5bMafxcQkW10cjpmIG7J0gtdFtFvyZZj7iYdhxvXQWm1nIq1eLfu1qh
6w1mfNAvIHvPUTY0UvtAIYHy7dK01kZnstTi4+Hk/HbqrtVu1WCS4XXAPdjjhGkZnCl83fv6zUeA
NFoHPov03h5mHLlCirRWrvHajp8DtQAwx3xnBxJdfzA8Lof5nhqnfiBXCM00mJpKIj5Y6PFZPhyu
VQe+xdky97YfjYDZi+/wu6IZGjehmgp7e+iq+As4CfIe4pqWUaONiN7ZEeda51DefjmgZywBAu5A
+g5DtdsnojshOJAUZI8ekVpK9KHtWavi1G+ya4CIFbF1qUsomyjVQqnBiJzpuA0NeUoktVCTb/ar
VfU/dSSLSB7f1S4BKmaWxYM+smoJOG8qKtCjZ4Vh10Zr4SAgHjnmDdbTzjNnH7QKtw2Oe9W/E80y
Hm32KLSSJzC02zYTe3UAp0bKnolqGaZQbXzsBCR1EW8mBgVOQmTsRl60rioKW1U1rhVawyfp2FH9
2wnDYKNJw9yzfsdzWDlu5uI15+ZBvbylNGVEAxlJR5tzRSMoKr+C377Mq19m6owi1nHj3GJ+O1gF
rpIfRCgmlxbH35oyqCALol6DGv1mfVeUT4MY2QjaWeX7bjICLtLzlXe56j63786M4b/Ng756NPyh
6g1nmE+fVM5zpfkcXEEz0ltDWStHDw1ojTuWRC70m1tqe18WEfVo6YBDJ8BFQ9ajQ768X7FsxJ+d
kIjHZHTP43gAYDyPmaNm9Ua0wVfi0s/IeaeOTu5+0VcKfGk+1stoKZSUdjiPU5tFIA3qWKY1jmdm
xhFCK6Pl5QgkNPitJswn+iQIW02n1LE4dScIsi87ySXBAjwAODSIPQPM72/WzqKopiXxP3oyIORo
hHJ4u70Hi5SnSvY+aZczgUHt4+/7ge7OL4rYWdeJc5edQZcoQaCnmqFVpHycb4/pVpf91oLHbhzy
SzUIhHA4Si2JuEdhfu33XlsBCwf4Um4u4QD/JL2Fe7lJ1I6sA853X1Z499lDAmFdfRPhYmLEwRuh
sn/KEQ/3+joY+w+CQnZ9Dk+NuMpMbJVv4VNR5MK9poBqcI2OTk7XtOkVTQLvQjgWh3e3Q07x2u67
W+KjsRVhKc2gtWk4DQ3pXR7JQxbDBJxrN1sKSng5pAz5IMF1Zsnw2TKX/u+lnq4eXNr9CSvBrlpZ
m65IXkd/um/mteefohGfWwrY1IBbCzrUVpulTfrTzGJdA1IPVMBHmYZcYqnda8rzhssPGxayg+2t
ajzuioC5T8QhrnYiYf3mwRWXYCIKCfGWDDqZSEsbSkmrturv78RFImdxohd0y35TCVkOXJjJW1iy
Yh86oQ1BQYZJO4nVfDdGdSh87LVWiyKLk3ad/4OcT2H8uovEQPOeL4ZiTlD8PFUwPcCUT9rLQ6uG
40ZbgrYtj6r6v6fEUM7/fiJB/uU7QoG0seMSWXDYuJZOLK8LMj2y8Q4WzFFPXiIW1o/rUaVWixG/
DbvY48rcdBx1E7t/dy92sel+ddDfmUiYoKalrxvF10EiP8OddYjUJxmPUOnhnsYoUl7HICvlCDEi
GWB4FkaEdiUt0wIqkTKju297scPx++OZFOW79gkubaiKZa7ye7O/CJu0jzKPe2CCBEOChhuzEV4I
g9l/u0vetc4woJXt3Xvjm9aV2pLL+E5ZD77sjZ1/hc845qhymsyf05gOkpFnlwsZ756ahgq630h5
oGiiyV6k2q5bNXWJfyWUQEM+obMhL+wXYgewGOObwYOFjGRrT9+qUUZFWSqN6MIUAzljS63vU4SA
3SpPjdwQKX1Wh85Bt3cX0s5UbDQOCHZdTEavY9KeZD5uIRTBfD19GYPqFLKHGSW14WDB5/KayO1D
667CpiDNakM+o2rcNGL0QJuqN2mRN53GcQ+aOPU0wIGiPWQYsXACd1lLaVASVP1Igp1sHQnDuGCM
QjIRpxJeRYNGTeBETfo+FzcXD6uoyL9ShyqJlgluYy0KRJw24KnePKJo0GGcaJhxvxe2wr8Mx67q
YI7/2d/FV/rV6YT73RevFZQBdigYfrtxU5sIWkiWUNdwY4Ph/rSZVH6x5BsO5vyqX+/NcaFovUmh
QxyIuT62Ef0HOAvZG2wULy/UDYO/KEG8vAObbt3MZw8EYjTNlPFC6FTjf5W9TtihQDUc+JM50BZi
nwsabo269QNCXulzyKMUoiRml4dZMi6VAKv+wFtaneR6beoij/qA/exd9dYDG/7n8osoKK5KV88w
ZtUC/RD/PavRZBEhKvf9x6LJcCgCZxHVp17xkT/6R8xMqm1VZgNhdMUJkK5h2+yMyRl+rQyTqClm
ZQEClew3olz2kidEmKpY0dDksqphBJuUhMyvMoBp2evrsFbXs72wwtUoPra2WWtlrEDpfDm2oSKE
eiygncyo9+PN122Vu26ff9nGrIcoGfKHvx6sjcCuvv+CStuC+KIcvfSOCJCYzGo+R7DE7aQI+nKX
tZAv5gp9JtTJrzyc/Migj/qV85DSwCKoikYx9IsVryAb4QIvYv+qB+19t+HWk/anj37g+MPE8zF5
6B/izbstdDZBBSrBNWL120ATkhEYW3DbGD0yhym1bW+em508IJL9voFkhE7iJb3a/bYbsrds2kN6
2aIvho6W60B3anZUAiEDY6v6cHP+wiNai3dWYrwxm9xpQSDC82pJQWJgcNlRDaFxqshpjg0HCkjm
YgVi0N8C8s9nSiaCqzYrmPX1jPEbJR3Vfy9mu5tL7XLLyBjeNub14QhvS19UhC/0ttD74NAwzK1b
jbsAKJo39WX75EmUfq+q8PiaVs+i0kuP2ewJ7ZZKEHfLb9RrUYfsCxRhNLjfojLBwilSQfndta4d
B5JorqjKmcAvcqRWZqqmC6UdCQsfrshINkYtWcTy1/PMVtWzwlREjw5xNVW0u7WLCJj5BhXHy+PA
PinHHIwn+w8Sx2hsxdoATzAoPK3LLZj7BEwZKAal6PdX1/fQFs44LTaWbUIChfuwjAgdyPVniIIJ
apOOletHj9QiQ60DzNtFRZjEKElN6UHbJAUCDNFqMF/dYvqe3Mb/vPiG+I+tYl3qaXfiquLV2Zh2
BDtL1BqLYsx2eCH4dxyRyPy5hTwxpq4lT3IN74tlsq9VStQ39js8bXx0Lq69R920VQtGR0CqxU0P
mhxLyAp6/fmNiDvY6M4AZhNbrqGJzVoqpaqgl8vl+Q3JhCoxLbEM8mAgQv/b2+s3irbXKy9EEC4A
rJz6uUmph8ssU2Xgoc8apUEBqoCbxsCucBRTcpVzFO0NzR+Ptm5Q6qUS7m3aHlVd6/lul3XzIpzg
YIcVZYchY2L/H5y+R7/azMprwoYjBvOMPh/7tgKgLQuPzjUh5XKWF4DOs0DqiKxIPMqMTbJUJEjw
UAYoKanup6Zq3+9wA/oVXr9gCDgcdfiQ8ubZ3q27MK2lSV2QNXIgg9V3h/WElMuM5oobYQyOzPQ0
Mpa91Re/OEWJC7FajAQFjK2txsnQFckgdS4MMkI0xyVkAO0DXwPoPZY0lpN4uKr4W75UjyzE8kLt
P7gBnimjyRN8Xfbo5OiZokCSdYnOikkzDr9xBhKn4/4zE8Jhisv232jDhLwBJjPQbIHjPCp+tYbo
bg9Pw2Cr2R777Zsx3EUmJTvRq138iqAFLIwxV2cObcwvnaI4GDNhdksOlheXfatsYO4o6AiXslyZ
sqwEtafgkexwr6pb58KOivcGaczSNeCoAuXZ2nMqmmwExwP9XdHEyeqWzqkETbWURtZrjT3Znh97
CMBxGZfAoNRfb/txIkcowUVpV8lpWgtu8R092vfp+Vc9tv9GyqnXvl7rx74hRt/V74luqQU0egc6
/lalyRkdr23kBotuuVZzYKabZLZIt59Og51DKBeVsKVUMjRbvzsEPuH1aQFr2bOenLhIemwQVQMo
6IB82ky9C4Qagol8U3LgdRjTH1mKgt936hF1PmpF28yinlq8QJIf4WPXBzMo9luyzGMI7uTcvAUG
D+I0qJ+UheX3LprRCJwQQO7ntLilPMFIGU7zVr4ut0dz9ww3PyUEESklPqLpPDJCo6lji+JnQrk3
gmGScmneDVT1WJ6B9E5LQheO9rnfdI4UyDn9OP8G/CkLr01RQieQ6r/7qy6yuLR7x9RJMh6UwvmX
Tg50pf7a2ofXk5RJoRC0TvV2WrgMUz+qmNR6wYPny3l6laewHKUKuE1zjQdqeaeieg/85MA6OBCX
EMhY7gzQhBCsOt0JEwxAgvgEHXmWjWl3l5rrDyjj3vHOVqQCzIdYwyuSuMiskbceZTPSGZJoNxXA
thrt3DQuWNzk55dUX0uftM50jimnJkMLzZDF16zC7zhZqwkCIoK1ZrzyQ4htLOoeLBVl+Jp4YtFr
2wqRwxaY57GijHdxds0b3BWrzs9yQloHXr5stf8OFI73dJ9Q4m6jukGqYsPro9staXiRQAS1mnYY
NI4bkVQ+xYrECoMqAlSOulzT2YQ5liD6gFsVzGSJl81xxgtwLKe0S1oY8kkC+fW61w08rmqzbUBV
EaE2pYANquUk3mUh44qul80PlS6TndbXHh+/D0r/AKUI4nbv7YHunS800MHcbJ3GVU/+95npQgu5
AwF/QklSLaIjtNQ76fSnz+nkWYjZ3L/M5h+qcmkphUhZfVQUI5M7rqSEEZB1SrxzT3qWUBAQau6T
8XPtQurpkT0lt3K1NCY+3sw4GsRPShw8BrvRzo1C5BFUeiIMRwBgt1PKruGbVvhw2YriwpsArDhJ
x/HHqQ60+wJE0lDzRoeqc3yGOs5uoLr4kpnzZtL8ggy+m4es6k1HsArNKOPwalht2dMXsLSGqWzm
DntQZ+JiZx83L49bpBC/xyz1+ZnyKVhLHLGMhXoLQvkkctJ0PyXBhe2wU6++yxpVk1vnKaqoRDZ6
y+WHVRSyXaSarEaKznnoHK+i1T41cW8arxVTg5QqyMleqTssC1NJ+suDy+/yIacQcIlhU5eVKm6K
OCJ7zxIlI37TBtz94ZTwoe8g24N6DgrXkc6PS6q/XIeE/Ki1RiABbY1UJQhgckFgt2+q5rhWZbUN
tAQahlb96osDKKnjPL78nrSVr9/Uh2bBZxRmwJOK4QMP68H0phP9tLKXJ/ixHTzGgmM9YdKPlpQS
8Mo3xi3s9FUOhqPCgkrKrFAvxzEKD/k3+6MRD6chbBd3Jr17MzTf3zqYomb1F2F4gOvJ/4nKb/U0
lu+MiTGvtnE9n2Jud3IjRcSKknPYaLw5Prtg/KLgAh0Qzpoa0zQ4XAVianpfZMnwZhupDYkLBiOM
7BErZhKBoxZ13e25S8YRMx4Vw5l0bxaQAPC2Omim2v0y7XWNnkniqCrpoxr2rB6+2EOTPdo70Scx
cu1Gc3+STN02TI/r61Bv9qqCVhwNfTman69llQdtIi0GfiAds9r9zJgXeJbOLTr78znbOwI+6gkM
Z21d6zX0J9f+eZBEcs2SFkm4fGAMuGVYQSXeW7c3yoNFK6Rt33Dd+jpB//kYB9tf1hwAct/cZWBH
M0me3YAXe5T3RYdjLkb21n4dUS3cOvKV4TarKsikkLNUDi3KnOYRXCWq+C/qq4aFJ4VBd9DhTPKL
4gTn6+hqQXr7db2rW7hLYPazWnYti+Sh//YniDXi+bSciRS+ZtQqZuDl/oTm3l1djbqALR8Dlkf0
tsnT8iXzPLI6rrv1YQvNolRy7bz1WEq8p0RPs8XrYcPJR2USgj4N3EjwpY+DfXi4wL4i69IJBq1i
FsXshO4XQSBTdEctyOv8Bs8XKlgHrlY6MxXENbVh70YhKqsQDe9oVoEVfzzZ200ZfcLwJxZDP2Dx
aa68T484OCRZFpr6VhjMS5c5NTZehdsrfKV28E1w0TKTxi+6j2ZzR1Ali1EtW6KuDzHI7IYIVNZL
9k7jakilL4l1ZMKM3cX2fJPlCQPqROz3eCJGlj84FbDz9xlcoXPPKzuc9IoenJJvaimz6g67t/9+
TMLL/5WaioQ7YN880E5tFAnGGPL0l4F+gQAmNpQdbF2qk2M1I3gLbyEcPSj1RvXdIJulOk4NAfyU
qGi4zc0HzkK07VMzsMynxJD0KaU+RqO3H8rnEqlAvBv/Bn9D+OCIqM5EeoKL62XcO9qKVCWjSqgY
HSlk+Vlhql5FnGKPcBLUNbaxm4moAHj0WDrvi60D13Zq41Bf5/i5Y317vw/jJiTz5CBzILXao7C2
TwDFpHMfLRq2jp+S/7l+tSVbmbP4sW4hlMf+cePWJ7wGIV1/0XFr+xopkIpUn2a6aK0E7xAS3+KQ
Indi+cYoA1VnVYjQVJ7Gklhmo6u4uWENFjow/oXa83ZYrjQKsg3L9Vfz0NnR+oJBP9znj1R6/5lB
MQR4L4h9kX2XbKMgy2suun0qeRtD9hwvv5O6I6M8wgP7kAx36CdSuzXuYWrvXhlzS7blDuqDb/OS
ne28InNk3cI3/j0g1IbgLYjb0to+9Ko4KXpHQr+888Chp7feB7kN2sN3zN+cU2111d12nXz/hp/C
ABr+pl+rZcfgwQJearNwGrLgiUAIAfOJFnG0zFQnKkF5NFevi4RO+vndVvjKRqvRsWwK5p/vQ6o0
h9kYkKrGvzCWRGNf7jCsA993O/gfafKNxoU+jOUwAy8ZZQvq6gLMdF7PWKM7836QhePf+I8JPTWV
mHgqu0XpNQFLkKjFeW2jU7L+j/IUIzBkVZqufBKbDYheHcmKEUWRjlggH1dhi+jvwey7rkogYvsA
NSbL7vC4e4pEclW26h+nlEYapkQV0n9X1X+U6kJOs/EmccxmZkJjzAh4N29BTnpTtf17oXKZWmrI
23r+1qYNTT0Dhew48Xa20VyCVssAK+4l/KuiFPu/EKsHwqOyX50SFtDiTp7ALhOJjcwATRdeLPPu
Hpu2vPN7qNblloXc0taA9zNUwFn5on+vRMlQIXJYF6CDynbSaX0hvqX0yC26O4HFNxVucQfaEii/
mYftr1JLOIWnTA+nViMfsQOJIfDbfqb6fG3Y3NQrjp7sRWO+ou8dDaeH0HOkimwNxFYMCGiWqp8p
4fnMWKnJuA8DWApv23+2f8zpSQQoQNYocxvc5eJ/GcDxo1VgaB3cyYLW36i1kfmbTxpydhqe5b1j
uz6iCQAQe6654QRJO/aDfJ1ZpsCx3P7gFmFdL6rpWwEq7s3iWcks08Dl/LcjRZdPnUKQTkoc09mn
wKeZNzt66y3T5hXxfUzc0c67IOW2IrCKikJVXA4tYZDessUqz4eRr6c5tloc2IveIS92lIzb6q/u
k+e7Ja6hw6VPfX2ZVt37ky24CgM75GjtUixeHLg4Hh07XhXTgCLBQPvgK1qIW15lb1NvFHfrQ7A+
r9aW5S/NFP2+2BqTHHwdP3lYxE+FJ3wzrMrHZC35n1YS1XN/fvaYp8+4I6rZXRjVhTg5cOxUoxPW
mbp1MIZ5VOzLelFCr6ipYp2AHBHFKY0AH722lUtKM2YScx0RhDqA6lljI52Aojql5HgHPHEUTdWQ
jWuCJO9CtK4APZVgULIekSJFhWE5AWtO/IJUqx8CFoKTHyaRISyTi/9E9sYTWNOhi9DcYWl2qnJU
+zm1rF8y8rHnyOfPWgbSn2uyVXnWxTpk0Uaya484x9dG5owR3S10DnHBf9ZZBm6369V1FGWIoezG
0JG16b7ry57BRtsU/gleYsqTxZqfqH9mutzr8+Ucj8ToZ6+ujJV7LJbPV6tVhhvMJmA4GmqECUys
RjnBSdsHbII8g2307HWGqAO4SvZ/OVfCRltLOtKsqdt60HFZhB3SMur6CK88Sc4V8LaoKlipyBFR
9myN1CYyQYWGNk3l0IgusTb8SeRfDQuMxB4VxdFo9CUBri2e4ZAUuQEyCYaXHPGYl4vBV98tfYVQ
vgJhzXxp8rFG/phIaR0/FiStYi7jVNcezgoHS1iQaGqN6bHWX+bc4skN6/mmynCvUawpJ+grWVpl
Dp6FqhsXF0fX8mL5Jgd251CRcmK4kwSkg0hEqLlgZUhbC0Fr56H9s1LW+d2fEk+RqZ0DwxlbIoCa
1uvtFlt1ic2flnTzy2Jcs2P0lqhhhgvibixYynw26LNRNxR/GU57ZY9KhgDE9S2/swkqx3Ynf17C
cCBbX9w1/w3fnFnPmWpAEVxC5k4idHERMEYoKhikGFZl3S1UvTtSRSaswovVLA6rHOLtIL6uQEIx
fl3Mx4PVxYVk1oA0cV0F13QNqXym7063GQ5cP6faKSqOI6IBAWcTwYx+77kXfWeyTK2Teu5lg2zc
Bbd2o/6VxW7U+ARX3c4VY3YvvizwAPIHY0DYbe3xLcwf+CI42vdr+XD3fYDhziDOJpGyzRM2gr13
FY4MzJb8Vkl6x0DxO/qYFXn+51ASi9Eojkq2cT94vSR3kNeoWLEmTpmu3NQn1Fok/YdNJrUcAOxZ
rlTzbAfQrMtn4rw5MvoCn6TljhKMu3mLm2CvZeH6h157tg06ZWJmastrBa67nnduRdl9FOfVFVUg
muklimYFeeHT1g9IsdzdGrbOFRSs7CLaE9uiiFL1glhCzU5Sr0gvSumsi/EcuC5bZ119u+5UXN4S
S88aXS1TxCSMgBwdpYI0bNUXJw8nPaA0rXNVUBlWlg2pBMcMrka4j6eQQwZodZ322hSxdhVgCJ90
0EdODINKZ14I3/oPsBk9PPTsgHiGmPf6bgtAuCFIfh9SIEdQpYWI4hh7gwqdp1abRC/RqZTlm3Oq
S1WflKh13E3OLa0zA4bXc8aH9amJhs9y5tLtdb8cBesJSHaObcRHVbB0unZgY+V9nXYjxm2M5c+Q
gCAlwX+UuMIKWv3IlIYIUnG9C79xKkjTx6LByrW/is4nw3kVJqE83Lj7wP7Txix3s4V+IRhqqivQ
xQb6N8dfXa75Yx/Fu8cO6jVOuIEAOZTziZdSRQXctFxfzKs+y4+9yTZbO7OphOMJjg3rUPe4TfGR
kGTepnKN3paWRnPqSwKdrX5jM5xFBOf0tTtPV5O0D6icPvoByopWd1iL5yjM3KtQHuEGdnsKX21t
2qcx1Qzt7qSfnrZpnyRE024NMxz7iXDQljCHiKpfouuagNpuLIL9snedvoKhipfnaADTUc+xYItX
Q3vu4qS4uweovfteBRB2JyU5lThur74XqAXoX/4VeLe1Ltz3Xf/KtBgHwq4kZRyreBq1mdTocvKV
XmngmpNFfRgXRhNdiJLtcKjZ6bo/zA/kyjbGIDa3UFav3iU7XUKis3FCIRZhtprordALuUtuLKjb
+gpbS+2ZelKgqkKxRI/NIsMVnRUvlZbHozexwX//oHZ/GJrAVtzBXzfLXfej1j94URP4+AREt89E
S/fcPIK6jkLgtryXlJAaX9SaEgV4i88JvaRFz9evyc/9CKWILsO+wsRAKJDMQMWeqNxusv1auG8S
KAJ90EUvSz2+f0L0nk630aq7TQSxd2H6GnHnRpdw0fc504OLDQsnWrJFe29VOa8A+D9X4JjzJjJD
puTRTb5K3kfl/Nw3slfTMwSwoUHb9dWQXgW49TvGWkhiRShAIWZxhfjQsIHC4/ocLIAXRlJTS61O
jttocn2RCB62jy+fl9lIN0iqRHP3Loh336dd6x6MXmVXltXpCkYG3qVMqQZRjz3uRGuX+PJRULLb
eB4w6lYOlpfFFkWDbCxrtJ+/OlxVgwYMBUzyZayns805BjXGivmG8cmIrCuG08aICnEyscwm5Hpy
8NgfCf+fZfqINkI+x6svaZCAGsHpJ5kWqPl2DZxglWU2Rpl+EBTVuyvv4pY/Ln3URUx0dto27rlf
FBenQ9hUTPEkXdI2L+XvM65NVDWizkKp9K1oaSrgbEYhyxyopTlUa5LTP6fmZtKpCdlnKA3XiIDc
9JgwBC3S9TT4rzR+HcDXHGf1pg28I2n0NNLe6D+oWXwoaQogM62YnhagZv3ra+4mtTzskC3UOHES
OkkSvK9gglxjTf1myqCjtOV2iOiH8cZaOUpD2oEl53eFxjXqG08yxdCTJVoCjarxDZedjDXxkNzF
5ilSpmPR5kLskipbHQbGAn6CQwLCVYJM6Y4ofXRFtNrRb7wAVfDtJVznLYtENO4PwYAc1elEtYnj
HR6+CP7GgM1RmLP5qBm4ajRn/ngHtXcPlcejFELDhImRjUX+VZV3w52s3zJ/xPq9x2xptZpgbJ17
+vpWiEq/USsESpRWs7aZxc95fENfMYIbth3xhq0GjoTt92MFpB8n2I2Qco8ddojlVmOkO8H/0CA9
bI7VmIXO5qRGzyBMVIxcBJLv0wQqPJaScPGjc8hoSzf0Bs0THrVL/FBnc9EC/CoiH3sgydvepvVY
n6nmbOWhTGcbRpPvfaFg3t9QZ6TXSvaB12U9L8pr5hJQssyOtt0TMLWKz1lfn+vMo36TkmNXSTyy
tufRi1eQfNe3d6aMAD/rb1JRGKs9ozISejCYvH2zbalNJikpGMX4LhH5g+LdWqLl7cF1gznXSkCP
ezlCdvVJaUaEkwPyBMKT1nb20TVy/Pk28c2q94gLGPHDynSDj+9GwFv2AcdYM/jNjQDfjxK1ZaS8
WDlg6Z0VLcl7hbcWL7sTfA9teasfESwn/PMWHazJAxwd66nmSbEazl1HfNay/mc4uO7AO/UEiUY2
m6D0HWQxz+xgMIch9m9xsc9oUxrjgyaClse0LhaSis8ovDCkfdAYo2Yts7NEXD/5JK5zK5trkrGR
SEz6/bNsQR5AaAis5IOaHJWR7fZoHZF1iAHdiIQ7iNkaNiaKpUd79ftVg/g+7ec/yQIe4pWBh2UO
AzbZoGcdlRQXhuK7PrlHcBWwlm4p6bwn5S3gdSjixN7iQtwbfr9gqhUek9ZvPj34ZLiKy5kjuCXD
VBHaCKcFTNJovqSzk03ySzUeT+49pQFjSxn4PMzXoGIOqZFUD7WuL6qZ/+BWGGOeGQaXOQdpxxKg
yWbsB7Nhl2xPypaC7d1vzZPoF2g5CDxBgMbsGdM6NRT7LP7usYDJqwDE0LUQG1pEYGOiiDe2q6Sk
XZfxj3BWryKiZ+LMc2l/VU9xYY0O1tuRLuojpW9ex0SSXf7IOCr/mX+Dn/w80jxb+wdKZ60+yCx0
RTRtbI1nzi87kbQVi/SaIZXy+ySwtcq6zcMGbuw3MS2vulkZ8IYg/8V1Jbb7zLtf0UxUMmA3qFPu
VMy2TIJm1s7AfSvtu30UxZrF1x5Q2Ge4SYwcRqwCsX6+SKYGUQtwjj1ABVczQ5l1dWII8Pib7VQd
n3JC/d6MPCkURA/lcWuqmGztCeNTEQZJ5kci09MIIlkTgPury5iFKdCI75bfW3uuy7+pfm6ASUsb
vcTtG52za5lU83j2JGj9ZqJ1Yj+TTHKEwhTrga9C1XWE3WItbg0wFSXV0hTwkK1zd9qsuVktQDfb
mQ1jBLizfN2kkRXGiyVOsm5HZyvATouxO0eMO4yzG7OMmKKyxdPh0/qM+WGWSrsg3ETkmEFQyehU
qqV+9ynxYXqhXMI+1V1GUtU5/Q4Gaf9j6D4u0xthP7bDdBuBVDpLS7VacH1fStI3UTMk4Fj8OWgC
r+6WXTGGfmly0RvI8Oe7h9XhAbQM5SFnHOS4PcHwMA65/j02ylkEcCQSD9LewftcxU+fKLSmuktQ
OReGJKu1VvPOGv5v5MjHxoKEbzDAeV1K8vbpYxmPq4QOU5wTJjPhW268qyn1KqzBMCzVEVT4cDhO
s7j5Yu/WpQmbeTDowypZiWQPN1QfHX0wrL6Ktu+rS/LJudE8OVzmDZ/qUdLpVuMO9CD0l9mTlc9P
u5tV+7+ko4V0VDXR+xFOwtsqNFUieo+ER9nIvUL9WNZCOJMiBlmFWTmDwqs8gjLcyp7m2ekhZahL
16461VQGGbUQSU3OGqnxRHdRUEYV9c6aLzmcXywy+WqKxE4VxuowIgjQ/zwSmw24IL97jdtRSHzt
q9K/ofKSfFWUPckMxpO+lnpT569VkvD2XkgNEVNQYJ5y2biivt6rzYOHsgHpLWCMbvgkp9MrmUKn
IgvCRGaaT79NcAWB5rhyMS+cKnABVM7IURKDXnELhEg2iHDRiLQhaMgpc54j49nQMkWXSG49biRA
pDB8w6EVwMPGMuN7g6b1x6EPP9ApfWciKp49WHOKjqHgfpLSDMS8RZrGzjSOpPwS+A49LekQfHFD
zwNjbWIgbUwCZNsWhov4i9H0G/XfvupcLO2XKFlMNCCfTKEqvZ0QOZ5PgqemDUqplVX2B2BfvUwI
ISm+CzEYK55bpHi1Xk+Z3gubWhY/J4UtXuBhSadtz/4h0eEcqSFmX8Pzst1SyR1KyQGHcH40QaeE
KrThxLJUeqIZ9M3bEJu6oUnyqJrqcSFRLvlgp/ddd3dWoKXx7aGo6EJGokX2YB3/TOWwIAD4FUcU
yn4akqg5749zREUkhtpF9sURPmY8zDYS+qKJzWExiKjYPlGEcqrNPz9s8mE7uacdP89sCTMR1Uia
QMOE8aYkfkLUpq8bT/m+4ZTCClM7x24/r/yMLt99lMB+1CGwWR47/5WOf4a0IlPeFzZZj9Kxy5AO
BTc3mvSRMM5uNHZWevvrvNnUyh4RyZPfHgihdkt2aF7JrrOnSJIC5cNy6Z8sxAAmZ6AgV6hfY1QP
1yy3yFRSgidgHNCjhixlwd5aAuhZfXMWg8xM2t6NIUvB3rKfHDUuSPzNEETuEDa1ut8Zs7Pn6KLO
b1cAmGh/AHmqtbLgtg5t9rGGurzArC3L3byhRCnQVmiWVXC61VPZakiM5ns55IBoV27utH/sRzwr
nubsE12z/PuYS2dLo5P6vCaFKJ35hEPmwHfWmyMt9o1xC1h873a6MbvXWpacyS+9FUrILXIH45JQ
Xlhyo1mFQ4Yqupze/9VsHRq+WIH1Oxsmij5CRM7w77ZvIrSht6K5txjJuCnb6EHG8W8c5XSrEVc5
zejgVkrVOFrrW8XTVcAkT8kdRjh7FjHmIANdhXrcYNDzM1/q8YZ1rsT3vvn7J1eEw5ladr5OsDvW
T9HCQ5H9jVb8G2+u//jT2NbMDdyDJ1FqC0f+sGcWTdWSXta3s3JGGxiwOdJmb5wsPzyUyLyaZeyV
40OU+0zYVVGF4cLpsmwu+R6myejOdedxyBFw8ySzTVI6mOks3v4TGtV+cB2aWAvxJ5odb/Y9Uxhs
lOoR9DitjzXwCZJgrnHbu3+E4eeYwDztHXy+DRZPBqxguV2fQwCp3eGVKNYdsRtbb4UaZMQd7vvG
GDM+KIDYzjmmkoQGV90Kn45D9PampqDbTu33p+jVhM84HHzd87Ly1f/sjvBqHEyY04SuWX46bP79
b1+4cMrYWwIVjgRzrEPw8qAmP35hN8btlHaa0h3oeUQTYQGHmSosmsIYJ3sLLlbg8RyD2ILHXNrU
Ze3PS7pxhXQ89rVTMNAvnCc7taL4GxPTCgSu3H4NFKPGxG2eE1QorH79cngqHxxCP/T0HJnOb0O1
yJsF+UuoLLEngVJHdJEiRBLwJUbtI0Rh+U3EzLbHeSUvq6UI3gONt+P4HkUYvVGMZN8HJfq7cO2+
NzrOr9AZFdpcZOx67n3UQ9wFjV40eYhNq+qRkLj96vRSiIPnOBJSkBETPNNCXJo64iq1Y28QMuqP
t5PgHQdFs1UBCgjK8YQDBkLRSubqTzyxeYF2W0BFC72GrbkB7JD/qztMBnGxL4PGQptCO+LLxoPm
VYj3SxrKtZILPKMU75zPXDDiP3lDrju6rFHrR2O4V1G8JktxO79tpgDe6nQg5XCbP+xjwsAkp6tT
0LfJv7vGD8XRUTpnPCG4yqS9/LtBkvJ2HfpOYNEG8e4ndhNKWGkOj8sEo6gaC8sYAmjoP+uS/63M
2D6aa+yn5uG64y/oU+ja47EDf3WitQ/O400JyQ9H/HpwrQIdnWXZvnbM47usZuf6puh5V6oK67on
EkazlpYJxvXtoCDXG0nmraWRZxLMWRFlZZSU3HlFQ5Z1q3tFkO/LLxlMG3YsQXWqgAb6KmUIfEAx
781Q9CMTUmDcTsuyhBFM876eC5oEOewllp43cqvdjM+wUJ/VUWh2CspXgUMjn0uZx9iSMCFdizKb
POrAzaTipSfcZI5j993a1Qa5Y9HM0Y9cLrGs8A+dLvdkcTgVCRPppItsOT7j+zYp1wOUscR4mtGL
z8QYTqy77oW9RAY0i3/0MMt44NiW45+fevUmmqim22yOCHnURVS/uTvJP7xYzSpVWC2idg7okG2P
CUkKnPy6Ilkle24cxRezwDhSx3LUeqUDGAU+uakRca/wvd0eKGIf16V/H3V4V7wqFAJOwLgjht2F
CvbLsdy+T+9CfTKveJyemUZoPeHSwwuPd1F/EeZpZQCoa5Rn34u6m5nqaufXMFE1pYheFqdCN3S9
VvIeOZxjMsioVUQmL0Z8VXvwAlhKL6f4HNLlfagE3I7Ysxy5rtZyv8l6x6DQDcEgNfd3tjsNhjUf
s21nzM1bLavDUBcCLbWxZsg2pSVZd9HhR2tHDylyalJW1nbb9cxwm3wdfrBB5sU0mXtq08l4A7Ak
Z7H1SH+F4uIxSWOj8SL9cxv7LlHngKSgdDMLwRoj6NOV9HOzVMRhW3aiNuMoZLlLw4OcuFmaW2SN
sFOb6MubHvSg4J4wc6Hfakxecl3F0/XriugANVGqi52xzkGlC41iyqrVp7/TfJ5gco3+fWY+TCf6
bpqusHA5zS/LE338yqUNnnmOrSUXYmEJbHcBtK4efEA2X28x+FgGsJZAbCaamvINLMdq9SDTmo/Y
tAJJBKPaypqT2UsA9Mb7Ayegcp0SZOt2WV2mvvPTXG0s/h9HHq5P6MZ/ulqUbkQ3DCjjwUK6erlf
CK0IVpkSA3lBevKAS/x5u+P4h3lcMGYfgBvZTWXozW1lsN4fxpXoco3EqvUoeTUeO1kI0G3QpfZ0
5mTF7zK5L7DUy5HPasOmCcJAie/lmM2ozhBzxsuGfsYAMGNmfXjYfW3oqjr/8FlBGimTSmxdaCwN
0hSVpTLlNsv4s1w7zGW4sq6k9lNRVhqgvldifcmKpMuHxKs+BwREZ9ufKbYSkLuGNYMMp5OC33TO
tcVHPQZot0QSq/XjgJEGr4rL/iDn9yUis3MXTZMrz99jcUtKx7LMGmUA+BdvsxnbGUi1gowvgXz8
8PYXfpMBEa+zoG0bmHW5kWsG7B4rgq8lMREb35Bc0qT9dTgEObcbCDolZbSz6T420u8EzLTAYZn3
v+k9d0PjA52Ncjhw7GGfLTeC13YIsRUw4f7tXKJK95YMhQsvTDTovoEmTK5mKzPoCkfQgq7oXFn0
Qgn/gNFwy8etstz070y7L6l1t6Y2+jK60sXORfr7gnxKivtvMbrX3wE5KaXuEI+46Hi3LQstyBu4
hAnORyfZv1vGb43xcRBKOW13Tc2N/YwX1ywrVOcLAmqgErUx4Pg122ziWHB7IUjcOffiSVMm9S36
p8w8TnjOfYOp0vOw9tnFbXrQj4Dl6fJgnjuJuyE1XcR9XWp7+DtaP0JnxfCEmRhHZ1lE3NBjJbc7
ouD5ZsoGFvaLdzXnlQmer2yDQxpEQMp7DRFnUP1cQmVKrRJX4RlKevCfxkk9BCoAW1hsNLbgfUS9
ZoQBScyif/5KRQk1qxuB5QCNZbIVM4tZ7jTMnJOziCKmyH7E+We3KlUC8FXqSFrOa02PlaQOhsX+
jZm1i2Dm8kK8jBAgFDB6PityAjsWqpLvMNKn6Hi5Yo+OHy3K9BSL5ItLvV62ZMwxTCKjjt3iLsi8
ZvIr0gG7jJCu+IxAXIbnz+m1ZHrmusEEOHt01wO/5sEoogiSDwRkrbhUSI0PCGwIp1648Unv4Fpo
eamBE0nDhF+QTFROsOFhTUPCs09yUmXHPkyQkHqLGWuNkTtArfLjlXIHtH0g9DcDkgvOwJC5EVDi
th20uFSaDVeluTKmVuBQh1sn1w5TCGslMSJM04hmTnTJYUQoGqWTgGrtVb2xO8RK4Gz2lZdL3Dhs
lzE22dgcHrQ0W+/kMsO1k0MNuKFDh/bxUu0lWAS1Jfyl0sB+uv/FQmX7bSdQ3cHUsXC9/e64U3g6
xt2YymcW8daZcdWvT6+LQUE3NhXKxXYtL8FWQjXBUc9quj9vRg7ksCBceQR8GTAjqZnYxaSUc9qb
3MNkMg6QHeqEfGXIl3njMReI41CT+xKKc651MOmHxqDbn8TBrineGswYTJbgOMjAsiTXlSRQ+O8i
hnkoQs+JEEg9mUkDxPvRPgEPmQjAY6SQXPtXyMDn59DOMngss64mNKhCy+Ld+H5x/AO7NCUj5eY5
ZMY9uYd5w7RUppZYJaMR7+U7BiwIw97JFLwn4hc51KKXsBuFDoCJ52amMwfiHHml0J1ThDyxJuUR
bSg+5JIhNMFeT7y752zhvEIL7nByOkzm/8svwV5mSTA8AD+KOfx68972FFqgXvB+vfzr1tLCiE8v
sG3HZiOT2cP8qC1JSnQyaAXtA/Rq0z5JFVm6S3k3GKM93+t2B7hfuPJbm/sLRg47onHW25f/+z0M
dGmEwJOISNBRO3ylSdbGyin7RGdldvChbX16xrvQIybI0eDuty5MlTb/MZ7c9Yg0URTCKfdNEGRM
QYoaf0AVFGBjehXbIAoiPjjaUou9sAJI2X8hXZDZ/WiP+bNo4zFdgZINmiyxydTow1RliDJ6c/Mx
vvQ1Z+cMEr5zCVb/Vs0nOSRZyD3wqQ3kZpe3zovpJ5VIfP2rzGG63YId0VCTNwN2vSdOT5Ox5u6A
88FyQUVC3Bg6S3uBLvjs/VRjcf7/62li7rgkmOThYo7Ex2C9b/KOlsoj7+bKgub2/vEruXaiEorZ
tuh7RoMza3leySkXaQPeiAccsOdObS5UO6fUn4qeQafHf9S4eGv4z+Nt1jI3HMkhgPuUwlZHOCVl
RaxkvZ18rFdpBcgeHtBkngQxbXDj3Cc+8BJ+I5JbWWPjsMORyeHljA0c/5YPyXzluYIaw+XuqGR/
AmOSvXRtEr4/gsZwoh99FP0jm4sprtlpR68KfJFWLvSncI/OPb7ZK52YMXSudFVKr9q2T52ZeEgS
iDmpMFwAsgKcTEGaMidDyR0oude8gcF0mez5DVdWYiAS0DyRd7/LNAOyCzlswYaXtgzcNYPsDhPC
Oj3U5iBLWPgl0umwX0HImWsQH5CQZXHMupIJPW9oFVXbUIp1Ajwm020UnePHxrkIkDiOiZvHfmtj
PhOKsH1W6XhTm7oOz0CpRBSPZWZ0cIk3RvGcYUee5tIM1JGBckUpBNGzdfdwIS4GSgJDetJ0kGjs
lhJXg4sGZ7511zjrzpCJ0BL6SUPuN6E20ZO+sbe4JnqMBSKd9kyESuJ5R5eGeJW/rjEFL4n4pIug
0aSSGpUvx39myT0YSIHLevON5/IEsesCC4OyvGIpCI0x4db6wXetNy6Ez6BIJ2ZbF2vgooYrflhq
VDxwvJRxjuEZZbe+DwSVx9/2URaNS1MJlLgDk1dHMnLpoio935JdvkCMo0bY6pjY7PcA/5t7ixQ2
tOYi2SWN+dCD9+Ah0yY3pP4ueY+ob+Hz9XwngyZYntz5zabvxnio2nbIZJvqMZyCKm5suK7MTImU
JXMCuKsyLfDy6c7KdzI1U3UveCWeM8yviJijB/Q4uueoFL16Yyh5VGnzN15N2/sLGe0Fxl1+4p3e
MWB45+R0dYnimuZ/H7Q/C5jaEZvg1a6a93aIhV0InYrArManHXySyUl6hFbaUKiSMLfBm8S1phYH
BkhcfujroMa3r28O1gfUCMGQ+7FAAuuf/ZuR4nFBBEGAqt7VkevqYOCKafB8IJHM3H0m3SM1Mz/H
uDC6r/g7w8oWWxjJV4AcYLu1gzbkYjz/8HoFOWSXDCFUjBHU/B7zIkGAO8aZCTHIUAgU9Yp9lr0n
aLbVeJ0oWIa1OUrosBsaWXxZ5caVIf/1zmNuApN2EdH9TQiVrELWCm79TmvqfMXOR6qgtoWA1CPc
moUKpVidaDpQuiqT+q+cF1jRAYxGTUGwZt76xMSiOfGh/IB6dkP7GqW49L8wbqJwE0/peGTmQ25b
oKtXPUtaory7hIPL4KFpNgX8LbuBBryTee3seSRkr/wS9D92+WNuh9pRde0KmCZZIQRqF3cnIq+9
X4dBk9djL17PSE6pKCMlxarrt4JxFEwzJ04M5IkxgV+O3b3NoS3bgkgtzUL4P+lWRdinQDBczyfU
TMOeMU6H2nWulcXijd9you5hGK4OQK/iVtSFJkqN45b8kOrttFRPQYjK/h0W15GmwbRJxdmk9M2k
pf1/8vfhqglMycxtKs1ZDfAJkesoyGvaszakDmookCYpHmATEsL3aw2r3VBQMJX8xOT57UUUWhPB
oXu4Uv1TACxBMruj39pSSYPH18ltUaD0BcrAN9FtHxBQuYn7Uazit8xpsYbxse35ZrjEcAAkpnzM
jCnr+Dnrjm4ootRDnr3/gO0hX/kwymeS7GXHDGeLTIf40/8qkuKxe9SLmQrxlGBRyeejrDU70Quh
oT/rOmQ8ZrH6CY1hVTxgZP1x4lp82qgpISk8Mi9anhwCs4oqP46TfYlz3LmH04N+JksXMHtKLbt8
cVHiCkvSFDyiz0HFp/3JiN65yu2BZrr4myecxdGy3oKVLVCYR7QE+g543aVZXneY84P00R9rbvip
0UV/4OP3qocoG9/MYtIkvkhKSJcNL910FixUPMz0M5dF+ZOr/DLncyXgjXKsVRATt/mW3G3xPNRN
07GOLHNrekBV6/d7lR48PMWutqt5dxf3YsZabMV2iHNnK15oZFDZ6cnlMpdBtsaYw/9zBYtahhLE
cdREkeqDacnuLl2uQ7tVs5pRpg3cjnSHlXM4SXiFispoklYpWGW7JBXxFpVnNU9OFVkSGiaw/sva
frsSE+Xt7oyvIGycF1inLJdI9s3x2dJPITn8yreemcKxXyD77gjQDKLFsd3GbPNlTwh/8nnkH1F0
hp/vWQpSJEbe/dP/0e4LV4BfqJRLN82f6tql/ZvxNy/ViaYE7GPPA0V+H7Yu4BMtpARgWSxCreh0
l4tPJPtRZDz3nHQ5kwm8XayXcAR8x5cB8bP6u9iIwnBO15kdIddTf1Fd502jJrKxj3gvUfJcCb4l
7prhuzu7UE6pTWeVYbtHM/0XWNuCcDCQIsxwupvpRmJ5mW8y6mNJIWQ2LrNCxlR1skfPe+5Qb1Ul
hdqTZFfMjZ9Rpm7i3maROL0eIardQ/y/HMK4XmBKFpQc4iXaWeTOw3pZKGWUWmBoyF/y6AvF6DnU
+dsR/1Gh1BwFQKuUkCy6a8QWG/s9sJR3pFiVosbte4cgQzJFqq6ipzPdelPz9B2d+ZakQwRbBp7u
Fvt6xiSX5wKyHCELWMtOmOPEiU8E9740aP8AQ50GV18sq40Z/nBp6SK5qmDD59WV88Ol9ZsB8ijC
HfGVVfdsNaAKDTHSp0vvV0ATU+SaZ/Uh/IWJKFEAa1dc/yeEuYBlqJp/sxKPSetdt5+e+1ouVdti
lRmb3FTDWEzJV44Qs3da27gZqCcD8H5t2Iwgg0eMTH9zhdrg5dg5BJtRktU6Y+/lmEatBnpk5Ro8
njScGrZN3+ZLmTZ5vJgDtEVOz5VKbIRFxswVdkzqWPcgViUOG7o1yDP3Yt5dVXTXRweqwfeeTCBL
uXituL9cfJL6KmvfYNKvjymSPTf78+R85xOjT2xMzs1GJgrf9Uf33xCXL/9uwub+zSFV7GgShaiV
yLt95fJ50nfZFeRCeFw7u8nmQ7JUdCGGyt+D/bBWXscKIBLC1v3I5C5mqsDh3VvuK4gsbhQSeQWr
121yV5+O03sid052AS9Oe76Yplovnfqy2/cY94zpR5Q7eCnbfX+ITHeVXu8y1Vw9gPXBZL6OWkCm
yDnWUhTQ/DrGmEt241N55fKnYYPus/TAGGgQZzs2l/ZCuaNXh/VAoA/6im49Ny8DavLVKPZuQzto
1M7w3b15uvfkZfrKk7wGzlEMJ1AykQXvfiOgS7Q9CpiKqlzdb5Ltnt9S3y5Oe8fNFmSzjTpKOqFC
xtmaP4cEcbsco18QymrtBNgyNACqWqkH1y4RjMPlWlBMHFOTwpUp0KleDPSoIihifCSOZf7Rac70
f+9RM/NRAuPfA5MZCdT5A6KPWoU95SbhxjoIAUWAgQZaeXWGJHNY71X0Lo+FrC7j6sp/TZJ1CCRr
tP97AtyikXiv9jKl3Uwo5pComvTcr82dGp5eO7sXCCTRr4Gi8Vu2HslD2ANj1Mfp8pb6uaXqvJRf
ag3DOR+GR+PHn5/UdYM2DzeUy+Ttg8qcy4FOGoK9BZBh7iCeqbC/EQg7MqQla182gi1A/2VM6+7K
/t4oQnFV8pycOZlHuY3vatDzoHE2UigynRYcw5m1vo7a3hHEvv1lJKuZ/+t5wZgu9Bip3IRhL01u
jHsGdNbGrgSG7eRB+E5lLga3dL8t08J9JVaiplKS+4PLSWC0eOYCS0ahzlQRy+5rKyMrjLNUJUtr
zp8vEDNUtDXKfIISUg5+6Tod6tm78nJLjBDOUO/h6A0YrwbR2BX5lV8XhZVzDukN+uBK6k1ORSrv
yvjS4irnmic3WmU7iK7rszFmvhHU5pW3LzV9Rs+aurWiX4mNjqGy2RJH8LC+cWqZw/Xd0IMI7wTX
Ew49YWlgXo+HSj1kDmcjiLxxhehwHwzRYdCRJETAZHN7wEhqOZeO9dRY8+I+3xHou/v3EfXAorT/
tQMBMjJFA4sWgvYN1NJIlIuYG9/+6+J2v6bnrQC1MXRXrYdAgIFuETCWaNQmsX4a0RUC7JefXzBW
jcBvWJafdIfFm/fSFM+aTUTXZVFV2iPSSlMx3yqDA8ok0V0R6Y2J83nq5axn1vPxtTEdYnComxOi
cgcCK1ANsOzqKCEYMxTOa+pgbqju8EFFJEL2Ya7c2pNO3DfczTKoMs2bLK611YwdvJImLNOxXChs
k3jPaxEX/krlLU6RqwdcI0W44NJxwsfMKtkcGGA1fmPbnLSKsXqPlc4IhMVBetssAoIv5bOvvJjY
FUkr6VTrdCoRzKoPTdOTa9bfKv91NUBFoWQSONcdWR+Eb1MYMJ+Zbogfw7UYNkJ1rcLVfRgfTkI8
aeeaqJswKA+i3RTQUmEgbAxhGj+AvzLZNL1YnrzADCZP/XElId1vaQvcZW+m0dvyc+Yb4styayHJ
R1Tkl6fcXfCYmmYkv3v16eFkKmid/DSnW4cUh9OfvCh7QmTJzE4aEXP+i3PqisFaW6JuYxF22q1d
KRGwum/GwMHXBP8+mFQDUmD3ll7kvH5aE7ShcVMkI7AdUeSUTecRQAahLmesMcvLm1RJRDQYR5n9
/hRv7mnxF1zYofqC5mw0jPC1VItPX1DvFFg23Kdk2zhf5wiSs/8UZzMmGO5i3o0XSLvPyz1bBuCD
Gbs4PtvAqjc1sarW6KIJkJfPdERTy+QZ9nNFXrFZGLqxrRMDhDKIhufBcPxLdnVd1M5iZh8ecBqq
v4iIc6G2v7VXWvyBlJhonqIBW2+rkvhww58IiUEqHErqSzFlJ5I6/km9VMQ1zasJ/VQ/hAcG9zCc
oyJaVrF8aSWjmU1RGp648L6Q/pLYnLJ3uHih5fP5ta8CBX8I41r5+ScgRU05GVoKEbDXw33rChI2
nWyWepjrHSxQGzAuAMydpheg4qMzme7GTI9fBUkYp2gWkn7sUgaXjZFY7qawcITO0uDrED4ptlGU
nCQFs9P+LiaHPP72lgdCHBMMAhIQZY27nE1GdngnfbqjgFrijU2DKgRK2zcg65prO4GxW1wXvstM
cPc2TgBY1Zgn5OgnGDSBsvFQ9zEM4njHZXD7R7buoHfRBvAqUZTlSM+mzi5mdrwZPrCqdPxKgfHc
sfGa2dqZnkoQ/8kBDmuAulvCVscBSfj8SA8ZSyaS0KtXiFApOoAObWBczZkc4Bn1cHrINBpVzyu1
2yPpGShd6kCjeFt2cAGQ3ldk9XlggMCA/pK3w396HJeDkmvO/wlCjh+X7A1khzKB7rGmtZAuGelR
9KOcSEGvckiHCBLkDV1cVwHWD5rPjAHrJ94be5lQ16t+7WUUh9VcTOL4m5S50WF/M1qyNBMuo6So
8IjIBzdzRfr1JDB5GDdVhfNpmFJsiCBY3m4HWbnhEJJ+EbKiDcKWyifDygqSMfXSo0ojnMc8qP7y
iDb8Nn3RiW3hETamjTu8et9EEzj309nViHmKSwVFjsLnfXybgz0nxx4b0sRyykqxxLRS5xcOl+em
JmW8BDQv75KQDp3M7Qy+XT5iRr4Pw5zzBzq/6X3Py5tCvXoBu1LCrOPlR4uBBB4fla4P22Dz4s/q
CkzdhSPaUj9w9sV9eRqQrMaCfoQmtpL9Kv5/vr6SsiJcNgk8713MJ3oFAJLfII3tS8xvziIneYiV
kBTjp2zaZ/PiChoiw0/m1cua1sP5Dsrk9cQteqXe0YAl6rqRVs32wnXPpCOqb2b4eo9+WmUZECSI
TM5IOVJi5Ub6GS3yGgw5k+kZJY6wWUz7LnIomIyveMS188dQdF4cNlTWcUHt8TVUN2I5wN6BjCGO
D4tjIDiByHpHglJEPn+X39v3vBEvcR/wHnOpERuBDkG5sQxdx18fOv3mbQXaMESEYW3KNa2vQiJH
SQ8eDtBqR0jggPdkOL42Se4w+rhMdCO+ctW0umIJIVMX/WHVuuD98N0CIHUNuCNVQ2Ba5RVv1wnZ
PysGOX1jd/80uLtPvvqzOXP8MsNGGFd01VTQQseEzgJ7N1ehvpdD8rLDSJG3YOIW8U6pJlcbTDo/
AXoaMZPv/50r7pSBZ9J8epq0H+m3RR+crkYhJwzoCz4UFnj9VGvYosRTj2lAkSL/L+6MIlQxAxSb
h3TOWQszWl9vjG87ksyIn2FJM8ATxC7qHQ2YJLp9XqA0oaT5OWzMK9KeQktiWP4+33HIZhTu8EB9
tfA2OBnTLMiqeP/975yq/JapjUb2yzCOr1VLz3KpcNrhjGbdyjSRguggmyDEhFUBN/Oo0z3mmEYA
v5/lNBVfqyFeA89RbXxNkX+p2nQosbNNxXfMU973JvDK3oykrE5pFFhsWDJMe07/8CanS2a5gjR6
Xdnq2Qs8v6Sw9ub52sIVo8TMEnjH2kVlMd2EypEmT0yuKbhqaA7tIPxSPMqGnTlco1KRuRMzJnkN
hHI7UyBTmVBw3W7itGsvOOa/7ARS6RFCPs3i/f/Heoa2KVijj9PAcb53+96TA1L14FXNdQSkqT6P
R727h/0IJVs9E3puSTV0gDwVqF+C0emMU87LgZphq7PPtfRDecu4wJwEE3nqVmzFvU04Ut5qos2l
7RrslkYH/vPKGP0aaPyHSZYB+SWr5b2NGl+fhxNq/0jMnngzjH1bAKED+3TPm9ZTeuaNNqkhZe/9
8MhnhKsUO4tEDgQUyVA9giw33pJNki+JS4AhQedsydZ9sH+29ERH3aPYf7e3wVJa0J8GLi+4J6bt
i7yLzf6lX2feHRu1dFr6yPwFbK1QBAjMVl1gpC/HMvNtoeB8/SuqVnu2jJbMLLCXM8Utv7/P+Dns
voxVAGljDkDDvD4dEKAMpYVDB7u2gesRIMXZnSadIToJG3XwrorCzDgVkCkKMVcN0eJb5iY8ucTM
Nj15fMc2JGR1znSdkwTbZCAA9OEvGZ+B0/8Gx01I4erkT10J4DZur25t0gTqrXVYnrEVjqDay2+U
oxey5SrIV63/f16esw7pcdtKwD+woYd/ZBmgoozQl8FtgmqenesN7S/e+ySk8tWfe6AOQwb5Uzg9
qzCK/xDUiToEe7dhSCRRgLPKup2QhQVMENvbQoCCk2y1Lp3uLJwnLZRndN+8Pw4ju1cazimStUYJ
uEn8+gNqVU6SZ8Ib0v+YEpm4c3JTF3pVdsmewz+VJnUa0t9iDFFpAcSkgkdkD6LZQnWxmrK3Wrzq
i4J6ZIEM0RS+wwAAUC/f0rTNggejkeHevcWCGL94z/5uY/Vj8NsMhqjmgzAftCQ9khMKFq1Mj+m8
WWhbpIX1Ds4rq9WrbdmeYhPrzbawltUAA7USMgZl4X1EyO1DXMeBHzY6ag5Z6b4xBC2HevpnXBSt
nVohaYnM5G51aWeNEmEL4BAEntvvGtmO5Y5otpwBDTNfY4lgoexEHiD8+yzTERv3Il8zzkTEucwt
rnWNKeT2WPJTutyNpmyGVKuCGdch7Re3OFavmpTgyxs+B7yUvwT3GJALJGG/yey8fYVdmznGbEjN
T9qS1qCaAMya3zW0PxszTbBZiZJF+zkuo2gHxfVUUb24bP0uwPPoVNvDJ7AII8VrZ9VaEgCdXC7Q
F4VC3AAXEtEL52g27Cu0Ss6sarBR12vLX4HXvg/eCOpdkl8QCE/ats+QPeo9uDo2l1SDlmfs/4o9
a0f27lcLT5iuy7piEp9FefQEaZBJOhCoWbPboI7xZeP59DMypL5cWptNXpdOLDp4E8Jxbc9NVQBw
pk06Q4mLY0SVgm5Du+oiVMfJHEr3CjD1P235k6PN28zATPGkm/iBMt4YD4+HisTVG+HcfdsJiDr/
RDr0+FhZl+kU0OlWwBELGwAP7HZK9o8KlZ9YKFEpBbCvk5aLOOeIoCRBu8QDu77e2HF87VnpEnGy
ZxBFvP+xzRIaUEIsYlg7Q2SqzKDCr8wGEIyCnevZK/X6gQkvgOpPvQdGONxAExzjG77LvYb6jqMH
kTLZb9Y6PyJtV/wiBDMqxYhvmor33uok6ZSGudAs4YWoW63siCMxwrwYj9cuzK54xt+kgh+itn95
Lrv6hVEVKvQ4ShUTrL/416IRbAtjLi/LFjvxnzIn5YQreCGn3IZOwW924H1wK9ik5khc0Ckuo0S3
ETLYtLu2QlM2P74H9QVtD6JKVpK6en8iLNk7HSYm5dK8xSgMg6NyCZ0Pru0DKTxHpEFsfKv+BIL7
fpErSnm1/6q8Iu/321Gdpr5t8MQVt0xnzApnsPA9VnaZBJmqRFo3hr6A/THEBsrZslxBHvRFDRIN
OVIo9DllPKugFwKjvTBS6sZhUeyTsR0ka80NzkcP8CAcgY7IrYVYjpXigIQcGopPV+kyR1YvgomQ
tJAEkO2GGHI6/EsiNt4+YXqaiAw1JaTLFlIVLqpQNFtwqgueHCmrxhHrv0JfIDL5mWCrbYei7Mu1
30ZaAsQ2kUPFzAJ1A80/nIhhjLn1s//Fv8p7nGhRsGHQmRnEfzs90xB0bAWKGByHQpTzm+gZU3Ix
vAMG3dlT9yIzn8SA7ahWtGPFVg0eQye6z3bLctIoAXZXDIrODWEqoDfNROzmfb/varjF80CIFfjr
1EATfiQg99rC7LdE/5qaWXB1if6sdWVnDSJwOTH8wl2PuIY1w8MVUJ+rkX8WJO+f6MIo/cL9Jo/V
nz3FjNZCjqXT+uTrk5XZeiNX2UVU/9fT3lu2tobgl5SJ02dYGHCAJjOhubWFZqSfGE9/hMytaA1G
8uTQ+2W9KpYb2NJpben6ZClPP1ff9QBzx+0moM9yupHDoF/uRbC+t8F13aa2SQh4w2AT61vxNo6i
NyoUawlvk14Q3ie1tZjHQu9pp9ePe0iVfSavT2Dq7qIjB8bJl8NZOFqQXeRwl+Q7kWe1j6ay7YWt
q/eHIfa/SrwtR99Nev87MAF758qFYNeoM8cC6+6YpHt7LoNHKY1GkT3PXUWF1g1MH3x8176iRtRw
7ypSvZiepY970pGfZsP48Wqmg1hDsPEbmXlWsl6lX+a4S1VoSVoEtRL159C5lZdM5Plf5uL49s8j
GqayUK5IjYyDOoiDk++cPJ+TpekMIkA+fvkVlygY8p89ze+Tv//M+e38scfAsegNKRuYrnlFrdz1
dnH2TJj6kDAQscT2NGOC0+P7YBQRNj2sBbLZ6mmsRpNtoN+65TF/uKAh2Ht+VvSVM3LEWzPpkCWw
E4nyYqQXaY+BNlxe32WFep6rXCYs0AmhVCGVphVX/v6tJwQtGqTf7p1vzJ0dBMW51vEa1lN36Sah
RzFFBeQa7CSieK4Skec9jJnlHlF2BdB54RKSXrz6hTd/s2SEF8ejNzZXS1iuZiWH2sUk8R64VwzH
xlq90NyuGGlMOc3rcP13YSglrd0MPN9H01r3fT018vXKxSXYX6yg0syOctP4aj1eUW/e6ri26CvV
Y/65mW5gqoM7M4KL9lrxKszuJdzmVO6liB5MSFLc9New9uhX7UNmbDI8s9AScK/C65mFAauYOfJE
7cT2ecjdXYQiuX/IyoG8vaB5MVj9Mrk5xi2VYo65j6UrwbF6bkgd4nShUlT3Lwdi+clua9Q7ROQ4
MwVcd8t75sLM+4TM2/KYRwpNZcW73REb8XDralqo1peFBU+jh/OPFJKCsLyuDNmAOSIEbFuQupz8
4uH0RfDz0mMRm1vKMtkHgd3g3vXwDJyXex44qpUEKMIGrvPk0VZ2jbTuT66o/5QzNQ3AvhyG9txR
z5hSQTMOfTqYqbYWxgaXuwzzchcORI4a4iUHNgpzxZBhIyH4UtQMcH6+9WvkE1HR9mxkSQZNtlHu
gSOBWErydYMllUuA1M6LGapVUeSrN1KsuLyP6/K5Ojx5O3XNH9hIdFTkEd8hzsGutMgvgssZ6dX5
B4s2B5w2BcRSlgfGQPHld0xt3Zf0bMPEcEcertMPPie2cAv7t6PQUxATiY32H13ZpxXQcwanOd4o
OZam9V957267vK5KzaFcFC6Edu0hgCEPpsfXucP6I+/HpnwkqQYosd2b/XILNQTT7Wiq+TSWZASg
0d/gicw+kgtbAhY41ogK8pSF5c4piBNFv5HrJ2s3+U/o5pLie3zT344xb3EoVBqNxaf07XDXPDvh
kGx55Ow9ANnHegqPnHjnXjEeTz0PS1O246D5Y7IPx0syE076QeASZYbUka3zMxcOvKWvLO98atzJ
8uFaVrXJP04BsYHDQQ7ZNwMJltBwVgs9r2lo7q583o35O3ahqR/7VAuYniMFrUa2zdTgA+rMA6Id
wvc5pZpMM9a8QIPcFzB5ilU4Vt4kiU6+RR/MfyBhDfaAyiEqCHEJJH6q+OIxhg3Lz6JrO7inRCCO
83vdDzzncU27KAqlgYVXzAYAQ/+40cFpUMf1HGnsHyIzve2yEnh6MG2gBBHWguIK+dLmOp73VpXs
0tVliX9buPkgNaoVwHos/fUXFRAiZv7SFykvtky4mK1vFA6Iqz6hkJhVZLiYX9aqkg2lmYVNgju3
mPkbF0/DGylHWEV60SweqZDFTk2w1ExLyY4oy8PgxTQcrxi1EeQJWUvY8+Eqjd8jTpMUnw7fiqjV
RWOeXSZmnsJtMKlsl4GWjYM5ZnsaUvi/O5GlIyADP8W0M+qghSL7eb6/Q9Oe+1/hmyFdSTNVCvbn
0jyVSrmLmCz+bn586sCfuzCjOxlM2xbuqFWIgsbbJ8SXOLWsGAyG55GpNwqJSx8F9LWnSjg86fGd
j06anDrtpv0TOrEvvXy9p5XD60nMIgUAXB/eLqgT3IRUR9icPaUQh28lP6xxu20HaBtUZubAryzz
4+kZbvCEie7F4fj3d09W1exfAvNNVNuv8HA/yF5Kc/awjRLxLtgiJjA281FLarY2ADyslIUVGO2t
H6gfE1/yR/jXc+kELDpmwoUKNGN78rIyeN6GmbIqoB9OtgbvMAhF4Be4IRQ8UHjOAYnXDVP3/QZm
IEIPZUtic/QHiIjCP8zwUxqEGP6Iipcrc85ybuiuv90VA3VZt03D3aOn1K0V++8Hl8uMxP4lvrSY
sSvMc0zju0vxcrvhOLgpkVUm2pX7iPCrs2SMCQm5zABp2s44mH3x3SP339+g6PXBfCV6I0X11ejz
zr5/jWkkDlFKR5YZr21yO/832LDwrz7QIJR55EsIeUBh0aOnip6N6++j9bAgFwrVwYfVgT3cWayA
K++abGHKTcDuL/XkmYmOoiK8kit3gs34jdlGiCdhVy75QanX+Dprb4HKv2W5z6EZlvCv1jUxU1pj
r1Zm80dLXOXcmYLq5kJiiDL2067og/BRtZa0HPLor7I/nTGi4vAW28XIjs/76xOKne3ZHvQPeCkQ
3dvFIcgoVjkK4mJcWcC/o3xk/9Z2x3//lxrThpq8kOZKgUkQsgo05B0bnDeMILqH67eA4fM+CgUt
1eM26LMRSXez+NtUESMsDvXmggccHoE+Wvkolw/5DaduHkUG1OnReWOoXO4Y8YbDvUmqhhVAS809
usHzz/PaKw/f/g0jPA0IcZ7zyKjq5d0VVLtLptBnVISeuoiUPqLfJofua9jNB5hvikL9ig8u1bTd
i00h2Nb7c7nLjlaUHdwWrsnImaIHsEQjdtzM4Jcdf2IxFBVOucFNgXPXp4ujdoszuFayW2VGHfNv
FAcVE28ulrWfbhuK2b1vs2qow5F9ruYwMawmlhsJA8713xz7mwiuwuAuWxUWIyH6umOxDVhUEwKp
sJUfR7nXCF4P5E0i17yao5QPiCOqeJN4bOjPvXpw2Ao7IlVfR40q/fPNmHd3Xn0CRN1dkZCQSUCl
kP717XCNpUHOYsJ2Kqd2wzsDVUHfWphkyFKMryzht2Kru3NvMoQfnwJJX8IZ/mU9I8yiZ5kRcbYE
7q54kjnNcsTFtnQ7IQgobNOvFpPljIvFBDu2eC4lCxQk0y7sund5pPkXBX8kXTxeq727aen3qsIt
oIaLSa/zqRXp7rWam6sosVWmE5VP02MAh99PPkRnvXI7peud+ncAWk3ZlrPyv3eNkh52tqxJe1Dc
Y/XusEyEmuqvDX4T0IkIVCMAp6MfSySlNuqE0vDx1sR+FKU06veCRw1745jzYc8D+9ragM51Aht4
4AfO87vFi+YLf7Y7A1LK/Axi/ImsHEO9CaNFcyKNjfQPiZ83Bkjhxfv8hV2a4lJJorlmYyaUib9l
RuMdLJQijPkHbFnQs3UsX3Qm1kBpry9GODFPg1s1ZfkdlzaySI2/dc9zljLQl/jBn4HqX9dKiZqh
w+farmGtPuAGA2mPjFL1hwq0PJYTrTU00V3LqHGwLM5clkAtemvEUR5XAl8JalY+oQv4ZBw+UQbT
QJZwK3aBUbGohecC+qp334sp1U+Ua6eFsKLcZt5cGshlUMGJSK0t+CWeio5NF/oq+0iXd9+1E0Ap
xwNfzpjWXMR7byzcRP67/f5s/KD9QKL02LJzVQVKniG1JhkFzSxcBhYcrY99rbybxS6u6I4FhGip
7vBo1lNCtrc+NIgJPtU54NihfhwLvW9SXg+7h8XK/P9S/EoKPIuv3Bek1GucF2M758wg8J+EsonU
vRIoyHXPL/tbWB6KZzjMFAqoGk52wBfZSI5t2BBBuaV7C1W4jaoTxlSkiVzfuU8bxaAtDeeZvmHT
9QsPX0vVkMYAG4RWggc5LbO53TPKsf6CrDiOQ7tgIQ3DOkMltLZlA6fkLMYZn3ohXWBF5oKuWZK6
4QNzWHIlwQ06VnsipPsOWCy/VYVicnvvbD1ZGnGvatqSNygwV+cT6RYY3WQJyU4tZnaKWR7eNAds
vtbdi/BjXQG0bfNqqy+UfkoMsBomYRVzy4TeRdys5P8Z56K7D/GXSqfDrOYDhmmFx+IqoTnSNRm+
YVmDShZq5IQcD1e3IHYJw3eKlmUg6W/smPRqJyMMd0TnlC9BxVT/i+h56pxbOvWWm58j1P0zSbsA
Znlk17k/SAcUKAb/w5NHwp7jDFFemucFTMeuNXDCIGPoa8TGmU9soXRl38J0eUUF1W9OM5evP1dF
2yMeP9D0eOhsh3Q8Uz8CxZdOg7Hfw970+8TV6p3Q5aYO8EEW6QWmNYdQCwtltSWPym4KE3UPoQtw
1N2cmEnBnihtbPc5V/kKtD1W9kWbLtkitUnqFUlaJO948Cg9TTk/Tvqdj3RFzZ2L5W5TdEws6C5r
vJS6Su2jFN59pG/C4uXTs2MXvF/43kRQeLKuKh2zi68YrA50vV1VIE4sQJPpe1bcH0I09/fk+lsY
IFExGL6YLzrJYKznHfXqkdhRuu/xhON4tue/rI3bMWOWpFRySmuVTPYhVef3hkD+ECWF2Bk7KDRx
ilChkDq796nVuZEcr9keKcAdFUT++QXlxwx2rik2Dc3eB38WnZs/d02M97KNDm1/fwLlLY+hu+S5
0WqOTpW++loLypWI7+4c6Vzg8yKFm6viLK97b777900iHKTG/ONgsica9hfFVXg0mIhQqioi2nYy
b60OLzLZWd7323flovAglxNR4n7UN+hy7gjNHHwHJZi03IkNYdg5T4y60IIRdNyAGpwbQDPjhmdV
tkRpqABOuyoapvhiXL6X1V+9bBMpDJDNJtW+/WQcrhq+enlM/AvBMSdVXgps2blBTe3//18Suxyx
H74Vmo1JcNeP+LAIEZ3UlBT55ieQPMswChP996+6p/5XPLM1anSMKMgbUe2SHFZvIyGID+8N9AW4
Vh/Qn2Xt+Rptrr0Et3uIJEPkmuXqfXh25A+rCBFPWSSlpChXAPK3aHg423puaLQbkMJ6W3GQ5YQ2
s0OPz5F5L564PGD9l9d1hs+LDW3h7B3ziZT4W3yRlBG49wFHIGCy8kOGE7VPeVMtsfeQMJQWso8a
37kPotHFW2BZZcfDUo0mIR2yGaF/Dmxdyj3HkdUY+y06dy7l0+mEKdek4Oyp8EuIQHWKQHkHLiJg
jEgczVRZCOt34AbqrGed2hbCGCVn3tJC7lLzTr9+8GWTwbxhlEMZV3hPLiiQt7FxEzvjUNgsCMo4
x3rzy8ZBb9U3rF7cF7ZSYeqQPNbXr/bNnxuvJabTHkcO43Wh9pfAv5LbWnWgJg26m8BZaz6il2PN
/yVyb4FddOuoP4a6Icn5k+yr2cUAY5TrgdPCNACKT+fVgBws7L9oZNCNv6QjqlEUmP7ztph89bO+
rWXain9C5sxakjl+FVDkNLDP09XmI0AttLzCUiW7ICyzy3aFwIAPXlfV9ZoYB5TQsmpklYMSHo/R
7mpm6NK54/yNIsxNOR6n6OLU0+c/l60VrzQLloKXR2NohwIXtGmkc1wFgh0TG/RnCq6j2ShJt4+A
tkDXDfnjVy+TrMVeyAk5O1Y9ju3fMgZ0c+vA3v7uHTsr3r0HhhgzkF/orS0QlxFt4aJToOR5DpOG
u/z9ht457YapDr+RHTCQIYgD2l9WAxAdPfcqLPwXHOUTCHlis7m4/QB6rEEX70HCHFFyHaVY9OmU
DKknyso89xjXxJrNr6Q72s6GNhglzHI7ROjL6LECa9toT89RanKwzQxNETO3uJdALTJWeSKVDKvl
vTywB3iM4eKPTfbHTRJTztclcRDsw5tCX8D8BlSoxAPw+2xWX5m+s72vwJGAMQ6qAjE4F69t+rnm
1XRTvCRl0IiVXOiRfLpb3eF03/Dfqk7n3JK32IzduRFbGH4SJypK+daUajSpkolrS0Tj6YUfJY6o
29qoP6o1XAh3hQIUNm5XIF+688mrs0jcDOeZ15MEbcPkYjXX0ERKdkjp5gQJQIcYwKt9HqSneobm
+ChPGY+qruT6yVG07+26XkkDjq3XmdnWoExUirBEGrqahVyjFqFxY0G5dXlAK6f9rHus92wSlNLo
UgDx+peGM6pElBnsiTMmj3uTPUpaUVJZsT1xfIe8dFtNXwZPfjt9P3vcn0O8OrYDuw4TlYqVhvA1
j5iwcaM/AfVGcs2Yqvtk7C8HnY5xYtYp39DHzUURe3VyZa7t2IKZbEp37zSDy8FbKlYgEvKD8z/0
94V7qRlt+RkAQH3zIBgyQn0lZ6ckVQeqlEM16xmhn83zq6lY2LewE6aWrS3Y/XCqW1fFOP+uqact
hVZee3ly8XpriW93uA5M3gEJTQHGhpF5UJkBISfAs5dMv1ZiVHf/QbjOuLjvvAsJ7LHg8hR3SW8B
KLKoKeq5CcF4W2boMtNsq/fO9MbTckfzUiAv+9/BVTJKd/J+5ZHxt5R49wD4F+EXm/GqZ1r8lID8
mEiHDsRck8GeE934Q3PAbjdibsE1KeDRIl6SYAzFw0LOhETDO2oFOYD8i08dC9IbBPzaNOClWXFD
qRiuglIj0RqBdgFpWsuJS5HzjkPWaOB+uaVfkSaQKekb5r+SzWq0fTdHkNhXEx9SGTRAnhqc0+++
MBBR08tSpDFwRS8IA1QtjCsZhSEyiC1eNRH9t73ODdvBExU1skScKGG0/EG8+MwUiyEgRIAF1DOZ
R4j3gAbGYFwZZXfjaowaCBB4kv/TAPkFafGnLoVo019cRfp1es9rBGcaKOWBQVfAO8In8MYTwUGI
3ybZrlPtWqzg2+BzdawLnfAsY72IqpH5OU6kWyPjalOl6OwXzZYnKckdcUrN5xqzdHndzhLIN7cY
BFfd5thu5boaJhMQQOHeTLdMQDR4ZbhBYjyEJkU7d8lFUoVyYW6xudBrh5Gf46PJQDz71zsOHk/Z
tptBodmTdA1bFAOrIDzVFcdnMzxg0Q7oG07EtfGVWKpwWD24yvalRq3iPhEYLwIp6hX8qQlrLdCv
/g4I3bHU52MnlANNFDcyzMyMuTyVThaoJ7RNcHi3SmNJ6C5cLJsPmmTReSOO5wxVZw98Gf0DTjdB
7/2c8zF+WZgrRnDUTRmyT1Hgyyl7EU6GEuWV3kkr8qO3OOx99jLCosBm9Gn+wVD5Z8UjoqRUMquH
SGzJatOP/pDL4eXcishzZfwudfC5UO4jTSIhTtqC6tHs3a8/XTPt1UCu3XAStKGk3pNcrByDAAxE
PWIdbUT/ASoK2Uk6mGst04wE09HgQgecWD4s1cPON926lkrannxspKs8dT0jSiul9kn+Hg2faBVn
iaG/VxqA/xtpxDbyx1WjfBmSf3vXp5bIxpd0v73MYdJBQ2uhHQ3ZdJmRzUQqlUa2QAGiyFHKIrzm
4/6mdJie2OJmmBeZJi4LRykAuQVw1F32UT23ItSW77cdHpqwP5b4EKFQ+QzAR9imntna+ImT/h6e
k78Oeq3mav+EevEZ9t3Vdgt4KP7sX8lgf3rzzBVsiqKYgCvf6zZ/zELN+RZDL/dQOBMBBcvihHqM
V2j/ySS9sCYdZdwFJIKKvcF8riSrM3lZvXziJPFRQZx5jNvdeRnGPyvXJI3Y1RlcVl1tijNqlSq+
XOB/T44Lsk9/IKDOSj6e9n+HyYGPisVjgmqUlnYSRPOy1hiygjN7nrdCfxSR+1Gew9MJQ03RBKeT
e8zcwhuN7z+/KaEOY2Qac0YIYnYTJ1dCeAx1Jn/iaaz5YdFQJboy5fUoE+N9R8lqiv3jG6euJ7Z8
+wg3ySXBD5ahhLIDxz+OJzCNTHKsehfeEo6cidJ2bIsVQBXJ2K2emzTCDpCie5BfqRTLC6hnO4NE
ScM9gswHOn0NR9xgcb0F/OhNddoOuRZaRn+PTwLE8NMmbhUcgOxK1W6m3EpojJIKG2EAlCVkMbaD
4oVdXbdexeHIF8T1FzYn4KVphjEWqXdC+M/9m+GxjSw4OzST6e5MmdiPayEoS7Urhje1hMyGVG3z
rU3cdIevmpAnAtSpKsgPosYWvitVXTS/hJA1xYlcjRKzeq2Rls85g4E9EAdjVdiFDBLov1WrOx0W
SuTIIEbHmnsXJB7nagP2/Purq6r5NWQRgGcwAbM1JeBT8kVvlRYQ+BrZc1vJ2BYlRy7+p/7fDB3/
VI/Q4t7J526fd41QTRNhqsWpqRfXqjfz5dsrsfQ4tjvgsr6iRhb6Nq21Dhd5ZpTOXAeaaYayEMBG
VR1mdF6jWxkV9vhPbQljsH2DerjfHR68qhgaJUqKBYQW4L+neSUoAFSpga1f2TIcebc3uzSp3i/d
DC0E7LgwFKOQGxXB5MUo/C2tVxm3Ah0mftbjMfZ49/GJZ6JlYjWhjOLOIz/NWrDOovY5CEfp/ux2
SsA9cB6GLgmG1DIbnZ4tZl/eGckOadbizgNXLvofIcN+6wnitlX33qIRFgxN3qYkr2JimHeubAUN
p+TJfMl2c37rS1oGEpMXpYlPVKWwKIDZEPNrj0k5oWrYwJiDLesYxvyVdi3VRapr//wF3Qc6yYKN
5Jhj3BPqXymuUM991aCs7kfuRTCxyjHxTwVMcjdVkXLk/hHqj1PqwwdAbm9u3CcBtsxMcJfs90M7
SqyeNt1uPRMMqTnPdLfYnWOHatmu9BezLx8le6AH66BoYTX3ekblof+TVCF0YMHuw9L8lnB7EEdO
YwAU+namaTEAx/IqgS1tE401feCAdocJMB0621COd+eDudI4hkAG8QNeoAmJHxjeLRcaJeR0gahn
sY2P73BP1g+seoiZlACmZXQiOt9SrjSGvvXLdp9kNdYwQ0wC6g/bQGbG1Oao0jvWGN80MCIIlref
3d2TmhDF6RzFkzmYH9ET6pnzAxIMdGyuOtDOe27e4DJwtCX7+5LYiGfkl3oI/51JtOV/nuSqai9Y
S4DvOWJbuhSDlwCs+JuvnyKgHxhzSXrnT34eGN9cBDUkTclppe7olJ5DekfL3//2ctY95fL0DHwz
7zH0BBNfv67IXfpWP1ETkriwW/ERf9jojv+2Qo+Wf25ICBrLY/wXavsZordMCZ+HrQJEhYPcMHHm
sH38kP1HObsXUFJZY62lTMKT6ZAglFEXqqiducotUPvykrcp5B4cz7Bw4PyQrhOkwMJ+Avk9CJ8a
Ncz5J9QU4zrpgXcwUfGa6GCEjFn6O5pB8l/qssIDYXpIieH7P8+hXmUKwWQpNaLj0CTwN8nA9efB
leMng3KWimeHN5BNZB4IQZpS5IfJ8QZ7NXeRxJqIrg2tVJ7ze54HH8Kj1qekxES3NpVFfjhboNN+
MxSmsiUbMPo5vAE6cd4yRdYtZ++hfJVZP/G/0OZVo2ehdv4CwZMxMb4aw7hbHr1+jPk2Kjw4b3nE
OyswaqxzR2aFBi5d0B8srBlXNziqmnXYWS0dDb2z/mmTYbHKzTaVo9oo9GX0Zz0m+7PPmBxzWBbN
bgPajwQD/FsQf+VkTifU38RJZCE/gPZ77/tDLhMOXXiEMiSwXo+6TN2+cO6YFaF4zBjR7DkN7Coh
YyD7lSyxA+Q8zcavfPlikqexcr0LNMMM6rEzqR64bw03QqkBf0YOrHIjEODxMDmLKstJ7NnLdnIH
ErE6AXuyLfmTi5CCSVHlt7kWheveGphdYWreI0PwtLSYycJuFb2Xwqhgi+td8Fiazus2oxb/2IsN
b1rdvB7cO0/eBmFBpO/ICGcPz3XKPphgvrBXuQeACJDMhoul8mTSnxWD4vuAoLzRQRhiL1TKl2N1
p7sHzNwrrY0clKESfLTxLa/wR6nu9DWg/Y9eW5uR/6cSFTLqOIMXbzZpVd1IFH8+KngWgN91B8D/
FoOlzQIOm3e6ayppRh6o8UX+COiooHQht9Kw5/L5n3IE30KDhobjwruMHmi1jNF+J2iqQ+X2pVHh
tML6d/5oEFesNX3xLNnB9EsyFyJeqzMagim8rc9reQKuAiy1f3gI5r7AmhY0dnTp9LKRZXKTP2Gg
OsdyLRt1suCTJr/Bxg0fXQYdg0JIMBzaicDwTs5PdZrrxYXS3VFsDw03BgfxGB7M944V7/TujcGS
DPE9m5Lr590FAVE3zil52paQdvg9wqcTpXpbE7oyOz2b5vm+46ddV+g61V06D47JzPQ+BdxzYO+6
Q7ZA45n7iiWEUxkwEjY+hRHFuECtfFbjVsxF1ELRLw0SIq1t71aUYbvH/fFs/uNw1Smxr234eI4c
pzpX+XlET8upTYPUTq6AE2dAuq6rY7jd+vxQN1xjs3xEP5c2kjKvpAZTw6byiGAs9povPlt6kaEK
mzSPBLmYVMum2PGOPWir3GLUYkfh17MtfvQ7dIPOe0zFIbMD59PFvOANa7PWSbOc5WEjh3/v5Ybz
awpnYPD1kjM92zl1jag2nzh9J5CjnWOy9qLI2N1/WzekHfNTayh9WSlusMxXClUlwvRu5eDXxn21
IB3kvl2ZdYAVuVGj9bzxXLx9O3ppFrVGZbFd7MIqMiLzP4hY5OKWfiz7L85L4SIHEWfYCbhiXX1U
czsxkohWjHTO3gaNc1tfJocnJNFyCc/mxbSuEPLVOEAR9q5k2K9o+x7zADgPLnMq7i6zRlUUiM72
0e9EAc8pGu9WWsU/ybnSSpd6TFBu83kbUGa3dREiCy7xC/Q0PgkfEPjdKucHxYuxKWbV+vcWnfTx
ev2DZWeEKmD8bgWdUXht/1i/uACkwmYkCr8M93XSR3C6CaOcwcAkd+3vnmPPNlz4u3x9oIKwI7bP
dxQDJ8qB7LgUDsrHR6PwHeObejIgfPE8yFaxr3PPiANjtFTZ0a/BaO5qRG/wWRl+loasxsrXp/lT
psnso/iIV2Zp51OXgMhOR5fCGb58vEUpibdsm0Ek2GbSt+0qxO6dxrmhyQv/L4I7zuNfQveNuRRl
3601kkSUFGvkCEBI3IojGB9A8Jnmmw4lItt+kd1ST/tzdewqVyQIT/xPHwxrnuMTP+mDPCMwtzLY
8ExD/tLMXAAin3atiG4hn+dOVbyT+cZ8pOuYMlIGiw6J+JpBJ70aexEG6S5VzM2JSBUqU29twP9H
BkGTPFxKHfSRYFLujBLxSPuqRFOO71ULcbIrhsJi8LdMIUEbeJmW17wFi3qsPuc/04cFhUcGy+wE
+d/LmkJ3UN8GF2gayKIgI1XD2uVVgOgly0WoXe/DT8Snwcmj5FcM3FHY48CEt8h76I/kt0M3KQHu
opA83yccRUc1GH2IhY90c8vQPZkTiFwE1ZrCUz/58P8jkyDG/tiSZE6A/0/gtct80p24yDfC0TLV
cL7VRuNsno4+nAY+ZwTg0Xs2OOiPbnMFEk/Z8576YJ4zs9ytD/9u2jkBlGhfY/tp3H2oNOSNFKLY
hLPV0XQwchK4rw+iou/ckv7HEySvLCxp1Ok9LAuN3hN3hE+248DrixdZstj35odxwMLzWmfMGa7J
CEnqAreEDOhku9RYOJD4JmYW4JPIo0eL/BuGhq2EdyTmVuFE7MwNZ+k2qcIP0RGMEF1bTL5/RIJL
JWXZofRIhxZMyNT+nzueReUtrhkgvd5OsHPp6xnqTqQETaKwXhto7l7K8a+OSDMQ+7IyDlSXbYvL
peRthse+REK89Q9QDudNAPvSR93LMjVnjX/z55QyCJT2CfS+owLcaVED5krvVx/X02ZS1SqgxtDb
3KuSqII/kqXx0cIH+CIG5kjst6OmHeeeWFKejpVdWntQ/0uKZxuSiUcUAC3IchiNkPTjzq4N4+YT
cGjCCwAF9g25KDyO47pPilwC4mIBC+JoxfnUYKYcuget3aVo8NC/6PvGVXP/RyP5KNvOWwf1zj2y
mYGPbXjhSp8k1IrUPkODjUNKwvicj4iz0EbTQO/dH+Xe7Nss4SdByiXfBEDyhRCyKuhjLAwnBF1w
VziE8oqJFx/3FMGDCe/nuW4p0GuagWkjGJnP4GY5b5lyXZaEbltFQjfAUFZiYGaz2QHc/kwlDB22
UYNP8J5LsFcVdXMEL5vGyJinyYSRB5veZdwT53Uel3ijCOclA4eYB7Y8vablCNABOZafwvJAU5hW
y9n3O2CvihsRw7hohVWG/+pbICczRAreT68NG+WFVZf4mbRlZMjAcXtabQZA5IxTTRdxkXDIedvc
Os4dIEO5u9kvN8gHX/4WAt4x0eZRxHabu6IgpUV7l/+FkCLCfRRsB2xskHLyPixPhxMB3Ff5/b4p
j+3OEjlzzyRM36YcYPi6EFHg8ePhnZBBAdmAxTMZNmCPWoOEX4+vy34cq0kh6snJRmH9qak5T3jU
ssy+OGzTPjnOg7rTVt6o3mhnotdo7mCgYRmVgmQ0uCt2tvPmhvWM0FfQTPN4Jgi34afZLzEoZ0ce
AkskTOH56sLkQpHT1eJROh86JbtIap181KZA7NgsrrzRupbONuqnSQtgV9wW7B9gtDDeBm0Lcq/C
n7cH3Trz84QzbEI5ZcahDHRag/HmiJPJKprtTZ51htEGmoCCeAS8PBYj7jyUPza782H+XmAyyrma
QPPyBhmNZgQaaFUGoC+g6uW5BHI4247MOq5V/O/epZe0FGwMOt9JonZUBp8M/k0IofzUDUwHWowY
Oi4VUj4BWzOYo+od4yU7we8meI27rEkF2aTgdfV5AVFuoZL/6pwBPNKU5NiD/rps6xt8//NUKUub
TlR5T7uSJ9Mjj+EbbovxpxGyWIjR6JpCv2WTRt73pe2i6KfY0hRi93MSPKnlzxIzeqObTBFBZaov
84G55SvskemHOA4KlnY7z6yA26pl6Md15BYYYT+9j5+laZ5L5AvYamrLex8mY2rT39Fk8J8N+nG/
5dQNYgpvaphYTh1Y52yLJEmE3JUAyGH/ft3BLGYRYSkv2+3zSulqnasHLUZ3gJIpneBGmAVDRkX0
K7+8BnrAeox5pMWljBrFmVamppn03bcgBZTF9nMFyCknHlE6Qk92eeS0m2/T+/KJE6BoFvAtfKGS
heVrpCLOD48XnMmDnz4ilm6TZOmrR6X5ig2PH5PhVKUploo/bQ5nNcLAYLbuQLH4BiRoBG/J+nX8
eJdRKP3pgq97kgBPe+CKk4m9auoDAcBL3T/c+dC4CNIFjBDEMiwJ75NbmUd0lZ05g6qHN4swgVno
MCLcUlFdqbmm+n3HJ50jVjRToLYdIqaI3ugyAjtwmUCDd+WGc+0ZaMb/wKMAVXuaiUiboQom7rC1
b+ZTGHWMY4LSeFfHbrNcpgM1IQF5TTdR05S0iObbGV1am01LiYQLgXjf5HePfIoufgVuM8LxTPmJ
gnS2E+lFik24NDMSi2AFBujs9yFcrb1J1CaJ1jF0Ojcfi4yw9jthqOAFGdDSfZAbGST2Edl0IPYQ
8+BTTm8iUiKlTgqFgXPr4PVDqPW/hK5iK8bCrrRIRyWa4diXRKVs7gepWg4/S65Guo1hvbLhUiR/
iX8SvSujxUXdFGwGpMmpGlkkgb3KF8f39hWQvdWFZQI1EPbu4wy93Yu71bDbI2HyRT0CJGSSwMIO
K7JuWZqyAOW+E7bFLIhVLzGIFWRUR3/EtmexdSYe3uJ6adZ1mLthydb6NWF5iMsp9Ufvh9YbV6eX
Ay1qxNGjVf/eg35KZ46WsnZogOXz+KBG/uRtP0favtKf7//2u79WebEUim8So55itk0okhvHi0F3
JzNcJgqUyNqPcHSdJeyk8SfzturdnmaAmf+RRXPmu5YhSedG8GqYaE7AfCBMPR1oyEVx13v4xA+V
4KxvY54oXVnjTMbUCUPmuJqzg8xHqfYBHNBx/AvQdV+hK+V1rU42c7mGY8upo3PMQLZcWXLQAcaR
08cYwGceytpMLwazMzIZ/7KJeEB0Z8iDwFewKVkDhghMA94ulH8vIefu4o6YG021cz8jVNKwW5aB
Eyfj1P9TddOrPKdbD6vyTx8NCdDQUrQAeo18J9ijSSWZQ5Er0rz/2Tc5EWmknVglfoNf/clbwXKg
fGItzkvt1oXsDqfqMCflLqsTKVIs/8fTAVUGofGFIcFe6ayEKwNVj/QTineGihZH+sT/Qejw9/7a
MYPRkBnCbwj1vG9BDK8K0SDMCRcyimt4s2BOHgqH+8mEhJKSCoX6xoUTtaF0aE0KGZHH/2pCx5XB
3KLVV5XPRZzTVQB3nj2TC/qZ3XK6Ff3pG7OCLpXMISpmiTGVcA/WfmzVebH+D90k/pO9nzB+K55g
/Az5sydjpEJXc7d0AflivRpozK2xcARoJ8+zkTsPf9lQ+JdUW90lBmFVrovwzgIKsUly6f9bPZNR
m7ljGDLSIHfle90C4/Wx3bryMmoDddTbaeVaVwYoomxNtYpCAi6G+Cciw7eaday8DhxKry9ocXqV
BC4r7RR8Gupz9vSfjbL3q5a4WBfOsAXuD2EfY7EC6ELOmFXV2M/myMa3sRFRGeZ3JNu2dNx0Zeer
4va9EvChb9MT3Q63belWcNexTS5S6bP3Uqj9l9EH4DSAB2boUPtfF24XESBVKZFYppzt8c7IFxo+
qjL0MyxizmBIpqV2EyAw44xIM6/scEFgMaheHhqeB4xOW8O2HChBnogGN2/YbfzfuIEg9peFHNvM
CkMGa5faYyyathXNXB7oYZQaiF3qRNkXCjjZq7dKbzjy4ox7era7eEIwRnf712+SDU+zuV6Nh6Sm
lub7hplOyFkCGvfLsvedE5qyhjBaBOZh/USPuDsxGz9t63AwJ//8LsNsmWV+epJUhkpQhLmylcLU
/gxxi65I8I2MsI9DRRGKr1LgBssLms6BFUe7/4l6c1HWtkXAfsyihdemMAHH55KmfmdlUGrf476o
YYLi4qlpn9FLyO2+c5zDep3I/5wTpoEE/Z+olEHPHmNAx71wBgj6v3S/NawaGS712TEoXsePx7Ik
lCvTQbRdwvwxebimgU9IrDYbmlHiQsF9s+ix51CAERwl1ciW3y029TtS6aVPuvf6mzGsyb6NwPNz
qBYjfGRqVYMCSRcNm2u13s8+md0W6uB7bOJRylikJzil7gLxa2rCG26sT1WVC1tFwyTSjZVSUwOy
/rnSNRYkXV8o2shzPSRutqQddLYFpO6Eh4LbMZk8RPiXVy1Sjp5ww43p2cbwePSKppodKCGIaeaR
/xBAxjiybOIwo1pjWFn4C04CCTYYa5YMkhR1bpeIyJD//FL6mlpzLAtRq9LK8KejDteTYyCgxtdd
Hs/NHUfM9anGC5fJuWNUpp3KWs0nbFIKnWOGhKuuF/KvInomKVkOsAadyqZTMPzgpoxZ/zvITW/9
x5o1KwA4tRcrakPDaZGGbAlzDOja+lgkUQSqokl1WhbqZ0jFS3ZssiO4zHrqv/DXu6WXB5RhQTU1
b9n9kK2OD26s+2evo4NoPXkjDEDy3QeEcbJbtoYJvUOzZLa14AIkhOad+7FXRys3TRwvEery+/T4
qVc7mMoe5wJw1SukqckNDJk18dQlUTL4T+mUxJEXgjUF7TwVEasc+q1mpx/KyQhqzrrZReslV1gj
lf0aqyKUVvgxzEdcRfmWty2TFyKKk2I7RvmjR19zJYn/xeMUB8CDZ6yCHu/01m176T98ohndpGM9
Al5R+oag9kH79GdeewRvO4JVFkIZSeZcdoEu3fev7qld+8snBYzv0VobhgHTXQ4PsKky/8KTF0v+
zYzbZES+mCVv7fU9vuOWrhMMNfVNc4HaeBoB1WaydXnyTFM3cshKTxLEcCRF3KbJHKT6FFFL6CnT
eCn/l0xpWaKOwsvIUVyGRNwHLbspWptTe1TPIJt6FPyqnnsh95hDgEk9zbA9Yfu6MOhMH60toD1Z
Xc+4lN2uyfvYadgpVpa9C06N/GN3b8+I00cVjs6ZoY08QioPTJp5FySSfMe4GRCWUzQvLBvY8mvL
JjJ/K5rFkckObgumZkZfW1faXLTnN8K8sjo6+rV5BbRA7SqaWWl/DDRB529QfReakEDfp9T5Zuq8
B0J9pLg8xV7ATeM8LZMXsa4IKoK97O61JLeBSlzRy0irOHC1HQ+O72HDbG0bI5oxAaBpGjKs7He5
nZTANDdtBh6OwELjI2iN6A8igECt9bDHo+ZUoUFRGfcjgSC6rPVovWMDlbxmwshezEdqDjpwVAic
sXaodTZK4zN+cSdkwPS5cpIKU6Ba3ZrDJkfbEysmCfVu7eVaNr3xrWvIGWf0RINB7wOCBE08NKbj
c5NcGTeXdOzI28KhmfLKAXO+owuVQyx0o6CcKYvfQyFyTEo+4fvW2RD7W4CIApZQ8FjwTgAWjO8b
AnU6XPkmGOr9fN+8Y/HETMd1FHM8b8rihcucOvW3+IiPH5flYCViC+35/cNmHeFJSOix6RXMhEaJ
QnDRfyi2oN344sQN9Xov0npDEj2mmMW6KlF2nhn6iawan+mTSOYUcDXAxsH64I1EH+3Y4oz8k21D
20NO13gQU0PQ2Ak6VG6b+Yo3+s1AsJbd5wCL2RbCl91tq+M6Ki5DvZH90s7V3Z8I64MjyyD78Oyh
TL8URYgz4BCQaEoW3RQHqc33cqQIBzYMLDxiAmJpGaFEih3rEMklZ9rfnZIAH6xOXlKQ0QUrMzAR
1QiGXoCH8l2rqzzFQBfgzlXKTR08tEzrrwQtT5ZZFSvAPYTEIQJZnUMyxtz1O7eSbNI15u5AMo2k
riUJVNcjQV4YmB01SwhsIDCu2XtQlaj168rO2lNypyurLKcOzQSapDwl8CCrgBrX+/8KCZC5yrq0
zYyAbPPIFWsDug43xz//aEu3ZrKWcFdSMS3AE9FZhKEtx0eQvry1de+aZGuUnn2hW0+FtWvxcKBE
j/k+5bmf4gRdFagHSlt5FKlkFxoav7mLMSASihTaC/9EZN60EYSn5tQEbuIxN8P96cXIl228wpgt
hhqpykxPN3/2d2WP+oJtUPVtoZFdz+P6VvcyTR9riAs7tADueyP7VnY1Ygqyuc3uiBjyaNNxTIPO
+nAwZMuECoCsASAJ8N4pWzE1tg+5QtuN14T7cpQDghmyWnqAlWElg8XUJN/vz8yXedIQ7nL+Qz5/
ybLXmaHPdRvRGe6/ASn3kKxumuT9BZ/uom9ZtJGZ+hrF4FClTv9DXo5VVGSPuRsespJ3qXCpNWhd
67rF8z0Wd+sFw7w9Iwjx/ttglWdSwMtCT7SO26Fl+Nc8jlfnd1yrjFQBvsYpCBgTM0mh1r7D9hGm
geFkKQ5n1IsqeFw8LMQR/GBNW9esqq+7gpMd8zdKQkXzfNt2RmhqhlXiLQsD286Jrf4+wcDFvIMo
Thva5XRQwdAgpv9V8ReokXYAtVS6TH2eCrpO/ySRea7lmnNEj2htg3MQSwbQawm8VkS/vWCEckla
Pz5/2VxL7d4aLrO33CklKdMSc6gK7X4ef/pNHKqOzP/bF2NPlvc+klfjfrHvqJYRKNXHLPLM0U97
aVJEjwmX4jOsRJjIHe6byOoPHRgMnPAMOzQtF9oSQ9451+gHuSDwd0RYv7fnfnEVoFPMpmAueUAG
p1f7WijfQr0sIc1+IoI8DBc2HQTRAMcDhVaGaMIWQHCOntEnz/ISMjrOcsjs1yFyo8qc6t723kG8
FLgIA4x4tzu8kL3DmREuzTIKnaSJV/joqwnELaXbIhrZFC4JC2aIpx3fWJnJO69HOHS0PDO65TaV
/4GN63qS9Sw/MCUEexvSDYwcZwLXKZ2d5LnB1Wc76fP5uaqTYPxBQfTEdquyiubGqOunI7lsb1Wu
pB8giaAqoCe2LI4Wax5X9cYiJF82Os+VlX8YmqhFcBwt9PpwaCQsmzmP4xJYl9tQRtLQ9HsALTAr
F8VwOepOVs0vwHEjHDRJJd/Vbd9W+7pEvuadtn7lQMY62OnH1Gg1gBJrO6lHR6l8eOv5X2E2IZ0P
hNWCWg0uGgpRzqjNfAoZVEnqKk2SO0EE0q1ha4aR3/uAFkHhl1c9cwUaq7n93W802FlVXjwez7jm
xhqcDtWtjuaMTY7cxjJ56b9dTLe/6qdd2G3t8/2eJnjZibJH7fgUedkHjEgVXieJPVslHRaow7dE
D1QQhlWuU4Jm9JzSpj02/MIiRnjNeMyPNbYFQBB4Lr+pac8U7rTaxRnjl9DYcF3JPTdUtaRWbQF8
mg5TjRLRbob7wddBghftu4U4hTv/dmF2j8NErXd+sSnRJUt6+uJN2wPoXn9Jj4eWEBHZO1xXnAJN
TsVkxmL8XRkpl2O7jVysT7MjuEEGyAnSsGjkTw6fhMT4EVLF98EpEyC4pov/whU0azOF6iLc4c6x
6Zw257i8rP6LW3MhDUFsWDi74r8asM3Rb9fTeZKV5omS+NgIzIbbl5thezrqneCMDBCRiQonJrjA
HOiMqxXb/KYuVAOxsaBcAEvLH4HhFob3ef5gBLdd8SGxJRcNPGvw5IZpHyABbS8xkbtyBLinrgAa
BG4537KQeOv6PkfWfEeS8RzwlmTKvy6NiidHwKxsOh4T+7RXwhyxuyPLD+vdIvfntE5GkMKAlcJm
ZVs+3TSHdyIPC5QxmdmXMypxSoC9CEqVpEx6ALwyfrBldHS5TgpmbWZDtGeoC/wFpI0OuIXyrwlM
3KueuCb1+F78SUW8lyxHPQp1fnqNwCQoem5YdI3QjYJFlvh2cN3IPYVrq3xdu9mNtcbqh8g1JPcC
EkZedCeQsfFyDvctLs28MP1cH5/QF2/552le2aUkjENYkK4l96LGG52DSiO5/QDMwljHzJk11+Nd
SYD2LodiOlZid6JshL0Ou3cdbXFJeWpnJjsnLlsmItP8LVBTdRy+1J8b2voq+RCcqtekZArwv80D
Ac8dDD5NyYfJRL9W4Wl31GlVGFAd80yRusPYPAgFZPqi3gbLfnwi4MPhjQkHhk8G83F4NSI/rlP5
RNfoDzXI8/PVUwFJpF4vZK2johBqNFP93NhsFPAP2b0DwDIu8PHC8pg+79JmEOrAYAlJLZlXNKKr
HC7pXCoZShkUkibDanLDnzMMFPZ06KQ29sYhPO+rmglquitjNtdnO3sGokA2UnF7ccvAixI2Jxgq
qghlrxDgFLrcnESSxYJsKnoq6voblEBQMrXIl9gUYVhQk0PNCG9I1ahCL51rD4i2Q84Vy6JA9cKp
w7bMtPiIB11lvCVj3TXQNdo5MK83II+/Oq6WzNJE50B+/XG0RxxYY78OHey8OCLLlYDpWJhkfkaF
QakpABCOCLzxGsKN8HVTDALrJ3macLRjBcIneQ5zZZJYhqMojEOihjZPcSXvxZCItFlCZSY69xdS
6aRQoxk3kgZLPV42zzhyrjrHJSdRlxbgVlROgMl0HWYF3s5yTRC3+i5B7Qubv/VMkkX5nenBIneF
E8agn1hILzfGQAZnQqMFPNUB9nLUEulJF7KjFR7qHstZOt+dvo8vS/2PcLzVNslvGyZDsobzCFyi
QplLbnwrQklMIXpWXK8KcdZKpZ1TjiuI3lJrjbTEbcqvV4GOGhEAGpjFM8X377njh6JdoKMrQcKt
K1zqkvgzRm6Tn9YOpqjCNDMtchCmBfMVoO5MgRsPJ+lgFg2fWpfADXyb17tNX6TFAVUrHmEZlJdt
Nz4BNS9OnqecToe5qub5rDxAhMx4yOzNUJs3zcUuQPh0BbYR03pnvWCA2zlCozbmP9xvI9Vo0deS
w1BU8HXYyY4Ii0LEBA/EvEpFFnMML0VqafRHy3QFVEy+Rs0g/UVyMhSVmlCBaddU423NEgn9bm7R
hQAqB9Hn9rHt2AV6DnJPKDhP0Tsvgy5/Mo6SeiJ0dlILaVM6hPxtO9//8OGvy4cUOxl2oRUrUrUP
QGgznArf8bZ69tg5fw1L4t6OYCpGZHZbl90DXwJG0cwZCEIV+IW//BwyunhCcJ8eFDkaWrkzgr+1
Ktwn54KrVttIlDiNcH2PeAULQEJIPtvywLbLerj+4KJVxuDwOSIy59/RtmZ3J27pxOg4km81OVyg
NVGlxx8V71bR8+ZNYztUzemXsnpWojjxZhWa+2ooDpFv8cIfRYf13/PNin9m3TXxxIz2aMPA0OLw
rOft/UInbTk11q0fJAzj9IvR1TBZAVPjXYvrtxx5mQfwEqNHO5qWo7r/MTUmzfgJF5muVVZn0jWb
MUn8eM+ejwkvvyKHUEHVRV7RMo/PlsbEXyqVoQEiV4IKokhGn4/yLcPq0Db0eMrSqsgBUQYTuv8k
Pa95GdXVP1AKc8H0m1YyP+z8KvpWVjOtPeOtLycrcXMJpeLSPjDAMKHQ0K9EvMKGYVpDdmg4yDNl
KwgSxhZSN2CpfYsIvM4MWPjA44/k0hp0El51Qy14Na1MjIrtmBz/Bdc4xld6l3OKr0LgkBIcR/up
NLqBXn9tKaWZ6fvg/DY8RagOiz64eMNNEQOCBoOCT9PxzH9rI8QYD/RZ9M2XIWdkgxTWWGG0qiUA
xwHU4TqqhMy0OIERDjlC24IlY/m2YyqSSCUYV9Sm3L4ltkWj+YSfqZ2fzH8gNxqZcb4JOjHzLZEf
1w8BWnXlIsyDrpkMytXnns+HjSadQrO7guZPZ40RC5bEgND1/S+cYxQdjPVs5It+aSTndVKg+dfK
92A36eg/+vJtFVfNfjaUCPHobFIJ38CF864GUMsWE/0hJ/NTkFfnxXDtXxsiCOCivEKckmVp9Yud
mG391ox4kH4h2HIWELhYAOlhubkSfyWFsFujyfzALSvdVjTxMh4WvqPirjUZVqBonXGv1mJVYgPR
1+xan4m+7dq33wMosJECsV6LBNtA7D+gMAzkcuS8/WJ5mewbV01nUoyC9hahBfhtR9A49QW5qSos
02vYKueMuu+zkkJeqKpQ32H+63q+pEZRgVp+aQeLBECrJ4C5sFVVEwwWBcAFsVtcpaPKUZlMxX1+
X8PqoU5R/NS5DjP2JXKUVvUFLMNU28xm0oSLXbcZ0QBR/9ei2ql6T3tDqgd8ISSCmKydvKzVZ0ph
l/KQ2m6LllBVKLRk/Yepng/ZJxCxi5ZfzCQ+nAEqzdRRxzlT0vVl3SG4KTXMIrT/QSsestXSm6wA
6q3sIPb/kM17LK8LLESK5gruH1X3MvnqztSc1Jnqmh/vHnsZm6Ikqtvmz8Y02hYgnk1SDBBvacll
2CKeLC4UIBPhO+/eZn1snOKEeJ9GRIsqrLK9/pv4eSdAVv616Lr/6k8MLzOZ+rp5Cn5U5uApF1bI
qFJTm6maf8T7G8N/F06lkKtG/ErUduOBsN8XRyyQl/A1PXWmqVgMCA0CzredyI734y/5mCsCp6Xi
0maTOI9HW1KjoUCkY7hMeEx/3FyAUssqqHhubL4Z4JoKx0hTpjZScuvSwKAxJ7vAhA6VdbSU/obL
n4xMTi8CY0T4ks2cOfMXRkk7NPXHkruIOGdO+TWU7+GBGmWzInbreEGaQjy5eRojtRs/1igLZ4Vc
4OC6lgjKSazFL5VCVtjPAlqTSRW9M+QkTRHHHSc3uYyiCBivmVc/AMLVPZ7hrKHhWjh7Q6dUJug+
FQTfmBIIfBoz+TmRTEx8o2zk+S28x/3OSFs/HpIl3h7ECmE7wORI+pkrsbE+yH9lKJZ08LnuX500
+foKiw04KXj1BsQa1/wTZFS4DVJ4MZ5AKzSiU1U2XwyR5boXvkzgzWKB/59R3js7WLzyTTWBQDs6
OL/eUZOXVu+/MFx0Zs7jd7mfcORmi8TuiA/h3WyFQ0pOtwQrDWe/2Ao+rSxafeEv++BqJXaa+toS
F10RR2OIQGw3EqBr93uxLY7Qno8GAKfLemDXjHzn44zkgP+JOTsjMe8ycYq175sq4tiEpidvpzWR
0nRwsjrObNfkbhYvanzXgte+qSeg5RHu6rOEal5bxhD8l7Zs07zOsNLJAEYUPvPVX4AW9eFcSCJ4
o4OYYk9hgejK8x/1g0F3TEq5qrwXfZrELzxUlCqoW1ZRWvPKQuJ7nIFVWvAmTIZ52GvqND70vC4z
tF6gMqy+t+nWO6fDH+NWCE1UyEO1zakCzYGnOs4Rh6afjYYVJvzrRZHCpInrFY05zCgQX8rXGXpH
1AVb/7/pHQ4xG0kNFk6bSz+su1PUHhLwEOK8WF+yHoUVG8NFpNg/4CqSie6pcx6G26eLFCt5Z0aa
dNK4ybxn9kEH1s9J4qImSb9uqR/TDYtp5JufaPFEgteLFDxtsygMw66U2GuJ9k6RWB2dMuMO2Din
6mu9zME6hVaXe1gzz3tQlfS6lYjatx+cf0fvTgJ/m27iEXsKEO0XvbTJ9elAqXtJec+/JNBamK+N
buCIrYW9oWzZ8Jm7aXiq/AXkGiK4CoygExq2pefuX7uVn+GxiM3qHabQpq7/ZXUrQvIybfK+IEEY
dIYru++z8TvLep87CrjX8412VDXsVAFp5k9vNoJnQvyoVLhQ/cVJGSVNWqKrrnMYJXS9rtt6aruy
r+sEiFUJxc/DAZNxWnx0tgjuqH6BMaSRldIH8dDRH76hH+vFCP1CVE9WubdWy+g5OWp0iBXgRQ4R
nJ3ln3WQ33RYx7ybH7SXyAP21Ix0BR2qcINrTaDjiBWuvPu7a2L93Bv/n0w3gqegFvfw264bLlOB
9rrBWpX/WWvV/nZUDPRmyngQDoADQ7tptk2PcrG5Ty2VAGgevY6MGZCNar7HXdULlCuJpdVe3ZRP
f4nlnD1o/HtX9CEdQFHgz2bCtTKKsk0h4ApTuIAM4QSeEBHMsyu9xYjUx5pi1igjwHuKP9yEy/tC
cS+TA7NT7eV+UU2wqBCktL2XGMglkOeNl87Xrzq14QS8P0wwKlAOdEPWwV6e/HQAzK7sZ/MSBoDD
VPTFv66oda9lsms9nzcc3N/snbT1IC4+DyCXYP9Ff5RQC4JAcmTiIDb9sSjMyxNae9qDjeqL8tIr
DoaBS/TAGq780ffuDFEAbn8Ch7RiVCbMx5DqK4FUR9MvbJfY5DjK563d8FTh5R9cD9Ayw+lhxIcY
iesYe1jwwZ5tG0E91Kl/gRXXobsh++oG38pWHcSXH22Pv6blKBdNY777tHtyQISIF7aCdmpraevA
qYM6ebI+fWiTYPUN5f0/QRRKnZdFvXMBtpkWUG9YRH0trG6B9ydDcVXBkZ03/WA62q7PIaYZ0Kg1
V628PBy7OmEBOVPxgo99sJvTB9QV8K9nPF6e1vONnNzwTNdopgMU2j9LhMrzVfr3KXMjLBg/ETzs
mS/yPaI++4jJVMuszfsXO8Kmtm9ZL9gYMF7wHoKl+uP0Gy+9/xWSSmwy5nniMmyXjHSK6rwiD9Lm
iFngP5IIWMM5+uqXiwHHk9aXKMHKCK5c93+hH9KW350QYdzBAAP+J2cCkHGt7V4LkAegHNvA84Fz
Ukw0JxcoHvpl93HTTZnYdaZxBJ9LAi5O1ySbithyixemn8cIECl35hfG0hYkW/+H5/49ba0XapUn
xeykI/MYE72PpAmBv+8kuNDlHnIeeHk4MZjMOye7e1THAWFCl0zPnEatjX4YNi3LwC30iXAFJ3xr
jFQ+QsMkQNaShrz/zb5Jl7kutxI2JuGlzd9vnreyRTmEboN+TwX0CRnHxwQ4MdKc0fqd0yLCEHpY
NOehUaAX8LHjKDJX2m5+CXL2UzHfiyrNrvbqjFOmgredPqghNOdZhgXjTMFJdYlKTQDU3WluGxnn
SHz7JP83KDKD7p7JUxu3Fbg6yRONCBGiOaX2xfYVUZO6VlVBfEFBBbADtBvRp/82MgJzbuIOW9x5
1sdf+xpZ1ZxKQN2T8TmYyvTvQai/t31SVOMaddL0vuV02c1leRxvTbtudPJzgAMC68RNUbzEiccE
1HSe3PIsIoouSdm3XNLv6it/VP3Y1uQZ7Ny9hYUtH5FrMpOnFv5wl/3cspCWKB3Qls5PrX7Y06AD
HGNeiIw0e4SvrhQ2tn3axcQCviMv6UQiMGI2y2ujVQWIbK3XiUQwllQzu60a+/pjfb73tmaHLgtR
PyRFIVjHz1wTNPRyecLCtdO7Fs915Rq1mJc6X4Pi5e+uobmRKNKh97v4H7nvtnihBcqffar3ym9l
ABJyV+HdXdlqlzl8x8Zprney7kaSndLFIQxAqkwtof+GGbi3UT8M2btskGaYRruGEiTZep/fxsE7
55wrgjzDqepnMmf4AgebDS2DZ+x1Zwfb1iwyNFCwdKcnKJ8p113gynA1AOV6Yjw2KRI0SvuogN9m
cY4VXHQ+O3sis1zInoLSHSFzvyNTppVnI7/OW33iVMU3uL4qdy5Fg7OCHXtsaRunNfdxYO7CzB76
KElL1OipZDWbkOHWyXNxGxpt9Xy31p5xsTfe5h1H3obmcD1oKHRyTFPiqhWMB/mUyUsv119nzqeJ
tThjcjLzF4E0KpZ0H0Guhmrq6CGBCQ1k0jlGnAzbttu5TtEockW0c9sF2tYRFMyw+ojiF5g5JmOI
U5rGyb/B4qgSO58f8d65gIWoe4LrUY5SNojdsFcjcjHVdftLRSZPOhK++cIkm7x6U3BSe4C2dnjL
dexJAygEC5JS93oj45QAXe+11Ku5Yi4FK+2bSQcz/rwhkKXcqdTVAIOARy7jyJJT74cKk8USSKfx
yR5FMl2EKRoVCxLXEoc3VvKtZ3S98v6QwmNTwMkCZVH8EWMGCFd3oNZ9+dbA56f2WtCcbk6e/SYR
4MHQeX9ZByykfLxRD271kjPZgld1+8XPh8yx/2J4sRRuRh37qBTUPbNxR1RWTNYWUAWHoWpl1AU0
rLqQzXwt610OvkWgU07m3N1ecPoNvBjhiByxnvv3iAZdVI9ZGeEteHtuW4Fo6gemXEozDb5lRrb2
G2kAW5a6CsObHr0t1Ga1rpzpMPgh3fbrbCa8ZYQY2S6+uO/kS8fittrtMZiDnU+v10NMn7hU9hal
+GZSJ0ob1ToTT6Sy5JIYe3d1qjPKyZcfxl9B4zmbdEeUaFLrZg+xGCPH9qEYNqnSBWp/VVB0d+Hz
P3VWzJmqNq/C14eRKlkMVXHJCWFgm4WH/95dLg5HicWEYOxDbq0rcII+fc7PR49QwLHv8/RVAO0M
7AuYueWj13bis+dsJI0NqmzcOTrICstFBHNfKBbSg42MbKcVeb24TyrGFKi4IeRQWq9bx73eRRue
fawnbNOVH/r9dxAwUHCAVJOXjy6/Chbt2eYJl8LlW0iWThSjzWahhyJqi5yVCebgaiEfOLHIKXux
uAxp2WVVYHxRJ1nQWRkw25Q3QRkboBKoDaSlvfi99gucDxpZ9bIWwIppij1OWewa3Osxl82dpopa
fXxcmKkFAmO/4gvIYblT0FW22AHzlJrReNFhroTKVhax5655l1fdnd8JNYowsI5c0t1BWQHuKxbR
y85VAmvY6d1HAypk4IFlF6o9TjeTLkXCKWBj+VQkUMpCUR+A7QjwLumT0MsIMX+Rn+e5YDRViuOx
dG43gjPB0FKcP9oZ8hegKKAfKYvr8YfsuKtxtmAA1VOe1bna35qdekzAOHKf9x0xgwOyKXuXrw9B
9RinvrkgiL3zfFvPMC6ds5vwa/Eeaw9Ar7HbrCTrSypLYbqvkZ8x5usrkkr1oDlKkTDKKe+qYPr/
CnkkEYP7maoakcNTMjYDJMUM7TSPEa7iJ8uRnKSX48wfjVSpL+Fi4uldaNxf6EEreiDYECbqLkiD
ioH1xwgff4Vd5aCK1O+v8jhtIgjSxAZxtlxorj1+ChShft4D7xP+syOBzxE91IXunz9v2w9YjuQ7
KLx1I4rI6Cr4GneNDrbpcb0rGjEpRImMcl85YTAY97D4kcOtIEkoEs1/86PQeDPRlU1Xci1SDoHq
VyouFTP8CGam0qJIaD1uMjIaX99T4kUIYGJqT8LmPtkdOKFeyx2OqllhG6WklvQXbmuj2bOZaue8
UJVawal3rB7LMKE6C4hzvBXDGWYNaYkLun+H7cIuIQo7zyMA7EiknCQs+C1MLodPFSSQLjTQDaul
Kq89un9/QI+GO7kus3X42F3EpnRnE0/9FvbVL+eSzXMvfH9z1HwQGaSXHQ3eaY8La2CtBaoQu+bz
6Y9OKKTsNreStrDEiNTlV2gKecCxWJwE/Zumz/Sxkh4CC7PYTHNomU8bw7XIG4A0dr7j4w2mKwP7
/fjOkm9+KyxFklZlqiPHAlYnnFxF0ofERWyMHSF5vk3C9sLJxRhsFRLOpUVboKXd/XO4vCe6Afz5
+q4uHlQTHTt59ZOxkNzPK8aKRVbkWHiN+ql2+mX7/YHH80XEVfZbkJu0l76TR1yW08Ti3I4Samql
kXmBo/hFOVp84VTvorzm8+XF5gb5jwHlglsLoDPuHquY/E2Dx/yDC7Zj6S4nExxxbE3wP9Q+xZ1l
trpHrMp5ovoyWiMbywrGJysG2L58sYMGVG8NMo/t41gqsb3WHyQyqoFLT97SjMK84flajpgkVIP1
e9mcc9QOhyFQusqsDMqJd2lCelbL4pGofKOYfmIBxeqPLUMi84R/SvDT1FEQY5vCY7ZxS2U2/heF
tN4uBebaWnxf0/RtIjD1WzCQnXCykDf3PaSdTd/fA4O5o0ayy01SwHFqAaQ1QuOx1ADftlEy6OTk
4YxKACrTU9QhbgDPz+IWQC3iPhxjuwgbnjr2p+rt7cHhL9sQLgwbTnCMk3Ueuo8gicpqF1ndOOLx
RKCzP/fm6R4/moMVlhEwI2Aj7MRbpd+CPv9AqL2gc+aySyIfwTP5m8uVvXTtwk73RpdZ5nJxH+36
nT7K+9BrO4JfvBCCYA3Dbfp4fr5ykmwc0oJeGZzrU9BxVUhDe2R17gmX6bkKSL9H2Hwzwcw4AA1z
h5adZzWY0INw7zithhIuLkSGv6OVyLw+eg7xNS8hl3FAuYFpKwc0lDoDBRsv45++jhwEZTz3O+Nk
kWLlG38IJ8fneydBysI/qmngK2eGkMfQcnl2oeO/Yh9CqjZKmz/kNP2RF3SNZckz97To5wZyFSbX
/id67HbeeNLela0qGN9K4sOxgpggHggH6o5Tj7XeSJOq8WLXDkVvSBJfyI+CoCb3ti1LalUVpQ5a
x1hO57oqJpWKyJjS7W/zdX5CQ2aCKjM+aG1kyU08Vdf/cTm1fXCb1rWWOhHn0gmnWKgI6t7NFLQt
bGypHL14+WrD2MEG1LeQ0IVfFgsnayMQ28yd54cwHUIkxZoseN7aDYQrzW8js42ZrQw649d/qW0z
usgaOAyt+H/LzkSpjxqZQL9jRfCdudVXzhFqhTr9cKWf32OFf20e8iCvVBDsC10U5JbQYYH0B6rT
hR5fArU9UwNbxnTjJ3v+w412gto7ilRD3OnsdmJ85BkmP1MHLmwcY17bKeZxok9oGZAD0dkRxQV+
Fr9qxTh89UtFcgJssay58voMYl6Zr62i/QrMtfy6wcJq6OfSSX7GIA4nmmgJx7EacKjRjMq4h+Lv
aUS5xxFgn76Fqtc0VCgEzE4gH6lcJPB0PQIIiEeErc/wOCsNuqHFva6bTKOAdsjVopqXmCV1NuPh
K7SHjsvOErx0B4gpBfhB5UocYOIacZh9VWxmMtMkeZQ42tRZ84qSanO69Th5sCl5UohIAz6Rt31d
fijLXQmFAeTdz5oncVKV33fxwJW1zZCyHhZPCOp0Y2HAnltht6cokFpvupcFrgyn1NYFKJ5a7rhU
j8sry7+XaJwuDSmuIUX0z/6JVsg3PQPPW4ew+USvJnAMWBOc2gWT9GlNCA+GwCjnnqhJuljVUhbo
ktHpDBY3bC5l7IVZ4oRl4zVNLzd1YkJOk6D5lnygFM5OSfYc+JaBviCZlby+DqQlZehsyBVbwbo6
bS2Ie6ZgJKN3yEsB+BaPWfis/yzFSeaifSDqCUpuk0y9rzd8z78GW+xBIpGEq3ouPtqRHo5chbN/
3jBy+YLXxpVP6DbMJLmGIYkjPhDVEavvLuIkuKivHOcPazHxUH6DV0ZOP1cBDuABJedOPsX48LfH
F5h5qtpIyNDZ+IdgiZsDK6lASvtr68GW+exjsAOcRlgwKGlmKRyUuKvR5Lw/5pcckrhu2SIzFZZh
icdqivyYZ1GNRt7Tis/3XmAQS7FSFsszGIVGWQG46TDnObqK623K7tvsUXFLdSyw6Nh50QaoguB/
2XSnIkLnCRPFkmjagkHlg3FePMtU+/fL6TfE47bllBqy9h61di8ZWxdEfOl0CqOvVk2P06nHCbRE
SZ3p+XY7g4w8AuPRcoQfqWVHqtvh+53dG94dTS+dl+znjKi1k0kBW1oMYQ34DkvC+d0DWkvlJ8qr
qtDzDtMkoFSTkRMvwU1E7A7K+OLq0nUz7PsScZFckP9B2v9OnusPzr6xH5l9ls+Ejup+34L7RV8o
a61fcsfusM6CJ8hTW2sYREP9yyWD7yghkc83GKM1lnHF8+l8neH2Ga9dcytFMosGeMBJIvyjqQU8
3P0RXjMq0XMhuzsIWKMT0F5P7lP9KHU7j454sujfjJvwCKgjl4Qlkoz3cnoZ8/J3zlQNV1V0ceWi
0gCcr6n9kn+BfxAhgtYEug49177VemWzLgDjcqweNrlBSOXQM3IoOIzS1MGGSBe0byJAl1UPKdyA
QR0gHz0bNGKJHutgCCwz49EKQXYRft8sKcOgMhXzqZiOICovHPEOdjN33KG2xDah9fbl3rTuJhSg
cI5xXVzXLXH/fM9VfzMEonLSUFIMVqViElybSrBNKi3xU9nBBgsGU/WRY8d9nw3HXCUykHHv0mcv
UMJSVSq1KGoBc8h5Keo07gg8qnmCLmVbg2NMocHoKAnJoaMk+Rh8wJIGMA/mruCIiKxYeqSXRkfD
qn6U+I4De7vXjvgCOikwDfxaabShng4INB3GOxHRDUHaPBX7S9BUCADoNsrU7+jrpnf98qEj032a
efg++ajNSUUgCY1CprOx9/i7bTq+IWfk7jnGGVPmeUxGJeUx33kTU2TthCiwqY2JNLRVve3puUpl
gZBnL7wMXnAToBgNWMeaZIvXrgthJEwcBDcvlUOliko61efipsymZhYR5FGcZ9d4jNqKt9C+5S8n
EMn6mSPXcqoB5Qdix6fDpZICG5nUW3BOR4Pju98US0uj3kjkli4p2O1ds4OpE3HRUXDv5Sie6b0x
OfxR/OyQmiaTmBl6xLwoYvbStrfO6X117W5JnsCtPr/9kTTwKU+6SMH1lv21iElfPTHDMLGEjdqe
z+khFQ1U8q0U7aJfI9GQ5UkLUDkXgQ03KDTEfCZmf+6etkndLDe3wgL/RkuDjsegxi1UxF01qaA6
nU38F5pOe6ebBOonD/mACQtlMrqlbYfsYBlUGX5JmXIgxC0StFhHxREOfObQJUVrkWOCJb7wa3uy
jgaIZHtg6M+F87frolHStJcTd1fuezy4cV4KNEYJdPmX0ggWo4f5NOKlpqewvfgggR7tW7PHVJAF
L1RlUX3x98GGJ9O1qaB+qc7q6x/xLgvY1DbHvsofIGsy8JVlVN5oobtbg1BBpGJ++0doJ2tkilvT
RyevuEOWy1ae8AjH6CDkOXydiozl6LThTCjMcFigiVfj+9Ya3+1aGYBe5SiuXuUUfSXjBu9SpdZ9
JZfCJKNEweNvFLp0eXled67d1vlPOszU1KT1AyON/l1vMb/qsGHkKvQOOlC2tNXpYiBjWki1CVgh
OzAD2BbcqHyaSYW4CMP72ZsCq7cpd5SuOCw1CbGP82wMEyQxtbOHkimOK/D6RR3C4Uy3cU3UK70U
jx4RfuwagUaJdIt+FKziqm8yfWa1xNBdhet6TkmtmS2/dRW7Jfu2XUmMaapfFJeAd4r0msEp3RyK
4JTblrJft1f5k6n9/lXq9tBbMuC/8yK5KIkH1J6Cs5ybcwt0/95PxzrmxXF1x737E1x8OXnW6+L4
TGmsqeWeTZ6Gt28duUsIOTrtBeiNI8H+7fphrSxlItbxbz8TH5I5X57rI/JmDB/wBZBqX0R7G2Pf
ltsCRr61RN7MHa5R120rmjCRrhPSprYv3kg3zsn3bf6NNEs55ylJLTfTkYetA5vQJL4w4gnRmbep
dZYilnmaAyOMgPn1oDelSxxufjwv75ST4bmQi9xQBTPpm0L2ZsZLXBCLiHazpOEn8Om70OTP9cfk
BWywfN22rR58pLNABXhNyNUaIyfjA9cGGlkWv3Vx0ilK2Z1mO5v5rpF9FWgPBS/Dwa1+F/YkLSC2
JPrI/cGddU8UH5/gBD7QTHWh0TD//4EGY/QSwS6ggF+zF+hXm0sTRjC75vXB9+4E017sK+BeOoYX
yp+ATwJrA2ZXg6Hk1erBO7IoHgSQ+pfFRNi4qSy6u9byum9HX8KuTRAf/v+mBDDBUxs4UW45UF1/
Ab6xsqYKm4J9VJr4yiOZ6F7vGAIZf2sGE1bDfVkfrQn17DuD9PgjS4ZmFmyXfAlo3YODW/My/mvk
yJggsYJLUhCSLIFXdLFm3/OWhcnkOLtqqx9eyW3051e48UEmbmu0KDnZFb2VqUOpwzmAwxJedoZ/
Ny1jlzfNnw+xrOYWcijgDiMSOoTiSrfRyEf9mzURDkR5cdYi+WbS8DLPp2SnnBPPyui25dXWEexg
Qy+Mton6L86kXvm+m04ZV9/8Nma+IdoNE0EZv4PES4YR/cASns+eTvN7GNAsxGnZQiIcx76Rehiu
XB5eFPZEQIfBPHXMBG9XdfP9X8/wtMMBkNI9YzGufxBBb9dsJ7rY5bPKa5fjfS3BOZ7Y1h1OAc4t
AJbh1IJ2hRiflmhrs1Ko0Rsafg+KEjwSU18nRxN5Rrn1Fd8XqxXuNDV7cSPIYIlHgnj78fonSR2T
EWTi3CIeLTAQ+DaRTJVxkvE6Uk7KINPIn8WxKlrdTyqGY1ml3pT7FKIesVAf2btdv7E2CRGWGDuA
eyt7pmQeDFpnMZHXbeyz5N5mLYSQNj76/x8jQHjTtAw0xc3crrEmZkNtScz56NjYlwX0wOT398Ez
Jqh6tO+821VVIq441SLfWDgn/GlpxrL4F6g8tr7FzZWBLzCzKQHYI3kkrOZvOWt6cXDbh/TbhxvT
ga5A9iw8KoAkSQmB/r81FIs1yndlhOWWViEPNN29ALcHuxeaB03gisvw6Ujyx/gdxdlPfNdycv14
RCsGJsUAb9dcVjELMPTOJjnpUviCz2Nmca724SgfMkCWsjh544qW+9kRj/CuobcU24YYGY40w2g0
TJ5CQgyTsOb6MR8ZMIZk6Unqd/JwX1Qu53saAfmIfMKk8lC7FNnkMvKxRJfaSAyVHJ8P3K12S8tz
Pzz+rkxFgTgQttwcDEMsa7Y5KIW6x47HRHj9msg9+ghXc7PyhUtMPdaNPQIqxHYO+D5kl59iMuRs
NkLLFiIAuUaMJeXtIR7mYpHdO6uqIfM/iNnobVzp6R06Z8qouCJsUIRi9vq/nns67l++klrOLGJM
krRcmhH30pFsl7Q1T8DiN1BEcRelj3cPv5Im9RLhChcOwzG2oQ6JmJFChotBvBG2GdJlhlAc3NN6
5Clnlq/tF2iBDtLWok4HIhT1dM67aWVi/2MRmNzlV6pQyp6oEGXIosUEL+8A5MSdIMbl2pMzLdWM
XBTchgiHK7po1Yr5pvsLtDeJzb8XEHvOFeGfX5qSt+GcIUkzadxbrvpV2AsWN24h9npHamW7MDgU
qiw9ZBcghfKYTRZfgorW0YeqZ1puJZdRBIeIkoIYvljGJwOIjbNZOIhkwlZMj9zvtU6Slm+mAd2C
3HZixpylUNCxDS0eioyBF+vJBhULRKUNIOxxhB2t+vWE6OfPVDlXwMsoli6tffwSmyljNzwJI8Ho
XL56FX+SrKmBXXshps2Ie+7O53X90/tytQBBsziS6fPyM731EO9QhITD/Pnn67rApE41AwkQifq6
mQallR0nZVlhdcfBqvRF6zsoOPQ/DxVM3tsfhPJIbepkm9jkk1m6laxg7V4H0STVDbLE+Sfnoc+T
Xs3YHp0KYXu7OXdqMBcDbDaBli5JTlDKPwkbq5kqk15Q7FB5x0FxThEepAaIQ51YygkC86vXXnaS
fA0jtD9D6IRz48fmbRnlmEeCpnoBkgblRyBFnW9XEb2OhO9FW3ghxfJSyfk/VM9Pbrj8C3lIEgS6
ci+YDr9bD7C+FCf0BgJII/V0+Lyk7Lf1xbmF2hvCc4qUFQwrXHrl1aYBHUdnXFCuM/5IplNkidwM
cWRzaXFKtoAwnFnuJniX+O/e2yFQWUsSgamC5P15geDw8p1Hk2TgP94li5F2DgbVbrpEtvM/ECDF
dsfdETJm9dgu03QzihiwLxpcZgAKxGIO/hAK28GW0rcD2CfXL1Yez9Pngecl/VyaCFF8FthV9YYk
zmlY+6w0B1V53P3ZeoZ6iTmDl6M03rqLTvEEqtw1HZlcdB6bQ3Hmr66w+8Na+XFQIlmGb/p3Amyo
ThD5V3CpfjBC5cknaL0yIXrKJ4A8j5dcGcNuE+rn3PQZ4HyvW4XlYiT2WJsGbg+afRSeZN0fxWRt
iYTtstCUIzeoVQrO2w0654lQ65YMo0xqso1JLyYU0dTjAvDT8RtYsigkOTSW9BM2A8UDF3eb8eXc
nH2j65v1jqyTLGBHRpvcurWpmmz82i4nIN7bkiyshpI4yk3+MxFJWiZHQgFf/J3u9yVMyPHz53rt
Vod/sSi0hD6j9q91XGhbzYi3px77C/biAFu4PkahikjEd/pC6SU8AReC3/8xZ4ImLlbC1P/JXVhv
0+veZ2chePJ5ffl2Xxdyqux42msZeu11qYvTmRIu0b8sDK9Rmu62Z4UqPqqIKHZyT0ZYCv6M8W8n
ui9mQys/cZ4Swuyu7YchSUIBrqlyenTcoK3qVZPCu1mHR4V9PqdwNNZwYJTnal9QO8/bUfbT+GLU
w/geWV+vuUxm3t/PVag3NfiV/a5QpAdgS9P0i7DPMuv0IRbo4tgFmRFrxe5Yqfdb/Z3K6EQnOUHZ
JfyfxAgt5YhNMLpSG6+SpAX+nYXTlX0sFgR3fvJ0ghVpM5ay03lHxKZjlrHQ+gU4pyAdYHw4ER4o
ekN23cTj/V4mIFI+G6OAM0rnGPBpI0sWXAzFYPWbLqX97w1gIJvQXRZRirbqlJ/MGn99Wyn0vHzi
8IZtCr5uC41pmfebbqWFENlpplO8s3n0ZiXdGkBBUYedkn0AIHP11B3wI3vWCvxm5fYV34cP9VzY
8nvTOKrcY0EW99nge6+zT9ULk42Bf6pbC3qTtfTFepMOv5ktetvgdwzy2DKQwoscxJg7+lXwOfQP
JU3Y72simkOVVHtQq/CuRF2Z1eBn1iYqWdTDNH3xjqJCbnumq8tjW5os0crwWeMpEPfNNeRndA1f
WgtxcE1p2Lrw0s0JAO8S5l42JTIWZW4OwYdhU5RExvVglFuK3ihxxOJ0IzruRKF0LBBTbik056my
EcK6OKpGz2reaktI70npFoM3B/ZLVmjjwg8iQWc+zNbyZQ3u1/K/JMzsrNkkx6KiHeBMtgdzcBXB
82DzNW0/HnzsxW+okw5MI7WaNOdkKwVj3hy3KGT8cwHQ9BxhyqXqbEkti/N3op6G4kdzuLUPxqgn
+4UPemski3mCxqCu6LhDSlLrA/vSk8tZ3b8ks6YYr0oLNFOkRmlYJIFUTD/9F5CvtHO8yqi3M7X2
Z8s9QLgHXTiML22E4gNkgim25mpgADMdusEVmfDmd8+oLomc+LWMIHIQaQcyOfZSY1D4bF4cSN/X
6zEVj6VMNNuQ8o5/1HwOm8q/uY2PRNOawNNFaKTv2XJ0ukYJDe1nn6IF6YcR6EfklZ6gqhIbJvf8
A/iXKFL9kk3aGYpplis5Stu/SHehJAkFnVM9En5ppX9GhfCMUifsThiPu40tm5uvIMowmRwzRoFF
XzE6xEQphndNcfjPdD8/GR8mqPKVBO3zJqilf5PonKAyBLx0/TSaQfPF9G2Kq+PWobn6JgNUjjIu
CLL1DZvfi5us0Xn8DCXHKtvkXSzU6ItWbr1tb83uU04b+7RZeAc6qSyGqcX03Yf1oll9y1ECdiaB
mSQnEWmYFsNPgeFkST+PRY+Jb3wYX0I2V4uuHL8aQuY1rEyeWubMWEiqLqrcTwcRezVaMR1xIU/z
UZ5YKyVkSTNWV1g5JBI+0qoAdZl+h3iJEGFdzIBs5Oe0a/Nhej1VCeu7FgS9vsFQs0QrzgR3Vrdt
tgmIU/HmKiRtLVsQum4XAFfekVq3Zs19n9WjEGOMjcDWpAzzpljy4DgycFfMQvRstnyAAQsJBkYx
gE0AqOPA5kSvon/fsZ4bJTfGtRXPDUEVjtl67D2aiF8DMlmEBw02VxMZLMt+Y2qp/CbwHnpR+xGX
K1moiZcpBY8rl8jkWg2CzHJzfE38VDu37DtWmBkA+57WMTlmS7Q9wNV6rKrLt92d3ng8CDcWGIcm
8ZX5YrGkDhtE5qQc8LBoGwyYJNzX+0NGI1MYPx9c8jbnIzpMvLbjq5sdeulnQ9ihxYsAYotFn5Eg
w6omhRMwYeVB2opaTOKk7z1K0BTlQd/l4gYV4MpAPz4cvSaJhsnf+OY/XSqa8GcGusI6O81R0i2R
XoeyG/wnvFB1Qgopm6qr4EqoEunngrCP9akMwSS+QY4yeok2RjzzU2KNPs2TShRc79XkoHqaUqGi
tiz27aYtL0RO2bp7H6Mn7Jfv7CpYYt3S1Boafw6I+Bzf5Cq8Dn3cC+49uZgAsDiRvz9Jd/QA02Ug
82apk41FMON6R4QpAFeYS0bicsym1Bd9lbJ5KNmL/QQQ7coQMqjNnKzWD8EuqTgaFYdYSw49wXxt
M8urjnduAheHbfETTT/+JNwG/xGMFQMKiay7vXnfrHt6ufmkIu5yvj/GASKWIqlJ4VzFien5naY5
mxWvYuwLtv+3CELMP5oHyc1LBji7tR9YQMoDMJQ1f0vLCKMzfsUUOdZnKIppohnjKgTn51QPIhrv
qXHtMlrTv1S/dyip1QEwb58iGIV4w/Mak1zfUEseupJkQ3C7tOAyvYNR1H6py8rDq9MsunUCTNau
aBne5STPIm7Q2R/sVQcUgFM38HNttVQtrejyWFzoXxB5g9ERKb3vTKYASMamp/H/B1i4nQQ3xfQd
9Ax7Wm8AKdT5lFSJT5pP6MavxjnOoy7g3OmocJSMalmT0bTvEF/EH1Ki5og0o57mN7XqvRwmYOCI
nSbel8DobF8knLwV6ntcPGfGnClTrB9S2GSJw6gx33Qa+d7sqbMmPO5K7L86frmFKUKkXj03sQIf
rh9NTZ3SBv0nMBk9Axm0qH2ocFoPz4WaEY77QCNPHGJHWHvVo6BeV61NM8jpwSoMkybhB9UIxxF4
6CSTZ3ViL8xZD5w7smrvQ5OBLxKAnJw8Wfp8rxIjG/jCwRZPmANUl3XvXhzt4olOFxXsv4sSDiVq
hn9zOqfW19ZgDPt9nKrBPnJFNft5LSZqe4u8zpWlIx5XfZEpdHWFbUOTxV0ezNvLObn2zAIxPhd2
uHVPMwjKBKATJBapyWoncaeBCFF4kIePW21k49DrL1mm0OaMXoxOPRE0cn/9qvrO+AlGFef3HBuD
L5qx4iYrqHxmvK27jAZcZo8MTTzNtZA08USlkpTIHyLOB+4xOJ9IbHk9Fpw18/YDpvxoG2B+JOFR
ERZmsYiGLVyfMc57zy4AxXfBPHgQnP1giNjERxYnX1ylIMHwYeyy358dsBkG0dWpMnq2AnWq4fDn
14YlmWJR95umJrp/Ts+q4LDHRCNwqt1i5rteI7tmHOWfpdaMwlS+8iX6GRNDmDbp6X0v8VDADFvF
9tChX94hwLSU2suByBpOiU1dPGWh5xLgSts7xucZWfrfFHkScvLlCeCW4+yEiYyLVVbc2hZMvrKZ
gEleoH4nxwpApdojUFtpUlldika5mUcpMCZatoFlPlpwm3OE+cbR1hSF8bxeaDUln+Ar3cpNXlSi
s8POZyWUQaya8T4wnIZMsdZKEeBce3TC8ACzcGQB24E55I/cS+Gi3BOASCNPJotM3XTjzQUGWI1p
rODL5It6vWP/RAM3pxVFRmeBkE7tJkru7q0OPoiQ1FsEBA3CaqBZBq90NFo05gmSdloDQm/OHxgU
I4QBw0ifnF5/U/hORTB4ycddvxmpRKsolfIRxF6JUXm0uLv6dbsZjI+Tl7VryafDHXvzii+W9oL0
zPEi7rpAGLDpCuA5OTTBH9ve7rqZNuAD2jSzpESt5RgOLgSBoFKBqWilDipqGXmLFXX1CbPNsvOK
t458ScPFhIQDzW7pEvcfsUS1EBgyF4E+IeyKJDszM/bMaOTxjV2d4H5VqB7/pIs2yPCZD8vvWLnK
/Q7S0bswGIggFDTKC47QXl+c046zK6OFbvYruh3GXkFhNdrABtd8SjtJBjHdxCQ8ds8efW/OdCG3
TunHQe1L6Lt/wxN42PhJX/LiHZ5N18rjN6KyeQbSgJGffXdmSfUriTZ9krR7XsW7h+3YXnAFmk2s
owN0NkfUFgGTlpF2EFfp85+EwNJk375qaxENJNFWD/or4IAVwzGce6NuwYfdwjkiKBEWUjkLdvi+
VHy2e4vbbLLLXmakIhLC8e2vEmLk4+65xKp4IZTF4802L5iSjx+nUb31L4UhPH1E/c4gF6vuHT/n
6exP0McMWq0wtQ5cganYSvLls0zm1owWXMfOss1TYchgl8b1d0vodRYA+yvV6tjbXSXzqzScDJYH
3QLsvjFCJrIUCThw92XhPELF2cMA1ZAQjWhKV+uMsDQwnwqkO8GyBPKbGnU4bF2E43709cxvT3ps
EL/YcdnppWPIVm0pjIPHaKYQve3l4T/hpZwiILQNNtMqTdWiv1rXe8DLapbeA1PEmRPtjNeF4Xv1
aqSIGkRww1MQ+51s+whyrc6DUE6IN+Py6qD2I6PnZG1aGBz7HRUpVMDbEw+yUBSBxVIcP9RoKFYM
nGtVgP94IKN4Yb1JoCozwmefVRGDt6W9XihaXJ+rZ6N/xLmSAnWcWB/trutF3FFe48BeReciVOAy
FoHuX7k67vyKtBt2Y55x7/Dg9jfE9EwJoi2nNxtwbW0dX1j2jvH/9pgTtK1C3LqF21Vpr+yRkAT3
28NJBb1YkediWUoYI7jSlEI1MR0gNSTix2vI+YAWZpHta1RsOo+HhDEujbTPgv55dPnngHONAcVD
VSCXfcqdRlnc3hrkkDmmW5XfGvRTraBdaNYv3twLGpVtgGAqP3POZgLuUuSBnkcbobMQK/9zqHOk
I21Wk7Ye4iRvPUaRom/16eepzWho/bnEdt7u7DPXMkx+heAVuvhThRbgBYhPmakO7EsGSRXPK9nc
6Pl+8dRH14GfBbGGObe3//N+HAzoTCgxOKg+Erx2v9IwcWqOwAfGwOTvY+e1vOFIbMJVkYYJtM2y
bCcDd0EFUUzUdi4lRfm7/a+8jYUP+1a32DyVCUXa8eNtsCajJsy8dM/Z4wz18ShV9/VrYwiVx/ss
JQXVCtSXM0F5/s3TTPkSvmT8CgFOUoBO+HTgMJ6spcNtfJtCxv3qkOueL2VoUIZ6m/zURQtB+WLd
7Ptx1Ui7jz1GBTwElt/ldnIheZTLjvOvbgvn49yJrka/3ShmOfm8Qu3TzCejW1n5eTr+0EMGKmso
iOET5LUyfFBw1FIb5QzzjR6OwowCi6aU2/3jweZn8ZNBquF4rWRPxgSca/btivMB58fj77LH8DPH
T3mnuAhPt1ykZkplgSvYvrbwEIomwNtWOk1/2LxH1Hi1ZTB7d1rODdIvt8LuCnogns2f5gwb9HEs
e7ob2F2poOEB9MHsbujNxQuJdnvON5hypi6BlTMTQb4iaen+UcyrwCdrKUeRri2wydTLbkhXiZ25
/LGt3hd7cm9qdxlF1kIu1PeX6qM3AQd0zxk3lf5h1dN2MtHLCrdEm3LbIJlCtq1gPcIPatdTkK2q
QyxEvg32K5eLncQkoBXH86uyPorR8A8KkMQ/6npWfF5fxHMASsn/ay0lm2qb1P3STq3sGNhJBEtq
KkLw9e9fzRG6iOcBcdN8fCQeE5E9iPy3gNeacyqwPGgLT3ytxS16CRRVEeEHsj5t6uQW4uIcXu22
jx51NmD08Xi8JBOUP0/9l38b0uQhfRyxCXt5u20WCLiCjzdUpISB35hAQG3RCImA2pmsMtD4TLOd
WPSA/WAWxz6C1t/uHffJN+cCeIZQ4L5LdDz4v2/HApwzVzvCwzKu4xnasaeW6H9NTFMZ70p2fxzU
jPikUpHWfBlgUjAHrmuyRk0Xk7Bu+6F5QQKcWU+8CYRy0sZC7muUqp3tMEPOsiLcDXfRQJfZzniq
u2naX3AVUFsxsbV+BpWax8PLKg6OTq5ZzjMHAr+7C2QlzQI3No9SG7iBDbFI8irG+qoEdSbyRgcI
BubeqA4DuOS0q6v7khrhq944vy397ynY0/Ueb7smnHt1WaXqRQsXCP7HePZKD50vW9rYoq2MYqGL
9mHqV2HhTolZnqkAia/baZS58Qo92vi8opRbkr5VcEhH5wKUWCPlm6Job6UIPYUMV13A6EVbQJZ/
PQmz8UzJnV8e/vB4zlL5XISbKt69A7PcKvZu395V0NPUrZwX+e7An1VxLCAk1LqNnO+8d39A8YOs
RvDWSXo2xfcRZ7AJQzBMDhLMIzoXEu6ytN03UFyv34jPo3l7ShWBhOYeCClfPrRwXs3t+h8SoAVz
Eg1C7Edb/SYhY/nANH+ghxQ5KJXDq3HMJF/Bem9F5UnI1e6F194VDVIjCVgEL8giAIIZTM1qFWwA
7W8ydDFwafs3jPGx6yi9Oo7M+Z5B3uG6s8v1Y2ciSZRkos3FswsRyxzpBLSU0BIieM8/S1/NO8Up
rIbgpYMMJV5u7E86Cx/hvEX+KQeRqorEsNafS+M78YIZ8qASzw2CFVszW5Qud+VPVz6/iKmPsK6a
YwCfNy0iiO+nkNiB9shpGqJZhBj9icpB3Al8I8B38qfLaHsH8XHjv+LEgg9pLFnP40jXAl9uYAEW
878lRPw4PEcSdxD6+F3/84QGKLP/oc9z5ay66y4/EG53ykIP2I+vxePYh2gGDckzynF5aiu0NcM8
OcK/uM4FcelhwYbhZsZ/w3vde8V7IwC847zKWRFzjr3HdmLKugAyo72ANmGmX+esY85hQ1TMWB8r
UkUpd0naRXhW24MdShfQN7gl7Nj6Lz/QKBPzS+UAeQja3AUN3wEgGheJA4t5oV7TwfD0/ut5Risn
oiugLy4OFQzVcBYu52/S9C2aU5D3E8tUt2NWqw0RqzOV7PHVdgx9frsSjOnB2R9+LwW5XuC7Wm6T
4sm0R9lDDuMNOO+iIHx7XjPkzKtotuf2C9hc32IOzRlFOafOQnsxFdgUtViZ+PC2awaDsasSwgHA
6U5MbSoEzAoEeecMWvhLkpA389HQUh3oOLtfEbIgC17NysFNH/OarIzXMys39qFWSntT9Q6bOsEh
CDsbFvKh668p6xJErh7vrQ8OoAdpXkerBwWscliwuUQUjRdM7XmdfNItDAk6tBZckXSe/oHH7ylv
LBamUaqI/uZiO3NsSGgrS6nTfX0hfNEVGbos50tHLjvnUrpvrJ+p9YQsWQyBMpYbxmSL+zdIpukQ
69iDohnmdBo/sI7in0PnHdWs/6REbAcwEh4qFB8cu4jrizlTERlIeLQS1Qs13LMGFka6V3AKD/R5
A56nriRmoryYYht+CJ1TivsmZpayemR64RtRYjyDwEiP0xhdAQhCRZA1uiBWEH3lFjct/hszt22P
yYh5tFbU82iQZV1aI0DUx8/a5DkfVpqVw/wx+1iZq0E20E+RFvtFz1PyXApZKKmjHQnblHyt07lC
uPDg1YMLa/Z9p8/n87Z0i39ezIGxcghf84uxdZpOmMNLBGp2uGHZullr3xouqHO1VitfIgER5Thn
nKYfSgfPx1xYroMB62Z/ki+GI20VztOj8XSvamHjNOiixwzr0X3LWlvCBv4185WH2c7B4byY7ISw
juNJNeKF4wmCT2g9mIQtil33VcxURL+Bs+lZl+Ah3o2BZzimyX2yXTN0H3XCecGbKOloZvtzdpgv
GJFp2VPjvFEtsowoS7OZ03Qe+F5BQgtUuCUcqYIqHBxEoFR1gJhOpQiLSx4ts9y47XYvn4nT7ceg
IIrgeKL1zwbjDuDwcYjd6Okq0J8b3XLjSH0LCpC9vbS8lZNU2aKN4RzKQjQ/ZlQc4cbCBhb4AsCe
FejUevjKabi/fBM0vuStVhsVEmgSvBPuq+4gMtIiuIdF7Ewjdn99gVqj0/XLgbJSH+pfgbWcQORb
ThYtbDPl0w3XC/zIHvolSd9w4dciytgo0beKij3uJx5/oF70ALtc2gdNiz3oCe7MygKX82YWuLHH
vK+9ZDtuVdNKWJOFboTEE1DwBF37exClPXL6gU0YgkadinF0LFL5RxhMLYTFSXV0CSX6txqNlm4q
6IPcFxmNLI+E0oiVya7emLdXnarwgAvqesG4jjkQnkaGtCSRktMRYrVfke8vNX5i6XNkoBqt0B3e
z/r8YKUlCNBiLJqbdaVQXE6B94Icxnq7ETSBtO/eBdYropgxlb6h9AnquX/B6JV1sQlppqIPDB6u
6yABNe49e82esPnITC/pb9Ww+F+0lODeJTpg9qqF0ODiMmTD/kcaJiPtikBptcFxUwI4NxBu/YBq
/2py5ZlysDtaIz9t/cWWKjwFrRZKEVKkpmEXC9/bOs2hu+4yZnMnD9ZCGWsXL/G8p1PvWISb6gc+
3oDn21eC/5Y0V7kuK/HZtjvo0Ht+kIdJ0Obe+MsJNghn9tlZxpFurDfs0NRJYZyhhqJSmwcDvvip
rxgk1UhihWTuUER23XOH+FzrPECXt6K0U+Y1Rly38tfjR1Amy2tXFHqDaaoXWxsdbpzPVi9xT1Pu
YSzg3D0ZtwTuHWeYUokQMbA1hGFZmGypJUNtAJBsDHTTxXltcwW8xZN3u9ZZF57i++qUB7Abm9Uq
Akcxk8Gu444aPxp8FHi5HcORYtMwYH3ohxCX/3mm+MSsKqxRsOZjX+hWSWOaNTSwpBtAtEykiudM
UFJxzrxlcmqOG2H1YFhlGp2Wt1coWHmZ0G9nINKJ0yZtsZ0yHNsv2sQ39nGC8VNYpkBnHTVJz8zU
/GvNkfJNXE8SdihwQxdxwSxUEHVOPImW30KuMhiovtIGFzwpQLm/tYD8PWmJtiv1G1vGqvJPwNKm
TYanj759pa4ZBnrkJY7xevenS0THky2RI9oJmibGKqmmADAGE+jysdBzKsrZApW5EyEK7qdSrsvA
NGvKBMoTSKbVo2IqslWy5ynl4lOBUhBGplJ91PPHsrTzJWviLbnc/TTblJiBEqS5Hhtv7IeLyrhB
aCzzGMxQKBZsXV5EQr1TTckV0nt87uXO4yNp/7hGTrvdSyUEv8zXG6WV49eGhgkrLYOf9aKTGyGA
iiIzh0Jrtyh+Ns+tUkrRIu996rgBOnvml2cQA2xxqjJdBJBPhng5k/0WFtvda5AzfklAKooyy5tI
XzFTFrUGsApiCTQlU3JX2lpCmS7lu1uA2S31A4jpV1umL1UjAZgr8OdYI9KaqIi2FBBENx/STSrl
Hcn8dKRaI5wXr4MZ/ZMwyQvdawKrVlzcRPXlDdru3zAD/uiioSvVxOS2U33AeWQ/1iT40Olikwnz
Wu9VaIVD4EFglC6oQe5A4NjFJLGfYitoAH4vu0xtLM9O2j1AbqEjUZ8rUW+DYQwCuuXrfgDAYOM7
DnyJYq30CbVwulan2ABg0R/6XCHRU47sQUZDaEFSBjNb2oLvitt5pbd7zQS9L3lVxqVAFrGEJJbJ
SMmaruppAX6DozegRTWkbT1dZ3poqigQcSRNnygJMwYTQLjxQFHIEHdwmLfkVzksRzpEU/y7To7E
AzyzuV/xMqBs5CoDf3za08wYmpmHu6boY45fub3dIEkcgosCn49tJGuMi0gNBQlIUUpjcdZU7BsM
ezFZQ+bEPCz+G/JWfz65PsamMcpuPTWip1FWx8SnvnDfVIFDgMwS1w3jD8IHfVZg3MASF7O0opZt
v+Rqusse9zI31hBLBMsiOx7m433LyPzw/UXWQ3E6Xh7cfs8sjMfx6rn2w15y+OufQQ1BsT86YUIc
hbdfI8WJrRMgLXx7giAIo63s0mBUcyClnq7auZabqIZYNyriKkFZ7q+yMuVfZ2U8iFMS8UrtxLbF
KlCF41bPJkx5r+9x6CElDsvC0l+KBynFDz/26+uilHaJDrcPiQtefGlOR6LG6IOM5MqzYc5DVsWO
rFupoUOptMNp4WVSxKGag/hGWd8WRSyoJl9REoPG59Qh81Wq96ni+BVojNfKjZc53etGJ7GalIka
AyNStPqrdnTHrC01vCYzL5sV+D8HmS4ptd+s7EKf4K/Y3+n6fwxz9HnyaCsoDNGgrjrl1oLYMpC0
SRJKM93VAWwU4CrQrHBN7a5EyY+tleffO0RyeB1rpjnO9Fu3MBR1O5YyFJHPRZeRYzM9QRWmPPEP
+q0M7pgeWP/GRA2RGRuqCITw6QThPZDD21ML39nce3WLwq2quB6+yKSdjrTPDtoeZ6B1Lix5fQ6n
b5itBeFrcrSCntunGbJddb2Rswi1yjsOPxmCXHktcdoAXmkSde1HBBbdRPwokRi0ilJSbk4TPc1Q
JY95uR5dW0Db/BW+Mr5edhOutcIR9t2F9ot8WMn3WErjhMi0Cyq1SUB/015xrELkckyHvPD9q/Eu
5h74OC9HeWz5TGpw0MI6Qy0GsTuOzd28DWx2ipketCIvuqRq+SHIvbKDxGuKFeHjP+qmwWlAdQ6V
h61J7woDtLuRDFZmXMdYlGwhTTn95ntfBAdfAZiNHBG14fs1zx5mpp6GdTvcAYpckOcVGwVq0cA6
dCMm6W+AcRKpDOvl20NuLcuXsU4oEeLDI4bhEW0oTqFuNBqdAtKx0/aqqgNPtRPWs5C9Ske3Arff
QO87APJB6hn1qr3zn9/04E3DGL14hSPnaONe4vANrouvz+9XFskqbGIy/84ArokyU6rbhqOxpi+7
9aoQdgFYKzI8vVaY7Mf5HrRtN5DD/48SB2sxKKg9ypeNQ0LBI6ruGqS+YX3WPfxsIX7u+58XVVGJ
Yzx7dSrcCpjUAUmY7qODgoZHo00yU5r/U6lQ1VEkHk6JHZkVgl2Z9tf3UPLpDz9603MbnQqovEeD
jYf9Jv+aGS044wE9LQJFfZ4RUMaGbum8/9XryRibCeevaWn4jtvKl2lLdvPkW1Dz8CX/VXYxnYNe
gviAMX7F//aGbGxEr11Y4ZwQXiZzunbfsZ/A4wvyOPl5IdchjsTv3DJAaPnvkJlw5B9otKZUPMOx
KI9WZ2m0qGo5gegOBkFbOIn+iF2K+OrurhtbeOXtoHBnClnoomxVnu3jUGu6WLQZDxiJ7zQkyeZS
bFqqqwG9ICOZR58s+zowBIOOdb9D4lGj4Wdc16MsMXuOKDC1GPiTYRXOMHJQV92k8UFo+LsTX70u
ygN1FsfVQTa/l+7/PPSNHZ7NpR4YlgC/pd18q+Asery0tp5DytjX7izyXXzxxl4WuKURmm8EOiQw
hlJzbyT7GyVkEHQpu45LMBycdEGx40M10A3xc5xwbCyc1Rerqmac6DC8C1FLtLvgZDdMCGdSRYqJ
P6+rKnkFyQYf8ky1VJ7gSpxn/rzKSSujrk4F7B9PLqnkHYy+/QE2s9Nx34+VHHG2iiP3mzmP0xiZ
mcBZWjxkOzsDfCB2xBD6C2TtgOvqWHDraeP5wZOpFq6fu57z+klPGRaqaFPCBMTkg2y3peel9egn
Yv5gQRwEtyyhuDSqcn/ZF2KFpoHirqAYVv+9Pfgh26e1CGtSWBo8qGOy5Nwg/MTRJ+qbynELpt9l
64idD+tU21Ks++khZO6sU7FL3pFUXGFNEb2AuHU9LxbOPwdktC1vER2Aah5PesZjJaYCra352IiX
eXozJP7LfaXQJh1YsAQLIJDZKmj/HlGjWdYzTUHy2A8ygDJswmk2oE/alU81ABGX+QZCy0kW51IY
yQLYln06XwtQ9v2ZtSmHbwpC3j6YSzlZ7DhR/9oav72oHB1K9A30ebO2CWU7Pp636uf7/bP7L63V
8zWKYqNXmpomMjTRx1GiWpgEmJ3xf8gDTflncSWic1VOqmGzbJEQ5L+ARk8KLPbDulC4V/bfznbN
/JFtOu5XXchHJ3cYGqIXvUAV5OakoB7uUzP+ZVTwCi01Z0ndO7pbojOkm+PVLty0LDzzYCWBg2aN
GDVP4g6IJMshkb4dXaN1JZhEkg2O2PvrgrCbj603Jnew0OBcoENqAk6fnFGFGEZtEMmfp3zRJjh9
0/iDNp8IIEnHCK/gRaGwLr/3jktiPdNoly1C9O14GDU5hAIIFC2gWdoigTSBMHNutshn9/0svm8T
6SF5y1rIleeNF1Vvm/mABDz0AGJRIxvmyi0euDKZnBzkJaYUFmrWNkxzIZwHcAZ3J5A6znnrr5Ge
OEpGe8Mvb73WNRuRor9zQC4flMlW/k2vd7SyI+F0syUabKiZfHEk0QtrJVjEvC7zmbTi+8poBrEZ
LeoxZEii3MOLU77VVOhpUapgZFv+q1xBA/yYmGOofTyGvNy4bUv+nxzT7nUcaOmqOe33VvswqdLK
G1OE00rtBzrSk0wvu4xLuuOh8nWaYpd/tBXUcizu/rDOTeAJGy28hJtrP+5RRA3amQlPm5qA+AYp
MyQc3tXS30SgvsavqebtCSxZ3yWzy4TbgNjuFgFLq9aKkCY7Zz8FOOJPHx+cQ/cHPRHQC/v8CwTk
/EQ+YpOSciu5cG2rbHo8nfP31lCwCieCr/5pr5l/9ypqU+JaChGOXZHfY/dY9Sv21fDywIM/vpk2
ZRUNgdZtYg1ThGSOeyWOa4J7YpJBHwSP/6kO+2CS7R6t422BZK77EBp4nORp4YXYj7e8YKbq56qJ
39vguq3h3traBqWcim5FD9+3UqRogbCraoX+jTYYzBxbEO+oIfb8L1rdDCAzEgZcbZAUH7X+XwQO
Y6Vf6vGHi3pppQfR6h6xK1m27tJJ9yPdn3OpGZecf9kcKuenqUtVVb3pvlhqHKRtNdgepOLrdRlv
5pQxNVanCB99pmY9UaXpf9u0F7WGq051SQxxvLSUytLoKn3i/48lKq2S1blrhSDI4ngYV4LMzqBW
oRk58j+l2e1vSxK5giD80W058rSXoUW+vAhfVqUZDW0dShJNlf8aodpmXh32TpIJl7jbhVnkt/AM
t9jVkY+Vv/b1h2QYoZE3QqR8sjjSax5j6/WJKofGhbCE2qNxZxLbp3W5AMJGnpcGWzGUVQt9scgu
GexJ487Z/pvr+AwU7epxhGrbOVsJVLQhp9kgzCph0elQZSTLo+CVfYsnUsMKHa075BXvjGYQOzrs
OT4mdbe9EYMGo+0+GJx1HEYZfpCNjydfICmDUXrdE7Ah/4YI+798vJxd+AMQby0kgQxgvdk0IgOd
C3MY8GwHlmEYaPGaX7+erszcSZGzDRq9Cl/OHTkcYWPzZQO2whaOaABeOOXVSZq9DLGbq54TYIqw
Rxo48VFKYaFbDT+gFIOWrDPzyB+sRwH3EkqWo21cuVsrYrE1kBCm3IBM7x7hSYTis+TStFi5hR2D
oWHkZgeo5cBvzjtANFesN9lRiDi3tDdhMMt9X4mkFe6arKQkCAKzTHjrD9ovwcJvgh6/rrtIbEUO
z+dilx4kZjSWD3Hcbsx4g3OXtmQr/V5Bb2K1vzcWgP0VeefwR6oHmqWN+PjavPFpMISHvg3hoYAB
cHZNn88Q/DMqx8qLj7h8ovMQ0kiAaWhLLqTtBIEnt7kyjfgRfK53CIPug06owyHdnw4o+/IbKwdC
Do3bdd5JZCgXl06nxSoTxEvCaerY1FlsYqB1QDmmfpKskkBETrHSySVso9YM2V8mrG3LgXVH/wXC
9/p0H+cu3rVEstmER6mbd5uIerMAzC3+3J0u8R9HJsrtdeThpTem+jPtI9aRvTKDyNvUBOG1K0xQ
dhXZ+gl52nbpr6kNPLXnDDb1xOZYy+t9yEmRS5SolMOcgrlTUr4Shx0TUvOrBgyCjctYFHWPGZ6k
UjXt0UsGWFVUt5G/MDovf4E7We4hirUkABh1G4IY/qc+GRTS0ypwJ1FqGWK1pbdtJpW93Jw9qYxI
va0hlfROpPX0papDQLYFy0+LZn2F6zUeVKMxDxa4uEv8MYlRNnw53PRCcLL9lDBr0G0766IDynC2
dT3AwZkcTI5qwnTpftJxwiq8+L6HygpV3ZBb7K/quO10tCbA1/ds7ZTjYxwBnNKYXBw7jppcvfga
2QlmzPkgberZ1QaYr8zpxEIUqOx4yZsZxf8fWn9ObDVucOh9c6Ke+ABbEW0Wnpfw3zPjV6ENoygB
tSYokaDXT9EXSBmKrkMhj3N/IeDBC9m9LORAKq1/How+8DZFzy/jsPEpG5Ye1ulax99/+UAB6lQC
57uUZH7lV5ygqlWmjO8fh6mkDKit70QREH/pXSUNUWiq3X9iuVBFj+T80OdyNHZa4kE8JzpES9l1
isYG5Yv1pScTevEqbpB7kYpZ7kIv2a8mAI9UbD4SXyG8TU1oCJw6b0nNFoG5ZrzKC4G8Q6/YPUXW
mBX+eDarAX/owLsThFUM1EfwNv+1jQExNnxLzpI9mSur7FExrroFpmE1LV60w3zDYuZ2xGbxNCsN
usq/PJKsEM5rLuwrUpAOj9U+3xTuDXrAPgCJwdHOwArpLdLdpEFCukxPJCwsCLsLKMTDgibTeMv2
zoMkkXYM1yfPPHipzkOxE3TYnRXyC2oTQt+4VJIgZUvOCYQH+s3Hz56N8gOwgB1HM+hBVmTuslCV
LISXiNOZnjqUu3ibciQ6Y8PqqGgViuOP9pXy0nNXysNfU6qJi1cNUMwiz1U/01PumZhtItyVhzJe
pud0Nv6YQBFOPTYIDJn1Wk93IClGkpsPEQ8m5aEbbf2VEiXX/mmb445vvXtxMSd8rxJTs7fXmjMH
gZ2ZhiC4LGNyusw3vKc6dlWE+cMdQiFdm5xdbXqLYbw6Ojoeb86R/QD6QRGxMGBHsmH+HiSfVXaU
v5VVl9b/u4jLbv+TlHBIi6JKixIs7fDgFSFSTwh1MQX+8vmEZ1W2AzocvqXy2/40Rh/e5BIkzyNf
aqiQ1qqEn7TqydckL4/6+xafFJqGffJltJabEn/JyRIRyyqrpJmpAUi/dnxcNZAjjj3AkFCqGiTa
BkJg/FLUXBYTfVDGD4PSQMcGp5vnhd1SRvaPyF8pr0Fl/3TKfcVpgwRyy2yPUJLL7KEVmFGnTFeI
TxPblD/FXb4BhHCA9zpazqVjD+qteMfEUUxXgWobbBqQvgvdMKghyYjMPfoMGKcOVE9331RkW9KK
qNwb4Jq4U85jWZ51jJCrRfS+ccwwQZRPY0ZZmKzw6ZbsYvwzpWZxhiogk3ASpr9TlwOYPZaE+T2x
b5Jy7SN7shcZnZmzmtMNlJyJUo98e4HpXEnRaRPYp8TfiYLwA6spU3+KLvtFvtq6tuFJuNQZe2cw
ITVoQSfxumsmrQDH6Qne6q593Lo3qrrmVHJkXv/MM3XHxj9ndjhTWtj3tqP61D54SmWnbXj6DePf
RS86S1GS0cEBAmTx5TKqhMBXNAeBaeDaV7MWSezYhrejfAOiy6459mrAsK5Qm81XhF1sohLjzLdw
OY8Yxs0zDSqPiS/gJDexpUJMKY9510QVl3uaCvG2usQGz1Wla7PIWDXs0iNFcMfajkYjclmv3wK/
mDiQTJzmJOOFnaWU9B2JnSeMpau8riWm9ppmgrc95MH/ldTXOwc8kehaqbxqixTidK8JBz3tmwQS
pxOQgE0bTId5lcOsHtaPwvlmjIZexU4WNKByDel9DMzIStKW1OrMf/hrTwJKzjQ0sn0uQQ8gGTsO
alvddQfI7hIQm8RHPzXVvxn+jsNIVqFv8k5KEONlAsffSfQxEcL6EZPtXGG7gOAa/ExFf720pys0
NrKpyIYoiNVkUj6wMhJmm91YrsQs1r9c2mRoBzCIF6H+dUYR3PP4dGZPTzSKNFcIJvIABTg0wbSG
OJWjaA84nuLkCMA9q1Xjg8A0pRB8aqVIGSXy9ZthHeF8IWYBHWMki9Y+t1NsTNq12RFRf4o9iNMF
6GGSl2JG4wv3Y+BF62CEycF00HP/NDGS52YsRMjYgi9dJ8sFtOIY6W8H82YKR6sYTfxwsvhCVsiw
1pa8CiZYrrOBDcufUvFHsFFP5uhn0ab14jdAU0N5u0F6LQEODv6p0g1LIxwc3hdas8Q/hLf5yFAZ
Qn0JXENf9QH1X0CgOFvd2HsL85nikSdyKyNwvKBKjVM/fuzYYHKwuQS9SFrAi86roxMz3tki+Qni
7wwgzsClTMTAZfihFX5kUv3uZuM4epAf/PQUhCLh5vT/CfeY3QH19NCTtJLh61Q3cn2rO0hanWkQ
rCvoXF//66nBl+xJxKClF0+/O7Fnn6yAr4tAzA+kGm75o0uLvHTyBvXABNtV2cYNmVMv+u4KT/MD
xrTb07E1yaW7AowQto+l/3sCs5UzMl8pdZVrP71KKB2g1kJYNiCl37k59MyaXLQmkt3oVuOhaF6o
C29oxQT88jmL6L/ed2q+F3hADRWmNbAHMk6nIzvNPCWsvwUGCxJ1zfH7sH4dGNM6oVv19FMH8WGP
XaQfRhLyRU6i2rXf/toBeF+0ywmnt0kW2pugc3U6LSYd1HmCTDSdRe8sTIqdVpp1vG97FTTWdoFT
wMEILQbYP44P3R0zE8u4BYXI8qGnAuywGPgu8ODZqHKZxPT7K+c2t1lz/pxjYb/4TtFvFVuEFKCY
CSh5XluyaPSzd2ekHOOtm3Yt67ERLozACmBOV3u0fmQ6wagcIVM6aAoViHmSL/Amcrxd5c5q6rUC
UKBquaIUBwC4FKhmE5rb418fizhzTxbgJ2MaDOetaco/6pJ6MxhGfA6B1OE7q3IHrv3VzIa3YB2z
3ZVDvKTqvH0nZAf18vaYyCjACBTYRKoXwMr4aivs+vtBILdPgRgoVIH+c1DW2htfmmXxBOaQyeeu
s6Pq1PScuSLIbQ+IrnCwu/nyDdms6qnZcdI703IdipmhavF8N9HH/++cQUCAl23WsoM3/Mm8Sg/k
hbyc0Vb1yx0xXzAlpbP734tzdk51/JmXc5gxnf+JTJ5E31X/njk8mNWe+k26wkW8CuJuxLJtUs8m
Qln9SJYAdK/noIK1YSTxxyNg882t5Q7PHJ7/c9EMXNcVxvu5VL1dX6MyDoyRGJZazPjcSq+Ib3i1
y/tgXCt1Lu0qYaM1FUJVxJZtxdpikCwOY3QzlQ772ox5gEZMhO9BReAeG4Op4uiaVptVj338cFRA
7bwRM5YiVOrwxXufj2LHgMw5+DG/jMyB5tJYJoi9YbwGoCA8yhiuuoH2xr31DA4DUOkvke2gX/3L
0kD24PAONZ3tuu51Ar2Wbuy/ieh5E5cAP0zYBuCD6HD8pOrhZiu1SM4YlqqPHIoTmldh55c6tx3R
puKjq/ZvORmJEqJD8UBbeqnaOCRrX/IOVcwH2Rx2vvmSDyB4Z2dGubdtpu3CDMD9kxufQUm0YFpR
hWTIvMJUrTO7wtdaHn2NX4Eni/uAwXF5EaGKAsR4B9EBQrBWNqRxmukObAJmGzS5aWJ1WriHdaEN
aHV06P6O5TEmyoUY72U/j0DYyCT8iY5LAmDy8BfBAQjH8slxTKCY7pj3FpU+HZPjaAzAeZgHHKG+
NF77U1Ll6ufGZqIxTjfMF1P2V4xS8hLb7aGKadUCwALHtBSnL0+yYtzDaNx/0zM/Bt4ksXWyoi8V
vG/9HK/9xDnU2srD41PfTUdnYG4vZMATucHnwtQyFm8ip9E5kM9VOVF8fDTUZyDewRAJGPdYckeR
qDYBOFIkT4C2mSx0rO0dYsS320GmxSlSl9QGXfysXfjuOfHMyCaDsAVwFGXdj4TivzyT65aLicPg
smMBaSRFvBFok5e3sRCjA5xvf5b09pyQGJwqLLDgSCzwXhVoHGHjCh01RZNCAukUOMBmyBABuoPs
XdnELC//daaNKnDnexjqVyVyhyL/AMlSPeNPNQezTQhSiXy92TNj0rsac0QNe6cs8AEDPgZqcMHo
oRau51MsPI7OOZnAZ61NecoIgW1Ba4JBxHtQF9LedvQdBE76u5ti9k5Q3d2r7zK8Cl6eCwVXhjjd
wX3djrnEsYSmXq0X8mL842W4kBWLP5MnZHwwC7tlt6XnyEgdyLvSCbkEiR080RsV4/Gbrlqcq8r7
EBQdLzCVJ/pCeSml6MXcXK8iSKZLEb46xlepkFuJesEm3YjnZMN/OCQl26qK4DjU4JYIxYv96YmK
uPu+PcalW/NAktFG057a1EW8RPFXMMyak3rA6oArIZCi5wFAsWVoBjaIMjYvpyVU5PcDwdxAZS5r
sDY93YqTMWMIJN32HR6g/w0oWHkyTmGG/Arr2swWIv9ZlO1mEiNQjZp8+9FMzGVbD0l6HauXh9dm
RlU0yuLlEaOzio4RzoWWfpM8I21mggSGyHBPZqIGXWv9+9h4YgpnrhMJH3bFVHrLMumAA637N7IQ
QV2wtxze8MXQ6RFoz6kr6dwggUAwP12GbSOcv/aMLViueQKWbO4Zrt/aE3bD2vAILMy44bwAETVn
xCZ/hDChaLElMK712p3ZSEF0hj1ZCx8IUL7zxOUQEhJDfdS4DAzYdBOkelFv7wHbrQ6fzqTSIToX
1eNWhaFrGnxJLLmGsTWq3lcISnWt58lqD7FxsPKTdDOaJBeB/OZSB/S3parYW/Y39yzCg0ibC/1x
08ZWRLTS55s7CkVpMEkYzNbEgVAz9soLJi7wwyhpQ8X8fPvqMsuGGExhriprKDYkceXKCT7x/m6i
teYHVj+XxXMFbiKhjW3+R4vLj4S+j5TKEfkiNlIZYN1f1OEerzrKbIeqpOfyYYPdF4LfY2oEFsSW
JAJY3j+wVKBRGi/raK3vuhSNgIQst+rRi3LSC5rFUozEZPLwhObU68s0r/ZsmmaGTQWCDLYV1PUK
5xUgJ0YO6eHCQ8rzDx/LOxLHbKXp8JWQF3q2c51jiUZcUamsh5eFl7UA6Mgx1eFCJ8IgkudfURP8
zpKammWy9hCseXdu6Uyp4vSkzYjQJBwiTv/lQQvXAMr/VV/juQ9VzzfEy5ZNWORNcJ5phqylJKal
bGuvJAubXusVOrxq8yKAZe5+YUwkHB6gEB0KjTxSTmKEqBOpun/mgwxbLzFvSVgVXYHd5WvHwbzC
0oVQ8dLU1b0OKc2F2FwEpG9kuKLO99V8ENPAucFI5mnPlod+hwmZMnm1aan1A2y3DAu69/yZ0B0/
Zcw53KXQOJbZ4pIoKnDAXlYoFFED/zP1wZj9MkGZchARd/JQY40H0ry9kvGzqyylgCRVCT5cgYut
q49NrI3XMUrfKo+5P2hMMrkaj0CqaJP1VF+JkZQzMNggFBuQk76zeGaWKyN9YPZsah5byt25eThT
1QChtSItwFso2YeDdDiBuCywAw6usuYErz2IAB3MQDFHPqkZVuJcQo7WMHfkxwbtuh128LtraYY9
79BW92d7VUsdx6gAmGPvyAmAJLNyi2isP212LpHck2dwUwJuw+D6ReZrN9uJ2NBi2xJWhyh+uLbp
2YGGns7Ax0Daz9Y6TraflFBfGHD1iVIvt59z0l8eYyanryaWfcd4KdV4H7VHxj7NGPrHzCcfwrRP
qg38UD0hN8gLT8lSAmkV1ShA0UdFpEZtlnqA3xJtBOvPVR9/PM7OWfK2YsSsbRAgWSl+zxKOHqZj
lkvbx9jEnKKBjzXdpTuXKfQULqE3m5+8DkSlulrJAtklHe+NpESDMzoPT7bKiPSvR7hiwRi7UNJY
ZiTc6GtOMIDa1gXVovJb4L6F3nAg3fFQwhCM4manwKj3QRKdzVj583IC0Y5cYpMWNHAvuqv/261I
PDPyq/lhJ0EiyyKZ1pQ/IcsXlifPSdYXpe812/z05USz7snOB08Szi1t7dYVYjOLxOkfH84w7MOs
mbV9orJMalvqZXuH8U08JJKwJfq78jH2fskD7+Jk7H1M1r/7iGtPCI1cRNem+IzgT0nz/wSjz6JB
f1C5K4wUR6MCFvAXLC8tBIWo1RDZ4wOhVAvuZ8JTF00jbjExY/wVX5M/yKe6I/OrKrpjEZlZFkcD
ASri95ffzxip0L+Ap6ihLurRbzfsSWRqVDZxbtYOo6ATVz0cY6zfN+81Nn6FBEGDpOyufR+NLYho
ckAW/3W+pzaGwgFWiz13wFJrFO6GxJq4XvYtDIkJPBFzJdcSLaynsqCgVm8rZzdl+6rFxUq7OqbE
ZxMxD8bhJReSXItphxe8VAyV9EtioAm305P+UhUilNrqhd66342Cjeo0UuN5qZHf/+8J3UOVu8Cd
gDEcpClgaLhtseRaLqJR4AqNKKETi1oRGuUoyBswnuJkst/MqeRPl8tz2FjM55ykYOsaZGSFGOLc
sAFLLi8mwn40wvDRTIraLMuwfI+8lcehAJAercb4YuTUGWV7QQJVdZsuibf/LSuvPB9VPU6/2ied
PoDV8OLDTDSywTpqMnamPK73Pg8Jrc6/gwBeuwV7nk2wTaRnPuKDBAnt8NGxJCipwEfijOHv02ih
xIVkjkJhmc0FJGDUI9jiLclh3uedwBrgpTze+Zg8jR6qU+bGlp81dTyIqXnP+UIDna6292Bcalhn
Kkjqxyu/JCRHf27Oa6eIO6O5udZFGZtkaphRnkf2md6oQELcex3hIVCqNXya0LC1VkUtDhqSz9j1
hXYTqZ+eXqC6L+Ht+VOykXvshsYluGDd6q2v3uCHEgO3WnX0PH4ALPU3aVgCZjkvjh588WFNQI/Y
DRz/PNfa4hXN3sdjgQmg6l6WbGFfCq7+OeMj3R6+JZcaiEchQgOaCZq6c0Qa6FDDkPZPNZWJGHGg
v0LHwd43o0nv3iR6Cg8U+9LTwtkGMW+4OULBZaHhxiHsVHBNdOM3+tWdYnuysmstnCf1UPhYO4/s
/zNmhqvif1IxrwAHUprSEHWnXVrdr1+2n91QkkKvvUGDkVo6+r1iwPkCAp5U3q9GhWJOS2bly+/P
Botv64fIkPfj0Eoi+THVL7woXTz6FcG0GDQvWntV0zztMYDEzL+eyMuWWMXCc7drjsCK22bAK4yO
dbhzWXYkG42Ld7AwUUAGSioeDceK9G7ygYIe9UHWoYJzHgUjA7p4qfUps9Vi2Qha2upWNFpxpaV0
WcGYwznHtqJYPgKf1uFmSv4Gp3MXbuL+TEh7e573Q7JUDxYPYK2cJ6j+iPulBYUcqtUzwvRMztFl
1Psxg1Os5SJxIUpCFUUH0AxuUthw9dbBcQfqryfiUZ+OaIyng3188oe7moGmLitMSbPzkw6IYwzQ
DFmr2EKL6sobMBG9zPh2wtzhWyX6RyvSc+ro9LPJp6JMgbjXP6ubMCqrRrZ8wcKKygRV9eiqYKz9
RgPEyAOqJZF+qCZNmA6Is2RXAKxBSh1VSW3K3lBhjJB4xC2Tp4sFOiE/zU2d4bMZL7y732kTKAyY
EzBjMFpYRJjnUb/Pac9eQcrVQkHeLxmToojnfF0jzT5yFRpFb1a822znmtEYhffawsKKU6vDpW0z
YitdX0w1SgDPjTxUxH+8mof2RLK5TQCDXCWR6XwPphnl+HRKrpqRNvT8LEq01RHuthPb5bv27xRU
vk+Grx04DX4NjK7HNv8GIG/cf15m+1I+vNMXJx6ThLei9swR88X4w38U/mU3fN3wRBkyFTPSBk+4
HWkEdgfOL5t+SNLlWBAl3RqzP0WSMhzG6gTlQFKy7C/7Cjdcsk0iKq8DLzc2hh6g2hcqlDuUq/gL
RrX/Ba6LQOw2QcXH4Gh2Eu7K+Q6gBnQKGTuog8W7WAb+lFA5ceykVieAjl6Eb1QzunAwe+/nv6Wx
kYLNsY4cxd0FgmX8w9n5CZPJ3nbOLzUfTWyCkdunk7PUXa0uYymTssBTGx/c//95MAJWPNMu7Ky/
g2wd4lsPVmftX2So11u1sKhgNju/mDovTJ8Q6673nNFBKojFmmFW1mpis8NO2ab0KPt9TNoqBndZ
usopdI898XbhX6kUQ/JjuirtEAZX0sdD1lQ/MnsR4mYufTJIw8u9UeiYr90rIPOoUv3f0s9s3Qlq
XKGT/cf/z9uXdzorMgZDAwf8OigkqseIh7QDXnJWmiTTic3ieY/ZsfKsLWj8+nHqpsaUR5wREmwg
ryTRS5WiUWtkqcbkVm8U8ISKLti3blTNnHoVB0xpAwW8AqBH8sj+Wh/ganGfn2UWlGwomKN6wW8U
iEWBOBExW+NIuVsYLLQw/hSasts2iODFbBrEs1ya9iy4R4WHT60pjs/cPmQ58hB0nfDljxmjYEe0
6iZgNVy5WQsZh6QZklv7SbFNb9EqIYjfbstIm1NvZq3DBk82I39W79BeBQoMGbSqOyITLxT1atC9
NHsI4pFDoYD4WahcycauL4evQ+dIIOluFwWJUrEzUxi5hsEu6S32JQqvKI3mWFEBPM6mjnph5iOY
lFmnLp4dGjMyJC7DHSG/KT6sK+1Rk2bBerK05DKEMnLiNMelq1x5OPqa96DTLGJ7E70pel6MANNW
YHvvNfBvrcWHsQFrh/mjJT8WRyn0IWhwpct/tP65JHD3ELv3lupoOncY8H0sVveJyBVXtlHxFsHr
10HJmfvlA1aiLZ7KMttl5TyNa2mNz9nMlBsfVOigzBzvywrtXpi0yoN4BiuphOBfeCWhSpmbdSoJ
BVi5ggWVKuxI7Ze9Npj4VY86ORsaTQx9OXxQ+rQ7k7htIMUIXThPLIDAOGgjX1C0fzPqlJP0uNfr
q0abTd7FdKdy+ivniL54xo7ffToxXedubXSUR7uxjUSJYCXxgRikeBttpm7zMrNPBLSb8prsSGue
KQHkjJHCo0J56BWghHY9tAtRyDMSk2e0l1A3BPig5+J8jedaiREEN7calcqO3DkhfzSt7SvoRoFE
Q2CYHe3NLCByCNIzFFJqm3qzHDIpOk+r+4keesfbJQn5wpbyjJ0bM9PhmN+DB2VP/NQ/1vbgjIww
XOQmm/AlyBefbZI9kRgJa9mHLn4kREvLZ0TGSRkcl6mGP0HDP4QIW0C3vywHAUULuEqohgHMJqMd
dlpPR5TlYEGVu5dDk75xIkeFxvnH5t2+WCTnsq4biKYlFRc6sEzUUmoBC61ET0hsqrPfw/XlYh25
ZbnBNPjp2oo6nyKacF+No9BvTDIogCPu9/107MgglukH3ndArbepvDgRPsB5dNIIcwOTZ6X59L8m
8VJg2G4XRJgupH+wK/ZtVtqfnNy96l57aufN5iax/HrhOcu0kM/3m/UhxanP74AZZq82gRFwp79W
r5kvfZXt3DaLSa/FiwbMo26Zs9b2jBNL4x5c2IkAjb0j3ZUVpohDY3NRVvHJixSA2k9kuT/qiPoN
lt8FF9OGHDXrlhUROIUqeXPHuyPbpOZQQcEHPdFMNpfZOZN5rNPv4NvfF2B5Fxbu0U/TDYWBzuD2
tzt7UAX7BdlUrO+LHyPTS657zqi3lpJOgoC6CJ/0BoPSbAJyrkMbO9RFu8dzsUGINitoxCehlUvQ
FDFgoXLZudU9XAVfL27NSk0/8HClRmAHsrQZJ1Fu/+thU3BhB1y0qTpju3DkA26icGweU9UIcx3S
QpLaLiPo+pkVImx48ArDibuPdHrb+54vZ2HfUBUMeQuWYkCkhQtzRY8hf11WpmoSyOvhohGkDW+A
Q8oDAm/LZS7LXS1fS+yDfDmlEGdEXZFTzxUyZXsjtSkB7Bp/6tb6ySvasw8W7g9nsIXLFO1zaBB1
mP0v5XeY5cLdZL2Cs0lKTHcPKpG6izVw5LhQdnE5ivJItE3/61U7aZ+7eV82X3fP0T+LY32OoHrE
T+sQNNdmRunuk47pKHeHCvfhhZLjTzSipT8ELIxlII/3ho6aN/N2P4cALAYK7KSY2jQ6w1Osf6XN
5uk3pfIQMVzSv1nHAt/at0bq8pLoh+pFrjmqlmkPQWt/NdoUE8SvZBxchqJEQDwlx10KaPKX5SyC
aasVc5ukoYhTpItKxiZHajSO1qGRf3dDOMgrLSooEbiUMKzx7L1+tRx+MN1k+qaXrAR2cey4+oSq
NKIrF4D6XKpIHlVuF2ZNSIvEXfVOLFfMNisrdKqmidBgsakVUIf5AEr8AtBZeFAS8bjpiEhFvTju
AhOHdoZiT//i/6yQv6tpImzKBIzgqr424QfSKZZZrHDyW+y27CeyLeE//2eEODSVU+pQA5095i7Y
2/dAPjcUatiujRXocXaClYFfKZsf3BI+9It7grff0NPMCzrqZhsG2qt4pUy99FAyRJLosGX9sBLH
3uMVhdZyusBY5+0FXWOqrUCgqI9VzG8LETBoJpmrDaNXJ/vybv9aMLmMVaRUUsw9Ad63RjkxL5Wd
7Q28cJN0BQEy1h3sNRrlW3go0ubr1zUz3R/SibPeIVLt/jhY1Xeawh8qrLiqwYRNZm4GhOJ4DVye
L4CBsiNWDiAMnk8wspssGv3482TYd17JNOlHzBCymXfFwiWd/Y4YHmen0n3ZQGICSBKR4s2dxb0Y
zItbNJhgqBRrFO00wlrnHFZL6q6T7A2B+QYDZs8XcOF5HilCIS3zeJEuuA3rhMxMSxWN7WV/pt7x
v8LpT9nUGwAa7/6Ec0e4yPBniDEHZKGpo08MAyDZYu+A3nTZ+vr23gCit5Oxkz3kEsLNj+JAUolN
6S3mMIBvQIMtkNDEyiHsTC0o3kzCU/tCA0vmytYp2cMUl1D/KPZHdYsg1cY3x4B9JEkCpKqodSz8
7TvzdPGwMW/VtO2mC0N7/oe5oQ9DkIYNgiLr4f/A8X9aTasy0Wn804t0Yo8noLyHMrKE0RmJ3ka+
vdU6ay4uw2D4M5yssQpEIpMmxyiS1M6UPrRkpDyJHCZkg3W1ekZdzezSzfcx3zlP7iihJZ84lBdQ
KD+6t7XBwMiYrU4UVzhto6ENBS6nAyGDVbrKTDma3izfm+8ymlGWC0cie+IwGQ1K7BHZekWFklKt
nlEMf5B6yh8byKuDcIQX9Fx2JinkSxAoSQVI/tLbSoGK2Wjcyp1gRd7MttRXZwVgWFXcqyKlUMJC
O68tsysg9FlPoaTpjMlHyesEK8bfL9O+NDh+HWlFo5Lz114zI6g2ToinaKcHpWQ6GkP2FOhAYnAo
MaMgBj2hBe96HxT5EKijWgKpZm8GqXOYj5DvyOVEd73O+UnKKj296j52SA3wS7AvNmbN3Rhajess
nnRZeeAF/bnYErATGSpnsAod7DxuRwmzEXY6Ubc5GMkb/vPWJdhKwt+eMjbx/N16Io6x87YGAJRe
HMLNyNsqujy+Q+bQo2D7chsSv2TuDj6NHLfeKsNfi8t+j0SL+8AsOaXy16rMj9e1Js0E2MyuEdH1
lju5kjUZdMsF08XuASDB0rk7Px59vBp0bMxvx5g7vomgvmdPipKmvkucWUHX/E5tiNUCdWRPBxd6
Rrl+zbjVR08Wrxuv4obJeIAqhYGawwZ5J3hNDr8ItKLog4Baj/ZkMIKedTHj3DUSh3Ib4asnEgVL
l/DVWN0EcjbLM3GtyY9SYSJulHzYl5kiIdvrC5zFJ0h+9vju3stzPnvDjqAF3FiyDwriyP0Rngvh
dg/Gxv5BxesR4JSQ/xYAThLuAMxUJ/pEPMtHMYux/y5nbk9NPDDV2Yu1EXto8N3qEoo1uXOgU6xn
VyGstegDsTUDAO3U5BjGObjaI86nVWKyipheaVAnOa1nNTVaK5tc3UdNzqtuFCZUxyTumA7eR1ZM
lkit7xz5v4gsis96cZYmdLYB3Tva1XdFGxGa0x0kjGuF2PkEMZ2/NxciD93X/s5KxoNqgPgEqAdS
cfwNfooSq0kanBHHtl3XljOMzYOi2fM+lUDTh9HcFVjsfYHC90Eyw0gJhz7FgtpiL8AV44A5JuwA
b8EGH0iRHf7QzmaWJPgWdPc3rN0fbeAxN7wb9X9xWEySSVz0NxkSmqKQf47IhTxmB/le35tqQrY9
J8r3uj/ojFDWg+a1ZVSLHcizrzfYQOVZ5H+NPmxWuncROzOFtgMEZOyAHB2XH7IUcVVrofMTF8cU
8mSzuyRfibY1W3zthPC3czF5sDhwyudIPI/tOB8ygwftErQTh+reKl0vrGJNa99Yip6I8pW203EC
rIW0DDTN2GC7A/ueWyQcSgbgSdAJcVPoxalpOP3Ylw0X0Qk+9qhyVwlVxTi1TWMQd4x67dDG0V5u
C6NDu5NTqFpDOlBLo/3ewQ2ubQy0abt06iIPL0l4sV8zzEBrIDJY4mWdh5QqLIaCC+HMevTx9gxA
416CtUcJ24673W9ALmGb2d8DlJUF4lWW9QGYv0F4gVxuOgFMt0ZQk9aV7ndgiK5FJO+MbTs+3BC3
aKd+uTGXldHZ7+lqUAbbpLEr9ewiGM2jAmoEqrm5Riw+e2m+DqUbvxQnsrc4AUl0runEAHBSOBPH
u6sppZPxubFcTOnoopMX9Se4jgv7gSXLrv6l74hvl+lvzEpTScEEJmF4GdEWmRV5IACLCxKeqmKi
RlXMHKKL51ejaBkpuE/CMrXetooUr/TaTk8r72u2znK7AWp0TiZP0HbogrH/16Pr2y4eQvzEfjNQ
jiYI9EddxnnYR2cu3Y+aa6+/iv7HTrZQflGoBM0EpdTyqPcZjOAM9iTk8g5OXSr1MkbIjDZvXr+8
LDDDimBKFrSGSqakW0R2LA4ylUxdj2zSrQLN7PFTAaE6XF3XhxybeH1AaiHSvzkC1mrLnOZ+kp/L
OFg5VyoGpo3/BhCWPivWAOkuKGVHoR6OPuEorGsBpJQBnqUkJYbJVkSFXSUZFBT4kRD1Ra9NJ22F
KWeYF8AVzuT77qpOQMR3EDsQTpG9dSivq5/h5yJKyrZCKdiHT/KJQPP+gGW5GnBDFbH//IL+TgBl
x9gyqyY21MCs3/NbXfoYJKgLHZk0Owm8cKmTF6IkU+xb3QdzugsmDA5ysa+W1N0fMaDp3FXoWmOa
q3WoEsDL/HhfQsZQBOBy90fu1xCqrcH7cis56YDAIjeiwtxv6lbTL2RC4THgCtR7BIxHv/xy5O3F
OA0Hi0kMDf/oDAPFgW+vfXdkrfJVi1UFwoQUPM3OVINEjnBA3XxsJ5P8k8Db8x5hOHmEovc+x/gy
u2TTeD+xPn28nnrja1mOW1Eyir4bmqN+T0hQUYLDlHWPpPGCKIc/A0GK/+b/kzdUXu9qd1CDyX6Z
PM/XPns7jOxx6JuarU3HuhPpCMGshSJgTZQF79GtOpsJdQ0OT0rnPN+wUNKJtl679rJWL1FLOZmD
hNN9UjJ7GaL3WqHpyG1ZxrHRQaW+Y4XqhPviL4fG0vwX4tV0K8nISt15xTkaama95LHIvKE2CVGy
jJOsGAZMKcZ+n7zyjVDghkHHMKaE8UH4QgbR/5aTAP/vWoUQPVBiPeuVGUlurSX1rtkv4FpH5UTH
M3Ks/MWm45WT/AqNONHN77PVyBB0inwX33SKK7dxbeQajJ28VxJVzG5uFMPYumMQ3rlcnoYJ9HEq
L0XlaJVnuOg2ycd14Y9QVUCAEPBsYkDIycl7q6BAErLuuhrmXswA+TQeX3+DgC9jRb0yyIEd79wf
VX2/tDRqrqyB5fcC94uFc47se3zlmN3y0PGMLc4qRN0ilo70QIT8bK08eU0o0jkHtpiBJAmCNECd
QKHGWOIFG9rYwQJBgLrxKq7ISLeVsSLAgbuV0vP63etYR3DO5bJ6mds0lvZFveg22+TAvXmTVRs+
goLzGwZpelW5XKtHcRLft5Oz1/NtZo+Jy/yFm4T9xbXVOnCVTrJOZW+OXW/4EcCbFQm8j6L58vgR
pO1onflB+H3TYBXkXEtfdozu2H7dUupO3Ls+bphCpRVpJ24iX88h2PPNjmk+MVTYsizg09VUNF7j
vIgT8vVAkwsZtWLSlduU91Xb6ZEbLJXd5NEDI9YPMYrqUjKpIt/MsWPRtj1zvIsgZ3YygbF6H1xn
GHLIE7z/p035Tr5c+1LS7IPfXCqewCrg609WdUhSRDfEH4nINsj71SQIwbxVr7KVYan7K5tOwd/A
CNBKXEx+uioGPNDX8eBHHiqv1uKYGGkKIsAEsh7x8/EgwdbTLDFK2aQUa8cQkwuKPZEmbulB57fE
Np4YOF59x2qtjjJs6FDKlpVSQC9PjTWS2EzU3vrKdBfkRe/qZVFIkYxWtg66BNAE914vJUEqHDzI
rlmDRXPU6aIaDjR1tvKdyAT6O3WyopDXfMxPHmSSfeiZc+bA33i5iRP9m0NORkkCCFAhGiPOOBBj
pR+VosjUYELWkjvKMpqr2l+6APA1GS6SyplR7hB9y+rRtl1a6IpiZFWCnSJQ+e4YNKGcmLr/ybEZ
3kaZDLAGV+BjxoROEzQU4A7EF7NYgLpE9IeOWsvSs3QjvFwqd5z23iOekNnwHMSKt+JWkEotASid
SGIfJbid8dIO6OGNJz7UNNF2rbXG4LW87mma/HmqrU2Tz3zU99RJz4d1HrdOshFrqLuNKWoE32x7
Gp21c753EEw6uV023cvQjafRUuds0k7ORpY3xCFlw5zz8l2p2ngnngG4oQ2lOzA5HrlPytiu8MQs
ArrL+5pMD/qAJaseKCj9xLMviQ7HH4XOE9HZv9JxuUWnhYYyKJ286yOHig8P0wLqs1EweWp+gRd8
vzAX5p9q5yfYKtKxOvyA0pWWtsdAafIDc5p34lh0uCta6tUhp6AhrvXgGJITPuD44IKVaeijK+r+
1E1A4vNAzNRrRPrJH6eZ5de2hwSww4BH3cXpvTFox303ZuxtXMMSK+bh648D8mRaJMg59GBauPEu
eJn1u3+jGbBuS9Zmv9dzRZWpM/bYDvbfaUMjeJmJpm5ZGLOgzIZAMl+LqjOuDIP0r8wXzqpDLPN+
fhe7SHUe8VI/M3d8Qdf1ArwOj/reX49Qb/nf2SfrJV9Je01ox9xuTtla6ArwhCAGCF6fTTwo5pqs
ISfTog9sDXJwVhZJyqw8rbz07EmQ149OmXKoAJWoTxPQlFT03c2kQSPL4xZdFHNMm8G6jnBJ7Ufo
bNyWlNcJegWrE1hsTP/qt5gm1bz76Ed5XjvS7AHaUmw8zq7vXdHjrE0jdyhGtWhIy7PMGERY2tdA
R0qQfM4pjvIEkHS7ReTnvPOLdEotRyd+w630Myk+10PxHJIKLYfvtN/GbklM6BBjE0u3ner6jvpG
iP/KYZuL5P53K7jbDkakrj04bM3ET0Z4kMKQMjm0kqDCbBUssWM5mO9Q/cBzMdDvC/EZjPjKMYL+
X4QvkYTLG5iO6qbeRTHYlfLPEPaVKwNFTWzKquFvmn+sYC1axXNyU6tnfF0+bLeeQN+rK1ola9GX
NptGlRv/bgsp8BszmQ/KwG+9p/5KsJcA8lpLYo+wfUaTjnuLO7CT6K0M5ZHIJ1n6OJoD8YXV1n1M
fc7u0MbOiO6d6NUgfZ4RtgeEYAa73e1hATyHivSxIVYS4XiBXLvlI7rr3mfdV1Qnxism1dg3+oZO
pDVVxa1c1F90lp2ETsRfePTmNv7r2zh2Tk/qqV+PGEo0m1UWWky7kXCJHv7CzDgNbWP4YZw4Ilo0
JHUVxoIApP6ohVC8BaR7qs1qRTjC+zU+hTnO9RcYE6SlI9l+H/fMvx/IhVFKAttEPrhXxXKbwOTw
oC0LTS8TbcTpQwYKq5U7R4eiBxiXVeDn8qOh8gJN6Gy8CSuwyuE69TKTsUnYuvxsdtD5DptBpQV8
Eal72z/5itpHgY33VPjdn/RxZ7dtvNItec+6UYT8/PUlPKZwhLXKY0hGneZzxRbfRdaD0LCCS8Gu
yI0BCbP8imXjWmBwaogSJzg09nWvRWcMcyqFNVBcMQeGONJg645nN4/zjrYzWDdWAgAyxbx9dYMI
xlDHMkXjdanjCfUp//orKOS6hCUboAatcyzVrA6T7/0+2cWrD6acdaDMebVc5UAHuKXxgkqQ1y7C
4LIVA1Ol+u4mkoLO6ubzdAeGdcqC6CmuhwFz24hykaUIYpw9bDMFn4ViVpqL9NQCJR3HhBJkvZoT
KMF5yXkYBBWP3bdK9Xa138TlaLIeHM0l8lX0tI7pKYrRdb2WQ7i0t5axCFNnH3IyE5wxMEyPUMSB
1KZVdOHcr0u9JDfRkrj19bnLAU0SRwvPXT8n6EwbWS5C/pMo5kfc7i1ustpBBhnQgVwkISD0y87X
F4vjrX2vsODiuN2HfTMCzVK/JwDVQ4JGJeg2Pn8DvJU73oiKWx76TeXjixJUVZdFBhiRHGemir0l
gS8nTfU3vLoJ6ipH/lWWITQpBtAw2rDt3ZvG4zfEA8MvOi1X/iud360Q+0ezQ6YxEfNDOTKb4wJ2
RvE/eJT6eqh+GGNrRpLCFrVUTPsCfG+qc8FpMNo3y+HO6fYfLSKDXB1o3BEk34Y6XmZepDbiKtMZ
2MLhcn8PelizFuxZ4qZ8zQodCJpqt3co3nNM0Uqg4gr2I8GehvCbAL5mB4OrmZODr6zLabLM/2hW
TEm3eJZR7047hr33oc/YWCo07kli2iFqm8JzUceNqYaFcvMsh5XxudTkbluODzwepAJDAzH1NXKW
hhrVYJ4FK4m3spdYRC0o4P8TzlrA1wIPuuQR5J7jatFShfDnnjfUwMBof2UlxmcM6t/4gR6a+3ho
ai7LR8mB7p/e/gIJh/nTbk7FPeBH7uADerdVFNARXE04N9dyfCGmRpq4XDFRYNOdLR10Ommz5WNw
YByMulzF8wSAKvX2JIXSgNk6nI2keCp3lFnhpv26me7ZtQV+OdDx+F4x+fCaJECDKVycbZvj5WEc
Mq+dFeUwcDBvQaE4htNeqNy99qTJMbuTNT2i/TvWGD6dIzPuyONzcBc8h6onfwZcnA007uS0neTU
SMBP/b7oPEGY5iC5HBEca3dUckB3WtUoo7y9M+eZyVVjL7v5Az4a3EiwWAAGjQdfAnQy4PbQaQ17
ACiGV+Wd00j89ZQ9fPb0N/399H6md2Z9UIuTwb336iSVAeZFDmq6jlq7gyo8ma/ajyaZ3xXYVtvD
5Z9KJLxjVMTmTns5YTKT65qGeR0D6Yq01uvHrD0PHK8w5VccAipFg43qN9muevj5+OAcpLhxzOVt
kYe1uNXgIjZ//H7RexvceviVTbFxv35vvIqxuW7Fs2/k/YujfrMyxvlGWhfdPnMQ2ICxcQADD6fp
cLlaM/N7kKr6UAu+Lo6QJ/x6FAHFVAdUK0+KBFAu43TF/nX4UhmqAE5EFTSpd8+4sWOTfV7KtTg7
P1Fl5QjZe2Y8EHSysI1Pt1wOjuOvIlsrOqp0euG9lmYgS7W0UuTFZop6wjTF1eAMOXjA7ogSfeRA
z2VhljcMgeFkJPzt6mfVZfGYtueU7b7B1hCOzZa6zhhnAMlYuBLJjgZRF8S7wLcptAXiH1BR8c5O
6WZkOPPqCOqa2aOHAQsAOvpZFvJGRxVLVHcfe0xLjafnQji6Y+UQ1bq/MFfjRYk0xghUI8J9xwTp
HQn66GqezjqDbgFwaVsnjRkJwtgc8t/p1vY80SuI7pS2aF83ecpI5TKZhXgzGYtv5RdOkBbmy9/X
rEgvwMcfgGarK2FD0MqcrzOIuZJEvnXu0r3L5H5w5ccVX2+jo1eTOnbHAp1zSbenot2lxjaxJRsB
9o9mED5nrVTypyaj1VLuAmIHNTcvOCGGzG62y0zLZlMh+BkkZSb/X6gA7jR68xSJhdVkJOTTajrX
7+U6RpdmKe2L/DhDA8+iv5B272xRL0gOgCjtySGeC/Osuy8RDAp4p1tppujogdECWJvT/M/RaB07
YlnMMZSW+AsE0GUWXnk4tB72rxHqFP6+m3WMAjUqq1zck979TYB0MLlftRtLr5fxwe+BufFtlFRL
tVGQz+h+hM5N+SAjfMO7TWMslAE1jwuHTHmkqD44cabes7zdzlZhLQxLzUPzUD3G47vHR/FHd1VF
WsgDUixmGQy+eIpg0UfOMe82jrx2iPD/tYOJGheFkiyMinEcIS0o+WTjJtYk9A+GHg/xke3Hb1nR
kjSLNIF6iUfrJ/VjlVxQFBMBYqWYAHj1JZ6s7beH/Ymy5Pm+aKS3PKzl096dhG3YPDaiF9PWmtv9
09CzUh6Ur5H9IdnEcNWrUxZHVHfqX4ICkxQ5LQdMwLlZQy6+VvVIw1treze0xbwKEFOF/S55DyBe
8BAwjZIxGW8eGj9c2l2M20twMrsN5nETSvmHQQPwchRHtCpI4HoMkLPFSgetp2tDl49P9NkAvYGF
6OoXfyZzR0gZb95WekeQetpWzdKFf6XcD6KLr7OaWIftoBWgHad9fNuBmb7qqYiA0qyiFoisGltI
B681en12PGNZ+ePiu28dfFpwMlL/PVluHzQ4/Bk6Zb0AzGMTgBv73IUQpF7CG9LzvfJBCgMGNC6l
7B/cfwcTQYArgLNZKL8iX/xE1W3gj1qdBaF0UBeJCgbDmUtvEL+lFVu+gZ/lveo4hAr3I4Wv3mNB
Hc0nKaB+nXkx3Ai5B513H60fyL8PWA98p+92v7JMg5NJNf6kYHK0BM4hJ5QOUVclOP88vAccUSvB
NNV0TJ4qPbEvu2S8jkPmLP1+rnttHwrrNHT1Ivl48suhU/xtZwQluFwJXg+iZwMccp0HfZ2LwNPt
iF1GmWBbuKbgqyq5RWgvnLQfew7dt0SQltrSEK8SC7VF1dTCWfISaT2UAMjXfbrLv0gT+GwT8maP
DYej2hXrH6HePLrfyDk9KKWCvhDM1BravacGeKYdDHs2VcJhIEn1GW5WOrxPKI2KfepbWziBzeAV
tHQE3VIL8qY2/jVALJY+hCBwB9aEGpF6u6V8gWRPkacMmQR3cI5rCM2gvZ2LVSdtBkp7JZRq+h1Y
8f0E1c5BOGKqcqGEOcCaFdo3EJroPy73vGTScdkYUTBispv6xhUj9SdMXZx3JxkeOYBzkV/dLvV3
DQlPwu0/CRYzbqhnal7/nUZafvcWo50gvaSI7oTPlo3knUaD0RVwsa0/pJPaavqaAoZ7dDcK3pl4
JAZlxoLLUL/nfwYsQs1fRgUmqYRhFAGuGAsIzCPWj2pZKhjfBx9pamMHIntL99a5mlDBXmeDW6f5
hU/Z7ohuyLtEAM5czg+jf++pEEe0b9JgV7gAXCg7Shdulf0n+GDONzWcc6bNfkMfP5yin7bo4vYA
UQW4XNMqAzhPTQTtlCHesKlGYkglyC632gsiensyaZzk+4wvrjrDg0RaSTl/uKQCyADWWGzXYYHo
n2wh6KpNYZwcgFIXhm0Upwplc4Mrk4V5ZLN+NpBktcDCd6/aWrvo4EDGGaEU9sQuwn6TJz/7kcwW
9otapHHqThOiAejJ8ZxvYQFjT3OaL3oO+pKzE3UUD96Obhd3g2+XJcbm0F/xjRpRqpF0WV/y2o92
dMeXI5gIo+y3mAEce+H0TcLdLK2s1bI7x5MaWhFzqTc+CQvg2P8ZoND+A2RBpo6gckuL4kM+c1q4
lVkGcgmXyeYglr2ff6I9cF2VPbGRCdl29X5hN79tvz6PnDem/rwAtmKIdqWdn0Y9r6D2hmAMSOqe
Wx0W9Z/hzZ1muTWV/vHZaqkrFReOrr37R0BypzNzCwkae3ZdPQJxOPMcfIjQDg4WqXgPfRf6R1t7
74PyhYKtuyU+lE062MJX9RFkBm+e92rjW6BrIY/5Q3oob5zyvz2OP7S+wWQ82ZuKNxaxd5xPtIeH
YVzdsLKtXrSvOA5tiQXU+eHDihPf3R/wgV0viw4yFXCY+65SfpbWsP1OXtNLWEKVw6jIPd6DxcUM
1+tJ+CehnQ3LhEKxk03L4M9QtJhi08r0DnsDwum9fFcVepJZ+dCosZ62c3J5UWV0UjCyrJWHTrKu
5aWxdcfwdk2AiKMh2wQ7uH57nO3YetUJowkQOfcB9RcFo6UJf7DQm9NKeBnAbwqjq9/O+o7XN8it
nptbWq3ekdUsgF+unGVY9zw8sggERjZ6PUNRXDbNlXTEFR5ey0hOpzdl7xrKFUCMhqM2DOsrmCYa
iqkOCm5xjZPbwHJ739lbhMsg6IBjlVcD7qrsPC5H5kNgt2jKCAzNVkdxnoJ4gQb01gC05mfxF1L/
Kuft/ShIrYnEqEpeeFAVfDHEOki1G1WcJzymXvcIu+Wgl9j/jcxwQ2EPZ+l9Tpwq/PPPTlJTRaPT
rwErHv6JunuwBmubuuz3e7v5Ye+UVRxz+BKOo/nBjANUi3Wo1Nw/M+aH3OTTqzc4ZDD5/QruUyUD
uxluDw7vG40xWGmdQmBjgERb8SpH6H7spG69yYP3oVn9PcoXQdthLj1LbBza/ccU8qaiab/PaTCm
+yBfS1u4RtXwrhTF2pt4aZCCc7IRGk15lUBTrbNHTErCrsr3OaUU7rQiFJfnQ+gYejIo3heQ1+30
M1SHB/cQWLmMOTusKki2mA3dwrWrGORoUdcSYkPEZQZOL0uaQQt6RUQInkaWp66drNSUCAcXbWa8
gKIyjAaiD/qPPX4y7fFY8/9rsMoIa6pEAJDlJC/4h7+WbjBXaa21MZ/wEG3SdNt/HCZs2Qr6w8p5
HiZmnn9TNRXhl0aT7TK+rXvCyNvwjaIWn+TIt3tKJamuBu71Bg2lUPiesTuD9IODb/VLgFxb1AXg
zkkqtMrohu9e/ezbPkAO9Pj1WCq5jIrxLI5pMenPnSHLTV4w7V8oSuw1PwIwGXQOwAD2tDou3Pnt
DIeU7D3fbDz80BE/pkNG2fmSearCf71sGGlWr5QJPYyriM158vJPslF4TEdpqV3QsMPUWlJj8/ps
dVklJcLl99rlocE32tooZSshoW1vkfG6nPGZntUOZavnFbE/f/d4FNxMUjY0qCv8a549+5rtrD6Y
W81MnuYzXU7UY5VCoidXBBOnZAI0enIXdh9yGEXTGd72YWxLXkPjPE36oAlpw1wNDG5jwkn4wb43
A3sZSsW1Arm0j/Xymw9MPhZxi+3EcUr2zavf50AU8Ao/woxFouC4aQVhLBrqeXZFADVYvE06I7mX
RT+NEUPqukncuhgj9FxH2LUfoeJuKMVmVAQ5iGPQ1T8iSxtLIX66BYze/YaWQxGCr4z1YgNJ/F7P
JUDyMpUBmaFsgdnj86L7/BKQRXoBUMw/FI8sN+Okt89zZdNj9rM4JLyv9PypdbPwEBglFf0ru7z3
urJGEzSEdL2lJmZIWpQd7wi5RhTZMsZx62JAJsgnmmVcv3NCRnQKAR5XfTGAYRHOU9Nqhw1uPy+H
h+jNnKePgKFMdtQyt8vjhfxI0V69fmCfesTiUIdzuPCXSom495Kn5h4pdA3Ou1AMo33ATNY94kGU
FBpNdNC53qNZlAW5wFiYRHm6fWpHiEOhjVig2sdyma7Dv4g+dpOE8PjKWiTQCGJ2FdhI7AVBZyhs
bPmdJ7PjJ5n0dUyLWgk9gAbMAchGmnnye/zcopGBzXkNQKAEwkioNe/RmZjVoLGt6Jyjx88khzKj
Y85YxhyqjGAnOvGygTsF6MjtkJPCsli/OH9r4MQJP7t1DuuH4McsQpMvDn5gURKNVZvxczNEIZ4Z
syz9I3WCqSlCDX8NJl8KWdcWgzzAuSA61G8I1IxaLqrAD/6IzcDlPgFSKH/mLJ1t5uBFcjOISYRB
u3xt+JljUI3t7e0Zf9je4ZpT7Izcic83qIS7X8HJo8GcA3Xk2YhGYAipovI1aEeIijoPqFw4Futa
QO3qf25NkMQt+mN6YOpuY7eC0AU58WndegSZzx7g+bzOZXf7aHSgZ1N0yf9xwjCDEAwcCtM1bPEV
HPZHUC5amvRSgx03PLCxqvAjedxpAbEc3uyHVv+0/q0Aewx4EJH5XJt0/L8IRk/EffXIoDeuoz0M
O3tVu0yfXm8i27qSj+hJpqeLE7ve8I4akwpyFvy4Nh3DRiwkQFEEyjkptv/XW6XnVZc2b+ubgIEZ
kzxhKhur/26tJ+lL49uEt0VT3XIjtCcW3W0IuUDcGfF11vw3CcsuT5JclJWmCHJDU68yyAQrfuIb
vQYE8Ufnyw5TI3QT9UftsXfUoeylM+LJ199BPKErpLWkL+d2l2CbzaIaRznVL/ep9G82pOAkWMwm
aoPJ/J0LPdz/cDPyowUH+ghnU9nYIXEaw8R3nAreWewvhVzKvV4NMVdSEwHK3FK1buKwlaDOd15r
/6hd97iOJWmCaZ5sQNZsgu3d2/zcV6tgnfmYAbKPv2fnHSW4JUyqZgJTPArQOxWxKq1r9i/39bpa
9wQh6jF9W2WxkMvtBz4gcDIRwbAZQ8YLc9jBc6lmaMC6f45EHHp+ML3EPhWtQI15F6iewxKl8Hn5
Cp/iiUffwjV8eJhsPXNrqWIx9mGz0fHgQE7M33nIJRrpZfU+tZLbPSQbkECUdl83Ur37p6mV5Fjz
/rtFcfJyVf0FwLxFJcWVvYmV8oZdc0OUFIcDATcP8nyIJJh9MMCY3NhXwKZd2wsEuvAr0nNDTSwj
3WJ9XoOzJIztoYyOaOYjMEZYqUPhqSLhA4Nyi5gH2YkptOop0Dc0uGvAR2vxwtBK62sNkuqA2E4O
2Tm8pYDz4/tD39ZIfzyJXnuhSM9Gp41eXqjKz2UpiTjCBmYZgAaJGW8avvy53+Xb9bL2T7FSghiD
/e+XJAdAGSLbWBnuCfU8MQ6rkimsUotzSDZYSx6hSap/WAqaTHAP1Al5dhmPCjdCN5Df41/BS3AN
UnR2+AAnp9M7dZQnBTGWdozP+xIB9feNagG4c67pYmIljJFX5U68AzR5Hs5dS70skesftIeXI26b
amo3c1I3e4HwXcBOQFfUyTd9Wyt9JmGab1eRKUzZ6brrpEJ77dQHujwcyQKwVwksd8tmT9y1yla/
0vNszl7Ge/8vbXJNHTpgqzylKcoXEPJGB37AT5fMVZW9tVmVgzo31DsgT8zDro1zwVFDGZD/gvn9
ueea+To5oXrA+NQMK8gI4YZd+5TyUz/GI5vRmoexxEEvr01A8LKNTITzRnsQmJY0vghSXgBJydgH
cQeIBD02ZTKsUkAsRUh5SR1k0zpm5TmHvnWHcfifFKZ3tSRilzhdAww1YHAHHL2S6xFjpjVYHOHM
s4PDFlO/wqYZ8ETMhCQs+znBdwa0pH/fim7gQxuUAdYnDqrNcubaiNG4QpjqSlNn9jMg+G/J897v
HTj0mh/llVx8NyHwtSEQobwglJ9PoTaeDRlzNfUHy4b24zaAR5JymmquECAU0DiTmVT9NBwcTHQv
89RCoK9GH2Fw33yK73ThqhEPdeqgfLSjHlelsdXsxNMLEa/sd5bWoHsnUebmLqId/skyxOw6PhzV
3xOG4plsuXwPmSoA/b+j/rXzLSyD7kxbztvu+CUdKf4TnsyvlZd3XnXQoUtqE5IZ0pVJ6M7QB91r
Lvg9rg4yEw0hzBTkTKoTKTGaMQHnqR/j7D+VQQuoIEkLueyBmlswQdTyR1m6PEzo+oaB9rciXxb7
1QNcHGAvcb+W6dKIsDNCxVf4SJy3aatyB/WSU4eQrFoXutOoNSYP5VVlY9v6tmcXHRDRfyL8rTvv
yE1VV6Bgnz4htwPYgyEm6LuhFLOpolWGsFFzYgMm+8aiV4Zj29YY2aIPBeICJhquN5XC3AMyqCsm
CZFSlm1gknl7/3j0/K50XtdqaENxMDQqAkMmPpGXJ5AMI3OtFyap8thEhXsd5PYLokFLop26+wIp
SmIMeYVuK9c8LJkLl8s+XX8gtmKyAE/K37ODYK04EWsyVF5a7K0zYPb7kcCa3OfeizICXfT0u+vD
PX9IcWcH4NRaCXLIs578o3Ou9YxQbsz2n6w21k88iUtnnLj1Ue0zGXCTDRyOQYEiSbfdUEBmqnAA
o4VmDXdDJ0J3Wfn1W6xoLBb/7jxbT62NVR8vqsawHUHGev8lIFYQpqm0TZuAV3FAnYqcUNI6HG/3
n6YRyOTOIiVGnyei3BT6NMLXMy5WYdiPfs+GmIgl2GXQdMswyvPBvtbQXgzV4ycH5dONWa+AMD9K
ezEmGnsJxIVgCtT4t/Xj6VNQAezXJEtODi1mXv0l7GwwzguEacKPXJWUZmrKZPreAtB21aEwUgaq
5lesAYKDiNzkqe2uMcfoafVsFwWyLNJxASDkyQcvVV2c2cnMkSOlS90iorEZuaNkLF7U+zlAd+ee
SKcLtPRZUVL2UTPS5p9SIbJbuDxHsBdEdMo4DvBaiYaQ9D6mLsWfSv8wf7DhvP2MEK8CdQAxNTKy
F9lBU/OsTMAQu1YxuGDfS9eFGZymwi88I5RFSsPToDsvBO01xAmPkgd2+UOvG/K0/3znW2IAPs4C
6ZC/oSYQXfgSvFtV3pS1fIADt47pQ7G3xf/4rjOnG3qPCE9xKK6CyTIk4JEZ91eRCIEP01OA3fIC
baUHaq1D0HydnclZ+amVE88maWR2D0bYmx8TJqy1Ih+gvN4HFFjuy5PPj0+DUeeKOriavyvA25fM
26uhXdP3wQdc0WPuEhGzxdWlH+VqAmrOcp4NGiNkw5eM8O/XIoAQ62Xdkm9LqLvp1j9A0eQq0wSx
Etz9I2kndGOdVBnEgJrW+RMgY3ZyXt9afWQUtB09BryfBJXI1c/E948pcf6ZmjTeXocYer/B5icN
SbS6Csnk7afnQGFJAwz8zBAbWuC7yO99ziQv9O4kSJ1csVRw1ASZ89zLVtdFuf9pdIYWUElLBwfx
qOb5BWYBkC9/xROuzzSrri9vn8GAsmlRcfOiLWFge0aCjdJmyUzbR5KM02t2DCR661Ro3GyVSHAT
IihBjR8huxihnD0O7PO7lKYvsx6zcmXfxOfuIV7D8+FT8RIbZkEGmsKPPWgL+cD3Jpls9dGhTyf4
bOjha56uNsakt9apE/6kZJoF2xnILZ4RKbfR2ezNZ8a6c9KzygtvrZxo0OryazgEuVm32SZQQbRp
rrtOYfFK18aqPNjf6VDOp2t16i7UT33MxfSFV+PNBhWhGZhRYsfwpDket6cZwqMBTYU2LxCTSmSs
pNcuQ9uaR6zlc2XCKddR9pPXElQn6jjcQF9PtifbWuMWLFD5KHsxxW041hkKC4AKyUb1aLbC2atT
HBLkPTGheQw3ft+lyT0DwSXDzteLXM2rloyVDXYeWAmBk/KFTImJFRBX7XYnRXKio4qhrNbVg8/4
eCJIht5qOjKYbM4q8Hfy8CXh5fqlB73fiKdnPYzRjvVlz/mHMIeGkjSVxwuKUijndRCGMJWqycnt
XaFbMqT8NtMk3LgHH3F5Cmpti7OmXHjI6iltUrklaQk6QwYcdv3DbhWWzF39eAYdaLrNTitC6QwR
CzsCavh6Vv/Zeq1S00m0UHn2RejxE34o2Uk93zPA8Oh6pNWT2S+4JVCuSvB2QoN7T9PCr0DiKn3p
JkIPHW/ZGmjfsKw5LClNsMMnY7hnsSXQQe70DSl2Uq5axegWlEstunTdhDvUcwE+fQkW47v/pxKH
cZXupKvNNWQ/IHC2qG23PqfqK+dWtW9iF+5egHh2OoHm8+9aIPEacQT/0Dnu0zmHCm7WdtxxQv9J
yyykAyMPqS5P5f1CK/MQW1b+n5PT6DtNl3Fk+uakyvwLM4gHmxzZwio0DSxXW2zvjF3ZSmDJ6L8G
EON8AInHq4cp5gTFvzbUxo6OMaWCvc74J2ENotjEMpRzjnefKYfzDalZ6KmwEXZDsTeHTOrEHIiq
G6JQUpZ0Xz8WqUcvLd5t9AS+uzr3gk8rfEsKuMj9as7+JIVhijxWmQuOyX42TrnI7alL674A+cKk
pMjxLrZFDeYEbbRtoQY7ZlGabOd998qbKYRYLe0yiK6fI/QNSvnvVQAhS3/2ualHUoQ2b6iB98jj
BOkLL7KCeDoQtbRL0Wx4wuM0eaq5FbhZnk7ZgmBe+Qhvs4Npa38Kjlbw2bhUhO46d8CMFIsnl6Lu
ECCy6JsRO0j2fRnkF60ph1dc40f9M9yzlf1dxugW1Mw92pvw6xz6mbWj0YXiKI3q+c5kA5pf84+e
jSAr+ARNLL20XN4Bq4CMktigvQMU9xdKQ3aWcK1VxMfUkVP7sxLJlQdLxIqUaUBIbQfoCEdrMse1
MKduhCs1TLHv7IhV8/ooClfepjk95wAw+ur1ULCvAKdkUx/0bUe+tLt2inyurcOP8nEcjFAT8o6V
8+bU6A+32hfk9P/aJzOVGJx1eddrjRQ3/6TQaDnu+OJjc9Eq5OrHBe5hEyxY8leZm5G8weZp4Gon
68koiFwVsgxvjpYoC7U4vdsDYweP/4LEnEnnWyQMDow2fzJ+w9AWoPIa346E6gdcLDUaZbe7h9sO
kAO1Zox4+GBsD8/MspddIGI7PsYdct60y58vyGYfPr+/JtgGd4DpO080lF+4dQOlVus7TN0ld9LX
bfoE80B3g/Cx9N24jes1BFNArY55aVK952gYPdQJKiJWrss8xmFw6rTGjA//m2D7o2dYDHYsT1UJ
g+b3yOPaj1/YF1pJnZaw4v/D1e5v6qol5U/kJAeZ//G+igUHhLPFCQR81Vyed38mpDo+6x7ReGfK
kaZ8T5RRhQpfzsV3qX6ViGKwYdee3ZCMTNpOWYlw88OxaKpKHyPOPJUwS46TC6N3lb6RdwSTLwa7
1XDv2CpYEqZwM5VYzcFQqn7fgqKhFkkT0eYTVxt/Y4VoyT8WLjUctH3uqvOzdtcuhCAh82UuUj3i
RqN/TxUU62FRSEBcugyR7eIyFWMn/L/OtimRn3SGedaM99YlvR/uzyjVYQrIQKude3vcVDq5hTUW
TRli8hGm2AcIfnwz//gGZ66wiQzXgAEtSRhBlsDZ2j34i6xY3eiiOQ3j0L7FpQH03u5ud6mLhBLX
OL5WqXg1Bxr1pnDrvRQWqra3+AZ6S5sD1aE8klkfNFyj296FFgN6Z2iuGYxw1mmwHVa5auTJxW2/
1ah6skAMhgu3Z1qghPtDLttc3nf8ZmGtYNiuwvPN9Nde+GpSzPmLi3CuW61U+SrdICeigqGcoH7W
qKEicJ4y3UVly7YZEBc2kxuMpLjh6LRZ2UJ4JOlufSsbQuKkiaNGG2yW57ykI+wSlkfPF0ye5i/l
2JoZAk7oKp+t9AlsQMbJL6KDN1tFtAGPMbSisQkT9pv/vHKdDGFXfQWhCK4Xci6hFZuPN6ARoNfB
a/lwG+qZ3cKGZMmxHXjdlHaPpOfvJx6wqx7GNcVl4T5+M3w2CvjXLVHru9yrCu8LarE7bniEJ1t+
fucruRMN/ab+n9WB/lVtImt/b3AaO2mWUCag/cD0bR0lU8djsbZCgrL0wVHgRx+3JdNGfc/sxaMV
8BPLHyBNqFo+t3fTVIQFEftqzxBF3KTVA6WDi/Upu2kduKcfDK14LYOGN8VfzHY+ndp+sSnzQCWK
ud5aZMDdRlHmQXM4hVErumVUR6nPVLgXOu5uEpk7bogPc+smSN2o09XJnZLC7MjfTMHbX4TnXnVT
yaNmPZqXwjoKxEYFQyKcEgUzx5dB8DyME0VKxUJdPmippBrjv9nDw2nRZbUF87kLmNieVD0BIRMx
ajRwvFvxCstSn7K8fLQQ9cvqe7mE0Iec3e6Ol34Y1rKtiHechKRMprOENW5O9UMVDlxcNbo17oD8
Dee0TW5ZmQAOnU/soXi1XnIRU6nLy1kIf3EX83ryVVU0l8aCs86l3ymdxDlsFmfmqN+HTlMrvmZ0
e4v5WtmER++ThVKKI4eMWd4EGDe4WHct8Gb66inmHws4EHaThBx0XqTnRkYItRUq0PUKHDyh/MtN
sXdQjawXQG3SSguPh3pHn9nNeA2QHORweQjUwFbdoV/byFVKHLeE6vC4S6EgLp4GvYwtD7slEoZ+
XoF6hKTy7kqYuxaiwnYZW1ug3nXS893SdiEIxj1AOPGPpIh4lCX/I17rBv0H7fRUhpAoQ4RWcQXl
7YvUDVyTXFFz330XKKKpDyCuwkXthjXJymZx6gENa+jBRxy54yeMfm2uQqJtzQNJfPXpTxm7Scll
xraNJzSmLv77Ebf9esjSqn5mV72qg4GGd92HaT/N5a+9qq9vOarhLqSBBzFmT6vwrBlLJ6rW+KKT
nG1stoGEBCtuBEwjg6im5svcDseqaDGmxejuMgHUPxCZvv5Pz0Y4xEB1Bl5Lu5h0eeOlpn0D5fvf
GY4bpPRVV0cs3NMllhoYeDxVhg50y/h/B3ZiIdponM4PPxWZlELZ83kxHGB3ezH143SYJ+Nq3J9O
epaNBW+qJdQbgmGeL+vLiQSl+HZ6mCsVmk9i4xLN5yVAFwvy+wqznCH4L5kGGXylTRRGjTIHA2z2
5sg0weP5iqmvhr0IXdRnrCmrbVwkcGrleCisQ0TAm0WSL2JW4gui8hGUIlSEQQ7f4lW+dhxFCOQQ
YyN30gbjeAt40u/cwiYGy9aHut3gajlWfYbJrxMmDzGpU0L9q8gfy6biPLqS2BjBXERqW/1U41TI
z0q4rHQikTo6I/Eubtju/8Q7PTw2I1Fi2MyCbnyqxAyFjEWA+Dx+SopqBgsCrXDbJo77xIDXIY8q
jagg6t4sI2nU8v2ed6bNuRb1lV3LVS/aWvMpD9emoL5s1/usVbt+sWnEHi3elbwaHZxpLgbvouaz
scGqJ4mbyZMey8yhLSyJGreg9nVpT8fNj67DZqY2RF0YkXWFfMxSNBKHAd4GAPe3dSc/BpTbOREO
dxsh4/Rbg4FnMSBt8qtNo68UwNP23dsrYRI+OYVczepGPl4Qd7IixRUcEfWHttxOW3nvJkOkaSHp
5dvvIDK9PkjbU6w5CpXIlbS9SXkzlaKakgdB8bcpwxy0LS2bnIXMp1BeKao7h+UIC9luZcXg4dIY
efEhhcqUf+BfwOgyCm0quiii2N9KjHqE5eRrE5Oo1064dUKNW2kl2TRErokcXNxXRhF/8T7nxS8F
3iMJpzlMBwyDKoQXCnDyYgTwLaBN77gj+L+OfPkjBIgsI+talZu7JwVmwKxTt/4H9e9YC4Iomced
YegJ4z3VBplTjQLWkJ4Lx8aiZnXTGtaiOSqBrVSPctaX9Nu1zRbS6u/DC7vBjQNbHzaYJLSuqeL5
6LuX8ROesgCCz/7Jxi1bkUUTskhIpDJH2YzNVCknWhFMbZKIMQC0jM5Nal8+ccTt7htMZy25iN83
6PsKlALwOuXy4hB8ZSCIYmkw4dHmgMrA3B13KKbo5uKmwn2GKc14QMkER+Ybc+S51q/koyjkD6f8
NzP2GqLHYV9V9dYbVNThEAggtbj6sMcASU9THsG8nbJfnO+tDkVYwcT4Uwz9iKR8N84RrvZpegFs
yGmZFFiVZU6rqZ7PErjMUmhzGr4AqrFlOpbG+OAbjmdfeOH/Krl7YNxpJqpgRNUA+heP3vcAIMgc
263sj0ah+p5WFeeuc5XL9jez93cWlAmi+rjFMDpxYLnf+TW9HTvknqvA/mw/uWICwtoiJJRddRs5
IyHtiOCU8gdjyL3ATj+QtjOg2kRsHEEqVw0hmI9jblAvdp8bzIX6Am6rcHD+qVVgcF+ynDOPrETr
u9S4FIINzQ4OdKKW+8VeJGeh4cDNWFjmiG8DUywOeFPY66PmdUPYL2vHEPu3W91P/a3KcDjyh8vl
FbBKb6FpP0hFrj7Bf5DvwLbKgS+Xuao1F2dkVP9crhwsNQZY85Kz0akEMXLIldSNrx9tH7vqcbCH
bQZMasgXqL+/OYPpaw+HJtSRd3lxVBcUeMqa4WPadEhEMpeRGIjJSYoAwdbJyDu3rLiZBMgqvtat
4dzwGpapoGUc0NZylPBMR6SLi7KvrO9LkwymkslUCf3n6Cztmlakr5phLkWcz/qItORUSEaBJH+l
r5sdlGNAicCC3lLh+QBngAEHH0zUFz18lQi0xXn1CYGfef4ig2DtV9D8qeVN+IDlfQ8OC07+HcG8
MapjFh+xFS904dWMUcILrcrcaqsNCwtZWRLofKT6fS7afMhsVbQKeax3HLpZHHZr3L+fVBn+3ATa
AfctBWV1qtPrTnfjdXE0VStFr53vwAw1K9Prsxoj8W61UeWlKKugJZSnVHwoGeFkHsj/zDnYRv++
yjEkgUv+4qyk5I4TroMCr74Z1k/UNZYT8Hnj7PCmbYm2woD6JAxh3c7fDLsrXJArUeNRUITPtgjt
psl7gxVkqrsaGnMu9QZaXjjKLeBKX+87urXoUBrHwQRNcodW+LEAqDZdEFt6tdWEHoGVs3b0Anh6
qmECKxEA/Dt3OtF8+kSgyPIEte7t0TRsGXYXTNGNGVM2TxGOxC5PNok+Tr4MXblk4GQt+4PUQfSa
giM/a7qMcL2lvJl8iBbbrzbNu43IXGcjzfASg/Jui/o54/5fVroc60VwbWpe8YY8ZKhByTN5QfjD
kBExxZwX4OFZ3fNfhyhG2VOGxrhftNMsg1Kg7FDnYUYQ2WkVGQKw8Vn/Kj07aGDzE7kzxxMWXQT/
P/+B3UKHnuqu0cR4xNLAVpdYmddRYsCMWdGgjjC6ZYVhKjjPd/Hazn+pHT2ikt/Pe12ojTM123tX
sTLMcjTFP7LyQw+uhdVZjGYKiTxX/uXAF+X2SAaGoWlNryxEpgtFQ/6PxvBtnt759rfqDMho/KWn
XsWFLryyDOaHptORs7amWCLtbOtw1u9Kfv+Bj89awYkZcPX1UfojPtYUdDOooRgoA5Z/54CA5ktL
aVEv1kqwcgR0ysS3RVZ0Cs8h8zkKnRTCz2tzcjzPWK+IJXzDb7yQc5jBWrYhLgaZUVmIiEwuC/ib
8e2S78cRfnyXKG56O5w9vUoiXAdZ9evMnK03vA0tJLkxhXKg3WL5zHi66e+FdyKaqE4b5wr99NZq
l1fUNNluhe+0x9YlfMALQVJbHzg4WI8seImTr+fdBfZUxStqzsUJmbhLijxNHJXG4aBAhrsUxJ94
6zorU1x9rR30O/M+OCK31vqI+VSYfi85JzA96ZZaeS2B0d+bYnyZAIpkzRCiRlaHLShvP1RlmNY2
3I/sFgMuoHqDz7pICY0nxErqfmOVOEag9nZO8XpT6KvGV5TDMoGNF4unsD93xsWIeOENd5AgXV6L
gYa7JAV12Y45BqPa0FS9+8gFnjAXdK98fY2ZzMhQfDa8Vwm1LKeLI8qP+Yy8zp7Xh58LUB4rodo9
UBcGFh/B4C8r7kpY9bEFwvlQ2COHnwXJZhchpPy5CHvLfjmW0wgEHg9DPO1T3429AJaazrwNP+pk
xW4Z1ONL5WrRQylsk8p9TkeYTS0DsSqWMFny1V4oivRO/uCW9Jjzh3IVjYvxChrYLxVjdONiYXTg
156hcMNQer/wjlB1e/KowLoiLjoLaHvt9fQpeDDHQN7kv49cIJmG1zyqWUE7srIUpRmy1NnmiQw1
NZJaMlhN7OE3SHN0j1HjmH/4BReYL9JQf4yZkRRrg+nwgHI3ERMQFyx2UuKBK8ITieYUNm+c5SWf
uTxcsyCHL79QDuGXRqY8Bd1qLoXdAJH8e5cxMJSyUbgBDB0SvlD1NgCRFt0WL1j3BHp6e3NhBAos
+8leAUfahyvsTrq8/F2t14N4xkaoexeuMWrrIXN76oSyBf3ucXp+OnGURcaiMKJg59C45CyxgNPW
AH7sEU7X/nyVQljh4dk2saUsPhWdLnmqp//iZC3Wp2ZBtI4mQvrhJwEBxFKZ+itemMwVAbEA21ha
CyEreQagJnNoB/RKPFawCrYa/mo4Eg65UxKBdiSFm9A0y3UyIoXueAoXcmwEz+RA8bm6LKkwnnHx
WtT8AblXW9hLEqrIWGqazIVM9PbGNZPJUCiFBaM63bCL+6b7qum46cy/A4oC+gTQiNYnP4vr+yG8
OQUICjAc4fEqNcPuAe1P+z4uQbcUj26eVbmn58yn9rxHpjxEnXup+mlS2CNWIocP+U0h8oM0JGET
na+0cmMBhb0vKpvsrRX2pu3uD1ZTVyPGIX8CROLHMHhKH2ieeRhGD5/ZJNmaERepBrVxkWZ9QuI7
C1km2GCstsrriiFI1wGiVP/vhKCh5QzIoT4lsOc/ieRXzxG510LrysVVdgtw6DzsAJRCAIQ9tHAi
jyq/LSQ5lfgRiKUepZrbDU6InXoYkJ3eW20lsoOv73bCV327JykistEINDC8irkHkTbs7UhoQMy9
MYSGKOqspUZOBeRxks+O/eVrV/qVzUny/KmZahfpAxmJcB0XgvhbTnkVOwQsknJvM43Q+3inCQv3
4ECWeJnyqUadkiTI8lphQhDasZ5QO+9m6krFZLzMN61hob+8K4G0fsaqhY5YXYJxD/afeK2eP1CW
OG9M6vcz8H1pYKUPGMLT/iAcurkDdIt+UMbP1AFulbOmO1KkKQWfdM2e+fwGRhkQs2404efscqVy
RD8+Y3IO8jW7nyOfyBpUhqtyHRocyNG4V3mxWyrXTNVbjeJbFeiUst6KCl4Xc0Dv0xJlGJRAA4Cw
JKNUWoAx+d9asitPO9ZOiUQtkAxwLi7Vf1axyKbxYbbvta+z0xvvNLmSDYpem/IW8zke1XIt8FIf
vmAHvZwRlXv602sVDmxKeNO24EIaUPszPlcUYQENRQ2UgJRMzTkS9uQ+vwiTAepY5mtCTv/JI42X
z1G5F6UNY31wKVxLyxmIpjdSWtLSwJNbVGH+Xk93qBf/gACoGX+TaeMv0VEULu+d0gA3jRMvgj/v
p/Rh6dwhlhcyA0k2Cq2+xhojStFTv5d7uhlsxark7joMMNKZT+p++CjknF5W7BpFdeQiVFcaGoXN
vKAFTz8B8FP1NtvLpxQuI6VwiTj7defK6rhhyDRJYKRqZvtA6x/ie6gVdZm6IKU9aYNJtuAlUwen
WmAuO1AJFgCv8Duze+K3vS6hGo0481R6FMHf7BUzWlu7Fc24edoTdhn/P65XB0P0JW6xyQ18dHIC
hwg2at2sIf58qLFuZg5z/yUjejNVAZzA4SUQHiECgw1OMe5Z6XVTIFid7lzW835UorNoxEobug1V
3U4e110dk/W3q29SPv6vWBpu4Tg7MoxS2XJN+pFk50udIRFe1FjiOQwgbzmHlDWS3umEygCmyGHF
2s3PfKvv8KdocDa2o+Mp8e44fA/61zHcV4Y7TGcsMrwb/AGyRlDjUE9K0zEuxvHO50ywRGCwTWb5
9QHJS7QK0jkYWKMmMwWWG5DcQXV3vMXfirvD9gss/7RCq7/8EhQMzpOekkdu8lq8b5SneTwdkEvr
4tArJIFzKVkwvi6RxRNQgQxwSA57NYSo+7qt67DEvL68+m3rCUwwsOBNCW1vqpNBy1Wc6jaTFirr
FUdECZZ79FBr193f2dmOGJAKqa+HyYiHqCxCY9pWomxjPfQNYvQ7hfpj6QIdd1b/c3lqYKreymIy
WFOXQX700qsGeBL3MDpWcdd1T/fkbION27sfzNtF8SAN+1ABw8KoJvS2zDEa7aIq7goFAhyl+88a
u9932UX1rj3+pk+zAD+6fQGGpskgIiDcTsLwr7XIbmzgy781V3mZ4ywRygmhlSBS5VAey4lN1loH
qF06g0ZQFdJ2z85Ko0LIOsPzF+x4WZlghGR+ZqH/c92v4sHpTilKKPow5sF5ZI12jLSpEtWWuxe6
6R/QpIpWxuSAZ1Wes7JNe26u4DH3K26gnFKjK8FdxIr+Eap+xvC2IHWQTUa7lgQCuPNohZvtX+zp
L44C9YgYOAY9wegWt+WIEDQvVvteATpINudWEJD15z8wCU+aX/k2fFysHXtWjES90czm4WQ1TvJk
Jae7dUIsDwcmAboi2F8fZHG8ccl6t3E2cca1HU2nlLmXYBp2uy16k5spMJ/uAsC6qLv4CoJFiX0y
a2Km0OGorAcPBY2xDySHp1N+jDX5H3FfDLOkTU5FuIN/NyZW/kgQX6kBAJPjggH0MAkSXjdzNLvC
Q/naELGIMaQWGYoWOiDtD1TxgOW5TM/qJZeXbVwgqDQEfHvo0d1BHcKL7eTiE8IFpXJkd9g2s807
U5SEuo49uokB/mpTngeh3Fso1mwz7LkFTvXM51Urk/VNLJcYs1sO7y66Jgpt4oe5HpA4aR0XdYG/
328+M1RMOGs61P1iBFr/s+IMePsgUcK6ivCHiwEtls2clj2zcQ/2m+TWyD9urkIo6ugiymbmIyjg
rp1JAd0sSa8c9zxvOlR3HHwXiflj4WMVJ7lIJmcN0sFyX+4m7KteIhoEtaHLumPQ1rdHrXPX1Dlk
DLCoB7/ivVEpIxcJ2azFMyfuRp1RMEvdBezedPyl7DhVBjJ+qAO/BzhyAmYdAO/JJw902v95gjTB
WN88L+fy6xSZX2PSL0++IWeZna6iZIFRcb7liRLvoMiTz3T5mK08XRrECkQShF3CDcsTVH9L4r+U
8eksEJieNTd10jjzLHdYt/U05zfPcBKfgHmDySHl1lVDCpTtWWW/JwkCyGyDkf5Hj8eMY2aEXFtT
2ju0q7ArEZdHlwblm02uFUw1PXa9wobEOTFvvhjl+CxbYJOx2Wjh7jxR1PRvvSC0PgKPex7RvX60
33M8ofoRaXTtK3gw+tRUuXCuxJVLPzjhlwAn2kNN/DTHM76yBnWEzVB7UPf1ilvp0YPXcYohujV7
aqLOnBNV4WTS75EIUEn8o/FtqW9fHjVP/2ozpITfOGl8bcvkvwFmvZwlCJCmvtpe10N3lBH42j23
1gCsB/6VKTdgfLjBFr7m/cRv1jc3ffM8Fi3f2KWYXXFkrAASQev81/c0v14HSLFIINQmyzuVMDzh
sgCsWu+6PrYaTrZ31yfLYLcz7uBPD91CCsoTcLXjYhTcKLCtLcEfyqTWqvR7/TkJWBKT94L7xnHT
XDpHek+WLDCeCNfdBXZVCoBBQ28tom6ZGkOKCJ/JIJHaF49PI/N0KkILXndeaDrpqifK8i4Arjbh
M3JczornybkceHJUZWN41FuQ55BhwIsscbrmaK9/V4cTNRh95gbbpk8QxheWEa1XvWmlKwzrDanr
nOdIqGtyi0+yIFQFzNUQRij2ovFYXzYrH685jl50Bzam9XFEpNm06jjpVVbZP4VclP7AMILJcDbQ
E/i3L8bIQ2T5+pbs+WWC/3ZSu0s2B3I9MVkr6mRhDSuBlFSz4jWHcocXJ7abSDr6K8wMqAHbq/g4
Xyxeg0LOZxy78sn/XpPrNeGW7KYQHdcugtgcHYHs6KWX9ppxRpN5NhsJy7mdBqTsQfqBUpoWTAgJ
qYKqe2CsDeAL7KwmNpx0HSW0DQ67Mksx25SVasJVG337IsysfNOzBCOYOKjcZql+3wAKUNqpFe2g
SEsLM20chanOwGmGRiA6NbU9y5KkNNzGDQeftuXHl4cWqfPQENG6KE/WbwJoXDI6m0JEfKLVdFT0
oWh1bIuXmQkIyhtQZ81lG0eECYMKMT+K0EJDhy+qAwPdOtp+ifZ/DXhNYBQwiDFybCsSgRFPfPIJ
xiT/qtT1gwJymwqcVgapXxU5hHv+SIF1hc1yHeCLNye2LxnkmtTSevMVSxjfgt/16oxp1uo3NpgW
l/qescTiavL3Vk8Ax7QdTmgFG9W/LBwNJXBFo9fwucd7NdzU8/MnxIvqmCrxWjAMXDQcSZCrnbkR
d2sCQtnzH+9WSzOFOaSW9sjmrQaPw9btCE9OK+IXKQ/LDYQES3xFjfIZ0hLgKWsWbAUyayu1IPFm
QjZijcYwPS5yQi5kP5gBzkCu1goeifRBMLajh2sHZ7k6Q5iYhzZF1f9ElcaN5cTM1R28yEw6LHKK
Bgl+uuf+GtIOkRXDQFE7KSvTOR/LTeC8oVq0QayYRP8hlVVQ4lYRH87PXtSBJYMTgothPpxqrONs
jZp+KT7yYN1xFLSGKwICxogtBqQ8WRP5RRhXGX9blCyZkhlyJke2SvTPYUd1BazNJBKybe0OgIef
Z8a8TUJB1KVktxmIobYfCOJZYrQlbaMdOOtB4aqwri8ljMjxM5Nh9gec4uaT4a1ccjbQbhYWgUcT
PLUsrB6YHsnBWclG35gMVdLynHlJDZL6GZYjqTFAtpa+Op9iwdPeiuRfuH4tGp6KMOE9XAesPyBW
9jCW2wS0FkJMAakRUWoXqh5K2YDJa4A4tsqwbSpuGDHRqZvCltSCGiesu/+EDF+KZMCggWTMm7X/
AzOpkppAZKvwVjvaLYqKN3FhApH7kBtMfV1FKhd/J9Dh5v/gWh0hjy8sfScL2xdPL19vH7p8ugFd
ZsIdD0XO6/6nNIGArMErACpqrHbUFYog+l67A2STXIB/xzNcC3DJx/cTTC1lZ1WI/bdh4QtvnZdV
gx9HujZ7LgfsGnQ0WkGfF+FrF/J6mgOkfjpCntxrjgf4ZLpGBOE1UhG9Ysq7wINcZu1/sf8lyFyt
E/t1tXSsEICxML6JJy+5ypurlyoyJlA6ZWmEkcvXFAz8/V0PDbpyLfWEsDXETMx5EsvTR4epNS6V
5v7zPUsixnlsb8oZ6s8chLo7VVl9q73JIZoiU+h5yWFvf8GSiwOKvYymloXaQbDMQZAvHDkgG6ks
jShb4ajy9JYS2brkV6BJ4/RRN6lhwap5bu2hP50OZ14SrP2Z4aGumKfnBpR2+9V2S3B0wHV8j/+m
jCDOd8qc47XeG8k+UwU9kA+VxdRkq+/EYRhcCqblNfkrOPkE2GZvqBl2OARqCZlx+w87M/Rh1yoM
cZTWXmzIxdQNqqvqQlGfxLQOhNbMxKhBKUGzi7+VOlrOdYjJpX0NyBZ870KCDjwagCwgoxWOXdiz
cCBBsIY73v5a7M9+a+iOme3cA0ggPy5CCsahGS0wmKBXQ2chjwyXaH0sX+gfV+/yIOpyVyxYTITl
cxwk/nXvNKg9vEQiMFa3Nvb36i89DgslxP4KGKEIK5QqOnp53xy82b6KuhUIsY7NWMuJc5oTbQTN
ud0wpvkvANpcGIIkYRQbPpqmgqBoFftPHnMJmQNx0x22ziHONbHzdT5xKuza07hY/hyq5bQN8Wxx
uMcvzalGbcEVPEHqRcVYjCJ6cl8J231s5OfJHr3eWUDFOGMw7OTqJQumxkeZnUWji2Tktbi2Qe20
mulpY9lBIKt4vC/zZQUfZM7MsjL4e1XE6pLPBHfRjDlazZTBB2Fw1STY5DrrVd5muvT7eB6hZXsr
k+QfoYwoMrTGcAiuIIxhcZAzWNxf0MEm3A9dNnZw2DFa2QVnaqmiC0s5UEN6wogBjvKpMjilpkOh
twAha7JinqO+OWCF4cKKoJ5eaVELUi+rEaeFGoasTIiEtUlDxRWoT5z+osl3ZTcqZj2mXDxum7S0
yq1cgVVYo4hwoo+zBbsI3Qq4q8d8TLwPAkIU/CtTt+pvo6ZFlGNKl7ixcCL8KVNa24ywy59y3DcX
EH6dwoDIIPauMQqPZgxneZBWFpd2P4AKMHNbiVhAHuRn6Znk3IX7jwj5Gcng2SCsJ//0w021i/zJ
TYDyRmSuwRN3B2jhnq5LVyJnWht/VIufad+0Yyd05xWQwqhvp20hrJq5rymJfOikPttviJGLlN6J
2BUsRRfNGm3nr515IiHIyrCF8/9PxsN/Z38DlWHQaZR+bpu/FB/tKt/1eUr2FnxeSJKx3XU8MHdK
NHwbYtIbCJ0MKTh7W5eKK9ll85XNkxsUnMwaQAN0579SPQyEUPxouHz0YW/Adgjqu6wrUDAhUQfx
DVK5ULS9osVGYg3Q4iRd2vtbZ1VGNJcFBJ1YW9xPV3tOofgjd79yrr143HRI5kIWixC7b49io6jB
bgcnW160SZwaT3ly/M+KMCn4vWD0x0PzewoASk7QAga5QU6cdoa98aQn5nJ93rz9ATJQP1fM3Ql/
a32+Dss2WWHvCuD+o+X/DGf9c57HJZObRfqqg/nVCZhZ82Tblp4sEXAh8gxxDGnopqAtCKf8ZdHM
5sKJZN9EsD1FyhmcTX+M04GacAGrtGxrf6rM2S3JjHQ6kH6PtZ6b0rFyXUBDf3CNMFEzjzFizyNy
ua8XHTcEhBXoz+bZvADLE2yBqOgq0fBkzhGOkGhHolVM1UTZSrFmZEY+97rEdvWnKiXUH42AlogJ
gpko9h+e044Y2s/w3OJfhgYgthQt6Bm50aVh0rawlxFXKdVwcbNiBZdV3f9XLvo4f7ZsKlXl1K2g
mHUiVtzei5Tb9eBwQz/F5ubwV77PNxtV/2y86Vb2Z0/7DvhMahPwQWW+7tBF48ILHUrRjthiWFNl
y2DqTZ47VKWVpS98PfljXs9bimqDvFI1VvmB3ziqaKH/lKlTLQiNB1An/DVeCrrsos7QJR0/5W+B
BOImIi5poRarPIu+YHnCUiLEuWIPkMYI/RKp/S5J1Iye7co7QVumbnQ9rKvfZN1f133kue9n/1D3
vgCGSDEEI1ljApGe0dIBqK2pphuHtslTgSPfO5WN5XkYKnPEWn9XVOtu2ANzUR3LxAi6TLv3Dfqq
bfSe33Cv/AEZ+VePO168WQ39a3HVedlXXkY5hmV5nSy0lzqL3igYjNdar6FjqWtxGSPivZ/ZEZ0o
TZdRxp6pqMzF9hAFyq5z65Uv1bxKoPORiiVhnVucc16g7vZRKCbQ2g2LzEjmbQnu+5hGbggmpA+p
njuUmUbvPQm2MdVyBazk1lOB+x5PDb64lpX3zD3QgXsHSdKAm7gOM0Qndm65veVdzfjS+6zboX+D
GYLOlFXFNo7m1HHY2dW2XOcC7LZ/1kRsYqm63PiAAhastxk6Cnmpt7i1S3d0P2CkkIYYXQZhLnaq
Y+xOfwnLs230189e03GgmTA7guZ4F9PSNyfAbvMk22C0n2T+WGDNNjxumQbqDBucGt9evqdPSbmc
aBBUx7dqvDEmajCBFc/QAG2sYc9W6LaGMmpzzl9aL5WpkG1v5CBim16Z63ixA+XbdOZ2tp9RXkr4
skcZTcE18j8vfPlqTXw/Is+/WRYmGfeaDK/SMLFpu5e7qepAgd3VObuw++QmIdcfsfRiz3TJ3OiI
3jColRPT3JeooSqacuTS2cQtdI/GE0/gtKl0nv+r18I7/n14q2syz3dY57QAZslli8titD4ffgf/
8SC1E2Noj7rIiuglkl0KY0T3yT0nNwy8Q0iGFkL3hsfuAO8uH1+DxyfLYp08qQKhuWKFk2PxVPTE
OVibjg1nnfeh2Sn235ZhxPjiLsbjJyJTUc3KTb0jp34aA/1dHvXNeHBtV00DMaMarPGUkJdu7xYw
7L6qbkBFr1NM/pA1M2u6shdtJ3CA2ZQ+PLt31eRQnwFreHsaaXkTnMjlzZkHC5jGSKXlE7ghZiDf
0luUO9HzTTclmTAELjwu8QdVPLVWszLYuZKlZ2mqu1MT9TFdy0aJOzWmXqmv8C/r05jh2/EQdNUP
LZ5a26PSsaEmWRxuNKEL6hL2k1f5pklaYmx3407zVMk2v8586rCz7JAxzau/pUx6w7Bh3KcdtCSv
+7JzqqJWPEJGW7EQpaJ0aqL6K5ZJt6s4v1u0+Zctv7yaxtSRecxxR+gRQjhul/rUINx7Nsl6dIOY
c1pLDrMKJR6B/+iBqBEDTjjqBT5VG3K+/px2HepQ98n3xSnIUPqEi6rZVj1W5Z6Lh1yBvHXaX96B
RHbzdlvnmLw6lWn8RnpEjCqiDT3XONz61nVosMV9JBMf5Twn4BFqPKwkFcVlgXooaqh+V2RYBVzE
wvV2rAyefK3wPW7IYsMby7DWef6Wh7QLuWGOFCwvutJgp6IhSh+OB7Y4iixcwo9jy3FPH4bxnFOB
h6R9yMAY/UQjwMS/2VEfl9/7Os4tij2a2TyyROMknzFr0dzGsoMnGGyv2h6jFc+mAVxmAlEBvWt+
VvhywCHBJ8BFamaEW39B2+5grQiSitl4NX0rcqfVItSDWVaDslSKK0RbYuTLH72q52tcnc6coAyr
RGrHZEsiFX6ONKPzufe3KRHmDdxTSl6UC1687wvhcFaOEsEf1iHdGLXiylcXwv0k+qe2I2cCIIr5
qch3cEBMyNx+fbX2xdeMy+Mcp3QNnrV7K3PyTNVGR86qW/WqDJjKaInrsMGyNJeRlekde3mKLlns
4wRHZ4LOKA17Ppx++Y4OxTXsDd2UCgJBS+Y4msrRG2OA0bmyJfG+ka+VGy1izLJUWXC2PFJwShmg
gn/PKMKpBhM1TbBJqBgKtlVZYyBuuJijPgr4PXJcNBNPCXSGu6kFCa6uPPn0g80YABIqIbkdjsvL
d3ItVIBR4N/wzBXZrF2lklwYcFCwknzZBZST3eTnpCobUrzaIewPFTLqoYZblJLC0P8fKXztu8PM
3JE5CTxn9nPyviA2U5WbgCX5sO1Uip4cV0Sdi2MJE6uGGEQr/OtG8rPI1d9Ap3jPGxBS3umdYyjv
Y6xyeRWKXOldz4RcQqbDxZ1R4jwWBZPoTTlEU3Aor22LfwAzy2avYo+CYrXhnl2HD23McyzQ0N05
DFJW+rn2tpR0pCYwzKtVHYQuKfjJaXf4XZNCaP/jVjELEXdTvu2KwMjIoJBFB6Zq0GLRwp8PWnFI
udt8pxAoceUp3f6RxXxrdcR4PD9kcvuM72nK8yx7xBDrgMfc7eNKOPj+Bt+uwGJVPHY1HNikgYL6
c40tjDFZBi3i50vVp0MQXWQMXe3/ila0jOZZLWhEJ76YoDk3TorOkjxggwY3JdpOZyfSpzXivGzt
gRAOD15ANg8jzQC+HWc4rLkXjLuSpeXw4xh/TYw46ZiAEylqqOoHbH37KELB7z9PVkkPAqrMcNHE
9OnZXGp0H/ylrg2IpcXb9Wub1DIsqQH6BiOE28QW8g8w/3EfAmMN5K5HCo8fWjWep54hGynb5kCR
JwaC5f5tQRutpl2zWuJJP1vwgQnVgDdYWy06gRey400lZmLaYzIS2y3xEm84AMZKco3UrOKA9p2M
zuAE8FIKPfFf8goUER6mhy1GR2TaLYXXqtKhWCD1sw8RfbcYgRNySWPpLxzFHR8ORsS5RMkA0wbu
sj0vfmwP3G7+ChCsPTgdCBLBR5a7LRzc4OtGQCpR2I6u5XPwdgUnG4rY/WyMacjTSSgnbfYCfm6L
TgIsAeJTD8y8u54c0sA6wbBVuj7S+i7zbY3YhjHl85Jhyr1FTyEd1iD7lmmjVvJpVQ7HnnyyBNAj
R3fBb3NyZsAERr656SeS0E2SviaNMxmzdARhXPJGJuDfdjpRqsjG2WAOueO5uVJ3a4tcMkwFGrHN
/oCqxraz7JUhGFiXMywbKp+9VVJN3dlQD/KSdaxkpNB1Yhr3F+D+KNIQU/nxOgMAdQPUQEBTbrV3
/MbKC54mwsRfkZsMEmMBdwJp78Tp8/G+7g1IAhKDY512RR2l/jFXss0MW8duTSlgIcbt/36HxMpo
Fv55WOy2DLe/rg+ZJ4k8WNIPzWU6LPme68f1ETLIV/T5Y5AMeC+IM7ITT82QvuE3ursQDPFQBN8/
cnPTPTISMBDHmr6X9J8thuEeJFEj0BF27YmytrJty5ysTZcZNLX+Ww64b6SbHF0lCrG5htAehQiZ
w+Ht92GfPkPT5kX/2BpxCv9FB0fYllv5TqLdshxoAy9R7N7MJyVTpHeOqB3IXCgSDoF56i+0kr3o
ufiaaMuiGJLuxyDAYPD4W1FuBqbwDDdHhTUg604MdWmC1jAlccOKLYoKyRJCtnuqs67nAon2th0l
v4EuqA/vYP7i7pL6bBhAeyNPoH1XlYfwoi6bup2aCL6Oa+XQs4rgEFHp8PzHiyxX4iyvtzzvPpyp
8U8ZuxfovJ1hsRhuPMIr1apyrLMyFhpDp2qU8u0esYAMSCpRAMT3QY2qoM8yWk9OJJrCRsVuA4ev
RHJJdmBcnbYZ2c9Ia7MZcDuPvUsmVC4QOdKfhVdrL9kv9HwvsnhUP4JM/YD8ueKmQadnA2GqATcM
yMO23dsFSY//kc9D2x6GsTJNsCNkT5fAMFCrIeKFoqSyM50w7bqjev5HmiMyPCEfyaWgXVxAy4Vm
6loOvEofdpvF5O8at2DbT/OzyerbaP20k598rxv7aEwpUWnEhQiz6zk8zTnvI0Aqo/Rtnq7PSGM1
zN7bSIv7w32XsuFhOZJ/PNyRtC1x3d8zMnrFp6v5zTZ5D3ECZ3NqL+acWnFASAK+pAMV1xXi+oMk
0FhqeqdfGJYZncmYRi3/9wMzIwh8z4OGoLk+xxiVvD4ymcWA3DuZscM0IpBomEWuA0NV8IOaYc+q
u7Hfw8KXhD0nSmPLEWqRil+iz6YQinJOSNijwgPZz6j7N9nQMV2ZN7ASrM31MBsMSxwyn8pOevPe
uThLIVyBx1mYcZHZWxS79RNJr/bLA4MGEOzsWZMarht5V5lj4KsC7VhVrDDSKybIT8AVQc2lpHZU
OfJOxD/CNv6rUr7Y06zSR3WcO+3G4FUsqL51sLEHBSwFWjsONqLjsSUyYe6fGu3dOSYfR7MNGp0j
3zDzaDBUb5WlhqFdo/lItDHRhbzVRKKiOuOGPp1qTY09diEAJKLuzs4M9R6/59rhAUpODqEhN5FZ
FCHXkWAeaYRHjwBknxXY/IotdUE19Jt4dd1TBByUMv3M3Vpo8IFe0QuLvViFDYTON7Rgwu4vJ/xr
WlYFHugYmPkpdv1oAC9+6qJCTIdTw6foLaigCeAkLBEjr+7nCyb03x1QDMr76GNBe6TLfmBMWIVG
iTL9XOhoKq6dE9lbLjLl7kCKv/K2E0YXMGl+7iJmfT4EOLDOG+yfYDf3fvqGIwlxlHrI1uc9lO/e
bAy5skLSw6jHaaCBqIHyV7FmR0y7MxVI60D30LjmfxE7PWc4xGj2dmPhyjfl4df/e5AoIMw1cGDy
p5C+20J6uw9FtFC5CjYw5uZoqgacRzdUMRw/OJnRRS/FDr4Ty+lpiN94uyR1cR8OnxKNXGyRa1M/
HegbJy15dvo+0SRa52sB9n79BbAGD88xainn9yu0eUxpIIYEfl8bLa16Xgvmplluc1Emk9m0Zt0O
eWRWMUDwGVrCL8OZt4nPBIfR0owdrayz0KqZyUhWaL0m7uE211t0/3hUgMQlvRastBGJ4udpyu9X
JN4n7SJFItJP3jm3ILvsZQDN7UWRdE0+HmFR2XNHveT97iGwmqY0Kh7nRPBaSdaBZBUmbtp5LHVI
PWfeuTmTMcwVy/LYrjldlIqplmZWuI3iqDGpELj+alZHY5MukHaGtZjdghlX5A0AI5dZD8+g7eZp
R0uqRaeJJpArmSXPXV9ocX2jC1d8fiRTcTvu8RnEhUJcM5NytT31GlW2ylsCIKDNvtX4eYZL9Fkg
Bg7Tc8mHRhWHK664ATumb+e7hxBESv3Og7h+fxbEwDMYEPr+bk2mnSpoV6bWpR7645bm6dvnciMw
gVUCA5gvC0qmsnH/WlZ7F9bELwkNrizosGON+PosUbFQlD2q8HAgOFHyaBECxypPYPwiF5H98hdE
5t30KUTXLS8258pTd5KEJ8qL5FqKVKKGCCAputiPED+R+u11pnz9Yc7yuCLtZgDJhzL85PibdVQ6
FlN6se0FJ9dw5Nhc7c3BCk3XN3+lXz46BI988lxUuHdZJ0hKlDkfgWHLRi2E8m2W4U8WNAHgPB8d
mpHi5suswfDJ1HoqqxEbsMwleD6zJkoTpeAqWaPcGr9jewf8s6brjtOluptXAGpIir6sbV73sdTi
22/mQYF8IzkHzCSBkTAVGFbxrRs9bnpHb4r/CbXEdNfOurnhWuqrWb3VFZ5RZ0/Pts/9TaVozRIu
8+A7HOKxXHGJ3NT8YfspVJk8Lpf1rAyvhdQOYR5D9nlIRnu1gTFid3n/X1C57YiguFkeRNP0zBZj
116BnrGv1zH5DoJl0NgWKLsa/8kxGedhdwNVPBAbAo+Hkw+Q3rvFptuh0tMEB6iIZB2J7zG1ckZk
oCqABo5NWfnQQ7yAjYUtEfatGCqD6lWL54LTZAjWq1weDbYJWsbM857xrFwvzEadNgYj20Vv0L2H
XIq7fXqjBJqrPYz5ty0xJwfVKDmBjkSVY9EiNEHafJR22cDmFOrlzol9rKgVStH5q9D6YjlpzDYA
+AVvmS7yqbFeJcaTZRG/roi8XjUH2O7NSilmyx2Hxw7cfvOAN3kbqFczuFVKaXDs6LZqm0xXrXrP
KXSuZSC7w5opxbQEQeD53bMrIlP+Pvgew/6Oqa3tQFso7GoC7YfwZdKqtKFLNaFFCLSbBDmLBXLg
Lsupr7gdrZ0LfXdNFfe3LXKtusESeOivbsn7ciy0V+sy5Tmno7BhA/x91uKGJ3iAM10hsOWaHfGS
K5olz9vcMHo0lXtwKkUwWhQGXx0pPa3/yJgYpbyjhaUfvycHFnqdjcJuUr2xvC0F/C97HEub66Wu
laboA3ArMi3xuvARfEFbzEbV4vzN9z0v9BP2RJSaNOzmQGgQJXUbuPn4JhhSYy1PTfC/vW0mnBPW
Zm8+odinwLQVDPavbDebnDhnETOFmdHpslCfM4psO86WOvabNpsN1D+z1++hfL6z409mTQxuOdGu
l7pgvL2JPImvQguWk0XO472AXvtb6X2ocTqxMAMeEiwOuB+2ebA2zi5DUN9a9RCxkmCQshU0GIrf
h6OWHStgDtj1uY7hBSEOoBmIl08vWzkNFwSA+1KuM2jD6UMOtpqXVdKYd4Je4o2gsR4vSvGlhC9W
+RpDrAB1fTw9fhieioT6lO0P20ggEXBpFviuOETjtWnxbjn6eHkJsAOO+l86PiyJKNFOJZAZtcbM
fP5paS1mc8HHVDYJ4QieSuZxRJjK/EaWpBwAEQGn0jJfoLY480mpHCn5Is/1FhGg6F2IeTD4muUF
5bBXT1ITqBS7C7ng3eyT3SVwGyZYQMAQv4lCsz9WnTwGGMezbrFYThGC5VwwGjQ6wUuNjDn7PqV7
EkCTUaBzIs++hn7hs20ixaMG0WJwg6dnKyeyOiF3DOoP008yuB4a96ULGheIVt0RVbrlekfq48Sv
wP3e+4lpR+skRt28aitRdGKLP5O6OovZ9Xng9JN1OlqqhqTWljAqQhhxfIEmXb4vVBnbCifOTmqd
8FVl5WfpwW+vjJ1dGTWf1k73f3+cLu++z5v15opHezr4URTAUMVUshuDYL99EAsD0d/XhBcB4XKH
rawhsabfysj1BKb/Byy8m0aEZEYWlrOfTLzujW6VizrePH2OfteidDkpp9oMx0U8sAv3erzZaEAx
3HjNGYKzeaRMIsyahb0y2T1AgGnu+V3F+3/7fRU64mdIXDdj2jlxNqvB5oGjBUCC0bUpFhO/QtR3
Ag0sk1Sk0+UvocLnlixgm04iuWIee/+ySYgOvdZm/LuNb91VJgEQ+CDQ78HgHZfnmAtOzko9ZgPA
zu5js4UgfhsiM4b0fZhwPQLbFeY4PVqSVTv2esckovFTaIemISYx6ZdYHp3PXRmOF0ISzaNUzJuT
L9iSJT49Js52/PJev1pS68DOiwbSL16nmOw3HhWNVFuhkEX8XTbrCHrsZcT+RIqTNsdDHeSeZRPh
nJM9SohH3AbFNw+dhzavKazqGmadOfbe5xQ9tY2GMNiL9SaIxZflg2UCsuPSMcJrH8TRXkhMYr94
NVklzbXS3eFpnfj4kR9ahol9m0OxmJgd3SZNMDd7BChGwY6xgoailRG6R56CZp5FV3NePGVSEmtq
2bCfXrD0+vBeaZesIo8oDvlGh92JJGvnnS9WjK16AV304FQMumzHFUD18QscIPi9D4ZYDgs5maeB
TsnfgjpfhmzC9UO4kEm7cHdPqwBz4kmTS6EhWOGIATS2JoiSdcZvAzS62AqFpu3s/vm863y6q3Pn
5ZDQG7S4Twl92zML6lMAbVL/3fl7H03hi11tw8Tl6j0qqEbWl/sP6447ayXk4gcwzwWEmgY9urFJ
5GuxIuHYYeSjJA4laCwaAshDsjjbL63zuk3xADEtJVTExn4GN3jtODNPct7kQvSgSW/lezlSU14U
ozxONRh1Olwlt/EWUjWa1hvNkMeVZfkNT5O25foKsWFevJHXLc07gM4CXYF+I42XixDaISKa5itT
yxDROEKSJTp74SviU8Mumy9rHh1JeDplolRLgi3YaCiVJEOL6hEZmW5BKP+yuXZPvjHscuDr2dcD
wX8m9BZraizahw92ycOqoGVi2f8Wyi0VtBWS73MvUQUnRPj9/nHVBLjhc2SOUYQc5cbfAskSIyv/
ZHmLe8Mcj8ssiplmxE3SsQkZbWA3uYbBOnvqAnuPv/nravxsEZZMUBpwYTcGGBVunkQ7BUuiXT+3
Ux/6NTGci9CHVsOwENXUPjbs1SjmaEaZjq6+H7/HzjlGVSbgpPPERJJ+2yGLIsIY0hSJQU0vRoNs
4JZ5RYmCHR+BJoCzQBomGFNfAaEg49k/65ugm8m8yOExiWP3Geky18/PI/PiM73Huma3KJxVGRTe
XETgrmlRg6sgNh4k55X63ArkrwG1cU5JHxww2a1g1eAVbB+KjjxIUwugePKbFytdPVpGrRIUCbHE
Hz6/dPY9OjEWDFoG9nlwNNZ8hTBeGDo9YYH+iXAKtDznqJ2ng4HlIIzgu5jzDRFRk2hgQdejuurJ
CiOG5xAx3Xv+9/da04B3vudu9B/40WtrZ+Mw9TIJvCITJ2fu3gU9PUJv1QTjouQMh6qVXJhPqQ27
vjF/G3ebp0mEr8DcdAe2TB6W3uLr1eNSBPm7Q4j0LgwJXwRVMj+m7d4YMorv9qewpcs51pXY3hkk
B27visAI4ygnaFxnGQbBWfeFfOJV1pLIXvUi678l2DH00pKnYrkwsCHxZGxmAGTh8plw6p1x9IFn
J5sVi5hA4d4hZnbIKWVzu6xv7DOQUUKujIrpW5oBXUjI6sXnYrIRz1V3XviCeqFYXh+fiLscuISX
7UgqIvxnJI71Tksd4a4qUyf1yhgaNTtsmRoZWonZKXI79HZKKAaQCLXc5ZT98vYoMlUEAm8U4o4O
eOuYY6RrWX7osFRl1siN55//ukmVTRFW0XCXJ0V+envGCeZ2fGSpWaAGlQkckosTTB6fOXgJJbHR
Ird2y5OzGwiPDkx2eeJhASPr+K7QxD8KQIZVuIbhVCN7uJSJix8SINJPssDciG8VJg1lpL2YzP9Y
cwymYrf46axR/Uk2dsQp/pmxQ3b7wle6NmtXrbBwb7F21Kq+XSlQ+WkF7RHzyHfpDc6wbZJcklQP
vgASxDzKxPyr9hp89xLl8Py3+z9IR2c+0SaO+B3ziSC/KN545L0B51oSWPNzMMOJLksRFJrjGpuj
2QiyVCVPYkQSMxKZGPxyaPSTzQvb38RKWiZAosQjfYRkp04WQKtVrqRdQ6rZt/5vj8HMpGy6xR3W
twauYALJVTsLH7GRtzs21ivcBrnA73mqIxiMjdEpSkQejP66jq0DcuW0UqIjuzxCS01OabEH4QEF
Dc+f35v2f5jIH8/gJ0l5+FjMuHXNUSHZeeQB8VBsQJ4etBbcSYqZzFigparHBQMqfPNbXXHcaF2L
8GyYysUbBmblmHUy0rdyFbY0x7/3NtfccoOHfx1dX3tANtXOMKcbhzyeUA/6gUezu16EhBLlFqD0
WPU8Z+Ytk+dhQRYAkC5JddBk2STaiggksllpLOcWy6J9Kd8j4B8yCJHTZQF03q44JRuvZwiilLAe
SMXu3ZQCmMGEdWt1EZ7i0DvUgzwaXeV5eWNUn/4+U++SECr4Bi7RyBB7K63dqkoyQ6VOQprcmuxN
DIZARGhKz0hpQYR1FGDAe0uUOrhxiQZpBQ5nFTM3LgkMWWFPmiFwKbTQzFWo2rv1JPVNkGRA1tA1
BXgYwN/2ZNqyQ82BEqxfWpu2IsTfty4xhA9sGJi8I7Q+tBvzWT5EXhg4HaRo48NSOiCHWub3FNoB
XzxC39t3+ttewGaQrXjo9ZZf2ZKHj+M3xKCRYgCmnC+ik7/BDHKDQA//dMhKVnDvc5rDQ3F/ql0O
v85rP1OaQrKv2ZISFkRaO76hASmCzCb6bszWLT9c51aLtXamrFf5hwrtJVg00Mw47Nc5J6UYLrtw
CJ+h5VqB48IwYtY22nKW1OHDcY9o/XZRqAM325jUtZTcye4bVNX+nS8g8eQZOeYi7YJSNxE2SIfC
rdj8vIXX6ZMo1TcV1rLmnr9JiT2QFVUNXtsV7jCUx9COoVYrUSjQTjeK0B2VbFkLp6Z1z9+CiOEI
OnxTCHl6zBCPGaPvD7/kPhIrBmQvLWhZAMaQiR1nzt8Jg42j6JJbyQmZ5AOQarNAdMel8M5GxgWU
hT02JUZo+S5uLPcPz6j8PEqQGX2qQmpS70Vmsj53/251oYRjjXOZWNa5dXRSFCw/73OWj8ZQTLMm
9t4U7eiJn0SPsPIta2mkLH80cJZxDOwKU/pGIHIbskRV49yXQmLSQl5OZeEGCKSHtGIGFke0U7Ej
tTDEFpm/QSpSH9NMXGlT2ZRLNLFA3T6iTuJ+xEAGTmFiISWzI2rH8qP/NX2KwOpnhIr/KvKvYCo/
BLZtsOUhWp6lWZnYLhZzwjzJUovhh0YNTAb+AicBpLS0JVypWvCEzvJV2xfkKMv8epAYbDyCZEr/
vaf2FumC9gWLEHZMM+Gex4jK0nWUcSMEvG82mnUxjTX64QncxdiOJLAbG39Z3QFAFN3f1rwhfjFj
3H458iIPS/U2aCPDBPBojRzBH1A4ClsNH4TRL5lHGVmPn8rNgioq/E2LUN5eNDqBrAs4usLcNFne
J3mUWfKkSDtD8zWTzBauwH/zo1F7+F8Dkebnqc4n0OhZfxJRph8ero/zqr+WIcW1V+5UPL1cT6bw
5XfFdcJ3/0TIe2WJlnzqvLIGd5e14EnZjNeTu/ZWmYPa87HBTMAkc0aVc1UxXZgGLdFBQQiWClL3
9DDpad16rv0cgkSXsXnDi2AniGMPmwWusvbDiHfRUpZcKqaPFKWwKjbSzP+Pp8i4ysaiBujcqbPd
Nmt5P5NzyC1eQFWeZg+B84rTvMZOkGNfXjKGE6aOTfSb9b8O5LFI59RT0TaGdYGJzCZ0OutCbnbe
ghixZPRDgedSQH9fu+Jr8HjF+HE4Aqa5Dag2FQ/YNWv2sSJlN+ZOgFZWixQDswce/o+jbBqEHvrP
0pLt39aa04ZwF9KPz8spby1SYKyd4JMhCuvux28x8DGlqDRrdlyRiGXq1PUpJbTgeMO6VjHW5TvZ
AYDjt0YeD2TgRNOSu3sKEsWBi27K/waEB5zu36/Vh5hRVeq0QpAQUY/TcVZqhHIYtL1VW7fmwR7u
0ymKgu+APJkviG181H5c37Xep9dr7zN0JqGKIVObfZkzJ5GmFZ3jRC/ySwxguqmaXNqFGRw0KhTY
HPs9MzR+CjS73xNjTFHUp1KpCbnd7tgmHEG8H+caogO8kXDE1B9MUR/QW4ESDPq7JLcYOjR5+ddc
Jl8dh4S8/Cd5sFW7VoEkyAhW5YBLSNqwmlPGuScUtywa0nmNGPklmGu4h7U/65+tlca6z4DYOlMq
GggO6Fjnit6k4sk4m2BSdbU33RDCmaIaSCPXvOtKj9fsoNRRtYTROCPaIOxYoEXbJQ59KF8zf7W6
geeNZKQ65HQmuqmZ/H9wEYzcnt7/ShVTxZ2auhAA7EEWRADD343+rPbhn/YahWX5N/KxRm0ae1Ze
PdW/YqqoBWx8bfrCtu6fbFjoGarrT6VhXUdbxzqfXQFalkkYp3RnZabMMhm4FNFWN+o7gw2c5eag
zQyFSvycoIGaWOaQl89jeyy+tlKEvSI7lblA9KZe9YJEEqvaBsBgnpdy/sKaTxA7ixW+0c9g8ps1
5w6Id6M6nz+mF9rcnBHdfpwM96DchoUaOU6lVkz5Agqd/ACLTqYpkMp7/vuJRyov9G40h5ezb+Pd
sOehd8QJnBXwdMpN1+8vV01A61TU5UNW9qUn+DAqgpkh1zvPag21SD13bTkEyzs8mq56+WSw59Yn
tOz4jDoaKaaw8IbiZ0nEZVnsbXQtLsRlbel22h7MmULKQ5goSHCB/g0WcaE9sD2zS+BOVHdhkB0d
C8S9fgcQpkRkvkUmOwazVX2t2brvmgZKx0uCkbCQ+oADJP/6NXxeQjMkYMeA5HEbl4EzxzXUQSzT
IhmxSjqGeLn1E45b5/uTDk6jNQXatBCe9h8kb+iB2SW28SmSq37T/altImp+G15zPinFa4/qz5/a
iCS7lh9LnubTSbvMDvt5WHCgJyOlwVzNkOtN7z8FYMm4cWV64pao0z2OvYcdGQD8Uwhhz+MtRoPF
sN4PRx6V9az4vcqt8J/+BwY/us662mz+w/Nld2YecQnOiZBt1czI+FJrTv9gusTFgtGyFKmTGNqk
xdbQI4MGeya+gnWtF2q6D9KKiVyQ8kwlYObXYQtVCdOQJKMOMkjNtRF8/DiruHjq12JZcOecscm4
WWJAJuzs+iVOByYBV37NwuX+H1dtONjOPkXXM0odpM4jPoWkddaVfAgBCRrjUJ18kL8GNt0Hlc2Y
MNHhbZAEL38V4kMyTmCyohMEIvTwTa9hrnQwtWWEtJfLWxaecSMpoH0ClOMfFaLNVhiLQQCh3hFS
OTfBmIHygUV5UZhmvsN74XSjZMElpiamzVscMmJB9KK7Kl7g1per1zs1bBCHJO7KZK5++IrPhwmw
7Z24zlFJJ5cJE1J/8j52cAmjxZ3KD/MPqXfXZ3IVY9nJvl8Mwxb8/WIrDcosDJoyPBRFGCI3HMGp
EtWGULgII2PIbf4fTerE5qbvuB6f0dgcJm5DoHq7aUkzOv2+F4Qt4BiRZyYYVHkFtpcefe5J5/NB
eDFER0mseHEu/1b7xbgXD1D07oZuyMn4wqEtEl5MWWr2aaOSjLAQMJ20MlYgisC5uq0TOsJMzy6Q
whYKSkQPZfIOfb7oTKR8SVw71+D/sbBWToKOGW4w+cP2sYTTqsWJ9L6zQkhpBqcRSVHaQjCYUrBz
AJij+D9wU0y4U2o3MA7KOArKqpvB888s9Pf7QA22w2iNI89vbzdqmF5M6c1GyxVNkG2UYxsqgAgh
hShUn0KTtwtTicthPG41q8PJ8gIob0I8dEzX4vkdfNkiiFLzbXIFB7paZlnNwKwWyO7P6j0cJjKz
H6t9PVl+k88mOR24UgwrFsr5ZbpcKCEv4UJkMOjXGpjWBsnS/duD6Ro+RgaULUpL7BLbKe6yGwE4
wvAemYMeHAzYRXo/+PvlLOfzgWEUdIZ/V+y7BMex36Mjj4GKfbgKzLETuofL7bhhHSBNtfFH4bxt
eejfyVKNUrxBTOQOUBHMp3n3SPTmgnzIpD9Bu1C5u0qx5yfFMQnVr7oH2xjCIJt8E3J2fpcvcai3
8huXj1H7V5zj+zToLDPK3ZUgXJ6+isGfPWDi4EEeTQVgQJNiDBDVQKGsTFvXWk3tCpHh6byCqDrQ
U+InKjYWbqzw3782JBrO3AB2jLp4VWBUbDx79UeW0CTRBHJL6re3AroBL49IBXVsoNRpbp9SLi3N
/s7SZl5pPH/alZtFw3jMkunjr4DozXLQI5/nCNWs8l0Ol6hmequ50FyjG+DTsGWLrTtgvwrRtXPj
INEpnXoCcBSwnE4YiAkpdCG9Gb3PDI4nBuMivnWOnT+KcBX0WkL/sD9F3C63ljo0FzmFU7yLIF6s
ipG5qnrpxHedSwXFlKOB+I1rDPvEEaYxOmm8IcOt+1jzJcAV5w4bAL3vdJw3yz0o05GbvVGW0+Y+
PoHN/axUiyiFUJ/DN65iK3RSo74kSwzhCi8edXmNnScLb5JlqZDzCOSpCs1RN50PP16Gsrajxzx1
HtSIGH/7/ca6nVbvkReJMsjt4TaBelF/tMjj8sa0sD1gs48oTZgK0+Nn8lgX1Xpie+Vt8SOjIHc9
r33wlluRGhlG9fkCqKUHxK1NaNlu7kpQhLLNnJX6vWqWYimgWBMCA00TuVm42PlfT9+ymioFKXYp
+FUI9VX0wHjwI524UN7kUP4A6zsUmZMVi9IyTl094mpn56SAj+MPuKb5qFZmQn1Qpr8IhGZlMfsi
xXWMGzHvjUdhf2jtlmjPBdXXAyep87QyZyeywXlKsnX1vCgDR6gQvObxaHYcSDTTcEun9dezVaGV
4n8JqF2eL3vzJqPgtQPa9a6NO/UT9otRI32vUsLkGhOZ6C+kqiN9/IgXdih2WiYh9FM5bbFgBjaV
SeO3Zls/d4oH8bs+YtOdpraXwqiIVLF1cw4aStP2zGqxDiIqKocRmzYebzlmG6AOe/6NbJ8MvVpR
dRiO6jA+T+ap3TM9F8R9aHw1uJpXGy8//kTdr/ewHcsI7I/z9pchJ1foYbT74u2ot4yWolgU9usp
v4HuCel+gTGEskVlf6MoCRElCTrJqNFWdll13DvBvUu8b0S1AsNfDFBK0+VEHJf2Tk5HRLek6zrf
s1/q4RNo6U1jys3ULWQoLRqj4fFmI2+IfzxNDDlt551Ufnf+EoGyCKDoFNvyX4mQe5eiqQAV5n9j
N4oCbp+rNkOQGj936oFR1PddZfleYIsZhjkj5ir6jUf/arpK2qE15lXB/BZ9OTQ9Hk+jbxGhBKlI
3MjGeNgBWTeo7hVG8UHdYJpxAYzfB95qF8tnCxXBJjFbawTHwnRB0D/c0hIo87HFe1QusmNsxH4Y
V+Bli9L25I+Z0zKi3zo2UA/nMhxtzF3XMnLUvs5fbuI8c4Oyn2SD9A7ssPWoA8xHbIMSyIEUgPIj
MAzCiEYix7IMQ1CGF4K6O8SK3Q3x9de7V0FXuK2o9cu/psuKEKOo7pGKKvY3BZkiVwWevBx9bknr
YPMbSUyOWEheQXmeocVME7GUPrr9aYQ7X4Lrhih/zk3b2KKoeA1QhJv7iXQ8h36SF6OEopzScgnC
WjfwENysmCGe49cvtao4mIZ/qMtKYBsEUe0X0I2GVsdKt2U5LIdYggsPLg7FEAr95171g99x+coF
H8mIWSdUNH6j5tV4d/r2P+Z918sVMKIyx6gCVsHIyjAhv8AtlVKy8DnVpy3i0YQohteIEHZpMDM0
Cg3ZQp5JR3URJ9dhbAuq8FE7LXATJ34l9gs8drSQ1QrnE5zzGoJ2AT25c/qGAQA3NwZ4H0eVK3M7
BwTpMPX0tSKsckcuSblSsskGpEPKECgilUBeWmKbzo2l4rNkVvw6vKllgPDC3g3Kder5JZXWtRD6
Y4Dy6kS0QTZRpWhBcHMyPiaISMSHKDn83qQbjpaiRO3N2NeMojqPlwvC6DDV2F1ly2yrKO4uS425
EIPNFMzHmI6VJbbE3/K15G7BcgKfiEEfaqBfPgBnek+likbTVHqL1z8J1CDQ1GUn7ZSVDDrNczOF
QfUsn0y3v/lT1HydlVe5v+cqGeHGtqiotF6PnGqP04anSSV3EoroTkwPbqaj9BiBJqzL70Ygl+eE
rzAqD6yYj2/Sf1yL7uuhViGD9gFj7hb2s/9+BIXg6/L0ZNVHpGYuqo3zNIUNU3Vc4bWBz0tE3tCz
zszhT6qOF4/DucyXRh3MEaxoqdO6nKYac2SgzsuFF3fCJoxmk76+SnUDy918acIy/XbQ8Z/sESx1
PJUNAblI0v4V4HnScJDFtxI5obw64BA5N/vPQZAyYCm4i8n13v3eAZwT/y2vxGJl3L3Ssx5vtSq3
t2qwYok9E27N2rp8T5UPfMqPEqNSn9cgBmPxJHLkIIrUVgVuayAwb4jEm2ZOp/CHnKpkh+wRHPA2
z43h847OVPfEO2FqHN04W+DWIQesx5Gl4nj3R5ROw/zqcdaUGXsCoSlSkk9Ns02r4wMKD9vNGkN+
NDFLrSn2mJ0jrPitTNQJ6XdrckRX/OixSbVlvuHfEVVR4AxgPo7TmI+kcPQAOP5jRc7P41er2h19
vF9s4f5eVugbp+MXlYdN2r6jCGdm4DAtvFGcnRWvQ3kbD/TIyswlT1Gumuv11MtEZrxxEWPaDI9p
hUkPaWeun8be8fNKYjBfyKvmoS4m6RwrHJcBrVmQaWpi4HYJWSd+v79oI0NEgv9+2g5J/+P8Qboo
0FofgREztwgf8vyBfM/vVdrw5miW0FtZApBtBSQcnkT1mhalvXvj87z8bb6XETP/v5WVUVBHadkO
gUb13+qmvVyHB9q1rX624EP3i1iGiDPwhMQcV5dz8tcs20DkxeRuon1ztSSY22tmQR/LUJ9y9d6o
5oAFsPKbb8ESCtHYWrn7zLWtvO7T+dmtSFQBCqszxL0hFJaBTE0toTGpM8sQceQuvL2JAEk9liwY
iIlpyfoznbz/s6ITg3XgQ3wL4xRa/HGsCGXJpWtSpRyCLMeJslMIVIUB7ttqqSAMCf82iWwe5FiP
Nhd2ID54G3G6Slc4n3hSjtsDkEmxqKYYLNgf5jgvp4PdpVzm9JOKMNfkUjhKSU5tZansQwaClibc
Uu8gdpgz1dQDdHjQGN4bone7HPLLSvq5VO/tkBtpitFxx27T5wZFnCjMIArErHv6osJFuPJnFAhI
SRUfUl+3vVBQXNX3Do4VgP09VDg4Ky26C0otNPFTrxYF0KwjEeB8HUrKZrNb9UaJRFXPhN+DIdnV
Hk1Wk+LHQVPf6GIrqwnaiZki231Lun0j4TlATzEHt1IGMt7wW0gZQL7wedI77hguOuibDQVhO6W4
8fRw4dM47qJTTFMfhFz9RajFok4Hcgkxqig4K6P1IwE7R47f4aUK5mlwuPv2pQtiNjP6cAmP+5Gd
MPFPx4R5I8VPvstHzO9nqPCNw8lUMcGw4CCim/fZ5Y7OpUF4cTLow34LugUo1ddJ+TW7n4C2+2Up
I3tNpIEL/EVMaIXc3/NaOLzaZa6P2kY+s1L9bV8/mav/hgtBCsyEsja/sQYKvr71yiL95avJtkwq
cdQxyUNmCLglPnkASzwvf+KAGgftYLB4YQ6PSPMLKyTnf1aT5nu1cfkyQcJ19p51OpIXKvvWIYU1
Ei7m+jwf+YAAWtSVPOJjsY4xt2okES+aGfKirpzSUulin0l4NiPP62WAHWEcIa2WrhE0Mg7YenwE
3J7eXRdPtCNvVtCtY/yOWpel4g0/EkM0pZSXw0jU5ZNEicdoHG4KDfmfndrxSMvGLMNOWZ1YAc+Q
AWXTBWDZJPe06HXbdBTECAq/9ZQ/uToXNWza/TupVS/KAdHt+D29+6DnI3FIhQW25l4wsi4BYOuu
nZawKlp1koIigAHZrwwPYZFFjbhGB2AkLjGqNdHBsQuqfM5Of+qQAyHGseURFr/4A7WAPzFv6R0j
ggSuyHwTbL62dlWZl7cjpvs1DGNFOqEi9aPP8rqNJXi+MsHPL5OxV/YSpOyP2+WQNB5i4Xfpx088
WCBeX4Cr65Bmiijzfooc33bHQ4Zfd+cxOD8qmtOTvuOqyM64/3B+7aduk9NIjvnmGctUcNeOdGXv
/d/yNRytKIdiTdJXtZEKdUSTm+tf22LgXoDPamA28HK8tior/qiQi9hqtEhkMpLFSsXZUpu7LWo+
V52bYR7jQ0yPdIu+OgbG1oRyT3C0zPDzGCMzi1BHvW4Sm8M9EUVfRjjmbRAPs/fExYbd6O/l1aO0
e+QVWcmc0XikcIq1rq6ESsClBCWYLhs8gNRQ8jYunXb0SRV36r8r9Ffr/JwuTCF3ofwKz20Av/2i
saaYVrr8yvEbHLQM10FOvCCe8DtiD6aUX4NydglM+69QdOgei6Yw6uvBfYw4MFA4QOcUluJBW1zZ
Pe9+PnL8Fpj00k3E2GpTA5GXCcNT2pk+OFOz3mIDJSWNPAT/lVz76IcKad4AXyGMBxBhaRd2A2eF
0R/F4Ky8HjBw0QDtHGxVoglIuT7FuBnK/XzFxV0+q3ncvMBhd64bt8I53HHdlcAXVX+BuGP9uacU
qlzOSZfqbwOo3x1YXTDxbzrig5BIxB+4p9bUYMdUKB8M602Xc2o75092CUTIlg1EnaD/nhYWozRH
ybt93rp8yIdg+qwTUHV3Kj2vYhn+d+k1IuCyfdigSBVgv5xeOM1URUr8O1mMbc7hnOam6qs1hsiE
xdE9TdTPyRoQY5/KgLZrcKWpEC44wtE1jjxkK1Lhauwz1c+dvcobVjplJStS8Ig1GCP9K4ohx+Xx
J4be5XSzbyNLqVZw3rhi2zM+SJDviUv8ztj90T5j9WEA+w4YW7xgxZeXP4YpLKwrK42nqpIHlFx/
uAY2/cPYPVnnf67bhc6owENansmULdK80mB+IRHOR9JUhwJjljFSDq6SWKjpeODt/tBmTHja9cU/
CPfL7EHa7Uxqo+q7lJ5+qGjYL5hqivcAABB84eMuhTqVmWLNEdtjAo97LYi/03raS0eivYAIL1YM
unk/4Iap49doOJ6sjnJ/higwS3JCSUqWt+JGhDwRkKzEbULuPGT5/3HrZi+oz/VBE84ZplU3Q/5S
V97veGSg9RyaozSwHA17l722Edre72aB4yrS6BxfvFE+LWQC4N4bUTNZHwrO/ivc6SM05eXQZiFR
/rzn+ADEACW8s2GNMP5AQBwd7lawjMM68EU6Ls4Tdpq3t6P3g1gpArNIusDhqYVre6yOOCHrQTf/
kjmWQ7tyfchXVWzGxEiSXgwEklwFTW8SjWwmUfeRe+JcyvAvjek5Zz0NoS6ya7M5QN6jnxaTJt/Z
pec5OTZ7GPyRTCMSUSU9hKCr1pouUcnR2K4doQkEYcM3LvMkpCvYdzroOtby/wsqbEkFeH+yr+pS
K0Z5eFPYRJnMs84//tUrIZQfwQDWQ8GeWLeMCO+IfnnLV1PpUwHV2+OPRXvXSYR6EpzRs8GMf1xx
rbWZqgV75sR61GezLFi3LkZKPla0VkrTAb66Q9grMuAF9c826zYnPfWlouuwF8ANrFWu+Loc8P9h
YF4BPfv5Qim3JTKucMdV8Y6sjMbnvwW7ZBUEv4SCY0nDBk3qmUcmiDP1eDAplnoggRmCXEh/LXuX
ugWzBa8CwIwB2+CCDSTcR88FsD1McM87mAxzvUQWjwg5vH2YhSZqbF5Z4BKfouCPfx8yVqmWXu5i
/tZpa7zJnLA6ep3jNg1Dm25H8KyqBhEyeS8uIM32yg56vJc36E79m3OXviS6OdDe326CMEBcn4PP
OA8BjaD1EGb0Q6cosQ+tqNF0dyWPx23KalnmpeAMztDXMwT8AOh0EBG0x/6/Ur8rKXqoKS7Mnac0
vL/LwQ9P59o/REGq4dDpw7is3DehuZ8u8UwrcOwCWb9it5x3MZwm3qgZ/7KyyT2UTPaDZEbIN0YP
vk5hiphqeHpu1d3qVjbcC2RbEN7QJMjhjqHkQ4ewf5c8x0rkmY1scpR8dwwRaePL/bD/seo8rSyh
wCVrL4RKQlI4sSc3ErMv1ZHijsGchXYulWqHHa9C8kKihujz4AlAW0MivOPELstwq6UcYspKzIHj
dkt7Y9mygjo6MjnhaYpWNiMHCfmuhZadowMuYH3gw4QhRk+GMPB+JFr6T+wbC5G2xBBimm/3d2Pm
0ft2ZM9K9TeQcImcGpks3ac2xA7ieQTPTJzGIho4yO4mpyT6fhpGzn03FT/OKy6UqaY/a2+NtxBs
lefrnKTnVmcV7K5gaoygeFBTSZFyE05Q5Il++6zLYBGovvG3sF06YPca2+lNUxTCNh/EkHeDK6G6
ddKY43qQeCTDcGn74SnD13IRP3Ob1k3ee8NsyxHqXcLd5a6LvKkgCMwpZcl3tCi6nRDuFgz8BpSM
QETXHIDBd/D6uLlVrC5DJG3Te3HLoXL9mZqs7LuMKG2lf2w0SYVmdYEe9YRtBu/3abegp8RTLD73
orKUUbogNua2H4IjtbsBvsO7vkMoj0bGPfpF6zlzkBAwOr0DHONQnLe4u3msGeaEfZhGWd/FxJXd
WwHKMomadx4UVOoGADqm1bI39tUbXbkGRAniGFaau7tJtQV1qqddc6QLWBzz1591Vf03xcbZJ9cX
ZX/bRVaI0KEPdCxLJkdha9P+BuJgee3z9CCvEtDtYcmWx5Liqhbl+fAESGJduNo8/Pbac251MdOe
KJPrN6BfXUr3MxPBmCYWyuDYAPHqR6vgZE21auDamhU/NX03GbRJ15KfD6i4UkVkKPTKnPLQ6FSz
49BlLIgGLK0tBpGR9pBdAfee9xYUOInudoYCYqk/pZG4StLUB0DhBymqgTK42+Ql565yuCCsxZ/g
sDc3NgKHqaPLjGDdnbviy+2eAnLL9tu1l9c1saJXpvxYXYtNTvIq5U9o920WWGgMkDSWTsFmnmCL
veYidPa7yfAuonJLuAkxr4w7YfNQLfdRlNFZEQVGw1g7f9JmVAoc4IyzZPWTIbYWFcIs7SiGMMQi
weRVaShZEi0LeqD84H2uDX5dva2rjllGTDa1GSzfVOLDirC3R4n4cUcNn3A7USd8arX8Cj4bK7TD
zTxYgzIyWBptfkGxg0KCUnIZg+QOTF5uqMbW1VgsVRpwpB9BxQ0BaeyXpAT7MmY2vXQI1USe7of7
Ma0rB+eelB9WSUlDFPYYLOcwRpTXLA0PcQgGNHL+4Z+E16TluHq4tDl4krHNM0bwIg4zyPuKnpzl
uEBwKM3x9VjpP3/cTZjO6UUA9u2HoTnxOYUbrX5W9QPcjlsA9kZbAzu+GND3dMvx616fKLT1mkEt
n7NQR53a1h/Sv5a3K8+CXzUzk7csyOLnbxJMt/VcIpbkVOwznCOqkUBeRZUQls9Rl81AKEqE9ixX
XnEF3aYBcwwUOMtWKit/vrkhIur1TN3cyRw4sMzYYktqi7EWYPr+78gaXGYVvq9q+6T/91hHB46P
W4SThhc+cYXIqKKrGHoSvhx7/ob4MnqXqMDXXKMeTcLuGrsqDHObDRq82uBvqn/7jWBHvJznsTVe
FWN3DWO+NxB6O/ZPoAhjj5IP69su2nmUXuJcP+5cWT5yYodWUp+xcy4V4E6pvTsMN+1N1Od/pl7b
oEXVwJEBfh7V05QXBbHLnskANIRrDLEUie5K1e8hnmo/P/gkmoGmlF5ouQ2Ks4X6H1R0pkUOq/pH
3a0EByYxakS2k0+y0+r6VfJHIC9UNN1vNUY38aaGXQ6DeqQkzagdNyURPks93N19o2vWRaLVSl93
PsHfJVqibOwIlixEbsNMQ2JU9Da8TTxeL33pG9CHqCCrLzx+fzsDcUqnOfng3kUtiLbPq0+gQ8mw
wvnAJ8S3KTFWmwR8I0/hHvSrvGinWRV3eZXlLPF8sttGH/2nD65/zGIMW2vJb4oaggquJtvvClMm
HDRiFXm76/79XsnscJyvqxm/j855aqHIFCM6xEl0m+mTfoWztNj8URPJhxBXRUPEf6WSTqo21ysH
noLAMnMc6WoSiTEC2S3TNPaMeHXaMldhsWOC8tZT3uVbx9ttidBkaUTZz1Zqn7pDud0enYHmYTg4
bTmBwrBYUxs9LXsnoTlGAhmm2Gw1Sq2ghRD4zERgd7wRqQLWXhBB41/fzy7ub6R5ZynIfbUpVBX6
xZGUQRqptEx7r2ri4XVuczwGl0m3VMrZH13ey863Txc51X0d2Hle3NkQ4bYIvM8CDLA6xcLqxbBd
y0PMP2d0YAvwNeUMUvcYHxtPhKmqs2R+gUKFs9GyvBYeSIt6cM7orX4w4ULNx9+VXuf1KYmXj62j
QXTKGvjTaF3XIKfznWiAzqY4op/2TTFQZ5RAK6MSZ4yH6RtT3v7IUbjV2ulzuYz7/FD8BZsDnS+u
7Nr9GWSFNU40RU8D/UDnv/gQsNtXzKPcSr0cFm/uDaPByn8WEHHK9hWBgnlTFThcqMMjMwNS61C4
ktITVrShPDQwd69tpe2ATddClZbmK+IUAEGwKQ+4FFRK86wDb5sT76bSHMb2sIKz0TXPlUboe56M
mpF01hA1LXaaASRhxXLtx9C+n2RIrfSoRsTbhJygsrhX8tTf6nPZu5T+mDrj3xdaI/cfS6QNkDye
Ib7U/u8p3HG7as885Cy0c2259z7T/DrNj1EBTaqDW5tHeQnSa2nk/9rzwMgoFAp6iVWF2oyag4oU
+bKIPw1AwBFHjycff47v1l9caV4uQyXWcyj2j9h9F5uTSRNmYVrnKL5ovfPyZ5wdoYMNKccIW82Z
2xeogohwUJstu2rx12kDVNqhITr7G4T8oWTJvUuRtdnBT8CnJBKMTbfiAChDzP7ZnC4zhBg0oetq
GRH7Ck2a+RvgCkgedATHx7XTW4Rk8Q5TTQRWHP16d16ZNHtzc9HTEQJnMTxUwAFF78HLUhlGJrau
pKW7M7CgdlO4wMhH8jdhibLwVQHLIUSc5zzphPAU4jI51YXwUk02tJDzubzWHyND/I74TEt223Xi
1qjxMhSnZwLVQQAzsTZIaShWrQyxxxQSopSK5zRXaIOG+X0nVAGJBzc4bOTEGAVHA44P3AnoE+YB
NuEoxOSnX3BkQ6qZIltSErloLJmC3bJsjlpEMWUO2ZkkPjIhq8vq4ihGxwhKuzADiBW+fAAFBzPF
/bLFf9puUCRAtxoPQQfl3U1xbzTfiPXyOeVglGrvlLo5WVDONgdYl06lA+Lq8ZBbg3n6CjJWam6I
0kVqz2/5iJ6ZKxF7cyA98NYA0XcqhhfZ/f1Jg79GLz1k3hUJi80JRpDncBGsj36im35cjLm1HH+J
efBwgKQ4jwjoLMZy1jPPf/g+6F9/2DtAi5scVwCxUVtdCaxbJK37u2IpFQy4LR2XpKRObrST0EUt
h0X4tdRCNOXSVLEX6LP2zpORBigkl52MDC6qo3tX8O0rpV6hZNQFTpZ6BDzL6666yGADspj9ZnWc
SR3/MtLthL21bkZh7uDYAZsHKx3iI2UKgEJO91qwabLxyxxwjoz1zT42jbZ4cXom+pKyxB8/UF/O
cnr+3vhuj/5ityoKIUY3iiI4YT1WY0sAHPFvaugCQ8cIgx+nUK5uG6eroBM7iyonyPD4/nuRWd9G
GzQF3V3m8PCsU/24Y0qiJMQlCxfFzOWSkO3TRGTNAwVsrpNQK3iXTf6bLxvkgXn+i9Bz12gQy3a5
SL/jlOMRYuKan+hEiT4Yrt1gfo5Xf+W12N7bh7MsriUSR3m+eMQ83rsiTF+/2KtnPp52ft9TavwX
7nzRQpVt2QWSdeZnCn+H9Dh8A7a/RsXWJBBCRUbB9K/KPLI/XGjpvtQ6PNNSgWejfvqRRUK18rvZ
mgrL459caJZKwc2qRGvuhGvDPskaPH4EXvJE79bEaz7/8k8QpDKsE8TIB16YGFpGpuR7JZcZT6aw
OR73q9lEq2eSFT8IMzzd4Gqx+hzKVxTKmM8jRCRX/mAMNUqGJWTeszFWhLjNz05oqTA+nUXSkBp8
VEViaUEpNwBiQE6u21ukL9XcGJEMNkIFCdVXFxy6wo4oK5OY4s820GZIcxD6mksUCvo9P611zvFU
pOmCK8pgtx+QwCQzuIE0gfCXRW7sxniNfBJ9gLMmNDJRoSnGcqKZXtHdUpoHr/SQW6/QMfOWr3zr
HPGaQAcil1KxTG82DRGar+WTk+9isV7iSLSqo10kmLuzDEfecK8mEeRCHzTnH19CHBais94G3fNx
cE8c6rTpQsvv7GZMWLaS/bTfrLCyT3kYJbZeKQVpoxDAKYNrPDe1oW+U/SqehQO40LdYK5ssJ6vs
FsjieCitm0tnPc4CPntEVOJzTzY1qzi3xl3xbFAA+/PzfDjjy8pWnlvCrlgOIgMcVii/3P4n7JqC
kaLxgzsQzCHpqbiRxSFiMTqo8o0qvFvewYOfkFpe23GRpwLmJbpS6zLnC+eUmgOnHXlcry2kehpM
5EhF6O9tnj952RZtCwB76BZ/RdxzgW5TdRJEV+izp4Zlv3pl9/GvzBNYbbBmREPl/lQ3c4L67zwu
29Qjp9zdHAUnuL9loZxbMVHsTEwPVLPNE5cptZ6Q4+5JoioaRh6gjRGITdpW/oNGB6v+aDJbg7l2
SWU1ZAhK9Preeo9gQfsoLEKLO/IW+3a1WKRnsuOHMs+4wtKYLVM9G5FFFT1pgIL2tUBtG5PDFbfJ
PsMCdKWJDwvbbSPVa2niKRVNsg38CLWQ/qX7vHWY4vvCEhkY38vmtlpIM1VI78WxTrBF0HSjt9uO
tM7qq58+0TxYAqDMRv3GPp8/aLKqF+KL/RZaBoZ4iBLvbdiYfuHjiDHG6ANKvDAssDkX6UqHzCaM
a6W/4x/ziEVisFkZwhq1jAF3M5HjTbJiwO8U+ruBkHKU09gKf0Zb4UIHaQnZzcEgeJUjd8rD9Puz
lvgwRClRCmloABikNxyjO4ep4MUuAdNe5eRtGwSYrUV05GMa4Fth9eJuMQYM3wUfw7DCnXH3zeXi
x5k9kxdbxbEnzYrnuewdf1vCeJ4gGHbHb1Uridx8u4zxQhhroOq6vMvnmGLsagOO8P+HEpWQNWx+
dFRG0lvegxKD+r5GGuCKhFYZOmmg3vBpwd61s8US3V4odYNOrSsPpTNRx+YfFrz8ZfziH+RXOI87
C2jULr9o2yW9BJz7FdWq2AO4vdG7zZ6WmNYw2Y0I4MnD69Hni/karvBXc5Nb5vjTbC0AUGRAAoRm
XTNAId1b8rFmRlgKmM5zeOd/iK1X8EsiKM54vUuGCJ8mxFNSxSSDusNs6RrOLo0G+E+JmPKjQRb3
iKifFSWD53wjvsyHbEnKGxoLNmVTkSytN6CoRUAEq6kJGpMcJwof/VNJeUA3JTNh3FPB2UBfCkxQ
Fw0nU5XcmWh+CxSZ8q4O//WsnMvPYTWk6F977iDrNUMRu99ifISKsdhGn5ozGy6ovDhsK4nWWIHB
x5v0WNVynSspJF4OTju/vMHKRGkoRIyj6pg/KLQsr3vRwimdbS7vtlnXk82kSr8Bnb5YlcHoa4II
tP62CqPqVpkfO+poHjm2Ii1GMI56lO4fp0n9bxxaXy7bXpkU7Dqff9bS86Ya/E0K2d/aL0fCmYMT
Xph+2YEhU0ByOp8pukgnigSjhFQ6ioGRUN55qJMIdrQmfa5dkbUJPFZOHmHRFa1NmsyXgspiDE5r
XkdUGDSh8cP4+a5txSKTnnHMywEJl7s31yLOeuE1QOsQmTZOdgApYBBMz0+bugH5kqGfPN7FlEly
9/zbHTAJta48R0Gi8sB7dEZR0jhFOK0z410I8MAVcRaNAoEXbXYgOQWEU9zMfmV4+5sM3Wxngk6a
P4p8vBq3O/i9vdAqMlfpZQ6vNBDDv+QnoiMOYoFsFGCjblBqxU3h1T01VwUDxr7f1i3vvKBHJ/7K
qD9WAPoO/M8e2V+Ppn9Pk1XIDqaA5GQTodWf5zWmtjpHMEzwN+i6C4y44oCutCcs1uMNRb8+ib0B
4xrazpnGI92j6swNmq4r95MWsNOIxugmS9I+PEnsY9c1dZCJsJ+Uyp+4I3hEddX8Mp/DugbA3w8o
f/jKJLY4ezfTIZ4aK0a8i/WewdvIvrdokEjnE9ZCkziYjI298URoJU7FhYBfK8IW+hbmHzKMz5Wa
XIaG5g51NjZbNupke4A5OXl6/0gXstcAj7VwYwnAOJK6E3Ur7xlJyfmiAxPOSVxYvbxZowqsgLwX
IgG48vCr7pZAy4twpZ+DjFlpLFzu05vAq77qirEVNSZ8FAdNJ6CaZIXl7q93m1IUMyjJiDcTeMNE
X6/zXRzNf7/SrjyDux5U8e9k7pPbDpKwJfH5SDM8xnckG2/0pNfxoD6YLPx4Ldnx+epnUyw4NN8Z
exq1Z57R6JEvxsl38q+JdHjXsXKCt1dp4Pc3ZOtqAj0VjrWGi1ZqSLX04ZzLVBARTZTgQ7ZsKV2H
Cp6AaWtuSrytqD5o/Pzzdy6Zh21xts3otObBMfxdFsUVytHi1IB8kmqpzJ8iP26IlXfOzNwD9FMX
JyqaPX/CUt5JDXlU1586LcGlSVecMPZWvHHCzOLbpO6lqNuYeRvaF4W3SmU4UO02+0LukEjzxUWH
TOuET8XNQjl2XYYP0qw6UvYdtsJF32vbpJLRSn4FkWwONOBzbZWacJ6o2wuvAa+foWdD4auj72DR
DQYlRfEO6XrMa1MNjZmZ7ps0pwNhfBqC/apYho/v/dIhYp3DPHFDqL09jqnBR6iFz009q2eKq0+q
c7rKW7tFGeGn4iIyHO+mBjzPGVgL3+RmQuYdXYMi0fVjA+mcruMRFnvxIO5bRWpAZp4hbsTP4Be8
4l2Q6V/LCPTK8pQF92mg+vmuW5zHl9/iMfeckT1OXFzZt+zAU8F1tgBULj9+DlreBST3zWbAeCd8
yDbrCRXqnUKaMOo6FCHDj+XzLwbIlkcaPLrai6fooTEjU05THpWIt+EWMPCjc+5ZyKhsPV0kyb5W
bUJcGasph1N0FwtFQnuCHgvHJvF0JLe53RkAuZ60rkx6igCVfDRovmCnCYHeeLWXFUVwCd1mt4ZO
21mn1FmnMBF3X5+Gemhhj+50iFK3fwNxx5CACAnE+73R1VbcX9q3Jiv6OwS2APHzW1BZjQvN4lC2
OXyJfJ3ne20mCjaXAn/CxzuuLvEF+7dTiqwyuGQyuP4ucHaDIbDqziir7FggH9zlBlu4uAf8HAxv
v84Vj1sloKlCCLbtjX6DYL/R3G3zKCA1uQsjLvh4fZ3xohYJAhI+/2N8MvLSKPq2EnMrzlDHmG2z
AHF9wj/MJKMGrOizA9oVQG2k2Vf1nSz9ZaZReRwjsp2jQn2tceZpR9dfoBi00uXiBXdzV2EP4agj
72uCb06ugtvfWcyVhTHCZyqBb5oL4PQvQBFtWCzKsDsRsTPc1zrzGhlx9GdzhxzveV+ABC1DRzH7
v8HrT4kUSswYWU0uZSaMDCEl0nYdHpfz7GeMii4SGRWhCmjiOZ0b4wJAD4s8JANc88QzWpFJs4kO
2Hjy1XjvfgHFMocngFfDV1taLtSUm/+RIbNh7kW/6c4eDHV6ekR8Tq7GQJUEPyyRaPzhlUAA5swS
TVk0OMGWDT+xXxQOyeGB69qtvjhS2214JjJkjPfBGUWb9Qj0Jx/M2kgs1ntfTW2mABbClbAHYh1T
ACS+/7tLaKdkN8K6zSOMDo/xa2bb7xJinUsZ6K5Jo3mFlEUvQsxsC/voYhzEFIaLFr7UZEL/fBFt
LKFJJ0PQewf3SF9IqixR7vmb0DjjWUnVJzHQ04zfSWMIy4nj2CyPwtfBqFC3OwxX8HYcqw981V4Z
5s4FK9yapscDKh/O8MA2IJaCjFFM9LzTcItZ11vYedlsFyY3xPmia8mil/Ea8lNiwP0itfJduRsp
+zcOCZ+qzqYsziylPhdALtmUUryKW4RQUanKLBmDNNBggwymJO8IhaC7Rj/JBMGtT/X2EfKXB5Rd
tVU0G2jEmJKRLLxPEIYhc8dchW6rbFUZxo+8LkC5aIqyU1dRBuxpikPf03RWurIRd2Wn+Vy1KObZ
XJH0fu2GdN9hN3v50kLnPLMXZVIJwD799vlg0bQn8X1m8xpoI8nQFBHeP/KurQTMDSqB1ZRgt0Rc
waQaKP32BbjEynqH0gsJXpfzDPduzivs2sf0JJBzAe1+/SBv0p1ZGBo3boI0fbDv8+tP2BQoaruj
KTiWmhhVijc7k0AYFNAPjFDFrJoRHhK2w/02SR7e7a01DtCExl6GcxD/u6EnUgdmw36p0bYpH+1V
WoauLH1BXHzhd1zbJyC3C37v43+6uAXBgI2eCNcGPv+mOKYYnlDctsTLLjVkTlGvI4vlz4bxncCS
+cezNlNobmxLSphatGrU/ilvEZLykGYF2X5iq+cc56dnNcT1m5EbaH3lLGWwwXzs55Q4uT6L5n3R
A3jLALHxmTBstupweH639K4Qo6VP7NvBsHyQHQ2xCOExmwcBRTA/eZcNJ6f301T2p7FA/uoNaH9U
IDnj1eSJZK082AjEW+1PNvXUn7OAl/Ktdn8feljw6C5X0JLMaf22HBk7XuAPUaCvOHKzhNC55wf1
1aSJ0Xo1oKWjznHOK4K17bG1AZTC9XD8C5uf3xsBVXM5M65fpx2otPMAoncyo5iAT8hytm9A7TpJ
L27MUjUyZwlwosbYydNFfQA4eWhlFYEwAiQ2o3DtEydRS4P2FkKeNiCbCShBc8LoNnb0kD5uSTJm
8fY3ELzxiyTA9MdxVM8ftk54glcJHqrhJkXKU360Uy5tC4ythcMl8UfNz8IK3MNC3ULBDxsApoZU
ru0mC5cYogx+f8SXbceggf0dsC7a3OfPwyItwooGuC65pSpupOl9K+Q4dGra0zUAsFZlhVarM0cd
Kg8A4ydjp3VVhhW8mrnHnhhvPAjw3ToOGdrS8tomA2Htjkgh7isG3KE+vzB2+uW5F+BU3eg07B9P
dP/9j4ZQDw1rq2NFesFTHBShFKdNuYnGe5ixGQavciQK6eVpm9NDBQTXe43rcYf0OQlCDCDaBqZh
VaIH5n3NrzT9/y3XxA0Y3M5MQ+6vQH4gSljc9jtvgrSQWd5CVJCZsjFniaXtK6Ro/sBh55galBRw
yPfIWGHcDl8vZC+Wh4JWM4/5hJ/Lna/wkhp7zt999J7LCCtQhUpchjVAP0zBuxKqU+nTScQ6ESgT
KmC1mJ++w5ANgYoZNFvIwAnlycWSQeokOz2RcrqiYsvLtWjYuf4qAkr8Oz9q8OV5Arly4/GeEwN7
8zVLkan/LZ+atl46nuEpuhlr32mdgWxMfaUb1bJMbBEvvMmEy4lw3gppKwR6gkndItxXnm2uxSPa
aStmESN/SL9PdFpODXPM9UEHH0FU6cFqMtol1sMgqh9tHFsvOA436gjpKG/2Lblso2uPePiSMDgi
0fn1ycf30zUCVYqQv3R42ZSB5rgG+GR6WzBF2fiyAW4IsH3/85gZl/P/oJnn+j6H5wkj0XIeeLzo
kYS/FDZIo6UzyBwRtaBYK2GlS5odmLT4xy4XI+e35ZxHIfMyL+H8j+3C3hsLzIJKZiPhsw4vC1Rg
HxzA4AASRA4u5K3HhCSUi/9TehLGVVYUfUAp87idaLqbmAg8X41SgqtX1vvoqN2bJap2NYAdV4al
1Cks3RZ94107XEuFKvXpWQvdBsAesLwcErTOAmR7EMvNGUABhO5aljAa2NyI+76uz8NCE2jD41+e
AmbtKjadmO0DAhK5N+/WZgehAmjw/PaQrbvhRLxQQs59lZei9MismKpr5pDHxGlAXtd/XuagDYwb
rZCNHHTx6bBrdBHqNMEQ/8vi4PWRP1VZGk162ZfUvEyotfxz/qe/4KwAlW6eGN7Ci5zBzeICVagN
Pf3RssnAAlvly1yoS+vx0GQGSX6f1tkjARWRjZ5yZJGe0Ycj0+j+33FgHxu4uDed5pp+DZG6i8Iu
Xrnw43ghVQIFXoJKhmQlbHAlnSF2TO0uGPGychDPujUnnb0dfC+AEX6AexBImSMM4+6myPfLPH2w
L83zAF4EOZ5EZYMLilZnfSe/jPjdcQ8lMszgByguZdUUTER3SU9rbWw0IztJyIMUPQd8EZp0U23X
xZfTO69AUR93AyMJzzp7MXWPdVIra9cc4tLvzjjL9lcK3E6YNR3oXvyYmdlOK9+HntZeBGGBaVpg
ppkG6pisxzHtqJez+ErWJHIRE89nK5tOFaKAeRZNFc8x1Hh0uYDtB7iV2i54YvjOGW72iyBCAbMQ
41am7sdyfFpldo8LMXmzKpIyv0cdyDM8bu8F1xZGpORMuej4E+Ia2kXtQ42aN+OvUMNPVKySXmX/
RziqkzWl9J49DxT+gznNYGtz4alaeWicvrjMagXYaIQiZvccjKb0Z9jG+mmF+XEgzui86+1tR4x3
N6T/RkWd/ubyJBfQpdrVmHi8T5LQ2g57qh2s8jBZltkDQKLFv8w/tu+bxjLx0MjrtVwrjecvGEbz
x4swD/+3QLBqvbpudcmliMBBdxRDB7HxiPFwgvDwAtm0oCy+vBEGbdt7dQuJdwhuYLfYfdfmATML
wFxl7OcHV5r1cAgEvORasFvRTG8O8YBhk00J6ANilur4Ar2wlcOw5gHtaKsn/GO/UNL5B5y3lfIM
tneNo4t1TgN3Ji9ctq1VIgybWKIL/5Iocecv79JjWczU52cFbrj7STp/5ixKWI89tTHj3QuXXpXC
JUj+AU90/OyUhT6cftko/8w5ABzdf76Xs2PpO2Qa79KOyRl47ct1LGXBsSqVQC0Hdzr+MRSmiWdb
YIpGafqC4p5FQTMwx8DrYGdzdhQTUeIEQiuwbJgBnXQzjhl7TlNU1WG92ZqGtPvDY04lRzO4yjps
yVr2tUl6dMOB/NEY/0zSxHzmyPyFUBVa7K9gg3IWxIoBNpL9a/kkDOnGhTBdc3oSwc/bJPzVkxKs
bjh21Fmee0YaJo5AF8VFAlbdnOf1PPd99yutVhZ7qGY6DWaJ5k8yhPUM0bGa5zKUL6JrBE+Mn/UL
obeWEGjeVfVM8RlsaI4s0UkFhR9DU4UDWroRDeRfzl1vqhUs2NLnDfReqXeQzfAdsd9Mde0gJFE0
cJra92r0q5i2QBeyycnhcldFOFPuSDspCb8g3xte1LfLMIDA/l5257a/p/BdM8BPtrltqULBA/M0
OleIRY6a49tMhwau8x8Jmbdh91X1KCQj6CSEj+lqqZjohn07kP0ZqGp30HZpmHkgqA2s2hDuqfjG
jBx4BTia00KrfPoSbBe5pTxyxUObXDmOJ+tJzqEI/k4BgW+8OteBhMNMuov75BsVFNR33Y7fhj5Q
VsD+ScSoOKOGOUTBrRI4/RvfIkKdSbIPWQNTIIKZvtHxLnOTVEHDR74ss8rJ/wI6Fkqg5tJQjpLS
sQjOMZM98EQwagiJfkIDAaZlhYPVMzGsEgtAkjpo0awQXW7gMOVbXQ683aElVwUmekMoU1vMccvk
jQeGBY3gptjg3IcuUozhJfFDGGKQm9pPtLl6M5u9No04MXs26lUi248RdPxzDdM6p5EFwXY71L9q
jFXW8LiGo+ZkIEAT74YqJKUxb7fTriINszjucKIgVR/c+vBd4g7xbIFxs4ajv54ebKEyeTTmXyS+
Pd+egA/aPfLVyigNP7sOxNxZ2z88Y87J8Tlf3Sqdp/PXvm9/rsjal/Qqy6lXOv2MD4ge7FKWeq2k
LsTEwviN6mEaX6kkszFaWcUod7O7np7SUricHb3y4/iRjnnGN+ecYDUeoBxAYY+uq1M0g6bEgQT3
q1eBrgbl6nKcGfw6RTiaQwbToaIEvm501q+p6QbhupN78lDLvVKWSHjMnmWb/WBcXVhVtju0s/9L
n+DuoO2V67KvkMBcPZqTCu26Lvncb1O1Qr5LAGTHmwLXtdke1t3XvccvdDZylVwCfEwdXcB+kz7K
wRh1mfTgbEQnQmvcftpTf3JqRm4k5P+INHBpirlPXi0TfDJu3a/oTkPBFWDP+NxuPYghpUxe8QZm
feP6seAcKk6t3Yc5rvHOxsJ56AJbt8HQaPzsRibQoDTdUxH8CXP63mD8qJ4JrT79aMijhzZxbGU6
XG6hARlUDuHekUkM/8J+wVVvhjBmvl0d8I9ABeq2Va0CKUiEHGhadnnKH9Ag3pIgc6PWEkd/GnTl
OXE9hKV/7bFlnpBrIgm1edM31Zake6CXbNgEPcMLPyqtVOU9amoHbrWTAO2W/SDvLFuWTOkgi0L+
srXit/3Hmw2EJmSpBPK4guOfvFIgBpiG1Us8s1lpgM6EI0rPik5J6i2/t0EAeIhdNL82QQspJEHC
+0VUsts912jWuCoHSptS5Vt6zhtDM4bnJjZSvQbLsXYh1bdY+2gfO5CZ/Wc0lxi8W+mABztjuVfM
gWGpw6d8FegKnBDYp4RIbFtRSo/XqkRtWpOMENC3dM0XzrF3Q+FyyP5NrIexzkCp8dbUgOuDbiVn
479bAfkzLaIu+U7fiSuyxiZrpGv9k+ImYTNdc9rtJZO98O/S618YCYfuqZPnyDKgFn1WUNHmMqjB
gsc31B/QkcORbRDWjYJUU7zaCFg550GvRIy8tRIykbVJoXpeQctpyosxwyFbyB/NOU/SQlZJy+zw
8+aiZSqBSYypCQcnZ28Qy8Zi3ZCel+5Xi8X84TYrWFEc1LOH4f7iFFKRem78KffKJ0Qb9U+fUDJ4
NTNjWoTfekRDTnwofDUXEm00tM9owecrl/2mg/4yrMfUA22Jf84AbL7K88PTa1UnG78lK3wigI+O
e07KWYoZ3xW6fS39s6MKub8PunFsKIuGAn2TYzx9dVfJw7VnL6yIo2+QObwFaK/LOZC1cnxakdPB
Ekk2aNyOkRjcQ0z79NYpCjFZBFRsk+AxW4PUztDuJqmYK8l4Z8zMXr4a4JrSsgzPnGZM/+Y0D+HD
f9DwzjTZVNSyla40X1MjJM/NVZ+v7/12Ki9ax4zM2vAVCUFdIy3wzVoe579B0fRjkNIuyGkuZJ99
ZhEq5m51phgqFJb6Z4d/XJwd8HGR2zTQwrrOabVerLzpyWEQwqIZ4hwyKSYD/XQNY5eOPZEF1X3T
4XzXfdyaJAvbWWy8NtdLoVtXFRoVCRO26cxaSK/ZXW9zpXpu60r5H1TUvTdq1xD2ZfawljbCGOCX
Mg667o3TABXSvW71Z4mJNeXrAK6/VouCNb4pYiS+KH81ViUqM5qBMQt4f1pxEK/ehdHDFjHIqccW
fLk+VBQSng9ewLDyhCcugDl8gtMA88FpKVU2J4Mlb5a/WhF/tKgy5kAhWy9Ov895WXQd1MBKj286
VnUDl3f1bVFwLUoenHq8M6Vt7OgL35CsepaSf4u7jDMEgxHZ8D3zVcKVm4KG1CFwnjwf5Ml6IRhP
GM0O9lOVo2WhnfeG8m2E7T3bkbo2Ajo64wv+2C1iK8ZSCyo51izAL5Wcz0Fe8xFzpghTg5RqVFdU
RdQV4K44maxzeaM1rKW4qain2Xi02HP0tRqH1dkzUMBxKMym0mr5fULDkU/FwM5zNesgQ4rNG5vt
kCTF+QAXGJfPZqjgUQj/svPpEp2+CA9K8QOJjmMT6tuUehQTvEYMxROS83ycr7EzhJYkgZzaTyNk
ryuwuHs34qoYA6lKqhlYGGUCet3rsiHHWbuLn7pc8SmAaHBryPmYrTY03gpavneZiv7tCbQkN0lo
sg2jHCKyY0b9Al0WV1w3SrWbKwfzkHJ0k7jDo3L/oyAfHYrHkYFF+RdSC1+1ZtgSTba5eV/WW35a
9JpXIe6qrow3TRt18TFPLynkeXq6V+N7nyfbeH5+vEI7ufmmM/TuU/ufqidJWHaxWMsyNKLhA1Me
LiVlrJsu7BJPpA5+fL2UQCUgAWp2wjzZl1BeCE72m5Ol32uECh5idK72qvJvELnnhGYQCZHhYoyX
Q+cPz629jtgx+rrEQ6CStfbVDgfDV782dv35qntlpcNhw0Vofr9mxmkmei2+y68+pX3Ac7glXK/6
sAh6Cr0g+HdDdLhNCuI5SDg0B5wqhiL6ym3YQYDMxJxhOodiWKJOJr/T5HJik018KUOhzPTbthvU
L3DQOOjwZJ7y7eyz0To4uzWPlioHY92wjfnQnB/HsOJ63656PuwhEVaaffkBJ1tuOui802N9yNIN
e6obNV2uLDQ7wIgwLaNN5ca/XzEDMYghBDrrxutl2AIrY3ZYL0MnTkawpww5iMcI61nNhQPNQVqO
EM9bed6CM45f0dMLLHDUaiRs1N2lEvwRoXKSjQZ1gVWgw+qHS6EvKKF0KaJ07h//O9ehzBTEa0rP
EScIEO+iBZZ9iKPN3E8XdkZ5BnBjObLKjEZxFwppEAgizGbzt9J7zC7t8ATxf7vdtjpU30BPyyE+
vGB+uirEzdVAINX1mTqE8AMrd0W69KDqyxb+oq6dGif4+Tch61FiUSyZ/LFn3o9Uq1oYBoYwRqoI
vHQ/oJh/feypBhGG750ygKMc6pgz4W9p3bPKOMW2+IFiJ8tS093NRNcYyyIAnDIz8IHRpT+Mnihd
QljqFGRADNV662IMaabK8IMgJIcrUcQXcCiJAiQM3Rrg2plfXVbAtjx3K47ULMh6oRm8JpKADPvF
qS3Z79EHLDLsS3NHUzY/L3HkhVD6cGO7EzFsS7vBJ4I4Syi5kI9zDyZJAsNNq7lH9bR/7QOhLruD
Cc4bADnPqGN10Nuq7SWqmlKcD+DgPVQgE6eMsKc4bX1zShcmZY/2eixs2x5SOCPV/S4GYYyk+Pt/
LEG7X58sKmTT48pfq4WDM5HWjflMupuKm2X9c8K/Hm72t+zOoIpPSwk2wbPFKoczaD9HveK8rgBw
KHdirnG8Ttxlo8lEQnSK+/tmNU2l/VbStH1JoGN6DjUVO++iFuGa9+V1bzJIjLKhzbPwIxGuUH25
+KK/QnKd26nioF+w+ciyqFE/1FsVADvix3MNi68GXrUmCKg1vZVZQ70mXMVkAK6Pmk0gzOUnblRq
DGRKojTMFNWIu2kohq/rA+H2twgFkI4Mw8WjhqK+V3ZoeqYWgr1ffVE/A5EjFabEhIqOCfrx7v7F
O0fiuBOaXyvZGdEy4qK+5X2ivjrjxUi8CqpdecwKxiV4f3lQCzSsTsgCsCIq/dSKsW2kdxV/Dfzi
CHW+RfEvC3xijvUqSkvBaaJsbToPABiX9/YSCzR9tf4WDXUvyn7GxWtJZLeEv68r513DkEIQxDiN
bq6gxxAy+Ia7FNYQxdFxB/Q6A5iTn5I40XyOscE6cWVkMHOgrhbODkMTaQg8GOtkAQpBI0d4OyNW
SjMpHxmr5Uff5EXdq/GMOnPl7f2ZrUfN+in/7RhcdUZ6dTu+mgarAYhAvbUW0F5CRMgO2YeSBKPx
Xa2d1sQzobgbnu9i+H4RTL/ZhuedO9ltg/xGwhkKu1cT7912WHzfIIWou0na8Pr24OtwMok8/zq0
7yZPTg3XARrm0O1fBy9sTIXRhc8k2p682jaE1uqX3ZuADNdysXXh8YkEtdtd2T3T1igsEjrLATk5
JBqXACL5eIv5l2Hvzl3R4Dzlb0KPA9+TW7ZebJjCNwUDpYYEpL8tLVG8lFj4B+EuAzu++MpHvs8Z
CNQThTvM+zr23Vk21sz65mlBeKMhu9dzf7su4P7shFB/eqel11wmiSQCOXzzJsjKRbpMLCT4mpER
HFWIirhO+yiBGCoZT4VmftnKjEYVgSMtC+NGnyCUu6vj/7U8t6Y2L+8NEdZRkdhBtLVVl24f3m1p
R/ZpbS57J5NwoSk3h931RMiRt/xAltyj2hFCSlqvmUL5cOjDZvIh58LVqiAKcT+saE/KaNrw0pDZ
Bu00oKrP0piEz8f6Z4Y5HoX1C6xfXYYKZIeSVThaNOu0zv/0nrCDbWYuexzO4OaMqsd5h+opd0fi
MiNKa9EhH3NA7RJWWzk/dpR2Nydxo1B2jFPMRVBTXRct/xbtwfX3FJKGbBPg1+X06+SBh75WsNBX
pld2BHhV1rIYe2UXXXxZ0RNQn7vJTDkBUzFLQtpa5JXYyWVaA38JK/gbjfJU3cbc3FZHpe5JRyeZ
shPZWbKSB0OLQWQLesTMFgctqbGIh/iZJ5bTHQrmDVks4EeGCUIsLm+Lcz7fRqElKJfJbqJttYzF
E1T+3uBT8IMsJfEmy1xXD/glCbrvcyAfX8W1X8CGMTeURSY+6r2SEmJ35xQ6j6oIVpK6ES3qC5PQ
zxCyqa0Ooa9i3ySB6YrQPSzY/3OvzYYXm8Gbe4PNVkbzdf7enhvLKPslmNWG8h+zeRs0xe0Zp4Da
CKstp0mmJMil76NdCGejdfZlNgFsvknKtdZhaWjwwVOv8DACaWGXvAb87WOR3+3WdF6YsX2A7O70
a3gJYpy3RO2o2LcPjKb2ggMOzVhqplKCpWq6GvmknmYo/5DdRUg3o61E7q65PpDFfYKEOopsyM4J
naqEj3EDZ0C7n0J6ixDJ4pRxa30jJhXyRoxHLdLKyAPOj7ffbggFZDEGfBysETQwMcW41UZgXnQN
f9qSkD7c514bQRPUmkfzrE1s0xG1jb8JBzG+Yhe4O31ieBPlvXt9W6aX4OEu7AdRbj4E2SSjFwv6
rBSYOtCE4G4FxqurPYnEicJXnmBCL2d4pcGbIu30dSVD3KE5jNbuOxhrCHEgeWCg+mGlAm7uTtz4
S3po36pf3VRdADImR86JGdSST+2ziIJWKlEhcpUnEHonbg56k0HGlxnxJkMzVH6MASt5ygFCcq55
6MRGs5RQhRDft5myuVunoe4YqXLEUp6iCi5/cokXOiJY3wZBS7qhr1hP6Z93x2vwuGRFvCXVxP06
Phjrk/VDSII8ZFxwO3zArOZAfvYp+Nwk/mL/w4rlp38bBod5oYqO9KT7t0h33JkN1Afo5pfer3GV
ZfNCmOcCzADHdCgYIybSLRAuM7fZFWJbWndjkecno9C7YLr1I5wX0O5zQd6CDdOiPHm/zYCGvD7o
5+TJ4jXrLIJzaMkDR9vADnIubpcMaICvuZHDNQwum3tYIIS/o/pit+2DUY503f7ynyVeKQRaALlG
PsqDjQA/KKFbFc43+SIu31sbSl6B6nJolnt1qO2R6F9usiR0aTuWhvRXRrpBlc7lZLRHdd9b2j31
HbCx66RmB6nR7H8qeAtD6Su0Bhljpba+L03uLs7p0iA84/WPMQjRseqOs4NKGLgZvTO8GevvRyOv
+LL4gQBhTLCudkhR9wTZu5sKLZrdcpLrWurqfkZZYTGsa4CFTm6vWTVzjBjUrvc8FoUgfXnoBbdI
JwOVQ0YWpNs7h+X1jCX8zQOz2QIZIv6+kcrD525XjRScbR8wtLnW1P/qKT5KspAOy4tR/Nd+yxCl
/Bnp3NzhuNA7vqfQ5xNutGMhVhIkVRpqCp4OH+clbc+RiPzZSw51orPXSx+pZUcs2l5qvsvb6CR3
EJYTeM88JxCg2mEx1jRt2FPtlJIgS3VwiUPz+BxRX6LfmXpNdiu6+6Drhf64oC3wM7LftfQzREd4
vKzzUucPZx45dRA3fOJiaf4SZsCEj7qt684h4DqvpSnLNtprYT9EbEbUzr9UMYwxgK4udoJqC44D
Jp1u9qTEQFU0Bdo9uE/9LkmqSpXXHnB7PoO9jWSex9qUSrQ0muMihfr8YlxWWGSOZkyoq7JeYSV8
FpRQagzf+GhfRoz7PZeA/JoyGscdf1Fjze33Kp9vWyUAO8KPmwX5N52rPy6AMOKa30aX3A5JZPXU
nulEtnDKho2VT5ZjmwSkIkO42Aul5IbvSP9jzwK2+6gVIqOn5t7Ih7jjLXcj6EAyTlwhiqJyQOjI
zpKYBe7PA5ihheWf1j/0le8m3LDiN4mvhB1slJ0zQAh4FwH11Yfn6rHU+bi4693bi7SzqBHYTCFv
Q3f0/1H3+Z9M0pI8Sm90CDAVkBNLAYPVQHyi+2d8x+OrXKrlaLaH3sD8P5xGWMCNJlP/Fl2WDEGo
GSsihR/X0zNCt+3b3sEIahiKUQa6/3i7qVIQjBfNujG3wgzn3o3ZbRBzB9HRwW9GdcMRznWgjnzV
YkIDJNRq6dDbk4XQIVjXuLeVHglHt9pWWFbdj7wU1cPOodrQrMFdRnGjLiUQ7KlMSDJH4J4QbrD6
bbamwnrFMYHT+vIqkilFNVA9Sp09KOW6U6nUFhRHLR95bwar23uCvmj32AmTB6u5UcqyKyM1TfBr
39cSLtwfW3jVI6AP2pTdM4EOvpURjXNsMrDhjUWJdz0N4YrOXWenk6dxWsQ2u3c9Ge0+JDYHu0Py
n/u2M2S0/y4H1y+f68kq501d7TPHxNOKM9wiXV9O43JNMPlJ36/gqqCPTBt8E07PuSYU6p7OFW0t
QiEiPgpjPAZbp16/gI+Fg6MgJBON4Aml/TIsuIMXlRNfwVpeKDAbB/Kr0Cco1hazJRdyUmRKxtnE
vEoSZbdeMzeSZtqA1+6YuuDeX3Q+WnbxEw6n3s+FMIXFYyZvhR3WF4d+6/xqpoW34gXvCZLjF+VU
VWpUKeQot6KAklOBCkDyZwxkppk22GCHqx+feCXZ5ewZerdXkWOIAFq/0GhCcD1VdU5CNpn6dnpT
/NorTrFxbBi43Rmcob9XfR/gHbCgt0xHVSA7C8txU5axMlxsvLpuL+UDBmQuIIDZ7jDyHwlUyVfH
mQ4+AeRdDeotbA7kBz9lQcKSa2jU5yORDwPesXllw/+5n3B5K1NKcOfXo7TeHO6r3kFPxOxtdk/H
K5thEQaVMhUJ0xiX+Bh1Onw1ziXbJeQY3r9vnrjTFwJgHpU3WZbUEwcLa5UQw98HSsZXURZQ3qBt
lZdvRvfvhhXpySHV99I/y+7DAZDIZxF9XGPbv2QOKF3Zyggv6kGgfGOwjXazhTMt2LePVGVnMY3f
yWyBFMt5RKxRPRIQDOrAmIItPAiEMMj7rJKiFKjrsgRxevULtBga7MtgxuCipF8xtFiV6/iyGyZn
MU07lyzOwHy1Hh0hLBVojSNLXiXzJhkN803ryeYVxlbXVH0WEl74pRctm9xt87a3eBNyfhilFFDZ
2edGzTAD49/U6RLGo6rugYWbHXIF+T03/Au48oNO1HqpdEe4GA58R8wzt91mVeOb7dVftTykyWjS
WTt775JtYtxg35L3xhoWzEBtLb6ZUIbBtPP465+Xt3gCg8cqiHeyEOeudGNkndLqQOAQZdvEN0qr
Hgcq3NDmrIo62ppIDE5tewZKbhyP4gLUNmHuMiBwp10axbUC0Jnn7gc/9PUGAutjoti5tK1wnru2
q6TAXOf54IUkEiQWf381SMWGBLKK238EzLI7UIUOiQn2Cj/TgXjNbsft60tjSFoKj78RmugKxfEQ
RJdNNmMEp7jwQPDksxvjwh1C3rLj/JqC7Nppl6lacHm0flOJZ/mmpiwdtmca/WZz1hk/sFgNMYff
XYEwP7++ekgt6CYn9t0r3bySf2X9jaS9hI7YzdrIh6NPHdtZgnbSPFdm4wx6AGFRabtgQq3xx54b
8LCtj9cTG5SOT2GRsGW9MBN3QuK/w9HHhNPzONhALNy5HsPpUdwLhvrFPAdrBrt4CP/rpW8xca8W
FHVcuFS7BvHU3mAMQXO0fDQYPU8uDsmKwfYPmqoi5eWdpl8f23BzE4+tU5ooTwpjbJNVTID1nC1K
C8U3NaluNVnDbMwyjfkfb0XkcYdsHWIDUos4jJJNly8CF3NDH30w86bE5AxhtZXet9MUqrhbTyBg
DzXIgokYogXkJ62SaW8ikLmO8W9gMcxI9xsXuzUGZDz47egNAGps4i+hzRURrb5Jl7DJekPaYHTs
L7fOBTmihPrVEjHfXnuyL4LpT7JzIevEkzI+WnI+ri0fQf5J4IGCjWfQ3mRQe0L7o6B6TtIgxI1h
TQgzfTJiGFyVTvmgnvDGauFgeIdTVCmkCnyTd9ydQbxX6oTxE9fnIMx3jPv8xfNJX1DF6K3gWcVH
v8G6mswm0cUt0tbA2fkZ5VSo4SzeiU+0qWwCrvf6stVdW3/snWSRCaPIa48IlZ3JauYbYaCcyfa7
CVlkuA99odmaxu9ZUclxZCjYqv+HRp3Yr/xmAlKO41G2lTK85Oxplg3q+p2dgfpzADVXcoddVbWs
JckKhKFZlU67ef5jp+ULRUg4rZ0WbEbOjjiANiJmGMgS53UvPX7NsG5BXzUovHNwQ5APE1+Hbr6N
ty0LI6nZBzRLQd/iNAugmb6QdtRmkblSf97IMpGNVaBrC66KIhFdbgsCt2YzzHd1zE6aF5dvV2RF
iatktOVd7SvhhqrjXbU3F9GsaXMUO1dOPSIfduEOuRlaB8BltrIuX5d/PaqMMbqZ6MezksT7mx9o
Vf/qr092JdumdmtYn2Z4hQS/il2gXFQXmsJ0bYQ/MNONvxlEtSonycuGe7iR+BYxrzLIhPP/ASAA
VgTN/0RJNFZpQjjoDXo466EIdVivWBIO6Geg782Xn5waDwr985pSvxlXEJLhfYg9LPzOqBTl9eXD
FRO9U7fUD0WciOT/vanjAw0DW5OTIjJeK0gP3i6aoZBc5/Fvqs6OTvRz9LZgNQZDcdZ5I9fxR70z
lPsfoiWcX0768aRGpvh9mrnPAfJjGGJ86Qbpmnh0qoWk+9/FqeAUIXh0d+E6GhbGhP0XBzmUQqox
KteG+VzS8p4MHuy6qu4lK8nsI0UET/0sg4borqXlsY4lx+3nfOETjxYNfinHQvJZljNG63ARXwNw
DszG0d4okgB+s9emZi2OBbGwQF30pkWIelKkCxn8OPoWzRJZxbSueBBARIFkC9QO2F0T08aT6tBJ
4DvAmYcJ8EK172PtUA/KeVJiAE5PfP6ytr+9mNCY8EVm3KuG4FMTD8rvJjJFVEls6xyaLAw/4Gz8
WSJew7JXZQeJPHJqSCQJbBZqTMa2HARshsQF7NA7ibsZ4ICPBuWvTXHGJwd6Zwcf2m+nH4N13FFo
toN07L7TdeHYmxXpG5hnCZ1DKfQlDeesYcheQgsOF4uoQhFkOWA8mBJ6i2j05sKbCFRWOvouLaLU
PEMXxTX/EJlsHrHK0lCUnvzLJJSdE1nkiyvfPMl0emRXGVfFYLe7OmCTNEn7vDwxrA4U61VLpwi3
/SjfElRNL2uNSoJ/B1pQYF/+Jarknu4hiynXDsEa/U8Z974xEBc/4iyj89mosDxhkcTDYnIbByVT
LwO3SIQ1HQvDmXKjwIgJIuSWewC/HyOSIubUux59GtBlv3OM6NfcxfnDtZofj2S2YM4emSaFSgt6
+D+IE8H95j8xYCs0xCo+L+xpx9eGFUR2QllG518JG9vBcNmbHPXuXosgvYAnigbfIRYY4B3ehdz3
w8UdqYVM0wUrYIJzI7I+AxXB4T5ByHETOre02XFzzuPG6IXRUZKCZ4wPMgZBXt9v74bVEGksF1Ml
KuOPH3C+A50luYeDe/qB5PcBJWUoL3wIk8/Pnt6eAFVJ5U4Th04QkqfgC92CEcc56rba98Zbs6EE
ZfoZM+6GruH4AiLgPSLXemJNQE1qctYyKA9bPpd77e/v1aWDSxLuHsGCqD86Lq33XCo6WBznhv43
Xsv3RjrBL+03Vv1OG8m3UOarWTBVoMIGvfhNl4SDOSjJ16LvCWtXYqjrMlMO2s3I+eibZOWwDK7Y
QRFV6wuo6KfEUbk7QYaBcwH1kgwlAaH3LO75VDDrGN+YvcVPIRjmM3ucqhetJGmMOAFM9buCik5G
1Wo4Nyhiix7rQyGECzrkBu1pGBkPFg6oiH2eDb62Y6awd+Lg+dr9NGizFdNccDDtr5lV+k2Yt2pT
nVxA0/yvEEgAJhbf1Sq9vjbgttbb1vpQpPOH/xsiD988HuwsTqV3KGCGjBa/PsIsZ3iiqauQorCe
69pjbgfHsxdIIvGzH+9lPRWjglpkofaVkM0p75qq/PZxhApEdr8+OzZafBvJoNETdUet5Mb0csop
r7bx6ZuvGJzXjRi4DonjTDFFz+vXmosAq8NbE1rZ7tur3FGZhtopr7Rkc6P8aESrYla1zlbRb4o3
eLRc1WeIpbrFG26dpoJ1hmtmYzP61VnnnRuo/MEM0vYo5QdefkPnJfyuTw0UmnMDMAMtuC+wOJlN
hAJ8LaATvb7BXDKaiauE1sZ9U/62bUS/1OixMFfkaQXGs2P67IZ7jUC4g4oZGwQvdbFSaPp3HlDq
ZUCmXu1UkohIDYd3Fr2Xpwq9rDNv/0xFFpybfv49Vtryuv+OxPvE++zwPVG54ynANAbUEWiq1neH
1BMfxE0ZhuOGUTd3SAGkBGttuKLI/PyNeYVTh3+SJOC6uF9T/J3NgqCIwyubP09S1gZ315SJ9CNr
gyrUBx4o1C22KCUNU0xqQGK/uOlXMsJofY3OVVnNyPAEqtPRsDUu+MeWvyA6RyZiLjJjE86XMyic
avMM6oCDU0a2+wOcOFqeVlv+LOR093NP1zXGHB9HXIWdbFrlIzZXpB8fdU9ypd+rWm09ZzZpMvJG
34xVDE8PemyHd8aSVPbcBPYRhKaASnkvV++GoeQM34aaWkWJD3LSFwr0ZH/oC0fSbL3uwqSnoks2
iDus8rndrKI6Nh36lfwqOHtTivJ5Q73d441GTcPk/sSR6gWFtdIeK2XM5rK21wB4+Wf70RChu3uN
CnKxdGBFMmQLpD0/nPAJ/OsQSMuJbLALJ9y/YIUIKi1bG6z44ilLqt2A2Tpm3Ha8m6udZ8kE0pi+
QXuKPxHc6xCmWIi+AX8MOMvmD0KFDf2E6HTioCIdPKOuwgb/VTCO91UUDbu2FuTuWAdoUw3u5USO
RHjCCIJadttOQAM8ecyXHJjQiqxaJjJgTrnrQi1hbRNsTAi+XvK05e0925zNDqlCFVnnRdgZ1kcJ
GgGtZwyZIfpgP7hdow20yluHh4ZYoBIpnJdrYqVdQbKVnO5wwFzXwxzYabydcdeEFir/iLrfGC/l
h5iflqw6WxT9XiWJY3Z5m6LJrf6mMJca/3dCbhNUsVU7aldfkJMf4MCg5y42Jz7Nja0bds5uI+6k
unUf3fhYjZsl517FjFVLg85/4HD6s5ta9iaZBw2Wh07KDA/Bii2WdUUaGtFf676bOADUEp2jxKJy
x+Owpu7HY5kgdPp/m7ZC6oM59kcELeXCyHe0qcyaGfiTrUd92MD/ODWba3bCVxNsoarEI3SxPdVw
gkdwQldoGg4FFDsP6S74Aj7z/Oy3b7FWifBWS0sqYpMmPXbZC1iXvfzNOxA9ACFqtSBk6P1AVDR7
jL+mH/VnOjWQFgvmdCfZVYPkurP8/pd4r3zlWPp9vv9fiPMvWcxYYWjsFLOV3SazuqUmyziyOUDN
t8chDNSo+pbSl6JhjQuXmlqU3o1jjlk+53DFnWTTPp8QHZkp4wG4+8WNvOXMpeIWSHSa5h/QQW9d
yhwdFmXUDSuy0kSm/Rc3TYjxc2SV8ciU5LZl+BQrDdPfEUlKTdVFPhFghW7LU0LqU+sUm45nfO9u
V/VFG9zkUiDjCyRUbwmmoDtacfwyXSJJeAg0dbQ4l1KgQxREe3/3lB5Gj21k9eygiKpwJXpYkXd+
oW3qYh2oqwCmvLYeUL/JON1RprbTDqqpHVUn2yQFPDlhbWlTZr00vszqnk7ChxspaHGtKL2fVJ0g
Rpcf6AohXB325cbGxvlki3sp0P7ofStXpwUWedVVHsqC4hc6onV4rjm+V8ld3MgvwJUiUytllH0i
phQJ3OBK3/JEiTEgTXfP2PIQ9KtBs3WwsWB4xgQ3vqL4jqsAoVx/olj/6EZjb3lmuwO67mHtv1NL
7f0hG4EmWZlgMjTdWIlLxBdYbBPJJ2Po1XSR9LhZ41ibsoJ61+jq563IKHOnMJngsoHI5C/guHqz
9LtsbLUbtaaUADsqh127/VAjhWmhFmpom0C6RkTzF80a+L62puo06DihaPHGFbCx82fvA7xAw/gD
gy+cclOvP2l67u23qVF4XHU9o8QYhoPh+axbMJ1SQ5OeOjhEsb5RslqlwOCEFtFttce2Vf1IIz5o
u5nk4X9P+Ts3xwTsD/RApWkHDMJL0yTn+xP7Amn9MF+MHoOrQhzaeA2alnL9OPA6+9Fu9GcpywnR
vcpNX9RfSsC12rw5M0T13Sq2pl2RZ2Mxvv9gm3PHKW6L1/paeIuvaK0HLAMuv3IRngQ92eCcgUzv
hFaf48XxYOSt6hCfI/6DCmFxMcc5qqutePpMvsyHOVif9Gzm3cOJuQXsVMI0eEZGzh+eCxUpjJ7S
3FCIVXJ8+uHcIqes3l9lLy9CDU4AMCzCUG5AYNpZPIcr44vNVxQFSR3SVo8+CbKqJsdjb3RbbLCs
x/Xc1bhW27qawuVqYFGCFdx9XcZicH/ijG/qO9fiY+y/NqX/fUGb//dzqf3Uo6uBGEwjnOTKtyvs
+Q8UUvf2qFrjObMLmzkPBn90n0j1stxNxtjvjnpZDvRJ5aCVqdu4iTeVJtUKgHgkuuNa4nvNkRXC
68IlRTFN3ap5UAQNOHugmzxAWAGFLfPoQlBmxRzJdxZK5l5yLd+LVVUqYaYGC8nru/tzPsBkVCwL
y7GuCbyKh8JnRRiw6lQCChGKDg8gKKW7UA4inGxOju1jLL/A3NhfOIEFHUMWBIH6jrcW9lWbG9jK
hnOXHjCvV5zjzY5RPu2ywxDs11M+g8xLF0O+nKQYFKZiRkfoRqyo+EYz1WplbfUVM8YsLFDl5/oS
E1LaPGkTH0I3b9r2DAoKaN+RHsUug5HqhMwXhR+aSYutn+y1dgNlTRbNEJ7jN9Qy5JmI2V8LS/8e
rdAUFE5VTyvr+5KcFd4QYt88gnZj78g73XETx1FxjnXpcnluSyn5jEYkMoM42P40oc5wplaDFYo4
28uNkaeyLnRntGAsH0QSDXrso86ejq//vHhNs/4UW6gelNFwiVOvebcd8EkHPfDnu+ISzXZ0icHG
QiOWg9AUgJibS6ONF1v3l6JcgXopf310xDqIRGNAy9B4pQDZ8DB4tUyMza56QYofjMrCxHRGMPQj
ET5o1P54tSG0onh0AV8fCJZ2spJtJEPirG0vkVLfQ9HnGK8NhW9+cxRolZne/duGdpidmucgrC+V
zzXGJnAJoj6IaXpGix+377uyYpjT3jbQutzVhJE5wALbm38VEQgytYZP83Fixggj9ye5NLmyPWhW
T/7MopMoeOlrI8btHu3XNzEKjbZbKJ2JxzolRYzEXEOMuve/aTgvkEXE2QZlS/rXc0Uke3xdCluk
9T7HtHGuxjPoOevZqsBgERnYMqIO+Gkmnxnp2+Wpu268n1yapYYJ1qf/Gl8094/8W+6swB7FQ2Vv
z2TCV27ImGHovAamAwYBgSakFmnHj0uz22VBk/+1ZrnAw7dcKx2EWQszkNnUkzoFG2lzGnwi17Ye
P/8Ao+a6ZDMKarOxaot1pzgGyiDZ5/n61Dr6RA21oPp9j9s4z72yX2HUR+N1QMq1BeW2IFe/DRZQ
FGy1Wpj8FSPmyXvakPVuQzXt/oJkxxwID/7bDNViLk4+G06qlW50i4S7QQDKJLrHE6pafigNdvzq
el26VdReSkd0LI95zdA9w+gCKxrYt6zlIPsemedyQIQh4FnrE0+YOUwetA7ENhhvjmnenmWI/p46
+tzbkq8Ip8nE6ywMCJi/AooaZvI7ChOwmiDcW2xjAn8wd2jyRzoiS91D6k0D/wyD4JOKEtpWdN08
RcWznFbTWZPHTkz2ePIb29NVGS43Y5m0mVJtknlnjOxhHyETdhOvZwWOfn98J09DQHVobQqZNZhw
FRhDh03jaCnxYuedT4Be8A8gTu8AeiqWny2Pzw+qEbMxtQ2sQO6VmHTCIYO+2YYvjd4yE6Fgx7q8
Mifxr9qu/4NQK7S0eD+NWzK8PVkrvJzMKHgCCkGQ/DBTXfycl0NZ02qfG0nmVXvb+9n6WZXSMlIi
4zQezf3XGs7JJLmp/8z8KZuZCTqg5nGC2SGUJf4GIglMEW/dq7rXeJThucb2ze97RY24T97bS5yr
jb8tcN5fJNBYHtkv72K0n64zueGzo/mavPrZn+gBK9jgBzGP4wtxUtv4hbk0FmtDRWtmIiKYfnO5
wD28POKPhMQwuTiesFODTUqds7If/8emgVsR5U0b7smdFQvCZzg0g9GLSzrFVsiiF0ekgsO0QFeY
8Xz0m4aMH2kR21Cv8GI7Bcg0LwPGdZCCIM1Q5jlFqoQtwckkhvzR5nAeQc/1WNJEybOu1ILFG0nj
4zAOd8J+rQWLtZJ2lu2sJtY4WdUpdgKjbmQpqAfCbSe7iJRvvUr52OUSNT9o/Nm8/90FofiyniEo
Vr2EPnNqaE1gImxnZOe19veA3x8wfPViJRH7TrPTJs4U5ZtF7tGgfiEOL8tqRPiCUEvobb2fsrAA
SXP2Ilpw1XQk7LTHrsg/Kt1mEKDSobLhDcpG4/FbAsyiqXBao9zF24O8raAec8vUYKT4ht0XMdpQ
byNrEf5U0gD6KWkh01TiiKGi7jW+c0uOs8lLJSJhjssPHuU4N0hhheN2Aw6wx0aX1boOEPW8f28D
8Wggeq1X/VBtZhj1eq+isN0bYGod/LD/A0VcMqsfN4Q0wChnp+s8C+aRTgDJBrCc6lUAtBEvx6VV
GYisCty+iP/GfT5pnJzuSFOZXLif1MyKrG22kf2r9SUvLFp4iVOSyzN7EKmW0jz5x9tOppp7fQGK
RSZSJBuiRteGmXOJnVswM6jyknI37/Tvw1Gxr5iAEIlxnKmNJoUdkBwkgrRC90Wr/xhH10PNIgaL
jbvH9cuaSEMbWzzMinDU+A2Xddfqap2bL+kWnBYos/s4Bv4O7oMRoUBfgbK7zbLdpRxPB2pRnshc
Wt/oAl2hUMyPHXjyrzvnDGsW4F6n1eJ6w/YUDxEzt/qeMzU6z+MD+sKIZn7mjRyDrVe5j+xldVJt
YDfunPU7TvYz8+ha1Sbh56ukbDHMQu0qIjQ4DYbWZfqcMOMxw6fquJHHEvHZPARW57uI9JZ/r5n9
5e9EPh5VvaSSSaC7qriaLcTwDf0c/nBqOmFjK8XHMu0isNx2QNFBypAMhjFe50zYEvf6mz0W3l2x
5nplcNjxmfzhedT6TuxVMQqOa7JLUL6pFDUPs03+CYbV4tUIMzr7PogId+wp9827H1oIqeDjASQ1
CJCu4Tt1v0g8rlQzFVm/7N0uZd1XjMTLiy2OWo+EoQaNv8IrIjStTIySlvgCSQzbYfNbgXArxv2U
+xoU+Ds7jyc8Dw1dCx7xAk3gSoi1SXMqJ8Y/1oM2JUvlbG3KVuPdsvwwrLQDy+eq1+HEV2gXCwiR
ym5Tf0ruuiIgsbeuRINmM4w5Wh77Mh4q8jj5QgArHpwS2QFtuFdMdVsotW5GiDHmxtJIq8csaf3i
KFyjGH4Lwz9FpS0HrUiz9fpQSrWRLNrSjelaFK0IbjkiDiRcKr9ZPNqP8DQX0FktWE6cTGeXVYTX
Axsm7LkyrXLDHsXUEiCeTOw4wUKtBnE5K1uS8qf9HONgsj83ShbAJA2sjXJL5qHK4zT+5Fc+ZpIS
h77reGzN77Jof1O1HcN+OJ0feNw214V3Hoonei0QXJF2kj3AVpt5SK/BH+6GuF77NF2YhkMUeFe0
3yYKyjTFnPqfliTJoa4UxUv+YTDFO/N1Lp8nKep4tKKrB2SN9WIzvQymteAN4snRtSZfdOyxw5Di
sVmETBc3eszzxTJMFR/IqtGDCi8IS6XWHT83IBlg/a/GYl0xwMoNjdR7YYaa5rfnJKDivREsG3sA
ErQo2ViHCotpO4n2yrVNnYbwrUzsleNzJGwGsog90APqJEP5z1gctoiBDJytdsUQEca/VVRkup93
a9BZrTQ6qHseQ1nlTlU0U19aMwLZgZr1ISZphMYZ9hA/3vSLdYW0lGQM4/iJdU0ifVrXezGT53Ip
yIEIU4umIFPOBHhmZvmlLnycGOMMsx7M73XjL24PwJisOwLLB1BlfQcNxA8bqPOepC4qADdz/lpq
6Ry03OIHmsa50yICLgNXUU/SbIJe6zc5IC8k/akS9NUVFbalPsOiLRb+6YDcjhADlDoTu2qeg1pc
YEwHq/jJj5deUgYOP363iN6DW9h9fBBXcliHKs+3nule6B74jFqUtHtvGNcKQFiH7NCn/dx7tN4V
PbRmuWa/S5AdCKh1SBb2c4jt35lRcSwJcfrAoboAISXP7P7Ejyh0HPV1xAPhtLcVj0JVfZ6/V4dX
4pwr6Ww3W233T2wYLRBGtV1O+I+jbcvoZ6ADq26NwcF7O5uyY3bmx4gbotPGneAa7UaTCk0ob9LN
rzB8cTOF4DR2dLtjn/bnLU6esCFDFIDIe+T52nm2Sz7ZedudubI1eRC0HsdGxnNw6sUBqHnZ/yh4
1MUaY/LZBB0a/hRR3gF5nKT0zOT/iC84Day+OTbg8zM+OtwUxgMUr7eAJbhUu8XwhAju15SY0Wz+
wdDWUFHFEBoNPp46wcTj0p6pZhaLKH0hC71ivvWPkHKxq3VZEUnao94HG3d2kLJrBh6GRHZt/GMn
fcRUDxRI8Wh/mBaZVEQJ0XO6f2jIvVXteCoa1DOnJrkW/+HV+8tca3FpLNnK/C8FAG7zKCx4DWC/
YbyfCB6kII4DHXNGBEMCTDi1rrPEdZRYrT04oLXCqUUivUbbVUas7LEIWrgBXqsEME2vyrgpiZ5R
rG9l2QzptB0SrKL2PiFbuBalKy7Ef3CD7RnLnZ0jvxrd1ABL8urWuCCbD9m6cRolJg8xzxgxY56G
qK9aPDNEHclB+oziEg2Rahu3c7eAy0wwKSD9/04+AwKDdyA+8yiFiUWNhx938V1Wp7nEVVRCzN5+
omG1y/NLco00XcYVVBl+/au6ErRtlv33G7LHtSiOp0N/oS11p5OztGgg68sRXsFELNt2c/HVJ/iF
ocPUrv/g9CNl/pvdhMxF8wDMEJQldXlSLItfHOGC2PuZg4kdkhKsJt37EhYNZpAqvzo9HwZb6lCT
nAvsdAgIJ2glpu9NRzOO3ohNTX/BDEoitjxFVNlwA5Vy7hpMzbtLGWq3gCWOCm4g7GNtnEr1YIPE
ZQRyDrjbKY0v9FUbp+oNb+PDbx1dBndCZSQJ/axtZlbEMe8JrVrY0J5mfKG9aJZTw7i898YVeEjD
GHGivhFB4rkNVzYi1ToPw1xvDlw5PlgIvzFGIuWAgmjsZeb84IULwvVboJ7JWlbgyyBt5XVh1lR/
qiK+QAGOTAfQxvfbctIb4Q+bDVAHcEqMzIlNEJmybMNs5A3cDTp+xRtMcBtIW/gklqZGtLukP1l0
HctuUVJpz8JbqqNbktZLsI9UbNB9LK1Bg05ZLVU9FUtp2pjNxRTwep8dXvOl8CFcz1RYwDbWfnkg
hLsWVenSd7IiRfAVltDPJgaaba/ax7Kkpd/7raA8wtQHjuOLlT3CEBEXoykKr04Rv9A0sXbK+ReC
e7wG6C2p4iS94aLVr4d+tit/w5jBoIDmBkd10aidgH170y8ArA1uIrz1deCF4Z4AG+7TvaKbyYMs
UigA4Z7wKOgSFOgqW2foqcF5ggGprDna1+OuZZv6o34OA0tfYJxQ1ZRrhsaCnm//IEWE8iMBch56
xs3YlS1osnAAbZ4lTXiNyEJvx/idscjO9pZ76QFjLxXYFFcGm6dYXgYUpR3WwDfG62gP5dVI/WTb
mto90COwQizCcfTjqefVzf3GHlmQAIXA84+5QR95+mB0Wf2S560kXuAa72ETjcQKGyTx5Ac8epTq
Qy8/SoNeLP8ImauVFLAtGVsHbZlwQ/5nwyTZpUysAC6tT9tVJwDwGmRRTQz8fOEfwtv18QSnFNhe
N2ZiFLGMWpL3AD7vEo2bY8oCI4LABe+376rdSXqSV7jeZhaBvoQ4HSJomFhHaPvy3KEnm0AgKSw9
R446AYj1VTEKtPdOIs75kDomlZxTCTYKQujwiTmF7I/nYiQLyD9ewg9zR2jYzjSYryQMoE2ifEBH
GHw+RDIJpHumw06APHD6XbNut+3T7q1IR2YpJnku3/GIk9JUJVIRWn+ljqNiIDas+n3Qv9ZKB2b1
zvMqR/KF0u5l2OJqsBtuHvMW1azG6/KDxLws1IP3waSNzgDjzpXpFl7cLpZzVOKC8IJznDkRyrzz
NqBav+4lSUHBvTJv0oCLU2QqF7Z4t9Tg8bkweR9k1VQo5BhMnBynbITeAxMM6vSyImYPw8My1rAs
XoW6W0CwvXkaB7dEk+2cm7uW4zkB/lc96bwSrXi7omvM6kMZhQNskbdoFdzVX8u1IbFya+gPyWZk
9wzzvavBnJe8DyixxXGjHwiDQ7F++l+bA5CjZeYPQfr6KuL33s68m9ZpnnUIZjPMjZU9INT5oDMh
lpv6qgSGwkLoLE29Jh8rRxgeF5ZDv3+2vWADC0Nz1l7g/WE8EU4sLFX19SvaZyAuWsTGCwxvcA1g
hFSdIxKS9rFHjkLi3Wa3ik6S/CDmZ4yjKAR6Fz5vTE8nND5Oar/dOc+pcdc875U+EkGd/sgIbmW2
64HKwtifhyecTQXOlAC+d6ndVY5p4KEQzoDWITC4by05g4mUkVattE+mPnxXPl0LrwzvddT+EFv9
2bTDqF7SCqYVOBPKguTF+Xp6qknAF9N5UTh7nR86jW/TCSdfAMJGwMQujT+bk8g5JZtEunRHojHs
gz4Y/ZCAqMSRJ3Xgk/yQSigWiqQvptbIj6ueKJu71BX5Tp9b/WSCwEGvv293F790Nw4g1nQVgNhM
gVwnG9YPAKtFfcnKbEfPZ/hyNqi7fVjHBjU+zeb3BWrOhg8MF9Xf23Abj3BHj0/Pc0ESAsEnvPFA
bvaoFfd8vsIxGZd9SFZMM3Mjd9BtuEpj4zxXePRkpCJJQWRINHA+wc0PmbYnepdJfEhRNqeaCOdp
kV63rowRU7/w5fItEEQmXJ6V8sC0mf3EjnLY37dsQvDyECxOe1zPSYTOFNXYjvBEP62+O/+WBtZT
AbHnPqP/7Gy73VRfAO7yxzOHmVsu8XFUdH4ngq+n8+nwJde9I9fr3BtAm5+sG2g0R8ycs+z4oSo4
RZPiHZGjPF+qpeOayBJAzYokrPQ7JxQKln/quzaE3dxyO9a0OfOfKCC7C+6iwQi89RZH+m5pkBib
jipToZN45IjB+CiumIfql1Det398WIEv3FCppUjZWKUrumy5ofjuqdcBuvPIkqOkW/PPfa/zXk7j
4iF1hgocRK4UP4mK7BHnH6Wz+24BSbzxeDYkF4CEh3yyQnb8G3jY5uIutklLJn9J948xdSkr7Vjt
E1VxkMaxUBnZBcKuPfar7yWmEbFeJlI+mZSCbGEvCU/yyBiX2Mc9RpOWvPhikY/Pef8TI3j72YvW
Jc0Mt84pc72dBr+W9RUqyKQcihK179upe6a2eMe+A4+V8SlnoBg1IxZQLyT/hUe0J3JHV/JxkBl2
C4083pVYZLiTjAWsKLPfpF1xJ78MHffgpnpKzjW4NIYw7SCAgcEjqkBYSXpdEaeFR436gYo7gCGq
kVNN+KB+8i9OGLGfMts1JyOtcZUoHWDn5PX/Y7IRuCqAiZUm5Fv8rfxaISQns1f8vYTb5Zp1YbEy
/gyiRWYZFUIdTPFi1MUUkpTxDcPF7e+D/uC4qIXTb69xwHoUFGa71BW+3G3kgyFGHHhqP85CiC6h
Beb0cvsfv0tZUxPkLy8/nGw3094sxCQX5X8FXBvxUaU0YUqfMOLejy7d4tLs0NL23h404g0D/AF0
KMnFLgekpr8P0GhzAQRcl2zS9SCndBIvTaXw0n0aW5cyybzpMAJaGchtW12+pKhG8LXFaGXWBIw+
p7bCLt2xxpJOVZOawiWBp18m+ZTKJSRL8uWn3q+TLZ4Vh8Pxi8MxilRmLooec4KMIsUMdDc5Z1ZQ
4lAv08qKLQ+saiqgWp4UshvBETdVaKfNhh5LVQGD+pHuXPaeA/Tqmk0xGh4GMkZgBVYv46Wb0MF1
GsyCsHdd967mpzj3d8hzOwL/Aiy2d5KYPf1t4+K/lw7uEaKPAD0UDTwl2mfcvCXAygcyutqWVFxi
NXr1xFGSWd0pX7dPJxKvEOzwDVfwTirdD7+07h6uTnZB2Rud0W0x7Gu8FeItUncEF9Gx+RQ5HNPR
p2dZRR438Bn6PBKEJD2lf1Yq52/czdkYm+H90pH+dzNyd3MRuESjSuVoA0HBCuTLPmV+anvc6lQo
j8U3wH3MA8pdPIwkW2uX7PXEXq0PgxjBEJY1zWnmnGNESU1HA8/bD7/tWHqFJLkEvvV1lLmiODte
c+QomlTYm64TU1TUwIuoFx5zaM3WGhVuXqiUfw1/xcJv/F7C8hBGlMmvcG48ZiQFMR4xviHXHFrR
c1m3RgSeBkAP9gv6gdd4X6Ap4h3tEYUoTMxKZRzE30JA2qHClp24unVmlMMI6W6/WppxgsAoZb5s
7LIm4gZwf4hf03MNq2ZYlJw9SazIDfx9auMJJh8PE1e0Yr/SOw2dQNJfvz0krOXPJEXEA6/eSk5q
Kz6YxcLwqshg3grZl2d1ptt9c1rpFaMRKqYiCF88vm1Ufw3e4xw+w6i4RSFNvvN6flAOzgGi1kFF
fOSkqd38Z69w/L2azB4as5IQKf9VquuCbGku/WgeNfkFS9Hrq0mgYW5crUvaWU2OkXO6aBhfJ7A7
+zTvgifIp4orPbpGXgLu5ESS/D+kc6g1w1Ue/oivTlUx9PkFJb/6RYcHSd1KieJEDei1xFw2iCAO
3I3+Ztw96bg2clw7urrJTXhs3J/sKTvyunG6gG5LyuICh4ypwSgEDokBgnOZbqBlHeK29Rf9+rLr
jyju3aGvAQetvsamMS+ZCwopeFdh+UdHNl5Y6E+FNJDqTCt7+yKQbzFLEYoqnw9juKssPrk4VZhR
oh6BV97W+fAQTSvj7+wjNQnKxFDb3wnTSFlzAtrEeKwpnnvEL9xGZop58Lm3sljSNaYHmg0mOCw9
SGZFmKqRWhi42+/dfxN9TLs7emZU4zfb1tN+2GcUvMR3mouJcUH7o3ttpgjkPz+BaHY2yQyLqlpF
4Oifupl+ViIdhN335TErMLHfM+We9rAoaXUChj0LrpCJTsqHKRHWMFyK1uY15QGs9n2pnU2jHxp4
4NLwYzY7WRyOAYpYke2gVsK83VRHizDdP0Bu5kXf38HvHLAAhL9yFexCwW+ZDsior4MQWxssoTZ1
MnrfkFk+qjEAcM+yR0/a5I5tDqkQ9Av1jbamGxZM/RG1Sz24rolX7wh1431XhWPqm8zBIejdDKGO
YtqYrHPhcZrhvFlkm2Jig4A0DEWktZZGwViueMukgfoS+WDFKysc2NXXZAOBrzYhucYK0PhkZMCL
24f+tV6DTILMcwRC4/ax+8inuKeifopBQspfWZQY8CBlvTzJIqDW83ptEltecwXMkgLG//wBqgGS
k6x8V8RzKpnX5XZO+uNHS9UUC02wCfRcDtzUUk/liB2dJo38s0es075XklEnM9K723MwStHP6BkM
hclJA4jk9uADfpBqunDEhjWvOov6zWXicibWjQ7G78wpu7feXzLDIdhDnEvYQCbNy6yy3MDfsFAe
WEWdadeXhammi3IFyB+kMR/fzxFU9OCoKT+l35QzQ8G3zoq92UXWWfSDvHAPG+Y6mRcLbZIeWui+
2+KJDb8Eji8Fkf5e9FPS+neHJd7oTjPG656c+MGwMTLkyjdkdv2Wi8G12WVgXJBZn4+OtVYNLS08
sGMk8n6jfkHU1EEugAq5B8DUyfcXt4KQrTiRr+B1dkO+uUloKs2peakHLG7dZ4b/nUawFXAZ99bv
ONwzrVy2khSHdGSD2riDLyYLlKbQYFjtgDT4G5PyxV0kcER4HND8PPtT+/W4zXWlfES4Of98UQRX
U8h4IL+TZo929ay4OHiV0ybawggqJT+bQkUpGiyJBg9PAwdjHPB2WZGUR3o0bf7eOzcmzckF9dkM
b7VothCE1mJVOV2fQ8/igsEmFfSUEEKXy594jKPGtk1/FxtPqmIvXRNDGNU8lLk2KNfR5LhpQbV6
HM+A5qCKrUOv0rOe8ovq+38HX7ujU5hqjXjoHhJYW9R1uDr7lvCReblZDgFPMjwbCBwmMewN/i7O
VtDgs7aJKvaAAZdcX4P1Ef5YOs8NlUJb1hwI393Mj7OBjOGZxgBP2twn84rqViu2e8IjL9SQLekl
LLbxff0yn2IyjERrjjjTb+Oo7wKlRxl3kQxIwT+Bs2PsDJW5QzZkgTDtvs3fCYGthmJcm15SD87H
XkKO23BgQeinu9CsP/Y4+Ftdq7bB8vkMPw/sSG/64vDuzK4ldnHzPgALAN5EAlDLqD88O0ar3MKh
crJfq8X4zaA5ttFTDYcDwgrGtkqlWmhGkAt8CwfGWW2cmV/9tJDZX243mRJ6jedwNDwPeuD5MaBT
vogRuQjPNp+hBC4dMLRvfG+X2yTF9RIHXEwmOfCiFWgbi0ESin+L5W9vHc0vl31rsRXILjPzGFbU
N8ptYoDydvI67NwaOAzC7U2DEeZB2yPPrOxIWb7dVNwp9NIHKmolXxkgPpXpOSdk9o3zkx4UhpWH
aBP8KeXA1v/Eej1F8VW00WyZ4GH4ftyXUFr1TqLxOrLz1E8exor3MGOGdGJc+ixpZD/mIX99fvOt
g2qpUXLyX3Lmrbk8Mu+WNY4asJB/tx3OrC8br5pBVsmPPqaFlaEGCaFkQChsvGod0+6HvBbqQqsP
tR8iYV1k56SXYiRTv7QsFjdY8a4NLysiVMiSfDwUNVzN8jq96GXefl87C6kvyNX7KdYRYxEJTtkH
DCjKkcUtNwzRnPVy18miNp3N83/F2oMCwazH0wQOviEdm0z5LNispvrove3ElHvzF0xQErwPggMD
6ZgQdggusgyafmzLqfnf8LpobRgmkkpxoXJwv7LBsWjPy00BKIAyTvOjR1LZAznUn9o3kxQKFOqg
n5y4hd/Y3yOvCqq0qa0A8nrog+5Jf64RdTTggCcVlBq+saHiXiGUY57WWypeCt9DfuG9ZhPe+e5p
6UEZQN19j+KA2vWnVWJPnWeKyn1Isxsc5dmO4yaJgH42vfDHdPzuCw00wDFha+N17oJINHyqm6J/
GsG/AwsaIolggc8LDqtXug71AIayrpnIAjxENfg9Vy510NObpd79lyNZg81oU45PlNr9SR7xI++6
+cp+niIYca4omxC4PeoRPHPbHwFaYJG4IFX8E7FuRF3jTlZcZKPsrcy4SI9Ae4DU3t25LIOI3rAI
vqdZQVKOP8gN+TRSowcPwix9SNmKFVkv26FaMa8mGGmB76ZkmuXsHAQe6TjCN5ZZuYRqScJrj0d4
GZvq0OzApAbOOPBpwBjb+81tZCNuW2wSHzoW++slelEub8WClqv02gHZJTNrv+D1fmHc57ulsN28
Cb5ZvO3DLH3IWSAfyTHIZU6QY9Yg8Cq0r20sPT+ibt4cg59xmKSoXnn+yIJ8lI0Bs1Q4TsUx7HSl
Tq+a+gpTZaStpdoTqFX/wJP11xnvxCvJixMBtxb71KaQVKxls4cNmwGpLrPLwsQVO5qIp3DPNo9v
tnHNZ0NdvUQiwi70nMy94g1na3uO8NwjEgaw96Mk8Ku/D/rktCUGpDXqDnkb1lDG68zNnFI5HY+m
DlaMJS7x3ZmnhBwimAk7Ywfcj2JMSw/513Na5sIzFQBCVpfB3iCbuwagcTZcVIovAOm9f9ks8ogj
sGidqvqnmF+vuaxkMat2f2+Sbu+FyMtAE4f5JQMtstra67mnwVHQ3koESrbeJThGwVwi8W6O4Jdz
4WSLyxfBjt40mGVg0cRo0EHpEb0+X6bvT7Il4PRXnhOphPPxltK5ewoTR9DJvbmqoyBwFGxzESg5
pQapzk/2FJ1CP1gP+jbA3KEj6vHI4jMae6AzmHIGgmkjHEMeaxI2AnAzhgVax9J11mlauwJnYObc
R+iqMcTceTqJk5XF4v3U7TWS7XhRuegBtjnIvH52cNXm45EmHhlRWVWeg7uB067vlwEdUSCTATX3
oVMU9+wG9S2KdsdFr7wbS1RqgV4exlCURgXLkv3kZnPvCXjdQj1PY7Ezfyr0gV7oRj3sRI82TpBr
fkY5Pu2yD7cGMWGdNxXcxZqcV+pCe6zXaFHAKt5OGbiVIbih5YgfXU15Jyu6Ase8cD7/O3hQI2Z1
goVJ8M6ixV/3LlOdf9hjcq635SvS3gibsvVoIGF1qeIOB8Je4RC7RLN9ozOF0fdpJuzcvXc2iqL2
XzqbhkrG9dAP51EBEfuN0YUkzql8g+zhRWbo2HE9mVsaApYOSuMRvgIwJup0zS3Dfg2lJy+Xu6FT
0lNUUAshfCdriuJ2OlMkidGrirzgOC88Fl+8p7x28IYdI3vC3DhXJgWYPvErwdK7Wv+J9atpJNFe
qVznO/3AzEbTTtVEwyMEdyKix91U4Oder94vGOLtcoZI5KdhXjIIVSZqd+pbutCCeCJ+05Dnp8Uj
YAc9Uoha8A1W9SGVIw3eejU9l48L7oZfKjR/uGDgVXneVrQ88+ZsuSPotrO+t8J0HVLAYEx0NMjg
jpG823uEgQsgHwtsFVKHGsizfyzbzWazRborrHbyp8KEruVkcbu8dWe2DbfyxsYaXoZUrlHSP7WR
B2r5h+L9SedexbvR5g4RV9xDSXlIHen1oxBXGViIYd7qV9fn+A+aNl4LgMOLnYmNJRs5ZUPSx8Bw
3lR9sfmKVU/eD4dd4wqguiWA7/NtG2SQxMY+xDlR30Wr0pKBpRUw+XOMv/NJUcoV/+VeIGbVNJXL
aPCIAmBXKxk2VdUf3JskFzMMV4pED70KpCt27KSQQS2qhzUkMwMy81EBYi+9QAfKHeQprPCIPsJG
3k10zc1LzKduocQSHm+VNmiAdUGEwx6zRyN4i6aqEORsiHpi2LxpqYZMdlnwht3o2tP6yax6hLtm
1eqoyQJs7Mpobu7IDgwVOIAljUcI8VpMRg/OdaD5g7xTnDQIxyEK2UIgT0YoKDwHLD58wOloUFTg
kSZBTNnSpyHBipWeLw3tl8pNlhJC1V/Fu+PSRtfTM/XL3QMPfIoX2MvjNMqLIcBM/z/21VkyDaES
zljWp5euDLczsD1jo9roB6pjkf0h97t4c0Fceo+HLvTEVaIUGb86VaK6Wujp/m0qYNsNilh5j5Qp
EjsV4lMtdHxKjfLRpQt0HsmFgceR2+kxQzmVLhoS/iJhlBd2HRqaafKIEMD+lJBl3x6fPI+ZZDbs
W9vveE64TDqUBffBbQl5mjmK+mgroJPRtNfyWsTawz7UWQWbTsu1+E2xxlfFWVIkWbVEqTmZI6tZ
HAJMj0A6BvXlgRms9xQyFrcBP9AqYs+ldVP9WOPh4YilPbCHE6Er3GYFulhvAKRupFKihLxjkvOA
bjfmWty0GuRWabdF4z1AF3j0tZ0gMv+kJAaqpqXChQsk6qHlVQc5qryAnw3KQEb2ufKkgm2ib+Di
esyd4Ib2GSethamf9Gsy3QPnRsB14XWu1jD6a8XCUC5AH7EZrodnidxRmieJ6hv0DmUEefpbC72w
nYSZahGF8YeIApOHrNRfu1HmWvwvYEELoS3TOCipX7FAO0MEtudUx/0QFmAvzxtjojrA0/cnSOlT
zGwKaNuxJ9kBxqESjika8uy3F0242ezyCm/EOTWmtGfPDqa/5xvglDxJ65pmmRpQz6Kl1SwZQEbW
DKt+0DqqElrmXst/WcQm7VsIM9WMv6bsV8irXtRsvK+/mXq9+DFcmJNpAgxOjm7m6giSBwcTRMb1
Kl1K7ljw/GFSWk20GymrC0hXLnysHZgWiRWrxJEvGxaQLyMIBS9bKpY2BnesSafuixllP7tBxP2t
HnD3QlufaQ22jNAwIhDtwGkYxwdH1ayyAzMp3jB0GYxGJp/uatWhsdgsKXBn5JsCe2oaNd5mOJat
tcoLOzTiEzAbLx1rqeOMlFaVOp7xX3Z4G6sIEhwFlXfVl/8OUNiroQSOYK1PEkXdqc8ste2r6V9W
jkbJzXv5yewCTEWgtwd1COtHKbQ9IqokVaVl9cfs01hH4bW9/krjLdUKU3cTqUWpIMUqyCQH++1H
uyCeJ7dED8zFY1yaPQfQo4idXx+3rjroLHUEiLjVBW/mZT4oO2RXAbkBpQoD35mCiXZIjwcyetIW
ist1K8Yq4SyqOxavHR/VbJGHiGlkjO2n82OJdr6VHilrSIhIyZhQ+lMlxy0tVxi5Bz+75HE5KjVJ
1mqMTox03WEW/3F49I14Uvsn1yCl2aDi0XHTmSUfLr6qhMoHrzdPcfDG8HuPvj16hpF/OhXavWVM
ZKFXHpK9Y4ENGSoxIMtrKLYTvkjhNE8x5FLY1HdjBJKA/sRdcOIsJ5TAML2o2wKOR1wDN4y/fuyW
w+VvA/yigNhwJvRi8HlQN8bg3dvMu433EqxDGlzBwuyt9mIFqFCo57poVNYdYxTNgKvh6Orzs853
vYBsllwIS4cIfaVpeS1A4A8IYnpr5YbHhooAR3W2SdaqMvl5g8gA6iBBXoQ9P6iAfe/BUu+0C+Q6
xy+1yikq37PQeQ/X2K1eDnL4iqDHTbXaZO1g3HtoMaKNAQhbOnyOTfMRGGvb2O6cQvM/bTVPtsAB
50hO5MU4u1DzUBaao+lAo2vZ2oOvzTleYrIPH23EPbuBVEa15LaXAoyR6x5I4U58dWAHXW55cywp
GcT0PXh85XyMtjIUaz3K+sC03dWrRZTf2PfkX8j5GFrw0J2ePQVRooJcHcdgIcQt0fQV6E77jD7y
Mf9CDdF3RgDS+I7n28k3AzTlUqZEh2UtgsuFIvoFhTSOyJgao611KBGcwvOoZqOdrTDXT7VTUKDs
Cfdvd4W7HAjsMFZaJWTF/f+P+MndUL6/fWZt5caMMorNMbCIH0NTMPcqIlUy32VnW68M7XMWTLfU
Lh0sFCaYP0Rs6LHur29CDSopIU0Rxc74qWhMq9ZNZ4vDpinS0X1Du4SRDgNnWNRCzNx1UonuohTX
Cx0zqyi77jCGVaBD6l9nAG/HnF+mLh7t3rVgjq+8FwBiwyuKBVjZe/P1VXTwsGM0P1nF1yX9Gc+6
h/I1r44RzJNWsVoVB1FBoqi+yGYCnJTsWmbWVtgTRqM7LWFDJfQh1/61HgjHDy5/m6aE6W0iMI16
qKKwYxmpoM5vge9NoQn5OCfwiulCecmu7rYd5HI0F41WxjhqyTxxsU4SYUU+cWu0A9ecEEL35/dC
nqEDcZkY2inMCSweC5Hnmz8Jdu/ez/zZgMyFWLPJTCFBAWrK+J+pN1DCQJe+mIeJsolX3m+gNWk7
7DmYIcjivQ70WqvzOhgdSbRUHXkVmUH25g6wu+wzU0SB2H2xmSMPsICGo/qG5xmKtQ6OaAco33Wp
W+cuVDJcWekL/uE1BS1Xq6yjhvQvRFUlbdIrVu5ahwmagEG+XflASSCUxiWcx2nO28CdIssCWYCQ
0WPYekEwYVxt9DmpnT9Wog32679FWDp67ZoU+EdBNGZig2Fko/yz3p5Vwxxd3PwqxMYDeqH+k8q7
phjfnMC/iLFxioCoDz2Xrj5PZpp+i5Ky8/LvVbprXk2AyCmhQo+qbwk/ztdP7sdF0YrnlNtYyEMI
hMK26cC03LoOUEaIFK+wjW6w7znvI2AsQLLpp/BAxSVM/3p6vHACeVNk2770ouWwdMe75LEboswd
M6sK14181D5L156wOg+h+LsEZdcY37YXWogtByVEmk8fOTzSGDCjbEoQBdX1FkXWJrPAW6rjOCws
3bDX1UWh7KDv5pV/lxCEB+SY9daEDTJCjxKrCMaFEpYO2e2tf3IlnASU742xv0CCgK1i585tGHtr
Lvy7sXPzBd2LnbsRcTK+e7txUHNzvXLacip77+6penKxXmJpDog+efMdCmtW+tfvgfdaDK4JFQZQ
7c6zpsW9pHKxUN+1lMKqlSKMqKARcoXNQjJwswizNNNpDyxlsUiZZEzQ4lGbboy4d8K9tOb0jiT3
VC+121GkmqwcR3v1fcojnyFTi7nh9YBWLt+wycDhmVuUnqPcMYXkDp0j8urIjPSlN5VN+tz6QSlo
JlNBT/q/a9kLm7VSPWEOh1dCHlACTgaWNY+K7rhh5/XUod2nBpE27izbUudbsuxQD6No4fEAiK5w
Z59EZ6lb6qoxIGLvv/o2YHjy+z+2AP4qry7S30hZaBvs8CDN0jJAo5JOfe276uTG67GrWR1Oe/5T
hE/P2mx4dsE2Y+CsLKFfXNRYXoOeDX2vDgzra89v+NgDSLeM1817fm7Lcr137D1zP8v/11dp/y3C
orU7p5eT0jS1zA1CP4ccNXf7ZrqIxNZCLRwCEC/2qBKFSUJRYDC5LaM91v5CnPflRYgoKVRPbFpL
YeJHU2hPOxlXRqL4VKbmCZ9YR4MirIL2QJiBze9lE0Y3M7kaNRo+DOyV07eF2ZW6+vp6L7kuTvBa
8AWYLstZk7bHu/f/krdpDQ0wP667NBSSIiJ+gDyoirxd9Wzn4ifQuaPdFmstkNgY/RszHvyMnzoM
mHK6P2PhHzoL0EFW96x+8AQkJPB7DP0YS8b1cP0Pfnm/lXdxRPHbVSTqvC/LLA25L2db6kR8PaJQ
szrU+/n9WkQRKEoeiyKyyq9uWWHrbMMhUxIqF+7hhDuqfe1xCvksI2kr52toZiEPDKsg99dBjfvr
OmFgn2wXiD6KNjjNQ1M2USnI55m8yM8NlPcZusnuAhEXg9yI8PG8RGaECv71EXPAM5wI0dDGM3OT
Tvl0CKRkyW8ijBSOFzvModf821vsGJZ4LT1WAoW7DJnpU8mkOIiy+8YDTWYy1uQXQ8cGGV3n7puh
7n9hV09nyFNXPWpXjhdsqMzP+VtjF7uzwy1i6mJIAIDH/bNsjw/dj26XSd7xAXkDsZRvUq2LUCpg
UUbDTVpADaFGWyaMJKYDBI/owy6j1TNmTu+7a6+MCGzia+1TVosOPNLg6KeF064cFBySuSRjLCTy
GCXJ7hOMWZeHdLXEIHkidvLym36NxzmlFfVdgqvtPQ8Qj4TMLIPwGd9Hdfc1o1/RGt9YFF52zdQD
fPh+LI2iAT5La0aUnPSYrr5GU7EsHWb8itbOZnxQQeuSxUh2bMU618+lAfYjqvhWPUeRatIwYPFx
q1/rsGuq7ldiHxgGqY9xBsjSrYZQ6HBpjJAn0jTr7vP8aYMnLotGCRPLBBbjuEsKKsY5jI/wXQCC
r9JSPSdHJOrESLksPuGAUxQrI9+m3yAoM1ZvI8q1LElvZI3BAxu/1z2drpRiLDZwwrBThnZV2b0n
WmJvBVM4bZDt+osPIyk/N3Kknzd9ZeSqVizIv8c0zU/j/ak5NozkO2Cl3kCa364KrFwNeOaqibIs
Nop7w0XErOHVfo8XXSEB/VpCvVvKbcNoh8HVms5g7CP5Hbr1xh7mRspM5kSMXArux6h09YE1sdpG
cQxltakWNSRMy7yaPjbQFJcm+O0kBry024T8X5ZBDubYtGsQN/wkdgtVG376XaJEjbiBBvhC+rdx
fHeGn62Cfmt2N3IKLakOSqGeIWYxtLQdQwWhwu2kPxHew4TfXIWXe/H1l6MZkZHh+iW8ymjzmU+k
qSBp52fTGmXfQSTUHDa4Y7XOkFNODeKfQCg6B+y/iouQvKA4+VFgBTOjevE5DBIcE+BNggLW4j9b
ifH4CJR3v5HzxbQLpHfwvkBcafYolWGHMOCKqWsty9Lk5TxKl8Xu9kj7rtDH+aHmnfWP8NsUBODG
TY4/pTCah6iwHNAfJhb+p+iv9pUZcXV74VsnNhi0kOpQ+c/wlP59sVmYrJe2mDh1g59PnnORzW8x
+GHyEe2M6/NddbFquxhQdFwuz6GY83tyhJnEDvrxwI/ZF5jA9gZz+zaOYSFmhPcc4iHfTdoOG2Pf
Pr2SXeHhGNLChc2mhfUp5dNxGgPVv2EjDLoWc4xd4TN/Ku/tQF3PUB2uMBWaKUDmBY/jF0MGcsy3
A54aavirlye8nZ2zMcOLLcZrfcTZuGYbcDQaSll2loIW3rkBYt2mvsPf9MXa+anu1J+gb+8qs2vr
aM55nS+WSybfiqSBhmTwim1aqZkfEx2P/zcTCp3Cfrf+/ovRVqkywhzdE/hqsXpQ0qDGDpny3sPr
SJXb01FMx8CnNz2izA+IaIjGsaEweJFatIap2eJcHEFFMi09ScSWMRFkZg/kR/VDvfUJ1BfcH/ds
nIpYgytWOYxNGsZU/YxLHNZEUivKjXAlKIKkJQF2tF6GS6Hwb30uIixazmyxKxVvdGjB6J0ialxL
1TQKVkTnlgatJ+DsnU10P7Fk9pyos/tSHOjJLPb0/YmyCx+f3tpnaB4n2V/4BJ3fx0fiUbWCTTX2
CmI0G13f1SiiaWYYDORogMf8m1gTW7OSKFIdn83g2DrbWsOYGF7aAfhQqzrI7yqsQgCopFG4SBdu
a2Fc3yR5UhXItZVasAxDLP722UdgH8v129fe2KjP6gjxOgzPZC1ueGt/v/6p3RBNsCfouyZ+LL3U
99rQWSVNhT9t9TGHJpckKFZ+V2+yxnfGhIDa+NMJMxsSSu0ZrnMrQaZOB6dryodHMcngzxW6f04g
WavasXJNCum5HCJD8eIXG9jNWxgL1e1Qpo6rulOk04o+Tdy7mQectLm6fFphtLmPwDruzToSrbuw
1OeCMdo57mXWcdkvr4Q0MQYlybb9CcBZG8WDAfzPdcCN8JpHaA1JSCp3iEdok/GnQg27QPfOTUkm
6AFQ/scWLuXpWeissB6/zTamBTc7olyHBTLh4OhkxOMr3d46r976Mq115np4TDVTuUdn2AxujU9h
QgCjS4a3ldkaeiBTjwcIYFIVJl/N5LYEpCfOhGCQhP/yJZreUrUkPMjpWC3XZUTYsfueH8IylpSC
MU+306CYtZceCkDQFSyg4AIa8YjZpPxEdQAn9ZunC+BjoXmjMsFNGbF+3wIAb3rFEem10i+DJDdk
58XxhdiEesvJ7kruZQvhHso326Eyr2yjvoU/kNFZarAP0I38mQzVzOdyBEUgTAZO0gGj6kQz3q7e
wpJiXagohufENK00/9PC/rbVhSUMrGSbnt1xsUU5iZuSpbT2C9V7ZnIW4q0cQMcW1oES7JyAaioL
W2fsITwRH1NlvR+zD8keHKFB53GonQfOaNJg6uQQ48Mb/NCncllpvEDv2kyHt1WPi3kDXA6eF/kv
WWwXMhlBvphDmlBsKEN23IuVN7yVAKuqe5+2GIjmz/zlWE9/oAjGqQH6zQwndWJ4fh+5rVim0vNO
hgjPSAt5ubVUF4gK6tntgTzBcv5xLQBEoy6ZYHyY7p+gfHWaFcfoVdfUw8ZCUaaALnF0usPjdwdF
QagGD2rdpAWFRhVXXkwgdty1Fi8ypEQLdr3s6uiBaIvHUn/ci2mDJnVJuQePVMcvZAAlSDUrXQ21
oJDsNOZAKlS1IlOHIomATG+dIYPt8ST+De3/hYsD3pQpLtuzwJWHvFFEQ8yqXQMZgiA5/9lLNasT
b5UmmbOi/Ofp3byZATRZsIDqdESNA+sg7QlLs/2nZxtRFSyT2RUO7Y+J9aJugvzSlwCiIWPQ1rZA
/mXpUklmghHDYgZL0jJq9z5ay6eSkQg7IcWAK+0R5uLtR5aCk+ACHG9IIwuyGzZ1udKdFSKcFY6w
qFds7nG/i/1bX6SVq7e3kBuc0uHvYTfouQpAoTNLoXGxsn5cDE/Isagd3cmozj339xk+SCC862eF
svcxCLeNi1N8zZic+Ntp9xwaDexxmcxqh7BRiia3I8mh/oI+Qi8XUlw2EokR0r2sRoVGoAZSYBl/
izBEtTifG4amkJhVc0qYZz7ciM0sc8fHxwjOZO13QKc0w16M3IjzmL+4+mlPibWt8SpzSQeNkZp7
YVXmUv89unr/aWRWWl94ilzU0DE7EU2XbkFcuT9zxNY09x+AkHdbjwARELAJThhL4MQdMp9919Fc
qMlItNZSGe0WU4bUPRWTJHxsvVcMMx2+rEaD/4VIPgjEzIN7/bPESETqrWDRc5S7koyW/jZpGM8Q
qySqm6kfzO2oMywwFggcBqWCqA8YBXXX2qdurFFlbJ5I4XS4MLuemH35JIs4h61kbEP4Ws3IruJr
b79Po/iw46jxWNdQHAMlpHDI5dzKMIJgIZmI0iwxfg9q6eYdgh61wQ8gA/3gSEVbBusEvMcEDhb/
7DYJIa00x2THAuIPYhdF3LS+KJT4EuzkqDM7t8bNaJ3RiwZe7EvIqap9Cd6sbk6ioHq0PrmUmOT4
uYHCPFDAeioRS5kvoLomdK0oSLkd+THg0T8KYNPSqa/sObpCkat8U6tuvz4e7GWUoXii9mnkui5q
CtQod906CfUGXYiMDEhFms5C52KrT/wZxJm2Bx3+Z8NhqNHyOIncbwRvj4K+Jm4EtE4TXMKzjIxR
tdXP+GyMV+LO3OMtA9eW7xu4mIRDLzdc7o6MCfTc2+xROwk0tk+KM0sBYncQ7mr3VkwAOS89aYAd
2rutBY8tbNCTkyI4A8+J+o5t2kXYUav5Tz6q+NVUHPY507xFKkJX4NhddgICCt5JKKunPQWLFiBQ
FSoCfVffR2Jxlrs+7WnN2Fez3D9cEwifNSdgg3GdB9mkRpEtbzs++MHyGJJoMpJJzLeaGkbrZANo
2FIPIN83jLwuEk6sVXpPtGGVKgAyxheGpay9PUtAGg3R7e08jEQFq79x/KAspckrr42QhuCJOPBN
tkgLNfCTAvGrPfAiN3WCAfp69e4620D1g02Eo6ncjb5GCNCzsr9sIZZv6o05QxuE1z23OsmTN67W
dnqB0mg6U6lzWeI2mUsHLdlfziWGVOaNmxbIGsjlgpVCbu5e4bbT2mbRn+FEZynMA1g6k7ed8fcD
WYoJA4xnwwrRG8vduEz9Hf2Q+D0DHtvjmz84x8wG3LQot2aln+UnjKIQfYhGLOJZXy4nNND7JRM+
gHHmNOf94CG4J+O+JxqjJnMz6f2xeDIHjOzf05LuCoov7fhZ52MitTlzjkfzFTAnonYGS1rfTX58
kWp/Y5F6CwlaPbYH4yf9J3Ok0grZYwZn8GDOHsg9fOcJSLH7vuRZNeSKmirLAcw23DqsbfRkWCtS
F0SoGTBPnCoO0gH0z55kCLyuaowZcg1gLxem/0W5PnYBpNN5Ju8ZrR/ZPoI4LSOzzxkpSJuBohBA
gUueiULTthPY8lZEWwtOVtSojmQWA7BoYIS6nMVij88jOA/xKqQXcmFs9HLvXZuJmiUlRhVqLEGV
TdADb5/EuwQl5eWuk0iKrBIr8Za7yKIekBbqMCE9dz8SHE4O1PY//t1L9XQvcjiwy7ZDf8yTcxcG
3OOhFzlfv9yb/FaUA5l+POTlWgg/jZvrlm5ZrCA7Qaj4LHREzvFInb786TCQsSa/SlOVyDKFVNyk
SdIcs5Pah7yz2A02ZBjScY05461hKygCAxm5auRXsO36WiFasJPCuyIOPr7PYbwv/4wFzRzn6MDa
MwZRQ1zpCYEvqMlICh3kCbsS9ivpQOi1e2LSHRcuGCP7sWcNumScqasjfMRg6apRQMUGL/KAYtdI
r974G+5xFKnWfIy9giw9T7QBMUtcLnY4S4X6+zF6kSSqYyhfQNlH7Ecfv7hajfrJTOpnYqCImYvI
LdbaT03EwoIqJOUnUMt2oEOo5Tf3VBkSEqOtr7SgisDSu9ZcC/3C/JZZ2Zl6pa2QfvLbcxlmul0H
M4jvMxCrNB3x5z8Q7viEVoc868RDWf4aRX/YHGDx0J6duLoBBqmz+iuA3QqbN8mtW0ckD1tdehvR
SdqpmMRw1dQV2hzefkjzYne1vGYbifzw35iZQPlWu9wDwCpo//YuVUhVFLgR4ZQOi+jcI1H4cGio
SEDfNgFJHY4ZXCj1I7bUZQttWgWUR6Or4UKTiw0c5H3fgvlPimviThystDuHTc4+MPhf40WVr+3/
hqs/yFMUKxGGCO4Et34edWoskdeBqiMKWCA88ivkKPPWM9S17UtSwK024p0mCNEEpC0RequwLqre
JfarEYzYcWrbZImg2aDqKAMCGI6nC2pYYYYk+e6rW7FDM5kQqdX1NEiL0qg2FCLJUlbd9VVzX0Lm
+113a2LDW6e2CFNlmgOCDnDkMRG9T6KApc2UG3TdiAA/nkFDGQc06lRyo+O1Sa8Mc1NI4MMIL3lP
JfAELV5R8iV2RWo/mHj0gY7eWT2DImAk7Q3XbBbscM+dklh5LzJZrouEaLomqr1K+nb2bKv/OJUV
zi6ZahwF+JsdwNZGo4cHfejs2m+947/X8s7d8wHkIznXdDQaHC3DATBCGYpYMQDgaDm7AgmG0UbH
zXKISPQyppAJrDQtMzr8jzrzXMqbVgSKgIP37lnqf4NEd3TN6f+lQOGNzyhxmLCuWt2VrNTMZN/B
pu/Z7q/z14n02VUnBvdaD5+v3nptThXaUeS17QswVSS+ZAtaSqjMKRh4Hx4M6xBD14s1znyd0vXc
3Z9WG+MZWzbm4LaqpvkMHx0OWrLZJdC8GYDsmf7CuJXJwP/AcU93Bk1yWZEgqEK9bGWCPhoG9sek
J6Tt/aRYKtlze3yu7uqlaPzA5LGoTln3rQ7GmDnqO984dN9KRrriOmgO+sQYneuvRIypjmEV5gKD
nzTcQnMhgv2jewdcKI/w/HK7K0oq5tORj4WJf+0XtN+Zm/+GH+M6bRbxMwPxT5vpuomauJq/GuvD
IEENN2z+DdiJtmL63SZMXWh+4RWEoeeU79vmPG8tXqROWhLiX96OkJQEiz1ng/4kfMcFeyo5Arms
O/X+62NbGjB3sk8ahBgtH+FCmknfKQcYYaR1b8jquOeznYqyzzmlpo85y7wWPTRKkqIeycl67I8z
IdsuUVphp20UNavBgh6ESRfQuspSLJ+7lCwiRaVy5ybe7zw2ccVWaKhZH7XpLnoqwt/zdeaJN5vU
b5u9XBEPyrCmGUU2nxNB79sBeBCfqLPdnMtIF/+TbaiGC1rCrLbL4Z/3fVb/A/eH9d9G4n0UevEo
vSGiMHmxFkiu9JngOSif1T0YHXgmRNHWGaVOyFUqz7ub/YkHvbRVcJbZ69SpdgMKH6QUDNNVTCzV
hXUsLyNYUWgmOgrc5img1cK1TMeG7WnNe4F/irT/QRVx44aFf3OvUddMwbSFp3VfOIQ7V5CHTthm
9nW/JHelKJ2n3E4YTXtjyPkEaLp+rYFdE7I4fiY4PxhZuwujnUxFMR3ICipoxW4XN+dR9X7EmCZx
8ErQvj+BCpVjNugoTrNCi1Wsy6NxuSsKqe5Hu0Nr2sf6lZlDaT1GbqVBz78rGIMaBXwnKHWk4x+J
ahUzk0+caYcx8wSxFU1TpaQThH/37MY+VvyNs2hyYtDqrrp/JBqM56Uu+fRlUY0xYJ4gDsGGGVGf
sHDblSTr4G4FG4R8kfaxgWrtU3aandEg2E+VamVvXQbgLfWkZ2AkzwWLSf9EetbIGQb7YX7thxjT
o9hMlsO1leEUNTPGG1hp4n0V6H7R/6N4IXd1zlJqxugOwn+zmKy5f7hu69ECufRZkre/Jt2jyFFv
qqHSr7I8ZJaqnuIZ+1gS/6NR7fPY0YuRUMJt7QHd0NL46UK41hJgwaglPXvf6xQHWAQC1hnUiqjw
NH5jX3NqevedUWQd4A02Dy/h2ucX8HR5lRdKJMs/e5KE2nTmXyg/hnk9/8nvAK6aQMR1QLUFKumi
NHC3mAWydym+Oy8R9tdlZ5y5IKobmSVKb6FtmoVTA33oMcC/0TDZ/qLD2KlYW4iObSoZAYleCZ6a
uY4Fe7LLI1CHNq3diMtLxKXgJXfngNKY5u7TSy38gxU2nJJ8ABUi+ZJNcSyVEXi4zplqti5x9zau
XVWmwsn8JLG9cf6N8ZhQ//JHdQWue3ZFA1+HfV9rkQ0h6h64ZYK3ZFVMHtqifeQp6m8NyPLPHbNe
HiHlCpQpnAoSE/oMSzLjCKslcqZKFqy09aRXyCXjcqd33Pd+yoONEkXGBNf8eFXlHnhlZjJuyTDg
6JHo6O+am8H+OE31VcnP8POkxOE4tKaKqLfQ978zYKTlWU9TlIug9HQaL9lTkrDUc0y1vO4aolpE
Ef7lXx4y0ttBsJTbM4ocRydRbEZ5tEieN7WHYF/pa+GFu4vK3T8ETkDT07kITZh6e7b1scb5UCeC
bhRSrmGyl9ycip+dxNJF37ZDb6yx2uBAoWLNjgsH1Bf99ai/BmW85OmDs07wurtDtjvcGAfilbKM
GG5QZ+T5yMuKZhthgQWW6IsO0NCPRAXmt8nk24QIscTUKp4b60bGbkkA0fgPJdOhtHuwr7GxgQEo
lruM1j6bzXBB/RemcxA2EqzpfXCSEc5Mop5w6T4guDJnzG6UNqTT87Y4qHxnq6MhlcriqQCYStWk
yFBe20UrQjLllq4ltxd0a7g++RZY015g8aHiBtIaNojvBBce2LqwKmLh939ySMAtY3U1a+oIUb7z
BZF0jIKWBL63m4O3zwbjRfzRhMiIb2zxn11SBDbmXlpQCDT6T6yHx2RtUFV1/bulTqxEFTU2g0kG
EQwH4diYATj2snz0Q3L3juOcSiStA0tiFrtxnGKMlFOPlXucMjAKj5+lL76t3pdCVnSH+/lLH0bk
uyFcWUkXvY+OrNa3NmTiRpldDK+pYjXmUq3wOt41L7a2P4M/WgJ3FtrzJd/Tjt1tZSNzYnYp8DdQ
pudiimBO3jE+dkg0zzB0OcOWxJK10fSy0/qu2uyQ44psctoE66z86693qgQCH0WRYLtPS+Nc06p8
bP9gCUv9xp5gJTZhx1x4DlrTrHPUiyTAv6m+UpgcRG02tmPNLC9ADNnNihA1p0d9kUygWMV6wmNA
3RBmCJRaFWj7kbz8p0Ff/yx5pmQcGtjhwRqZXdNaPHC6OQlxUsU+EUhVwQH/IEkBDznW9/+P5jSd
JzZ4XFnehcQj05b+MG1n3+OKx9dnv0j94gU0SFB1ZKGLB4IQ3m7lHWJ95yz6dvI2WxhNytf1tG3e
cwqfTEEVfyti47CfsUglxfti3oau53qaa4mbKFFBhFwWaoZKQOQNlPHP2QjX4hZ1vZIibG1NnkFr
HAfrXURbTGoCF3j45vby6KJDLIZI/Zqfd/CnsBGr2sgRHHljREF5Wlc9Ta01iCEcCDwk6E+MgAsB
fQ8qCVmmx8ggt9ppkFbWpGatAYK0h82DsHp/9yypvy5BYOEfjHxSpnc96pn5C6luazoHQQdVPAHd
PpHHfRrdQzrp1eIFHI7dRJDHUBMZWnab7gvUcXhRiFTiQEnqXM54VonTZ9x9JrQs8OPziGr1ncle
m4sn9dZgJtDWY+kUBHAmJtpZSb4H9om+Gpj2eXin3HckQBDeCAgMhECR9gnLaUavzGWT0Npb7o3Y
gP7RnJE3VkXeO1GSiPFwtay/NyaXu9R+rRyppzkHW5WfmLuyymPjLoMIKB558MNDpvf/u84iDhuY
nd01SAJ3pBtAGv8WwWzhQxatpuR95E+d8gRh8d1JvUAxkmeq7NuOGGawftWT4mQTVCc0Pz2vGBxE
TVUPsrcWVXyEtpZI9ykKb967C9FN8e93uYqqe3h9Zp7FJ0RnJBg1OHaYnEe6ov0+66x39zfWd1kX
wS6SJFow5NY4w/ecKlLdLCXqYIw+C/JN1GhNOT0UbraCfNPj/9s6pitl9VHveLqzW/3nq3dhYYfi
XKWxgI+9+kXS9S21QVSOH6T1hzBU2i3LnJpq6DmXofuNZqGsJ/PTMOs00AmH9IZ869LV1z2U2brG
ZfhioQx44WtvgQvJBL3TJ0PXvcn8/ZjTm2EtrbL7zte9FpL4eSoja/c4fdl7VfY/muhVg48Tct3v
YTPVQGF0elxtlJqdubmmluP/U6BP29qV3jlGplzHPMLQAK4sDQdaLFVu8O5Bkv+nbFQfkNPjKvpG
UIk3Nssr31t7TOOpQe+1EaNQIaHh4enlkAcPx+Wj5kh22mGkiAdUW2Sj6fEw+TDl6p3L9Aperyau
nrwIEMvHtQgzLcH4PvUxeloIJxiJLLjOyasaAj0IDAnbNLHQog0ZyuCqVF8AB4JU6ygCg8ijyCbX
fCIVg1L6YOhFkAZ60yFDo61JBvlEl2avufFUCuZPKo9x6UJdYP6geufcKLleDwVFuCakb+f7ivQ2
BR4QFEamRjQqMzyOwZkfCLjt9VmyA7BRN7isirSd2bL8/eR35eCvNuQ9wbQm9bc7r8hH28ytzdWp
ufXQvmNEV0dayXBAJqFJl6NB5zbhTTDE4dFRSbPWHoAsVraj5VNRRutRStPG/kWTtnvtOIVk1zWU
i97uBqQf10gOyDKfsK7hQvZ0eYIhWGzQOQAeIlXzFXI9LvBPMP3ut5ukMULWQDMfo7iIkk1fXpD8
sQtnajWJEFZVOvxV3WLuzyElHmOCJTz0eqyPxdngudtZNLrgXWuA4gWZgBCZxwqan+2BgearI+U8
qVJW/UeKOKUfGaQgvsyJGeFrNF/HlWSzWJN2SaTTWYAAi7e6HpKvVWAAByfUuzxTg+T2TWDAQieb
+fMRDf93HYu2t+ORG9H6H5taA0G1PjwFBrF5FldzMG4pQSIP0SLD6vSkPG69ON0O50eNJ3AS138x
og/LuRCklHKHVidPNEcUZBtyFypM7I9MON/d14dZPtg+MEzhCTQNX7QBCAglnLk7ve6qGsrQ1o/C
U4tEezpSTpUATiEAvIblrVQ0ql411x/duGp2vpHQ9G+McRGQyNRiSM/k7j/ggKs/noWCF9Fsbtr2
cM8jedqeUtHxpf4/1bnNuuQzHrcfzkuYsDhfc9mNXZMolZjJe1xDzlKNXmJLis4Ts0Ubn7Z5nFDB
cTIuy3t15+MIw59GmI9UmmMXkS+FV7rA9yB3BpW3NKTy3xKtMQEcZz3hH+mNeIh+lRu2/v6v+M9J
WfwP3emWbHlNDTdb1k78aTjNR76CTGuOKH8KFL/WZQSezEYe4KbvpXbpezS78+aA+1Qm649ajWZe
7rpxJbc1X7gezVp9eqbAhNkaR9heXjq7VK4UB4YtvYiMa/XJWjBCoaesZ/Jocm9I1+rbyv0zvYOc
XbimQmAjP2/dIawdePgerIGwBP3Z1Pgo4DAIolaZfqR20jtU2ZC2gHNjiT4qKhFrBXzpB0rO+Ux9
+k1xkZbgcee73+XB7BqyfxHsdEQHitbtF13jy6vGiG+ja62VnStuXlIZY56Ty4QJDozu2ZzH5LXH
JYPlE5LlrZSnEUvUGGzgAdDMrUjlM2gD26JpG+GcY5tQskQiMJdw4ttVk55wDa0pnEG7JlCEnj3A
VrCnnWpfiD1HBgcWevDRrEYIPQkiaxs6ZjL1IeW7/7sTNmkOHWyfsoMhCy1vyeYIeH6q2nGW5KFR
A9FUSVKyhjQ4s7xIEr6tSropg1YgCbGxs8eZld3Wb2m65ofywv4J+VAbjGvZOJMJzIriad73iuSE
jzAaNZS6iNmNEuUkPAReUsmOMkYNnF88XZ0GXiDXSxgRccG2ycguUP2w2cVNP1WwxGbAJtGNpoUx
lkq8z+S5k24BCZsngpO+FUen3QXsTqe4LFmo+TKsvWZnhn9t1B7OsXAKvhFQgo91QYhDBBELk1xO
WgpqxtWFpBBmDahhnbfuR1MCzmrHJ1fwa5zYTS4OUhXp8/j10bNeUdH57Vr1GLd9XNeu0TwGlKq7
/0GIE37kGl+vqlZikY9v+FIyBkLSH4pNctrPtu92oHk7M0v3xAf/1+La0nRFx+5R0vXjLksTE7AL
XoicpCp+sgtaz/b9HxeM+jJ+Umevi3wFuFz15S4m5WgCBGKyWxwDwpys3xZdRMY98v8Z4rxWHqh+
BiC8eZY5tERnwGk5DYDpq09OfX5xBcMvgXa28Nlu007BMgLkMVqEI9xjVf81w3i//E7NNGiNjlSK
sne+4rufhjM5E/Qa4osROoRBqDCLibBreQJgIwUbMf3rT9dzH3ycsJsmEmJBt/KDBY8Sd4LypzEW
hXhGn9r7kbqvK40BE+0vwZX0m218zPObwtjzdWxR2+1u8cpcJXkThqSTKYc0zMGoyINDIScoz/tT
8OjFF+EvSfmpkTWmHCdvoL+9rj6Dy5yS6GhHxmAwL6jCxJns+YIX7Yx3xECakxZ6Js/3X94vAiWt
0ruGu0FB9tKpauql1BD8Q/CewVd6roIFpyeXHR+0LH+gx9bhZWoWh37JpnS+vTIloAfttrqHy75L
S98oY3UVgqWCnkLayyr3ktd8cIkHk7XWY92Yy6Zy9I7HBKmZnHi19tieL1WSs3x2jvQcF1YNHwVK
zN1PM5X+T17WyxW9LulRYsxL7dZ2iihFRQmq2wpQvZ7Bl7kaFZurf+aDSdpmXGXe3b9q23sL41jN
QSx+7uLInuQw3TRoPgSCUvbZILPY1MZZ0vcUy9ypLUMzGq9j+VfdKZ911byrUOO29E3VgAkRUqMn
C3Wf84OvMs8svskHDMouWg9SZUrR5A2axcg5/fZZyMRbQ3+a2WSD+P8Un0PRN8QG9ygQLotEXa73
QLresH9AsYQLqCBaYogs3Fn8xew1R9yeiaQ+Fw16RjywkVHu9ZLWPD79OWaqAzxCD4cqIYR9nfK1
gMFfrLY2SZ0Ll0iT3VF2ARvvwSwtyTqUux246Whitfhxup9t2hu+CEJ12WmslYHnFxWWNsvzlNzI
knSkioZ++nT98sPWouYFhYuOiPm3D5qzSHKndJKxqvj1iu/Ga/1zFpWSD/JJBXipCNZueSAQmSWe
y/D5vF/qpGnBDXJlJYkReum5QM7iokcmn2Nd+EBFbeXl1tZb0FrWZkIYPgtoxNXyfiVvzlPQS2ta
jhe3GCIbE2h4vE8aatP4GXGmoTmBtbV93opGF/uy05DROB+qGeSNdfSJglYLHLKfY6x/FYvUgwrq
OhCx02Uf2/wUI2fkLq36VDb17Y+j4tGTGQyPiQ6KQ+OsL+jivp5yVAFVsu1TskVzB0bEekCKtp6j
kAAFu8epFbMg2OE+I1tz58sIBiZv5eTnoHsRLsxhGjIXiBJH/vnVPN7+krJazyDUEbprjquevnEZ
cK08SIUrsVstn5bjni65/tZ8TNvnQl65diLjHYBh2Jij9jKMQLopN9p1qCVfXTH8NC2uLoDwuFbF
lerBCxZBhNVURRA+1uiVvrwmSI/fBLnp2NOQV+si2LkZil7Qj1Fc8jpkzhzII9qC9WrMdPeA1zPq
kK6ZSwpAwBFuekoPWESNQoHSCvOWjbvpAn8CRL1sIYTUyCCsYOc7GZDwL3nZ94UhtUHRMWze5Ncq
4/gMzESZCnooCyw6TBUO4A9GFR2uf5sNkn4Cqo9MrJmOCWkRuy0Wdwk1NwXxyW+10fA4VSvFwrQ0
Go7QW7LHF048rBhDsobHx4NbZ0waEpO3oQ+yhlok5gP/deYPxK9quHpwZ23Cv/KRbgGKHL9tdMWL
rgW2baktHuQfaigKcgLnUwpmy7xaeQejv6IBPVK8hvGxLwANF/3JJ9L6G02bzGjun/3ovH+kwlVz
rDT3gP574VwkBlKeNEcbRN0EcyxZmbEWB3OCkxr//YpOp6D9ak0E+69x4kCfYLYhlxQqQ0x3w14c
+BxxizldDLuGaHnAcTAZpT7qz789rP0vv5GJL1qPI03i/UK87gIN5vtgg9w7FxsBvs3arQnYlA0l
+2Q0F/5sZ9/WZmv4Ka4HbsaARAC1MiQu3R4YSUB4snnSh3Z4lTKx22Wj+x126t5XVAURsQzhUUGG
nynWTZaTxA23Tjsj54tpkLyEXtUIaeVEYhwRMDkV/R1w/4ADIYghqZdrNSeEoEKAqX1wW3Xj7RL0
sXDIMqdOtx70NTuiWsXiLNeDU3UUSm0mWWZnawB8lz0rUu6Xe1yMQOtYFfip6GNfjehdpZ/O2lDy
8hqNYml8/6O5cHVmIGKzFLul4WwvWs3lT+9clbbFO+dy+xWDTI62uVPqgGTWF7cdh+6/E404p75E
t8YNC/zV/0CbbA6RkLXYvqU2j/712JjR1dFbuP6aoIC/dGKp9pt4XP6pkt4ld1Qmj7bTPF+U+ih5
mu1Lvpz97dWeLiSKdcThhje0Zg60yYGMjdSDQtSyWGr8I2KBc0KCuNOvqATFoSdCHVKeunZpB6dZ
+6u1rhO+FRjTYBc0xGb333qsn/I2jbo0Uic5hj6VQL2hBd6i9U3ln5Bbxl9pC4XLMrFHvwt5c6S0
WAupPltN1aJDMmDavEFYIObtWaLBASKlQvnw8vCHJVXZVHUKG0J1+Uw5ibeD8gMv372EReWYMQ0o
csmUQhb/Qr/hoZpbgoDOpyEYNVaW/X9s/wh5cGE02oYS3H21YULmSSmoII2WBJ+ILjXJOeHbqJrD
N1+vUHOorYrJ1bm3TVmj/AIEpi9tETo+oLdQ18wzmv5czDFCo5CEdt/I9v+UMOF2/BOpR4eRhkjV
9Ygc2L70H8LKgPR8dzK5HQUmQmH4bjC0/Z0MgooBvJD0dncs/wxVa3PyEtzy56Ok81/Py5QsbQo+
7OSDdl+4eFzHutCiDy8j7TZ/icaHe+bh+WCvPqlJ9I+4MjnGuTJeZ/IzF3uxOstPCZFDsBvUl+tt
hX5LifByHCeGIrKcrjwQ8aljvySQVp/uDNBwIugQ0bU6hDT1fscaF0gQJQLwUpQ2d0GTs3eCg4hJ
XQFKk1h0jmmDI2E+ziQq8w8aAEjTmVnzPWm+01xlQ/cYsMu5fhSF5VeNbrg37HoIcQiVYNiOUwLK
OeolgdCO23fJBpV3PXJQtBS4mP2NOh0OPVu6ogBOaXbiR+5stvr9zlnkHy534RCJgRWvsl5evJu/
Oe/4pxgHAy8Vo+fD1hHfzED3G3JnxMn9+4NXOGdVaXDRlG9dmX+qnBg+1sSwq2EOj/bMeMTD8QZV
O2qe+4LJYd3SKNpN+gn2zmFTV/8g/u8mVQXvrL87Zp5ZOSJ23cfhi8JPtW1S/Zzphm5+15ildOwP
KUEk80LuCCjI0OWUJJfNAx029Mjd45BYOH0853DqrDDqoTY79GOk5b/We9tyOdm/P5W3sLQxdD46
ybpuXk/uiNmhImW1AfeSeJ7aPuUrQl/0QJwr22pYtAjRWrA2WIGie0zjzIwP7FGGYk+M3TMKnOpq
5uYfXemF+s12J/HQcP25VxqQFejv0C3+5sGKuM1YIZR/oh3EIxgY7MZ7L/4A1GIyCU3pIN6dYwbe
qiE4sOdH/MtRa/ao9QtieaRO9QT8hosApgnS94hIUBXJdu1eBquWx8TnHY6+CDLSAX4E/64He3/k
PrY9TvbNa2PHqjYv/vtJbx1Kck1n597a1ScDPCRi7x+S3mQHPrj9ZLDVS8olykznrOQuSPgPuvpw
Puc6VF0wicMtJZac3dmLrBWt2CF2+2RvKN15azKkfVBHVPaiRPUfH7MDGCHXaBzaJWyHgbS5VOCP
E428FBYB/t50ZeVJzOle7evMp95d9wpoCW6Eh/FvIAKVWljPcPPdo4/VtSPwT1ACELU//I8fZacF
ZXrIkquS2i1yMBxDHSy2+mVR70qDVbGJL0eFOmc615os8nglHA31sWeniOynMEwC/CS1bS9fId2C
aUzMOtdHts2K7fa3i2CeW2YgoIDKtt+oUs9/uMpRC+elXnzhdkwLJ0Zd0w3lMJpokgqi0cnVYLjR
k+C+iqxZPcxsIN0V3jmU8dKASLlC1j6RhK+/xBnHj6ttLWia54Q4gzoWU+2EPjQ3xIi9HZiy4nzR
HP89skbeYbBghpnRepYWrvL52D+DHT0V7f3g02KKxnMrjtGjqT+HeJUFGcdTxTgil59uuhJ4VVZ7
RMMAhZv2LwsW1ShQaV/zRspoh4qPpEjcn0k0NxEM4yhNdZSQjdJFCdvbhAapY4Fm+VSwYJkq/XtQ
fC1Qj5qr+yyObs66KueQ1BT2d6jFyX6AQMjq2DWImezFLUJ54qjELtH/hVM6LzGH+LL/lNXGiEgY
NDTi4WzPtEDDJgBtCFx35ApeGuUIF8qEJozwQoq1M8MyvibegrMRpEPSzp8aesaNsOkLSe03Phio
mUpsNSgbNkoXbl0EEZT8Pfy/DG1k4vFoUKB/lKOYy2VjU+D/scerBP7HOs0BybbKvep6xzCx42RA
6KxQYbwrlIDRkqNNmSslgH1AYtmBkxq+jYdScJt63HXqHIovoRX2uE2kaU+uUZdtFs+HSgIznBPE
fqvX5NFqGbzTJlH2LEEQC/ApKXsOQriB7x92uvQQEdJNGijVkMbbuKBnQAfx5kXFw5w0vN+fUjSN
mcatnqO74ZcZ+M2+SeMBm4ze0GP8tlJ3pP1QVq9OCejhqCJyQ4e0scsjvrQW8zKSqcOTU74Dfwy1
LQhH4Z6U9al715oz0XgLGtItCaOn0i4MzamG/b38c+ZcMqSdjoPbkTdEtFmLN3AtqPl1LJBsB/kS
Nf3oFR1BVSJmMHL3XFosbGUtKpzElKwQEr3tro0EmwqTocIwTu+5Jk380rGxoezfYll+rOPICBvi
LFvvM8nQKOCBsjzVVktDzWGc2cljvOjT52PNaGScfLg4e5WVYf6TvUyGiEkvlGF7V0UY+AcbMQvN
3w1lmy2WwlmGuFtURawd1mnY0uZsF8d36u5Y0xrkoBdBeup1lZ6icZLruwwpU2O8CnRXHXs68HRX
wHL08MfChnAL+sS0Cv7nCRmIl+FsmLVU6XDCCEHukbtgJUtfriOCvOL2SYBD7WXUP11iyJctZCod
eTgy/wDC4R2XXqyIt0JJB8XS/awv+ecXVROsr1GFlZDfQaQA/jRaFyZF5S8ZTSORy6VUFvo1M1ZS
avbhcN/LJmbNSViMgCetQwqwwq4VXMFNgUOw8/A7ubxu248pNjskkUXKIxNl6AL9h3WxCQthRGN5
7Yu6zik4HR0iNdWWU2Z3tifHRWFoGN/YerOGNlIcyHmA74Xw2RnwliTAAhb5MTteu3MaBWaCl7xv
7Dp1+Jp+8Vjz/Wm060PbCdz0weqNXiuvnt4qznP9jTQcmueqOHIdd8o2kQAzCcmLX5U9wFg8rXg/
BdY8xASBDEfevPM/ERW4j1PXlmAqV8qcbrvzOm2DeCGDIXfwCut6af4lvvUaBKJSyrm5Zddp67M1
R84fKlNdwRiZdxG20Uwyai6z0zMcUA7WSMytmJ8/hH34kq5qVnVk2xvfK9uDPuyNfQdfVWU7Vldv
qzLPKVgqq1sOc8cZcpB/bzFO9mCPWc4W/rXyitAqv2ZevYj6OV8DhGXUxsOIOYKbvqwkhPWu6u3C
pubRHGEzjFcrLi/vcY/WTydmJE3WKbP6ULZU/AQoM75sLZ0rJX2I40G6KDiO2eNXSYCkvSnEFkSB
vrEx8dQWswk9UxJu5VX7Oy+KkQwM6py9Y4OJFAPPt7Udmcbnlgpmpvhf54yyPGKmXMRHgEVfR6Yi
cc7EVfdRGVUuR515JhzmlSdxWsAFBcEScCIk9e/hAnAeAl/px7cXZOjTlVha0NeOEh9SkTkLH+4J
EgBjJ2OZY2QCYQx0sl66OaXr0BV6OK+TfMEnWyXS+ogXDqj/Qpcec+9mH0GvkHfbmUTPY6Rxgm1w
VDwzhqBo2xThmd5BdC+aPMBElErL71mM90JhzQ3GTOA/yaCtIO6BPxxPlWpsD8ePzx4YvfzL+RKN
6SOZJ9hFio75qtBOOpl6X4gOhxTYeapvHF4m9izJKEvyROfIh3iN/QFGFqQm5aizL/hkA/VrHh8+
f4v/QI6b5lCeUQBpyPV1ya+PKLDLMuO/ThkosXchH16c6+R7SBAYvJLEv2obQl4U9HhFJD5CU5D0
hmaqAFb/+6r3yV0yHcdv0MhypgGfu65M3LQplnAaElIiSDRqen7FCJJIJnz4O+ugKhR/sZnAWK2p
3am3FhgJ4Y6Bi61Cm1jBmkpy7QW92ISO/26/0SwBEFOX6p93vBx6dM12T+DOwPEEBA0sDW7tVp1V
265PLa/qtOViqFKWSTFGGHlo1prsIYILxZzxEDDfSj7p7FKV/FUxDkIjnot35iy2q7B0+YP78PcC
lgr07oA05BW0gs17A6dCAllglEzbWy1GTdavYekPLjVB3yX6UArX851Bfg1KKEYAXoCF90Iw4KiA
Uq0q5WpHP4Rrtjr5bC+lZq3J7mq89dDG1RYPJV4pjQ9wMPUS9lSdBZiXOmPpM08Ymai/D9S0N85A
l3Sfrld716sIFWa6tKiLq44i+1AZv1JBKn64sHLZjzyca2AxWjHqLIEuhBXyDdEe/ulfZqd3FaXV
0awXL533P677Y6/vEAUtvl9pabLU9iFvLK6HROwHZlK03+I6uvxanwd2eUJWOkKDSzhty8Sq5JgX
iqDqxgYT01GATL9dBKYb/jGnyDSxHHNoqLTw69jREw0AHf0XM3DQ8ugSJRxR3+eYoQA7qgR1ehes
+cshrIqEHPlMin7+yEJzvnOBjqG0DLRevHdMbPzEyh49ASohmmZIEdbcYFPRDNmNdGfALkpEgZsV
nwlL2ufhTy687lv5REOmPN8IMyPPj5Vbd+b8r2jQUaoGnlQlVRFDNkNFm8CqDY5WT9l7W3vDLr1u
loETWk7HUQv3v7G/c6RJcz5T9434msRwEdQN3IHutNsDMo0h/cpa4T3LoDDqXoLAyrSDahK+nJZr
bd3i/QPFIiU1FZX46TzNFj13bBBGg/BPdg+lxBtzokEosKU8Nvrgp6a3jZD7Rhju2u97Oap66Hja
1OrjVXgXcH16p1BgOqAf+Z02fQk7SXevL7YYceclfUytnvTGwbZYCmC6buf0m59LY0oyGxHH9OrG
ICKXP0W83gLihsvqLPb4XsKpIx1cDGXZIHV/GOvQshlFNR1RzSS444UbW4WdT+ME9ic4MjP7ii4+
KbYSlq8aJJA5eALECKOCLNEXCA4MTyiHgmS50Om5nv5hPIH75bSOC+KDVSfbgZZGut0QbUtMAHsE
xkjajIUq2Okb1cAm1aAbtNRqN3NFf6evCmreFYtYzb5sTnkERkNJ8PEh3dabpvMwcAK0/kygVGO2
g23Thuf8yp+1+qcLultiTffjN1Pxp+1JyaidMb80ZqbIPVN+i+c/nbx3tMQe12x8md5V//U4022I
RPlIRQgJtajEPe4/QLolBHUHKDqemWEFJ6YzXGtIMXPCyHMz4FQ2QVv5yjLs+YykR6MlQi8cpwTZ
l43Ru6/g0zMD0HClh6ioEnCric3kY+5L5S88+3mIZGt8HkOBj6uDVj0y5thj9zu8qWsL8f14YDLr
Q9esnjSlDd16y2Ips1ZMyEz5EnXrC9rJxxQxyAhDPLou0crQ9YlUy6EwPPyeCl0O71NayIKYu3Q2
6zx5whMpIU0qMw7VqS2njJ8HDLULZ9FFr2iIsRKXaLeRu8uhDaGC15xT3bCJAgb+4+Z9NYKmQ7uv
5YM+ZgooeSF5LHZLNQsIMFkju9gHu9SNGTcpQZuLyPpZfhhKLrnZMc2me0WyWII3MduEm26JteBN
HPmovVSO+KRtTY9ZSLvvFtU9wynsCUNj+OyXOJ6F2zOsPCXel+80pmiN0vVHklvL6CU1RiW+QpFA
1gGVNZgCsuxQNmJTZESlBldexkIymWAMhG8OXV4DXVynkfJ1pSBZtGR8JiCi8kf6Umu+fL2y6tkW
dv48cHjd1Yi6jCqXmu/6G3V2Y1tqEZn512uy6y+O6/Ihkjf4qnzK192kjEGa79EkrFgaynmIP6K/
QWvsGp8BkD5qj++OXQnEcXuREK/1itBEw8/XuMtN8NNnIJgyj1W9YScLWAR5Mw7DmTLwyCfhFDar
n08PBFErvxxsJ552ertE04U+DQnEkUciFfOlztllkYQug2OQANnuL2ZZjTP8CSBDz/ePpKRkIGkE
O5ohXvCp32Huw+bCAQevydEB42N5OrvQ6wPoBsf0u9pRQ4INlwbQYEDyUB3DqkgQirQAEk+1QWwN
aXhILmutc96L635E7Q5ZshcwNMt7qQYDohu7VsVs+pTxEt+vmVFIqfU4nAo0u+k28UZOVMjFpOjz
wYPtpPFz0nNqh/h89Hr3cr/bZ8IgXNzo6nrmvLeK/cg/jw+wGNZKU8cgGlmNZVdZeDbo1EPBCLwf
YpKKnQUc1tsPKrJ0Cz+9YDq0o/OcIYdoP1WTA8LDoOjV7l34ixciSVQPhkfwnFkuV+KEYqn8fS0a
GA4yNs5KQXrQq6u0sUYKxBlW9jYrQUoX/KN7J5kTt9VrlVWJqEnd0avvzK7znoBuUQGO6B4dZoGt
30s2+swXvj5zPJeRS4as9C/uxEio8n314msugh62IlHBNAJggshK3QsuiqPtj/zSrTzuMOjuYcoB
tX4n7+siJ89Kk8zLdSTrj0h5i/4WRdgIltKa4HOy/9Uf19mE1jlGuU0zOgs8tWBuLgCa+6Fb4VfI
PkkCXCAA1H4GU6oHpEOSdwDEHJOB8V2m23RXdOc/CiHwDenfDjGzvxIq6LAJOlbZxtQeZCTelt0j
S7N9K+ACpESe5+M6WOZdRuDYm0B0IbVqjolGoC8ipd41KaGxdRRaRnHkS3FFqzs1WANmDIH161bH
TTM0xmkOqiEYGfhgJpzO28r8UduqFZDflFfoMABx96Sz6WakqIiYjcx3jbLqyvFrj0pvWZv6y41t
voRrZcQT7nTssMaMz3RCO5ZQl4L0zefFD1IapoaDT8BAPB1V/hChUIw/4qm4Im3TM7nNgNhi2ezS
ALNnueL9DbcTVW8nvf1tkPQXLuglWGh68U4gNl0gzb3ctg5/Ksr9LEVkeZBREwg1mjluPB29mKJs
0gaRcoPzHd5YiblaXqOdc0xZjfxKWkH3HNB13zlN7N1TPOlrUYwgmm+npz/Njubk0uZ0M+LGVJVu
kJSr+CS3zPosliqIK87vrW8DBoPICwPOsLYzCHsTqhhkrVep60R3KPkAvMmr/UsJuM2lUJ4kFsza
EBw5Kj3DwqcPSNphc3NpOXxs2XtX0ENkfyOL3WJYXozs+h1SnSikaD/8BiUnMCawNBIQ+VorPv7w
hGsH+Nc+vu1UsT1wCQqsOM6SfrKnj/xQ27irbS/LB3TdgJyYPFM0NUNOYN1QKzx/VON5R70eC3vq
42Sk4AGe2s8YLCXMUxgbzEfoeWdFXcV68UglHyl+qsptMyC+IIeXiWdq1HW4nRnFHtJaUdud1rFu
2IkNVW9iMsIp0kddtMzB2+R22DmNUWCZh2fD1ePVVmdxCCL2SJ1ZltcQgH+UL16StSElWghJ08XN
TPPszOtkvram9U+lm5b8pcrkANz5oMExYcPR7KCe0bTYbRiOE/8nhRCOKTDIXctGwIPx8B8A6tyu
eF6hVlG9XfqN+MZE+NDoN0PfxnfWe7eHKVTbrgaxj1QjCAIR3LOiTJ6wZc5/o0GzqUT1Y2ZDf1rU
YIfjwNL3ms6Vkx2llyyb8cUSm2DN3tPbQ+XY0SbE1+SeocTm766Xf1dNXdGg5p3iv6OcGMjLdfYv
u3ZmJD5aKoqALiNti64p9Vs7S1Bwe1xUKxl1IuymJYVVJouw/8CPDBJYmwcPjfTYu8XusXdCdLWL
hLV3h6faHPs5AJo/m/LxZIAVFo/AtV3P+slY0zpGC3qDHvj9IrLDAPXEJlxW5eJVRBAgHj8swbwe
nz/Qf2sogIT83BVzjR2N9xgEGFZ9eUOOfTKXbefJsRPiOELq3cdN5NWUbzbrTbIuk73P/MUgWtxn
J3Y+aGUoFKe6lKG4VLRvdbWnt0TH0TdPM97Uahs8v3YtlDydIQb1g/qnfwHrD7F/A6QBDxQx01JZ
llD7SotU82yI28mvNqtDrRXSW2wdKhaMuPmw3D5a4/eOubKGUWyAu5ypjIeeIs2mUrpMXZZL/vus
10mpo1tK8IB4gvckSbhWlYwP1gRRSFV8tzVuyyA1JEUArNejDcGd7MCDX6NDfQqes8fpNOo1DRQ+
US2xX+xfpy6ut2MO2HPEWgu9ykb1BZPuIT7UW2/kqfb35v2UvHkio/HAgDGBg7wDqwbkoAhqcj0w
3ER0pd1a7n3i9z/uwKe2aWLXe98BNSmO7OMyfhtEf8CxUNm96Ng8GvRgkelSXTYI6y7E4eoSVe31
PkTDnTXpRm/S6nG55YVvGmubia9qkl38VOzvcKvIlv+61EWia5hOO1utfU8tnRc6hPDDaAR+y+SW
c6r3oDYMZzcITbyfv82xg6XLl2hw7pxCC/rHDEAo9msK8rUzFghzfAUXN5V0VAd/eU9OQeGkr4+D
G/scrJCEyRGoMMrCYaxt7646f9H2vfwEbKfxk7Ndf8ogfQAoWWUDMw7hDtwBlTt1yzQQMHotl/pg
QQJ7JnY0eN+idIlqZE9DlXNIi0G3XSYc5bimsry18n4l7ARvrpfmZVQpXXqa5zrvltgbPc2IJD99
KSRrQAZpTjkJiV7peZpfbp6laabOvidzJ4ZvLHTEhZhMRv8wNPjsbFLBd1/lrmnk8u4o1qpWMshc
GM3F2OU8IWaC+BkERpJGeAqbqvfDMUoNjIdTV57xtxmVFBNhw9sCW61hqrCvYWlQuf2IPEevSoZX
+vssMsJEjNowm8K7cnFzMyuHMh2cJc+KJ1BhgDi4K9to9UfsSneHEYAjjLWEdvWk1GnqlbCqsE0t
/cO6teM6SPh9zE2vLgP4YVcKIiMrNb5gj7twwQkU+oYeMNf5FuYryLS82YpixSvM9W2s9LZ08vZq
asAiXD6rODc7dT5k21B6ekVW5dJ5StKvDi6vX0lpG09wp4KJ03hTRE1pUeIdQjhv/9jZI186JqkZ
oMHxWSzC5TKoPQkga9VyE/K0lNhu9lMsh/HqjE0qH3aJP56dHfmOgntOjfgQpkOn5yQY1DrKI/UJ
D4PU5j4xXIEkGNzPcc2Hlni7kiydK7vq7s7y3EOtrPeuV9iDvDv3tSxXgNRg+Tc4LYQBTTZ/JqBI
vVsjtiJ3rsxXWwMiwmiuulX2L1I+m9gGJY/KpoHIZ//Og1F8JP7TRyQp8LjPvbkVwLwsOwmzxgUV
hi04ow6rTAHeXWyA08x7OY0Nf1Na9b0BQ8yN82An4w5FaiMTkqK2aeCv3ayD2gtV5st0Qws5O+bm
YIHzG6/Mu+Fx3qC1kmJf/lHY+rhTmW+zNiaJemqfEBQiGY7YluJMSfv+nyctnPEun0yhDvhEGtpb
H/Yyp/OJAed8gPj9KPMmTTEQIKL/SOxYF1fRfiWBDVoujCNvtNQSVDzK+vMYIfy48PhuRIbfxPJn
sYnjzVI996nazGeEoAsqUgnX5aicxh+v7qgfrm90LcZVfNdINLydC9ZL0uMLSkFWmX7NSBq71hnR
OE7ugxDOG7BrIz3gtlslWTcZXNeQ7+Lf8q9M7fPX6lLVdZH+hL1t1vSF6swLqLM3HnJ5cnVx9+3q
N6ILdbBic83qrhmTFV7sFVSq5N6KJdwoRoO51GVteDQ0Kngsi9Ha2LHkSeFe20LDaBji/UNBm7Se
yn0IOIDXifR8SR2969cHjftZDBBljo3pgKn4fZB0ZB5fogeJivkq2LuDUn4mCXZ1K0ejt3XyWKOP
21z48xI19qvWVaZyI0g4W9e4FuqjMKGS288iG54jvzveVHOmeVSgdD3dmCWX3MMuvCmepZ11bchK
cw4ueSu3rBk5sc08K8oJBrWcj0Av4G4o5GnJwwIppc71k1dEbx7CoA7U6VxCPGJgirzqvTh2M59M
UrDuY48WTQMEyt0buZ3C5KcNX1UOCDgqJ4WlYOHYIDrhN0T4ugzZp14pWrg59dSuf778alWFGjgh
5ewgKAUvOmr20tzR8HFCOypoO88TKT4WpCt5gqEGoZ0/3dw5WskIK4OVnUhxdzi3vmG3h7aHzPr0
XLAWm6mW55YdD0W2RdFxga7hoqrFowg0DQrC2rmRc4nRNGcTEq5I8nGLDm4Br4yYAl7fD1iWODrF
AZuercpNcHJYV9CmWVGOXMSkUIoU2KSxgfv9G0iTN5smcO7ROLHFtnjUTZOFbJNbhkuztbhaDoGO
VsmVb759cFQ2ea0RY7NfUU+m2ZkggEVz48pwsrNtzxnjWU7JlFqVwNUEzEojFEwIYh81m4Ty0Ymp
3U2YHFDkWdoo7brgiWtSd2T4wIbYcORmvgCIVAPh2B8lU7zKpyRG99WCoujz/KYv3yKYn7/AfiaT
dIlVQMpoRTE1jomizNJeQdIaWHY30CWqmr40uJA8MA4EtQxf4FDMpNKtuRG+TrwL1NyQObFW861n
W+xGizvY1yMP64vtCPjVmUo/tqrby/+W54BTN6l+tNjuaQ4pU2N3wi2pLiL0zn4+KPalfgmejFYF
0q+ztHfHxeGGvrJma0/lcifihQ7lybtR3KQGtixiSYKuZBsf8Fcyefr4c6eN0AJWX6XZv4NqQhG/
f56QZAD9xHJhuFU2GYJPDKLKNdHdz2z66DGD/DLFxlA+YoIDqzEPJmKD6tjtd7Is5uv6LQlaH4er
wH/c1zRyUieuBhTfC8FSohxUlp1YNpGIcDiH7bdBifDdMdPjL1DJpjLKt+eO1LpdqsI9uRfJWAZ8
CL2qK976BzFUjtG2hAOg7qRv310sspXtk9ssnCLCrfk/clQJ4UbLArT+rqe+uguUgx3UIym1WnTo
0FcirLeYJrzp0SkA6n/KyREius3bcA9+hmu7Pl3EvVUBiYB7jQbj4gXt1W5hr47UL2gwsoWATnc3
9y41fQmac8NIwC5TfeA6yl7bhF2mORxTk1VADVg9+oLCGBjbfcbVioEFZ1rYkEoWKTv1Xn/wUAjK
NFKfgY6SiJYIM2S+LfqaCrM4d1V2aMmaQLbXAOJTiodFAH+9CxIca/Xzwtp58qIeXMNay15tujSb
zGIsZ4h+ejYvE7CfOvoS1M11aaqR+WEX7AJt/iZ6Ear8CK6JTGbFFEUUihNx1O0jfipLthLnxHvX
85MJX+M+gkcC9JuhZTwEXqsfbtF30w8o6SXSJ35ru4tlrI44YAVEHVTHAJ48PSYUXTejb49aS475
Ma3btsUwvSNJotMA30n3dBsNU7kjHid0fX1iDI/SMZWh7pPOc2ZvOjQZEqfKLpeS8h7iyWYAruFD
Es0XJZGw7vYykpIjiAYX0Sr0aPs0LE8/piQfn+trs6mTg5T0gjzX/YppnV4VHIMLOUk3gUP/YwiK
KvfsSnB6LcNgrkrozAxiPFAMqdACcUHSNoBkXhJ305g4QfRkrY4Ru2N9XCJexvIr3HdrFA0GdvUH
sOr9VcWjVSVY4/BLiy0CySDwtqlnSnB5wV7+Kg60N8416ewNoKN3D2JuPGA0/F2yQxE9CoVpjBK7
AI/gU1buKk8pLMYtjmsV6T9OxvQ2MFQPtlIcULpC6HQidaiyCanlF08SEGC1tKX7bK9utj7lrT4S
4gA/4rveNGzN+2SdvuZsFUWVscz/0TFUEW2E8b4afgwUPMj55bgID0WsKMprswS0JfL+W6YciN1M
gXYXUKDg+EG6KAokc6RHfHETOPPHCvCegBV8LtlSlneSOHELjZB+NUM4X4wWPWgFzCcI1patU+ET
5jXJu3JYtCN5zr4sYvKaydEX110WTpx/TpnHm+5mjQoiojsjLUBXFksazzFh1Fjtci3TGXy/Vmbr
LT2i8hEuuAWMhsqpnUZ5ZLogjddsNduXkoTW2f1NjlvUpTuRw0osBMs8vS5XkOzeYxC3dQIje/dr
H0HsO6C8gammO9aZWiwyRmAr3bEEafz/Gu2mKXpw9D0CFPa1LATF8BnpPlsPjfg8tx/HT28wnDZM
2paP31GU3j++gWapNIOAMctkCPOF649SGjWonl7yt8Ud61K4yuT6ComUHR/B4QxEZc2TQYW7olVf
IAfYyf0g0X1+1x3DbmhftCj3qg8+QKVf33lgicblI5cvFayLWrH0Zb4UIETD7m3r3eaL0qA5pvQf
voyJ0fOjqK0nODOg8ZVttzi5ByDhIIIXfrzit5aS2NeUyeff0Pzv0ZEuqxjAh3PWZ1fFNqBGJPL9
hqLwDqMcmBoqgh/W8KNkKi4MLTFL3N/2PzdQ9WFunfZ5wfWnozr/uid6cJ3e9IaQegE7+MP7fZfR
9tq4qR1Ru8VPLC4iRKp9U8Ibs3EOYrxPMeavHIFPSFrpuyCjTfOABm81XXdRPuAVTTMj8QM9brGd
640nc8NS/VVsvpZAUPI5qzIaz2PhmXT9cAsaUUSb0ZOchDyJ8+9JS3EDRmYRZS2iNmr+ITJ4Stdh
1CyBril5+OwFabdmGiMbOeJPQ1hTPxDTfk8BlHCv+IferCQCdwjd/fpCGuyRPa7ZVB77EGmsGra5
P4qte0mgSKtYEqpplVenMkxexeXZrAvepujNzfjW2d3TPxrv7C5MumVOcvXmQfEyjpqmOBqXBdx0
Sqtc7sLVbVqMN/jxlC6xT0ArHYvFRxAMfX81PLQ94kW2AnJyu4Qz6PJshRJ0RX7K6nSzyX57RHVi
gdbyFedu2iojn35Ic9KOJuYiUS6bPhbaJLFWD3KCMazUifrrl1xT7xoq/TsTUZNP+mczAhul6zcN
41bHqG38sqJ7147a+NGICM7EbJpSEwGo6nSzZwX+pbjFWDluyytQcnvRSt5hPwKxu2wi7Gl9XN/x
v418z3TAEzR+TqT4x+SYgiO7zqaGfdX9ZCJVjQJPGTQH1321QAVEwgpr4hKRTq/JYaLlgnvkcyYb
rpJueyv6DnMDq5r7jcyOjuLdFoEpT5RA0dfY1F+R+qwvLVeav0kFrQ0Wqbkgs0OA31eIRJPuPFsc
A9jeIhZO95p74Xc1vTl2maSojHoXghyjJdVjF/FCUJwl0QtdQj3APGoInvQ5Ze4bepBUr4eoIZtn
5hbDy66PGno/WMjGc8zKFdgPg0/W5n6bVmg5dFYruKAdjNXEmmcPQa3tzVQ4rN2E/97FBrOuQvfb
VxIbLHWAGqHSpDDzdr+VX4kH8LL18qDBIsF6o+lMykfAHXH2HKwX5qZcKtbIjgrcpofkQUdmuq85
Q4bwTYK1Zpg1TlnV0WdwsuFyASBJzZUTis/SLBZJkSvMW3DxfQd9gGwsT4kA70gb+OM2CoMPq76X
jyu6ExR9Sm79B7UrXGbPh0R/aDuVBBrRjwItWEZi89LaOPbJopoJAnLJT6lzSWerpsC35qTmN8nK
hff8o/iSFgDMD4NtDoyzVFTV7KiEl7vMe5FM0ZcJbDJMTd17ITEtpnGPGTKqq2VPJy9vyLGGH9+O
n6wGnha/5nz7qkzhIh+qcEr+7JI4Pw0IjZnJzoLslUsN2ltxAh6qr2d/vb2xh0F11ObnEWUa5FwA
iV1E8bAhC8lYggcSP+wQwdY5SpCcaV/bquPieYuKGxNvcQ0BzKmU5Ndj9evQPpLIJIxpm9ldmO51
fgfZzI0wWbqgb7J7KIPFGA7+5tf6CEFCS9Oe+S0QfFF7NZnZohuIxxLx6hUrZPPGGLINqCtlg+CB
RCRzSDlz7u7vTfidKO5m1ERLrkqPHYNrRaHdYNxPEfRWT4R+tKhGc6+jauAMFnfZraihOTtQI9cM
A2zjqyOqCkv3GG4noH22p4AjGoOs2oCVnRWhKAs5eGUE1V5F09HmsKokeEpiotzDhnUbsmdjTpJU
JrbJoioKPPKZUk21ZwhroGPuV5avz0YCSHYIMxtbpty+o99NyWkLcdIVLXjea/W+gjqaF8zH8UVP
XXm4SAxs4dVgiUl2Eraq/2IdaPPgs6QVqlL7P+ltbUFEUZ/tLhlQgkGCaufS7Wi9RZlojxlhx0HG
rJLv3vf0FtsEy+Ch2gwyJ/tsbbXga9zR61o5ZLXuOn5raXStF5Ws1lGMZPSWTDWjdGgXho40vPyI
lO2KM2tSREQlsu94fFErLEdiKOufsZmMQ8PlAZMIAT3TLS0bHBS7+/0VC+UjnGkgh3uZkWBwx0y6
R6TDzG8D5J9SggURz0tuFezVqRZCuAdARx0iNp76nuCSkj/rZlwbUly2P6r11STGxK74byFH2FSw
CkazpJXcjpJgYMB7ASyb36M3olGENbLA7pp5EdgZa/O0+02NqTEbnlXZ9tNqUpo29069Z0YHAhg2
QvujcMQm8MBk3o/PuNRS+x+z6dRjvzHUEq6nGpHMQ8996Gd8+y3Ur6q9Wcuc+y0BK7jm406XSXdD
9chgA+kodjKesamUA34MqACtmKWtR4rsrwHJsov7FRsSunBDIHUxndshU+XLp2mUezVb14lS9Atp
imgawr6r8a3HmVtlStZkOG0aWBlXyO+sQtz0yjksG09Z0DoPT1UPJO58jynR3EgNY+SrwIHDsHWx
ftTpkd8mmTvUEnVeQ/s2R0dMRuITzvjmYj/tmDN+dtxLKSpWvycrXJzcW/ceDfgf5xQiZSsOes9B
zZzrySJHkX3Ll4F4HPo1Lg1RmKHarBW55eu+oiX9TWIBxcfqj1hbwFOS99Oq0/MvVO2fgrFwvhw2
TtX6b3SK3ccnaOIdMy3/+Uc/AL9pQ9Yj5VFLTWIQB6XDw6lf0BQf3MjKF6yP0C1j4F74CNTXT+w+
zuCsdGQPbhKgeLrOsRfqVVcA6X7uXzFPef2d/jALlUArHWCiG7v/vHezBk3Xs8csslDJ7A51gvWR
31g8O2KTfvLCJPp9kjciKh3quVSJsqLHIYWh3M28CvGLVAlrjmBPdd7brYn/V06cuvXvF6wGLDD7
HLLkmEzYBvc/GNYUP2d+RgBRG7UwopKi4NdYPpb1g/zzGOR9ZTBnyKAduR76Hb36k12WrL9U8pzv
sHWLFieSIk5i6w430qXp7VubLVjFKV4sQEky+DsvL0d3que9ONAdlfR2wtyn61baSBxTq7iQ7KGa
5t0NnHFXjNB6QAOX0aRiIG/Y1SuwCemetDZ1z8DJ/ANbhlkq0eOpt38bxeK0f4Rodp5v1Uml/Bn9
ABoltbr102B/RMIgBGIjESR9IGjDoQZLk7f2rLCFlUU2ej2VtCraA9ROH8aXYyCUtYPy3i6YTBY4
ZRQcMrtM4kjyoJrLIkljMcG2aZuyVFsMs6UA3w6gSi+WhSw1NLOdhH80vAtZmIvkf2nbw+TgS5t/
kLvpSJ6J75GC9ZR8Hxy/nSwjKGp4QlTV8UcfE3NpCysO8g/Tsb8wLBwrDG8X2XhT+QrarhWQWcNe
iEyXv8kosAgub0b25MZ2nhZC5ttPdEFJMukkIHGQCi03iDZy5zgpTg8pnhw1rVMqD7D9dgPbX93a
XBhlvZJ3MeEX2JQ1yQKl5SHOSG44FVHFFPK6Wz/+nAG1eKMQLmUIJAE5xEVcoqrtVgWDcRCZ9t0q
LuufQM0EHj8gK+u+qQjPi8VuD/0pXJrT/vkPBaIF970WdK1uQJb33vbYK5/b9dy/+DP5qOy4o7xJ
AyxE4PL3u1jycVLTGFDGwW3lhB0uYyOjyBOZx9C8bvlWL9cYLjzxoz0h/DE+As+34TXxDVcdbalX
c/MqYx90PGM3QlQVBqG6sfcZUPtYenbd0Bot/RUIk8xGpvbT1FM7UO2R3YZsHj/HOuyZosOc6GPw
suxtJU4PNQ8aDvEmv3hem1bloNUGvm155VbEgzgmXyWkz2ywjhB8jA4f8ppGAX7IhN0MxpTxzmq8
FkCViJKM2VrXHIDCY4pj+sxhV/mSLqFIOTwjheRjSh/uScdDKfh6cPnMKceFzQL/Z7MJVeQjqgHq
k7JE/pulAPtUD1Dx4xgssDrvd0cQchuaXpWzaPhN31jHwqpkXYHjkpr4kj1RZIox+eLSpeI98Fl9
Ri0c9HkUWeHhhu8mvSFkHHaeCCtAtX1NlkZ+6rV/QdWG05r07BPgcqnFd+5/1LRV7vuvJB6d3Vtl
46lZz6Jw8U/kkPhwOPMmmHFkOjsE4xlTj5sgWmVNZO87oqliqYkmw9RVs27uFerWsB8jQDZPNUiy
l4+NYJ/bUq53CqSHbYbBnG99asRNVsRdxsxh0JEr+vSFS62EyfcUt7/NXcjI4/ihUlLxLvudDYUJ
8mCFeeUrw/VR3FlE6ngypM8zxn29rxlzEm7wUeQo4drATLsw36I8JcdC2RlKjXEUM/tYcN+6LiwM
YZFl/gZtR/Fr7/khNWFWVt3x0MogmI5oSfIJE7KHnsuB+0e20nXyeroEHSPplTSWa5jyr/AX+Kgn
df0Yb5i4wsZVzA/pwfzWxOU+tvD7SD+ubyilLhKyq52ekIBoCaRCKZxIjZ/7JN/IATrItsapIZA6
CJs8Q8z/RBwxr5j2ZjFVNHEDeFMMF+8Wap5g/reZ7WZNZXlu6CvxmLxC9xkLY9+0a7+mghwKmfgJ
D/J6i0mB2tqFyndV35QiWlBQLr4yqpQKzO5n7a/ewVIT54Nu0+hHUk/7hxKool5cDtCP42AgpOx2
EvwBEbxIg2IXhk1AwMG6FSct4I7CNZ2GeY23W/Ra2SQrLru2TjfGI1wxVKG2NU0tB286oz1inVS/
/OKKqjUqxr8tRQdkvDTE4Z+MlEBfZ2VzwOZnXUpbNmonoQq2f7G6RjTDe82BliSKrftX6qA66HFO
uYHcDGA9JkJNj0V0fvq+cywaFjQBsw8sCpLozbLZiiRZFLRkmXvT+PviWgSPtjJNf31Fo2oMEouI
0WsZmnM9SPMrQ3giCuLf3+nERhiw876WiiW8G5lLoQdDCfI/NvFW6/yDYOJu7LdbPIawBfSPho4W
EcUCC46y3y28TnxFVdpS8a/DbcSZN3sQ95qj7fPekFcioUgyyaz2+hXNvtdU/evI3BT7hhzNZXyn
RmoBnobyKzGt4OO6CM3eaf8wNLvgbxJQJbiRewP5vvtFBbUA5gbzt58Kui2Zgp/QvYCagpWfMwTH
Iw3+UuAAIETXOcuorsdhsbw7MQ3AkLtLE2Rz8KZti4mMeHbfhwGq3WuR1pV6UqB059BymFPzLrsr
egrft5bF88KKIZfaOF8jdk4OKy+VGwC2wEt9IRS9Sj+6g2USwC2OF81O3ETcc9yaEPNeEoSu8ryi
tLTFqUhFiMB5XgyEPNivMK77+X24i/DteJpla6BalKpDFDJeHhawgwGRp5EOonMW6Oo2m9h5lWRj
GkxCYXTTKabcDGEHTxMpVOWF61tKJVXlp6ra+hh3Iy7mu8fVVp6UTRV0rNqhFogz4ji0JnsZHRcY
n/K2mSiYuqr82hZl5g2i9bZoQ6Yz+7+YgcTeUiYRmk5D/ygKE+J7DK1t6GJPgukEwAiXQzzRc14u
uUZIZWefL0YjdqAqmFLMtyN4EoLs4tehYmXdTjrtsrXWJwq9twzZ2TPMvbWIDvJwwe54G67phu4X
pj/jwbLVmob+t0iJh7wbw9pduDvV8z+fmjsCEamEIbfz5CHylm0T7ACPWP5HC5Eef2zeU4F2Zd5p
gRYop9o9gCRDoRiSEoA068dVhvXnSixhOprwsyHkkTzCCSeLsBhfatFThYd2bHjAaHYFCL4Y5Liy
NZYcDTRmO+NzcRyBTQuJUhu/G6aaNpoyWR/mJl1SqmFqH8jKAYVpIhCSH79KUIfCreDjXJd4YptP
B8FSlNd58rNtaKvtox3fW84NDRDVFoyuiMRXD2cTYShHKRCGv0h6RKpTYK725wC4ajfS4b/yCL5L
aWz6YD4VVwiHjWFSnowqW1+JWCM/bWmiahZTF/0LtLph29IheZjxc4XG3Q9s+h5U9tCt3kh6tKrf
7hn03tU8G02Utau57dL/HOH/JXGvUGrlYe6fv3aH+1xI/Mfjq164nguGHXn7siFBpgTC6y0VbGx9
YhcEYpQZlymsK/Kb5lhCLMvXKXtRTPz2o7b6A+XnAxE/mEAwpe8XVP6xMGgompr20pTMAjnxtdp7
iSF9KHDjmD3ptu19CA+RAu4T7hNqhDj8TOXCeYu9fsQxBT1syTP6uWaV17jYpwI+xvxtp73CEH69
79IYvuVDhbRwGJk07wRo6JtEPFFusn5Q8E/DUC9Mg/K+zrvgCt/fPVrXK06moHne63aQMYGAJ5u6
dQewVC+qVJQJqUYNINJZVZVpW2HiG3zFi7fGZ3zM4Ud1SiHk2/b366k9Pnw0QLJ01wjlLKKkO6HU
y3wVBL2DBzHl3swxA8Oz/n052BXDfuUvC2jQktP9O+sqgvpZbs2f19DAXAh9Lb1KkyNQ2lviyhLy
SA2UWDmoxYBDxGMcpxG2AFTTjNMz5Ssbq8fSCyUPl8TnIa23/wjHWddFczMu6OyfEf/U9YHgL7hP
BtiA/KBHf1331J2wYoHKWcrjnN0MmezXSM4dPoxzJgTxxjuPUSILnBqw6YXB48xFCqoQXYIU8fvD
leUVOUKkeKamX4QoXNqfGT+gJc4S+WwGPax3eRBDm0loQ2LLEcfDwR7Sa6Ra7CtfiX1iHoKHjWrk
20lXKZHuzKYVAM2Zolk6LwX7X8aShBqNSll6JpZuowGzgBULOYEVat1fRRjWqnYlC12meyvdgI1S
iaXn1Duf51kjJvHO1Isl7xaXfLafAMK8JiVdKVckdk0dmhnQi1BRSS2h88WPHuU5shDIuP4u7hjh
ICPJs9ZXemIDyHAaDXYhgOAb5Lk1x61gDXQl10U8z9Dw3x63fVbRVJPcMfBPn3zUT2CFn9QjfRVd
9bADMX2QjK6LCFIzZK1bLSSkpu2hn7ttWQXL/euDAPrzw+mE4pla1yjz+xoxo9hFmgY7IpfC4Yfn
r9AHEn7MtB6TDyW1KsI8CQ3sPf6Zc14zjiJ/7W8+7o3tZo3q0HMA5VQajLb4a58RxlTnT4vS+rYs
zDa01h/HCdF9hLCzTFdyJPV4rC1ttjZBjZH49Cr8bXTXorfrw6CNeFNqKMUSgRkJMkGiGeQhXlVb
4dqmnbIwtj6PsBkdrOdSVtM2KJw6aEaD2xaX9EK1tBKVOe6glXHAMtqVnWOI/Fwk0eewJUvgFR7J
qBPBW7JMfWrY8S6nnqmdrZzpVSbJLceVlcAbrKDZujBPuojYu+TE1Orxy1i/DvVw2uNhRA/vNoSR
Tc9S/pLJuXH4jfYXir4rF62qtTtQc5m4ZgLjdYDWenmMyEIKio1j4+uNazUX3MqSBq4cSUHYskwH
tym30aTBZCVMZqx1vcKTu9QYb4X2dsaA2tn78/3IfgRGLfUkpsQxxr2uYhz8Uq+YQP5upqwJHQAq
ti8SSZWINV4Zp65SGpJ3fwL4GGwH0sSb1H+yJuOHMxX7mDVqc97fS5G4GOvxtPQK9gntg0sxLypK
eqkFljyPCLRnc+JPYmAOYAH7etIX3kwKE9qsfmkYJuUoYT45KoVDaZwdWvoOCp3CV9cLcHlZ9d5R
Jr4FR7/2lb5Lu91OVtXv38OAdSIAtD9D5LEGdf0h6KLOo1Mvs8ckrqclIZMLJ1BZiANY2t6lRuSH
7MDAHPc6VBmK7tRfUTr8hDb9JMqf26yimFA9+RA4S4RJtjZg02OjNTWEjesyna22zTUfWjUtjzHy
aR0j2Q+zlmq+Uhizr5WI77MHIIX0te/5kf5oaADKHfvDqEAp2Qblohxe2RVEIXu0vpj3LGRzYrdC
WkE4kFchD+ir9cDCG4tzW9MOL0InrD1h0WyhRVNOuely2svSqHS+YcIRQ4nzwUa3j2QacqFa30bt
t+uYLxjCBqgaUmqn/LdZmAQb8/DyjDlx7lD3JhzYeKmmUQgGe5MSqFya1WyJeTj6taDb3W2jLftr
abj9tnTfqY6Iv9qsfrvi7nlknNr7XQyzY5w9ITp23B2zs84EMKdNGKNzi3M7QE+jzX8dPnuyJ20X
5V1cWsdq9272ChZtnGo9nFq3d6i6VT+Aj6N98lKutp+V3FhRCjfw5KM9slndBSCNw9V/sflDWBwY
zMJ1FsNv86J2gA451tce0nPWGu/N3K7rTT41rrrmeSVhoSHv4Sn1BtbWT5PGSfzzp9KYYvRaJorw
IwxyRvov6GKDCkTker18hzrqXdkZLQ5qZNXwxjvqQYYOxKSZIg1YhfpM9crwAuZuDtBF0mWt1WbH
70AuG4MLdKi0R2ZjGT+gvUE4bXKh2OYxeL5Apq/uZhF3h79Td+eh7Z220NFN8AKbIsu+By8H+7U1
mu9BV0H2M7TUJgo0Oh1zfFZL4zcMr3lb0NOhlUxid7iUIzWvCD+2PINIWgNdM0aZk+5mea08cGYt
ixlrLUB3jgkWTWXOPgYn+DMYsqL9sYapB5nQT5L2+1KWxaqUY+GaRFkck8tDymJEgougC71asp2z
jQtyRlV4kKrYFKbikRquJLkytiwOJ64MrAe/qsGQ1GwE4u089F10varvyQvXIGQCgNclhK79vAWG
S7gYXby6fq0QnVI62c/QvW4IkzFKgYDPiKSbjDFFcyrwKsEOQX+VPCxVHqMSucIr0ETXx8q6PXsb
ZA+r0uSwCP8qK2Q+EN5YC8846x2ImEkotStINGRahAS6Rw3LE+IdBPbLRDF+9ThQX0IsytetjquI
3C3wegLMSqw06dNvGRB+O3+5HAwg6Cl7lU9rP1jYFnXtNXWH9MhyDRzvTsffwWpdCAOcJDyFoi94
jbA8hYSJrar+fJ6cyavC/sOu3qdyGFQDTpp+agNXpnUp1J2Gv7w7siz+IvJmQ0MKI7Ksq/GFK+zG
qX0YS9ViA+mSrniwwAxfccoBsYMj1XqxMSA9YMnCyaJ9WZIV+lkKvPTVLT7FErj5jgn6c+ovlUw4
nY5tfrJMsQdCJo7ckfyLGVGo28TSQpC4AVuP9XPsRLEv5Sm2ZFKJ21cXxfuSR5BwnavYdXM4d/bk
lGywI9i+jRIWF3RGnR4il3PFcAoItcn5vjzNcAZLKbrmOAkQ6q8ItAbkemSXe1UoWPziJF5VxEmF
7B2PsqOefOFfTuKTfPt29XPA8nV12CcnMywkycknNBqfb+Qq+vg+UCN52EDYyiXN75S9oKra5ofn
y8dC7CTTLkFqNWoSI3QXrzM9FvTP2Gyh0J40Qqx8N2CV6b8VCX2pahGHy9AbZBQz0b3Deg5OnhMR
E7G2pLe029axoWoFFcqiapIVFpeNSM3AXLdWPwHsT7QfQbvTU+djQYpHs6fJesvSuLayle/PiUFl
+82vEHE7vUMZX6hPs5qWmT16QMg7DDKpZZme275wVMYAnvF8QCzSy+7PEQQtCfGfV99Me9QRe5OB
Fit4Ir3RA5jSyhnP2lrrP0p7xV/Ssytep5GbV4B10acXLtwI4In0zrgdFffhoRulbJsQT3LcwNkF
ViRU5U45E09fqG5sTIwUN7czzTNdNC8xUsmtDjJ0Atoxe7UOVRvdcK/Pfz90Fx1CfOTV7uH69CMy
FHtHbkot8m4icAQxcv0khXFysctZ/bbz/V1tRbmMnOg0Du5izvrPXpi+6RBNXktwtpXi3eZrNzN/
NFYLF3RvQYN/t2wy1VbBZrPnr4M1Tg/wF4jna1xAcobBHq6DKVfvxDt8nL7lkGPPU5xKmkYn50ym
86DIBUsSOJNWmQMJl3tlR2iknYBUGd15c6NmEqyafBBHP8X2XuN2hRTAMeiBtNzJFkDNTFgzKgmR
hPfpdZHNZGZmUuv8dChp+IVxq1Dm+YWUBxpMAAgZKvgreBxEoAFwNFMtqohnpAFGakMSEMPX2meY
lFeqIqdYmHG5nRQj2Mx+T47B45HQLVTG7A+P9Z+dOsi9dh8LG0+uUUkcixax9Y8sWStG055/1wVw
2J+7PEeAkLj+RTbuQnZPnrCKA/WOu2viHd9J3f6AM0RTpBs15TaCKsV2xiFbZL6jNVPAmlV9KutZ
uCysv3xmWTLW+dI2lAK2YmD3wyw8yxwWPU7RyQtyiXXmxa12C5AGYF5o+j+53ZKho7rhcGguUS1v
t+688ql9gCkYxKK1lioGlKUqaLfAw+w/+NN1P0RPQDznh/Xy+ixAz2fRnP/Pz+Pau1g2jqVHMyw1
mPNcEwf/xiKLvvo4LTBGX1FEdZaabNfWxPaWFlmAbnsDumC8AOD7b4C0cImf8Qr6zssixTd17KdA
1woYRVuykR6DB1nfT9S++g34FH1cGv+8mqDc/pbWxVeEQT4wmwFyxGMM+1YfnjR0WGM79h15mVnq
dp/z4VW/qCXt4OvFoFJul8DW2NErqfINoxsRHFrpdrcofCZX6h2CL/zFKtLVPgPIM2wiNbfs5JMv
j81HG+zIJwfqVj9Myn7VfKli35+Tr0Z8YktcWCDUWwq8ALquTJ0r970GBdHqI6LuXMGktxV4NtSb
YXomCYyGnGyp+euP6JCPSh2Ulqg5wN50u0hWYoNM3lQ1uqLL5Ue809JrF36Q/fEkhfy+7gYIXOlW
Pmcy438Mosu8nehDB512QST3pXc4FaZ1K4oWKzQAT0aw1LlrMzTN5nG+Ck4+q/mc5zzlUWikY0EN
jyg9lH0yc810RBs+iqYJWvkI0nvbqk3t0vjOoYOG9XX2sXpNuLOFhkvrUV9foiHpnwH2CNeOd3DY
8GOEFVrknm3iqxmex+BnSuPT2jZkajQdb1ZcYxj7E728IG4uWP3C8lo/YLUm8YXqUA21w0f9wfO7
C8pY6xSEWuyKFiCw1x1qRdgsMlsFiHfTonFBzlqZeFP442UaXj6OV9myYxgSmewApP6XgtWrd9yh
J+4e6nCkYysiUmuGGOPKqKaJTQdGHfr/wBCYI5/njda/kQ/3QkArALQufqUztwLTFpUhFoCDjNEP
dgwh9bZTuJwdRg7uRfoUQAILl+g/Wi4aIiIOzzs0m4Bs+NWHwoROLMPA5iNWtWKw5sBxodRYBUIN
zrHhUXggWSRkIu3sh+qhueSXnxMLo/nk8C4XuEONQvWnWCRUGx9NIOWBTamrPwQWjEepNaFKQwn+
mw0ef0J6HQV/scLyHKMMO7cZRt4bukPE3f1qJEV1dRPTwKr2abVQQIEWePSpSMA5ikQkVOSbbdpM
WRaf4NA2QoY0Jl+A6JIi5/zAypAcIGIcZLvHtllwcm83yB+Znx23OJ+LjfItPbOFiZTwCOsT8npF
QhZY7vl7pVvlT14ht4/awNFOa31ecVr71/jTttCruOrKv9CkA9TBVrIPeg7Y55jsTGI+JKCKyvoL
v3tJ1KPf4bJt8gCaxYvOnfTGhVHBarckNi7HlZfNfpTwZkM5C5V86Jel0pSPEcMn3Ngq5cvfRRYt
NQA3FBEyk2rRqtyM9LVHLMdrl3W+2Lc/28dlJWPDusIZlKVVIHgn12Hkhj2k4pfU2XNVcKjFBOmx
Pjl/yYd6+gwFeQtb4iCmJj3Nk+IK919nKrw1w9aDXHR33z1n9/kY/4j+HfgI+F9BJ7LkCG9dLgIi
G56Vg0DrJfMnUpJgHJ96qDeJXjkC4CKKbiJeJqv4+8HWNtbdLFFPEO7n2+xs97QYYBHyrMZJCZZY
dAaTmqXoHryOfZpeMdpUeJ2phy6sT2So90XNRVXavAMKQnWqQkKnYD8stLdrtK+Q32vJXzkdsopx
9ZJuvDunOJeyTU8Hfq80K54ijhbDKvJ8frNRqMp0J2RuKDKcSl7+5t+PVlvM8NuQHopv8GzS/zO4
XZNYqygS+HWJV52D/Hbug9UHifJNFGXpJjQc+bp9hlaqwxrG/jPZqe4TBtns+C1GwSQRp+1gcEjv
72uqaLUl4dq9Bv2bZnBu0R1b4wLO/0G9kUbn3O8A9vmOHsYISmp+7j7wSQnRIIpHwgW8EXmsDNrF
NukZoR7zrGeXomYrPjb5fWk69fqQD8bsCE0zsLBA1eMuWFjsi7lyVsPRhauRn8w5yj/YQr+i5GAP
JWJJGeozGT4K5+Rg8FsJ1X5gtpWhvMvCx4fWzLNf9B7RR+TYieyoAPR6GmdBVP3l+n0EwiRtegrG
TSfJVTUnwdgGfgjlJwGL64A7sAbrhaq+DeNf+vea/HYiJi4sCtpf8Y43gPHR2AO8ILISLw1c1w+l
lwYgaIFjwZprocQ2TmmBHOVglPoEsPMkP4b1GqwasukoEOOiH1DYk9dkPnbLXnRCuWqwXy5YKD1B
2GQAjR6843fsv/v+kXWrtCrc5s+xZxVfYeT3Gt89aNRy6oBDrpJcIqUudEqOwWHC0AUQCoTbj1Fe
6mqOIgKjx3CLQ5R2qFYLm7+W9AtIcORMU5T5vlTTJnwjyfT8imyS7PWvfIEszWOrNSpEsyAaisUJ
h3Jhn17MTdcZ31dibdEI4KqCMjrdkIii4rwGR27KBMQSZe5q1NqN1S302dE6Zy2Whtw8mguPt63C
uVNyKZUXmL1QL/DTVpcDbIQUqo+8Qpd9s6g9z/w94bQZVI3T2QN1bfkMH1hDpY4lncV7b/F31cMr
qhcQSy1X16kmlBmQRDchSqSi3lL5MmbvxVE4BUOv0Oros1kART4CH/6LGt2QgQ/FPbcEsXOUfabV
gW27vQY37Q61ndqGqVwZIZ5aa5p+4nbVqavvr/T1VPs7P6V5E1uNwnoNRHIgil9jfBmdaPJPKvEd
NcHOwbCDfh8FxvsPel1MPy5uFphxn4/APWtww9NfL+Qrc3B9yXU+2A+glcIvqzmZfyskeg6/ErRi
vVdhvugYjcNypeqKZIaIHXLHttLWBT+8C8vWKKl2gF9mZPlrzITgf3tRVA+tdco3mj4Xr28kz27j
DqlYS3L+ohB9zpUzXOtzRBlRJFSUw+zCnBLP+gSvzVzoE2+UhxE/uu1T8ZCNhn1nU1+crpt3HOF9
P3OJOl0iQH0fJfdqS1MmwXkKepDz3dgkYPs8OVfwLB2Oh5SMIgc/f72/9DTMSITgWH3n/ZxU94r2
GsCaLXKnjEs9FjO+8Uf4Ttm3nVf7vn/XQy4h+qKJ30gUdAgTSrDiSFDMHiQRUv3juJXl+aOeLF82
E8BfgDTj8i/g7LV2SgIU47I3wdn529htbdhc4txE/G1RemEm+p6WoWzHb5r3ZcNk0I2+cr6gySsr
Awnk1oPbkop8xNe1Z0HCgm0LAjI3iA2AQ31h2HG7sDS03yAYmUQmwozVaLnTwUwOlh4s/sW67M2d
am5zfYRDll5M01/cWOaAne4f6o+829D2ylDA+QNMU/4vO0owykyKH8xTjT2ZMn6xV4AKAhsL46hp
G7JufkAl38BbdIOfgJcNXzzQaC8DMWnvmdrYGfWsFln2BIQCA1x0159Cq5ecDYIZtnOv4ynfL86G
PCVEQRbvFhHOZUnpI157xAF/acvAUF5VOk1yabo590n5V1k/Y4MllDngdBOj4MJGt+7TzocG+dXG
xIXttwUO50EVLjOw/MKM52FKcw5Xrwa6drTobI3LQFaMk6Zp6YNwFZnORc6oLtl1UIupTxeqrWSo
Dp5PEICwYlwveJRokGWbBaz2XyKIRsZ14Lm4syxOyFapzz7B6YvRKnelsHAOq/VIreEGtyJr6dF4
bP0NeLpsxQzokp7s9euv0BX0dFRYqgBQyqTti355zcMmeFjbsVBEel6sZ4Z9WWO4hVVShpZzhI8+
PqvfLogQHWN3Kb3N5MjEEcAcDVcSsXSkeTEBM9IOytz3Dmr2+P0A49zHY0L0MXhKvekuUNEV6Tph
r37EaSH3IOu5ww3E9kfzJ2Z1GQQ+N7GsFqxdFdN1FFgT9VaAjYvUsEfBsONIrASFBgZ7KDx/zUz/
0bq9cHN+bpNksGSS0rgd898DEfjlrSYOfUR4U/fvMLksIuL/EDYiIUbOd7KIyRNvEnHIUQ+n+xs3
crOiOKTVtIdLQ1t8yFPwrm+y4tR1/jfaN/EC1CJ+naRnyh7v5gu3W/TfyqZviR7+gwjJlYTQ0RNi
J/rSOcwt0X/rBuald6gAxCtHxpAU4luQC/qYaqoA8UVeirQ6hIYE1KP/C4rzddEnhHlNPmUZ/X6t
Osr083UJPqh/oVJIX6ihf11dqF1TEFkoxhR+U0M8Ma4KTcNLbdgzpfivjVnz36ZcDJ12No2p1O7L
SrM6WJBA9r1ILLDEFYN8PDxWp2yoTBAr0jCkr+orOXm3U8ooHHbt4sda+L2nfDXlfJGwgkhpIqRy
ip6Og6eW/T1nSiQCTw+b3QNc3NFYh8j8KYkxa2jf6mCciAbJBlEEUxK4x4zHFxfWCZln+GyBVPVc
c8141l9LkG7lPF9ufVH/Ztq2MH5hbiq38MKIayBLTc8baKDUiXViOuMhBKdV95NN38ItVzSSF+83
BOdpPCLnZT5/q/tTxQ632pIlk20hEdVxlP43xPtk6G4rPvTy6Bo7r8txR+zJO6flMatUwFLBHOP/
LfEYmP54ICKQjUPErg48Y1gNSXrzpwIyxuXYMlCAXw/uwfi5hRxL/rte6yV2so0HJasIV0xznqm8
VQCMV4ggXEFxedq/pAKC/xCr49d+r6X2Xy++ix1keo47KMzqdUNsPh+3FGSkLklP7DsUC6CRW8b9
FtWhAJhneOPkVSSeP8jfaEfDAJIYTltrdSYwCP6SVKDMY+Du7nE6h8Dc5A+l0aD2Cqi6nUJV+gP5
90qViFTngVq8Lb3uusQ91Y0DOQNlaFUNAF6bulA3WRm/VaL4PBwSOIGxA88zU/ikmTOcw1dPkhJl
UciK5G2qIgy2Lxamff0vbS1weYNTuPsH7klSsZTOi5DKLO26fdKWIx+x1PV9HZ8hSdFG983ceyTK
hFv+qCGevIfV3+355xlm2K+1p53H9HBjVd9/ATVWWSmomLY9YwCt4cEFAr28d7aQpSpoLstIlhT/
aqvZrP4gDV6XePDGt4XSuvOZhKzZITho7HBJh+bpcNDiDBLNcNy8B9rgEFv9G6YrxpUMJUUtkwh1
Sez0lbbhuKfNsFtBO34ylC5f+cdjpSEgv3/v3ArHGaq/8cUzha57zxdw1+TL/TVh0gSCjyQKJ9VL
yj1lGnFqSbI5/YVV/2lS1c8vUOq0i/dGngwxyXQATKNn8FIENNsQAh3qdMV4CXkQAO/V98sIkoJM
/Xx5upMeVQs6D5wp6CGrh1IoyYB1SAOrXLuh/9PRctmnFjG64alCS/mAkq2p8+WbjvXmf9qrvzf+
zHNo8ltQh2U6DC9T4VnRjqpJyNnobjr5E4Z1Zc4iHEQjrAMpG8mlvCf/mIXUMnt0WP/KkiJUqtg8
lTkcqGhBCv5fBDKuLYgVMlkuWuN8StkpIWijXof/tP7gCnlpkpqVhKFMlVFTT+NjXQ4YwsEDdKo5
T3Skn3Gjv7v1lB8bEE+6v0y4nOGK/XHpbQOWve8bSOYzVGvAHY5YQwtFJizItCnZRt4YgkMzvMJV
AAfiFqHswTlcuTw4SNGMyfrKlQ/Hhcy8rv0sAijXnfGFF6m+IAG9zC4k1hk3/1JeNnfYipbSNBSj
L3aY2GUhjuwpNynvWVlQuHBvcqnFZ0G+NIqDt4XArIPNqjYBKxBQwTq2H52Qf23z/fcrYQ3/dFkd
pmpxGbxP37iCUtKDgmZ7M2P4HhQeZxjHjNHFvWpz1CMoAey5t/bgcMfAOeLEDKpJ+st5Y6emtcOQ
uik7ViMvEpjdVq4g/gfZEHEP1f8P/7Nep2C436Y0GZDk2bs7fuTsMDd9ufOxIZNu5rMKKFq1wr7K
x4HATossfF6WpnT+AzbeEIzDslj1ySp3tAwwZi+KLb6TAfIStTwyAsOouiP1lY0NeUoebb1uKiOY
mdxSST+Z9CtOseSBBxzUkf61yl0/+V/TgT7jzTveQt4PLJ79uy+U+6xLw3QgTqbiXYnjB3c2TTGQ
MGqLS0HcTz6WFsPndGiNrVfNCN1dYxE4o+zFHhm1MzeeIGbGi7LdLgVBq/ITkxf6Jga8PHL83/Dd
OGk9lskpcwZko1CLdUoSrPdNbHrWwXAf1fr8AMDn2Pb8XbPAkkxrM7UJf92TxM4KWD4jQ6c4oJc5
ZspdPAcswh5KsiYASdttV+4DcZKg4boLvNMeKRo+xyYmAO7FM9QoKmHfScP7EZeLzNWVzePQxYqy
6NQPevLoQ4fLDokb9UQOYmtdxPl+KBYab4/EAuDCrTNXQRMftPQf3h+dgSjpn/AdGbNAT5SDpB8L
faNtCpC3wloUHfdjv4XXBjm8VYROnKnfynrO/vWfPFNXRfoFMdui4NyoAocZ6SFGJG2crfVLmuvF
hzngttIBg8dEsAjHRtIiHKfHmqlCbO3Ra7CXDH+lQnld+Z1e1xMnOpG6wPoWjxWagb8k2VPz8tn2
THGX4p2Jd7NWqaHpCtdZFo9UYIjXwpNAvxooN26aF0KmrUSqEoyo5rvgNfkqgVILpAqf4Qlh9Bsl
YU8dMXp00MEr5WjSbbrMW55nkHqUFC1k4s5AI7LgNO/AWsIidRDax1YzDl2otcaPbZ2qzGjXBkLt
xqffVtcAwFu1jaJPWoDbxNWcjBcv52AHau1pXTmZkHD+1TI9aHSbxj1DiyM5BieG4iKXgbM16yfU
ZrIr8j3fXkUgne3gznADfnIxabcvEUpoQ3TTkbS6yf5NWtCdad855COqp/FLoNSLq/XjiLibVMn2
iftj4QWXnXJnEIHiDqDF93lmW2GHGY8DwEXCxEs4aJWql0EAxCOev2Nz8z+29kHIQUV4CKC8tS+T
BRsctyWPtPMxxXloWoUN6RD579Ufkqq7EbBgE/lHSUv1Sfpcsad0eLMQn/Q6tNwjTMdgZf9Onv9t
zCvYer7poTBlhaeXWeL5uqV2WlOt3DFEma96ZOQs0nYYgTqHBouUN2RPQci34Wc6Vze2d88cNXOf
pcgr31C1gMbrZgaCd5MOa+7eaTJQcdSkB1j8R0/Dsfpdb+aG8GHKfRVikPeP3VNo53mSdEG+gVZa
Z/uRh1qi7pWKutGRYnfusNIasALcQtwttlMY56lwvIm/ct0BblYzu82Cgtro2nUHQmN9chx2Bhx0
JQ3eJ/EARhBvW5sulw/+eo1/Xj5MoxGB5sMFx/xjzHO0GWU2nz9MrsjyoRcajq9mi7tB9FyE+pMn
gCezvyfDxmJr7TyIDQUeTFp1UMTQe1tANHPNzFMoztDoaHR95TZwA+ROxD7GzFWuPbth2y/Y2bNB
eN5DQuszIk1F327vsrBU6fxBKUc21eKyGWcj5QLpEqum39cat8T2KX+nXEsOf42gppPjehGZSn8Y
7BN8HyNplf4BBozphJXoY0zTk9jmvre5xd/KXcfHhnic10+dgSflGbyGfbNcm4h2XQktYvHrLigR
vpmwpP+npGR0fqv7CGwbBBC0jI087FrjKa/vIYXIe17JweijboZv3+epBgsCDk5ZkS7XPWcNYzdl
0V2b5ZiMYiTqZdT6kKKmcmtZMIiHKYrKfjUc2tJo89VJWtUry54c1lcbE26ZyjLadFpXSVbFuF2R
4UH50xOMjk+jmOF0pK8Cq6i26X+VJyEvhmychE0uKWvnNvEAAMqO802LFOWxPJfv34f+QjV20FnT
GpmtdsFEYT5WRotOjC+e+dv4xC7JJpk+otTYiPkt6FU6RjKYTAgXbepLPSVfoZ6/I8ULK3S3gS8W
cZrD/Pu+XKdYhyzHV9QfN8saiqPpUOla5AgL7akXhiLRX/SoTXTqwSMvv0Ok3GX2eBzO+DfLB5UG
3OJc9BMxqlgfSa1uHcYDsiAEVNwM2I+Iwp32JEYFJhbEPSc+RGECfeKEFl2MhF+aZT+5Go6cL46w
YnSVFK372okreIQ4vpeR7tw/DISq0LYQmqI/Ll8VcCK6J70hjXJoZJ4VpCsaADoh3EQPvezjaCCt
DTkZjCL/FmG20HYZ6Kg3WSgphI+oZ4ZvkdoLU1scplERhV/lT1lYEeynb9fHdQIXKsIsLj0+tCsl
h3ekLdXlnu3f2nSg5njHMCQfB8o9J+L0ArZ6s8OzMOQoVWxmQ0Ap+jj4rTXV2CkgBrF23j9ZkCyb
xTM08j4lntKt79nu+VqPasDuMZ8cb4T+prC/dZ2GTARqzupZbsUKk55BL635V6xJHoePxec+wmdv
lCi59k5Zz6q1yyxccWFQvfTvL3uzAG1KTYAK0YxYMozm5a63iwf+2ElGYL2RCzLwcJIMLLdKWtp/
meor0jhNgjuw8B4A+xm5FEMZsUiPxfEXxal1YNhABzUxFENNIHK3ljnUqnaFL9VGo9R22QgTBLpb
OX/+7PT/2QSeLELsIDm+2WXPhJx4JMsYbsCpZ+SVCHGKrePYYbtVChLfCUyRcK6J+5xHSWHUYHeV
P/vTENMUZRziPY9kLIXAeHSOmBz+3vehFpQPQhjNjHaLizTc/fqoa/vWIUufVLRGWRIOia9Cmj6n
JDN/K/QZ+GRHlWe7fOiVEf9N2QeBGZJPfL1lniHukZhNzcWlrMJ1iuB9S/mSCo1KgbF2rsP6z370
LcTLJ3Y3CXr5ruDieWmJF6ueGzsIg9UxEwGVhlI1qGnT24TVGK8ktT/OT9LrVz0FeM/hr3yTMc78
/Ym0hdX3yjxpZUDRHeL0Zwo/oQ++Dc1bSydLKud0345ZCcKYfTo3NW+kO5TmB7J7kfVHY2ZNENu9
p1pI/Ssy+bYN73w4c3ram5XK5RN+vZL+MVnVqDYn3s3wemwbDKE1UMy/B28x458Rv+L/0Ap8YOgK
6ebcfD4dCqCZNzZQR6RngtatcQhnYgua6WO7DDCa+rKYyURMMdqqiHtC6+5t8OA9DZ5efzOz98Qk
9I2uZn3IoSB0HXDhWCSEv18ZYtV2UZx0jBDeLhZRhc7+kpY36LTpBRJoJ6Pf5KiYwW9aXmfqnZwP
V1zvXZvbE2AGGxPwYzTpZiSwW4scecJhTPZfbUw3ZchyHkx+64qfdCE1s+E92TNFqjc+8Ey8vRu2
Igi5lFmHPb/7MZd7V6o7qttQRl6kd7RP8eYEvu4oeb6AyEZSEVncCCP4e542Wg9cvCTGemq4lzNj
Lkg+YN6G7n56lXT28he3A+Uegf3gfS334LNTk2ePAzrFrPCQ5yi8x6qxyIrFzUqWezFZ8311aaUR
JVNfRrHNpanynG9dsVPnKhql9I/BZmogADUYNuXtEO6hqvkf4iuTMkHwStfe1ep5b44yR0B+a1Kd
bCn4ZAHX9zpzLIYNpGVA9Btg9Ufhm19GiZ/ndpErJCZM0Iv8Bwti7BNXxV4lCybRddB36GHpPEAw
uYmW4W2ZiLODfhjADwy3JcQ5IfBu3ZzAYTHfZYeD42jiRmbRCyK/rn8IkCXaIjKdQJUNI3wEDEgX
H+oIDVucLFTt1HVisBCtZPDqPvtsiuQc1OhhNfl3wxOhBaeovwk/9ePLLJvz9v8uUzpBKImESK6L
DDtBu0GKBL+Eq4DFmGl/pc2KOkQbxLoaCeKyoh4p4skCt7Qvo0KsjNwT1tWtEOiSHBV5OuH4OA9R
ZpmKLd7RyicVWh+IebUFRqwjqR/N0JRdMRJWQEsv5sVsDUWEQPAFe6rqM6wqU0H/2BdOuqFkpGjq
WzendlkGehFgL8YwbQXMO1r/6Dtl5+1GVy2OW53nLSsR6+VjF74IVszVP5SvRdzWalEokSdNcAx6
TWyfrOE4mSRQfnrNjaY/0StG53D0wZxJhWOLWci3e8F74CE/ygm+lygCWkfYBLWj0dbrPLDfY35r
DzpjzccWbil9TtStBzFV5bhixgnp3cSsUJ7taBB3jw7P3+oc5KUEUp6T06UHQf0KVZjWVm/VBHzl
cffgvpCt5EcnuhU15pROUDce6mmvLgthbUox9RZFiIpFyLe7wBZx1mNEkif9TzePQCP7mTby4cGK
ENPwk8J2hMOeid8OChcQ1q4W6oW2GfEra1NT3s/I2xVUYXJnpgHE+CZ64HqXz4tUyFCEFpXS8TMP
iJOL1lg1dMLIpPN1BpNYBEVUyASMCAwmKXTIOpjWsEgZhqgANmMx7Haw1tw2H9pmp9gPR9u0Gsji
g60aAYCDSp846t4GKg6TAbIDeyOu5tWzzkdfpTz7ibRqylr75pEpIU0rVIj88PYfFWIapXymVJEF
AsmCTU3PMm0nQ9lwmdGYcp+ssMtor0sDdWASMuzWAEGhi0QHy77AYdh+9tv3AAQKx9+TqtNxziCv
fu7A5SsSOGJxntgtxA5QQDWulSTpVFiVyrkCzqluZpZssT2Z8EPy6MAXtTzUc/oncmWByEbfD+7X
MpxSAs4PrvX7JwrPeOweogWVE4euOgpsfw3clK5XZYb7g74Y7i/eAw9XeIqWmIzEPp47nXaSIwCm
NNvPwqlXthsWhOglMou3r0eD69qXyW9eVTbcuVpGWqnSzEj3mYK4qX86KI2syu9WHumManwPMzzz
bHKT3ka6O+C004KhXkJwuBuWDx7qrNfBcl2PfARQSInQ8fbgit0+qZ6k43WnRQaZbumwJDfRqOyq
4EJZ3x119pTQoLm2D2K/RFqgTriAPUuw8S4qmVa81GsqE4N5ueROPXlLLm4+b6sUOJTVIzYK5jkY
DZnucD9FXsE+ruIHzpQPk57QLGW6cKjY35HipRFQpFLxBGnfPbJysAXDNPx6ZkfcecFnlYKKUo4/
qY6d6tNBQ5qweAwgSapj+PSdWrIECorMyI5GojI7s1xgsXieIBgcaCk4qvw1y9zbm16DW4SwgBd0
8t3djeaLhSt/6UpLDELt93aHcQZRDBujwoM7VMCzBuvKX2wq+fcq+8UJwMccOX97iuwAQggMoIZX
KSB0iZwWiCfcajBCAFN3uRx/MD2YikSQ/KmrdBoHeWq4IY2DF39XCszDQZEVtQf/3cbY0K1c+Fal
cMaeVEsmW53cOtHVnNS+lP34MuclNApuVcSqTFqadmvpQi9zR44K32WVoKmFqTf/LwyKVM1ur57I
Mc5BrgkXQofyDjrCN0C03b/UVO2oEiu0Ch0Yz4cD1SgrwmipDScZCOF6zRwyRzj9WUJIpxpPC+ss
/qjMpqKAsm9OmKE0x6a9IXo3rlIbKnyGBgnnsLyDwrseVG9WHt387iDggrkloi2tsUoX1oUwfzEz
OnGRStlKtlJvXgzmZC2RlClAlfqltwrkxaXtFiV0LSlxBtCh/FB7KVU8nn1m510+nW7E00eAqGq7
gIx7UAVznSOmLqTx2hiGSyztc7qdUVeKQs5RKP3FxZ1cEdfRwXRb42KIVoLmOTmWsmQI8nx64PU/
mYM6/9aNJVK9jhhEYe6XqhvBVEvIE9GpXYy/Y6S9kTYuNtaJby5OFpqvWD2RwaXc7mWOgbJGIuwN
UReIqdpMAKXqjyMVUF+5+SRx6w+RtnoxVicUTEpxy45OFFAelWWh0JUohnPUdbFTF2f4CYZACfBX
0for/kS/1Dui4i06XAZMZNXedBLJJ43kqZZUumXzlGXOyybPIWqzAGwPluGeoQwB+nqHYn3Q2LHd
1S5Hq2O7Qa9xTh6VXRUNNGt+V8/K/xrC0CbX97oC3U/pfdBNztb+hEjcoSs5oAoa6xB5DdqRDxFa
vKUuvgYSvFT6KWC8gQLl1J0ulsKd96DOHnbzq/ZcCKX1J69dxX9X+KTH/Y9FAdltaQoO4PPNbpFk
IFpMyEPhZ214hh9xR6RqEO81Ik2FU8l24AalXELKER4zsHIt/+SWlOQ1Z4npeEpvTL8BlBuVLX8k
1gbV78fkhBNBIsuETmRDTuzpGm08JtEWtF6eSlBCFHfL3mPVe221fNIEs3eXt12AFIBb/6Wzrb/D
WGllu/oJpzclFQgYD4AM2sP9t2xvwqA70JUvw1mOF5hNnZWOH4Ej4uVN6x2gQ9Fg/QHMVU9fIFVR
95FTvkoUQnxjYFTOEY66YySBRG6sPlnNJBhBcjSszEz+fqbe+mUgjrntP2vXs7iAghaCsT6K0aBO
jvuz6UUWViCSjzD/WJ3ipcMdVwD6EGyBNlEbxCJy3SBk27cYoeA9J7nx96CRlsWBkBAii0K0N/eT
vuySw7ZvPhT7X60F1M+wsRfDvMuwWwaIWkdfNfD1yGYPwTp3wThbi9AE8wYZczoZ8stoBN2gIm+J
5cb8HVQHCTgReG0EUE3OgFiuQv7DsMgmK9wJu648kkhDCgsUPeaYCFpK6amPe4zUXF/Ujj9Z3N+0
6iQ5+Mh3yLUSO9Nk69Sit24Hs3/p8JAVfe+WcjBF3epVJ7RHMW0CpcNhALZFORYj8pbSc/Kb4/5j
Q/pLPRowjZ9l88WeZRsTlliyB/oG0/uJzEDb0fdkYJqlZYBMnAA47IqIjyGW6aodCCmeyl0f7cHt
zwnNCt1n1ZHIjjWAE6pUL547WQpT+FjaJrYMPdhpmnqt66vWDdLeQdTCUKoPULwjt+LAqDIrMY1G
jO9ur9CsmAdwSpjfpnd8Pb966+9wCfXMGu47l8hdGrqPWuZ0Oqq34GCKrlzAsde9qhk1PRmhrHgI
oSyMNvg82KDgIH6r/Ca38/KzLVltkxsemEYNInvv5sfYWH5wTV+/RXA6p7ahmAucdtTOJagF/dry
WZHrjMCzuaG+IV8sEo3dTs5vVzoTHPhbC9/3HuFzbpm3P++xmv6qwhI82GYxdZWN+TR7M8Bo5Ei8
7YAV3sVQu6TO/f/75wQo3uytkhTZ9bYVYoUlUNo5v0GGpOtBbfcH06M5NEwpl6PH1/sxG8Z6e0oj
fgqrSSjaaGWf9EphmABGfuFycuFUtVQHoeEx2W/SjoeiybykhJddtgpST4jorFWHyQA53eItQSdJ
xvQxrEnOQ3fqQ+Ce2716MG/LPoxh7/oCS67Ql29OVbDcAt4yJUl4f7ckkVEApSDOhKyhRuvtfAwY
nkZ3E1na6tbsBDefEj2vbqJoklcv5lTvD/cDfjum8sUEZrIc1tjEdCq5AZiWmQS7nkfNtQRwsDiY
SllkqXSiZFibYxKZswEtqikfY8c8nraX7ud7LEFFn7V1U5Z4eVhOc6FgzsS84w2L1hF9Ugx9gAJ/
G6Xfw+sjBtjkjYDlAkfeNAZQlEt+XCHSGtZOGTYvZPk00gR2/CKjjiLH43ozG7wklV5VLlvkNLEh
t4bPHWkKQ67X7xwfQEEek9mDPwdRxgpQUFocqOVqNs/P+pPq/crbfrICoQvOPjo5RtKk2AQma7fO
M7q5af1tNmGX4m3JTquoGFnc/ttjJaOIHhF9UJV9iJvKi/12Ivm8ndTpvXgZEu4oGmnLz/Iv93ru
zyZ6gGtz3TC3JKs0BRTGjMAIDYm/MHpcM2bR1qQqDvhxF5TESAwPOG0TKHhAQYX9lzkwwxs89UKF
5poVU5+k/Q8KbNp5EAfmglui3rjvCtBX619FOv6kpjXiHHVZ/VDRXgdEXVEecoqp+6xtnL66HvlD
amQYzxbiz/LHhwRvawgE1qPELU55jAY0HninsD7Q/h15H742BtWFXC0r7+OXOP2qCc9yGQx9gA0p
sUob/SrNX+91R2Mg/sOnAvRch9RsQMIkXfDcD8hoySavvZ1rW2X79wtGj7Ym22gVNr9zn7FSF3ii
5EWz+yFg4jWUq3O1cLiqmkyTf7JSV8SuuiIq+UIjqCuD9KoyNV2RjPuwbzDujdcrQgGTtjmc2paw
EsGogt4hBSg5Kykfx2d1lCWKvOO4mqaJLnPMkZafLPj8CgiHorDQl85+td/hbhjnVTXyh9idsBw5
CVfLqe0aWsDeX/vPgMYg9R34y8pbjLezjTkqnDWKTsMU3kn9jqUCkABqvXzRY8pT8CYm4+Ivn0kN
X6lU6nPGurcgdsDaHOvDETgDeAYRNgr7/WRAN5JVKrH0ajSrzDyD0i0uX8lWxlX1HWTE01z1CgzQ
l+K9l9+fQHQIfupBi7J9FYZQ9h/eMRMYeOl4KV0AONUrZ7RuVhkc4v6XS1EDrkHPWnrVXeHzF79S
6xkMdkyTh/0Ftq+Cf24wQWce2I+P/I9ftPks5kaA3fcm//r9JPqth0UJCPb1O12jIOGQHT+SaMxS
aD2bYBW2a2dN19hbXjGlUJt7Edxl2G2VLJeRyuGvHVnCZkk0dVu+fzrkH6IHB6s/JbpOBXQbg/co
22t3g9fK+Fp2AcPJ3ePlpDlWGCkddvAIOUYGfSfcrWOTifu3zivARFFxZaHcDYx/TKPBTcg7YV7X
vIGGPEiZEQQspTn8o/+fwzZEeEEHzs9T/K34JlwlNHnLVDlEvGdfSUkYoLAEkIBIjb4qN4pQdJCr
XETZo72GqpGFZZbtuHQH+8sLSMbig0yevUBDSM4JRsWlWjgY7hpc/WHo6YvbPmB31BODuirkD4C7
fEiA5QhC/O2fdZhBSK1qtEe8/SfQoP0Hdi+mld3+yFcOInUvQKDTeCDGsMI7XJuHDacj9a0Q72uU
IiCnUcwM3Gvi9FjPurBslfueZLvZpZ4pbFccE7iDRBjLY0mBR7kg1Pk0EtlZN91GGQY6Pqs1X7aR
YK27mbAh/5waFkOyHBuON9Cfqxmjg0X9q79bB60YoIPPRO5Gmk5z6+ysfpJBz4l92DQIiy+qi4A1
ZaBUCpYGxPd3WZKdWvEOckOHOlaXdtGYWAhLjzv43atbE6AsU9zQMTGkLCh4ZB4bq0SJ79vX1Nq7
1vCSmdarh14RPYeYIGU6ivzdDJn3WfWCzMfHa0mk9KCnBk1mV1zBtHef1/xFoglBt6UjyR1ZlW3M
eYfARSi63B1XGLxSMZygD3aFBJU1alTtgIfD+9NeQv8vNjNCtoD+oczMxBiVLNiG4Ec8TJIBL5gr
a1EnWWYdKy7IOGyVZxipMqZ3FQYDZhXU6DxdYbhhVeDHaeeCH+M5yLvdon1KZZViFhXpjZsXy4hn
wvxvjkCdP9FM3a5E8oAxNS9xoTZPgpp7nd42lF80IlV4IdqyVwk352cXy+Rrmio8MLCfzUqMEUFQ
Sozv9mb6uSGkvmElhJfVQojiABjI5HCTOmsEKGkUGbvKQ795K7KoqydIAwf7oqOVe3dD34i1/zkq
npVygUTCCVONLADxyAybd243cZs1suQRXKoewl9eA7NLwcWbfNfFDHaMSUYihKMsAgUmMdoEepMT
aXF3ROe4Uemt/37qNkKuQQzlaWueCgb+P+VYy++fkkhQjFvVGq2ZuEOIYS8QzVFUNLy1jaLV0KwE
36buCRZ2bo+ynXoxQGoRgLObZqFMyah+yYdTmYw0gPRbTt02P17mElmfXl6PNwRj2YcvgW5EFSBg
7F2Pq4Gvs9HIY2Dgt2rq8OD6AbN4mEq0YtY8cSnwiYMyyRP+05NiEcPSKv/6ropcV5wuhS9zvc/Q
62OvVgY97mBOEleAjkkETq5KOy/xQaC/LfOrZaGpIh+EcAy/B0Tr3qx7LhwVPSDl6BQ7hkalYnBs
InYnC3VWZez672jiRTbb9YeTuOakbnZBcUIfVPsZ3vUyQsYQBGvp44DKd8pe0LBB2ywCorxXVOR4
ddN3c3rPZyyEwAqIJ3/zTokcyGM9NIdeb82Ktg7khGXD8bN+Purar4+gcc54RoUXLoKsKWKzmrOc
Txc++8nPBpMzpryg85wG6QbG5/+Nu/hJ6ttUGR1dX6OOQp5rSZxUxiWCXUDRrdxJUqXu9V7YwYwf
+BZqXtmnBzlRcvRYfN+qOo61+gXxeNKy57K/b10nP/83aBD3Fg5lMAlez494qbfG579jtaWh+WMy
SSYVr64QyFeWm7Rywn+tV0JA8rUDPZgtRi8rc3RJffWqemEtM667a+ECG28FUUN6WbbN+cwAScxE
IJw/xD8W6zanyGexLA9TU5Mrp0RnG6UbCz2xE4GD49hr7O/Rmt5RTaWJ9lUYgmnH+13B0eEZbndX
+zJ/I1dyq538Zw9JZ5voRZzUnF+UbXEqhP3oqye3+oE6szZ/Dk7cwx8Puz9R9so7y3su1YmR5L/X
jNU1BwU+LE787sjNTXFNMu7GXu6EViPrhSW2oGvw2dzZRC6Q7xITc/mkUqbuXlG2xvLMLW4aMDdR
UUA2TWkpvk4sLbxcSswGVgtacw9+cXee/r1Phkpk0zNbVnASmi6diQ94yxF4OKmgXhle2NFWfh9e
XvtHrgXZ1GbKUJm6wvyIwm7eCTUejje0QFeRmegMOGCLzCpTe0XjykDqANXRVHP2v2RDCcBA3g7q
ah4W+4VaMoS557rGnqgM6++XT4W0cYviccq4U7Yv9Q6cRwpT0E2PxhE8fA+L4Z/ttGWs1t+sa3y7
YFQuT0AAZYOvycTQKKOoVVB+nNERuv0N6V0bWUeAmdJLgvG1QM79l+Tzg47bzBtO5ABmpcdL56yz
ymTDkhMYrwF/fYMGiQAx6JQ0KIGly512f/rmneA00DGf+7izGm9NJIbKo96a4ALzC6mXG/SqvBVH
FfP78SkV6zUEAfJkR7t6XOvBj7Ny5e3yY9BrBBrOfvN4ahIvmXwawY+Y+XdMnMXOhVdWi348H128
xXjJpdTja6Kcz6yrwYIFgQsZoa2ymZbDv+AiLKsjnB9PGgYCLevNTxrDcrgi/OEo3XnzOefxP54L
w3W9B7eScY+2CdTkNdwmRyn61W+pitgb0L76NLibLlEp/udGvU437D7YG3CDrRJiCjNc8H7Lf6IQ
bzWQUUgP4RnHa+7XHfYib/TiiJTQtihHfl1iOD08ft9P69z3ZTDu0mmvmPde2J1ZPs7Cyc76UwVe
ybL6Z+/RgTDrTKGby9CvE+F5Pj0isUoyHU8IG3h17evhNo7Bh/Himh4BLoeDf1HSaxu3frk75Ssz
dA+t4opsEoXKnjb5XYPm+OBJM8EwOmWa/9P1rJO9wo5ZQTDvY21F7P46TgleSJNZ7+P3RyhHx0kz
OszGlFHCnrah33JqtK6t3PxoJLXcEIfRE+6Oeubpy4jfAb9yDclCoQ6UnV/QxDU3nq6qlFsqzria
thp+ec+mRuNYOqcWj7LrOwwbbp2JrKDQzSKSvqv8YYqKN93rjirChPSwR2SgEUrcQIROJ1gx6T3c
vthVzOEr+o+C4N4zYdvEq68o3BS9WZ79MsCpSwTVsRpdBLeuZ6py2uI0i/Yz9ildQHQuLdBpRbv+
qVmtB7SoBzI778KP/wwb6ibIG6L42G9fT8YKQLXw1lJuCN9QysaUNwfj3gsv8knNNy1wlMctDlyN
S8oDPjW1sreuoO0JpUVzLVyRRj1nv/rzhbD5gdxB+IX8e6b2gJpkWVRcF+cQDVOJP/naJiPD0q6V
mlzgyf4Wy1NJIhpoUCUIZ0nPj2l6/XB/6LFK85Rx+JMXLRDTO45AZAmgDsgu9WZX5+9czfz6Y09K
h6pkA/8qBb1Xnp79d48pXfRtc7g5xJiGed5Xg+XfB04bbxC+p1pgGBqj0VPiRWanrZSY8A39eihe
nIEDszl5172a2SYvE/FcvL+PILZiV9nnP0/q9kvT6NTND9xG4TbX58KxTo8Ou07QggNz8U5/SYjj
+TKS5lZKjOQSskuWb+gE81XB25oajfTl0TTmx1peHfaz7K1c2OMxE0ohgTjwOi8HHbDamLCzr3gm
NSba49q1T2tehr+IguuC0QGDxgJJlkrhYZjUQOWtXyN7WkePP74buybUZIewiI0554KfyxRn3yxD
7RXL9uNj8SC76kZQ7IVk2p6xyEAN4OGSdAqqkiDUb8Tbk3qdvNZ9colSubJoL1DVEC0pbtyRx1xr
IrwEYo2rEt+kratlrbruuw/Ig2fO0wvxcd6PIu+QH7kGb4HRQ/slK/Kzi8MofBXdoUMjIQe6i2iU
2uDSg9VhvCDHTlpXli9Foh0PBeVdDHFD4JzLhNJlBLFzlmMkKczTOaYDXXma44g8cEFWGKd2N3/2
XxFpuYhcG1eQj/iKzUslvrFFwvFWCZCd1h1lfvHUWZrblWifqAMZGh6Q9qmW2uykoFl0BmVtXBZd
H2OuAPgKgCszZIlXv7Ww8jA/3bnluBz71G9O4KQi1DiSJtweMOptyHQvAS2U1CzFJTRB6uKOa1NQ
4P7eC9ReQKgQHvpyY+htzJWphGYAqbYuJyeZSCHSLyFZ7foPq8tWQ7tu0XqiZPsWZOiZQ6SDuo2w
OnH+5Lmyz1JruNLe919fueMzCa/mEsYmqjYale836b8Gce9kKkzOrtP0e08Fj3yIvHdeCAyBnXZu
rxExtmvhHi/5lG/9EROPX4u4uftAh4y62Y4djCAmAFc+BK1MUKj8ouWz0aLaCawNQMhknGr2Pu68
RAILAxCl/Z13J489LEaezN7GQQR6EZS6SBiSHMSngdVTCHxiHnp6BRrlKSDSl3MP5nOXZrzY4nGd
DxyQ0TWiq5OrPiuQHAztnIzohvCN5yXSvt0eRwMPb9CkFoDZYRe+Sg49C7uE/jC0d4/4zIbf80Dt
JiW7He3vkjaOPOgboqzr9fLczy+lWKu+jHpBfmH/6wclkOYh6C58JVpiNT3h2w83tbwqQpByxXpP
jV+EpfMmbRTtz/bK6InziOdsmNRGyNvG4vrrirOEB6GP2yX/Yaho+p5iijWWU1ojZZwmuahswMx0
ScWYmdG3s/k0GkvaIpIQ108kFJb66d9/HFs54H8/HnDH2GUYMYJjysQ01/Sppdg4I3yn6NKcx3ej
BVuyjm0BVnfS0xXTitdfTuEyoHwl/pYXLGcVhbwLnTUNr7BMrEI0KklRxDV9DnxhmGGVVuXUD1Dj
H7Zsbk5fwVOfvbEr9zjfpJSU2xoe/jT55ZtZl3ubd0y3Ej0fkHSnCVZioE4vjjmkWTD3ZSA8Jfes
RqH7yTV+3Fy0jrEBG8h6VK9L5/Q0trQzOHlHJbCKhobNeLl0DVu/KsBf5SWvfFwgHWTeQZGysM7D
SSViEGJOS3B+JxN4aPXqxi3M5yoBhehWRFnIT+Oi/hNmsbR2djU8d7IAVBqaaHJPAvM4AdLh6xcB
1ZQQH2WAuchvOw+7y/27+D9CfKK0XMnLlixeZh7SinE5mjXfPcX5V4coPUWE0/4/foumWq7HezQo
ISzB/Sh6j6upu7IXvjo/Y3jgprSaJHFxPmlWKuHYMZ70iNeCvN+n1Ft35yQ3fWJyLrcJAsjt6fpO
3SHXod9QN5I0LHCntcughv6U7se5guCmpd0DI7iMOE96ktdcjCcg3MXjR4YN7gUIqQ803vu25v9P
hNGxX4AfAqqpl21mT4ej0sHTfQSVKIUH87uU1rMowkSw1CWdNd0VTatU+cd5bU9DLye1TBpkdtV/
7Hteq5m5HZcrcEp44ET23LBjQOi/wg1xndOEAuYI6vAM6+mXlvDXWt7o83pyMuD7TuTY3kg+eHE4
G91ZFTVBdyFvOVXOpDkhZ2mHPySrfb6yHduPUnYd0KUISIius+x0YFTNPXyXfqSFd4RtLOvRGg+r
Z3zxK8Ao2zkW1g6ZQiDgsGemjD++aMi8hfdF/JTtYAdTJ3t8KiEQSauvRtR85HezM9Bnywj0X+7i
2Ng3zFr22BCK3C4nD0XS+Z4iSf46Os3zD1BD9GlLqHtCZh4bNRxZU4kbtCmZU2w5buzIWp+VSJKw
w9/+24JJFYHwe8x0bx8Sw3ruUC4sO450ShABqbNQPpBtkS9pcZdbBttdeZw397qHKSIgbkxmhT12
0jkb0M+yNSc1jc3Im8yGCiTkNPjj3kfXvFie1P4ECk1STdwjMoh4SOrBDPSMl0r+4TQCjJS5c9E7
ty5nMN6mBMOwkWkSqC+JPVpaza6mJx1flVtLgQdrfF5Flo3bMoT1eD+NVsz1fcdsT1viAqdqNyij
TjJ+jqsNgeyNA4Xbq9u15h9MOe95DqRTlMH5DQiPmyic8rEuPoRFebwssRcj2W8EvCjGNdgrQDWE
54kP8bcwM/eUAapmWIhbxtr+A/nRdnq+LD9eZR+dFya2ikOKSDo6blAIBX5P7dAxcmHi1sa0jS48
Lqq92VGNhOk0tSDuTRKo/eLPYQRUTMr45P5xzYzEVx5PTq8XOZPL6YV6PpzAkhZeFGNI7jAsZv2F
tJfu5PDXTcJSINonI7Gg8KBP4nzExwL38k4Y/ytAzaMFFvEeXR4b9DioLSrYrH30N4KUTVqDrjis
U7ctYNXmN5+vvsnsOgBsyoLW8m53kJM0rPy68fb+QRe3Pkl36lKBA45WxSB+8c3PX1Z4vuk/1OOA
pkTn4/dJUPM0nIC0CJNcK2fZhsmviNmwrhV6nES9n002a5g2odQkp0UHxBXAwOwY57vjPG5y5TGL
2VDYtnZLuqEah3zpE98ecg2kk/JAuwt1oGivMBHGomVf2nMSkV5WDbOssiQuaEChYb9iS2qDvdS/
Fmghc/eKQYAz8ZCQ7AuL2AshJuDUGLWkx/UpYVvRK2W793ucYQwZJQjwkY728Hi9c+VQsyavwkdN
8dkTIvYjh8TPRIwItJBoHbokQWgUou38raZPsV03Oi8h9TKQiuPxIQ8YJ0M4apli80cmwtB8AJDY
OSZ3+XqV1E9W71rqMrxDbYz4DeQ6N4IV3L5dgTP/Rw0YFjeHC3lPTpzX5I6DJc2PzFB9aXs3hpDH
IokEPBYukHn17k3H53gPYH2AYZUrcaP5I4ss5la7xmyogeGSkhbsQmVYjEk77o6GtdjGkaUmyPsN
g2rqpKVm9St2GUPajrt7w9IIu80oN+3z5IxG5Hc6bj6spBbs8QvCGrCI47xs6LoCTAjPPKK0rqe/
QtSfjx2fOWwBld82kkHxTXq/KgugfjtdeCIW9GX47mQzIymaDk6m5XbgNFKmgPODRzxKMZopqBqB
L+J2cS3vDlSmS97isiSozHQBZxzsQguzoUaTH1YM3dQYnBO0iQWc1PFywEErlVOvtvi0JYnFjhrY
y6G2TU9rFbiB8bEINXpgV49H11w1G6BHJfuNMRfTdrbAeOgIGrbcBa6ocqGzl+13lHkELLUU9o6J
HWRfmo4qZd2yuEbHtNTFiWCmCeAklluqgH2WbxTt3FVpCA+PiE5YwGyaNAVTSKp8t3kkRvldMB+9
BcZMkjJRMyfyxip6JHjE7K4L+NvoYTGIO/cvvDnPUicQKX55ZcfJlI0yTWjk3nrbM32SYj7dUtuy
/HO0X2rswQNvSzjRc5gl+zMLAOlQv2cs6wwZZn47Eg/kvQvLQjzuZ6CIzk1QeJpHXx6ny6rQK+86
8iu4tegNzjALc5rZBVUq7xsqlkM00IEIJJdbA2G+IlU3o5ITcofBRZJe6wYOa4EvCEytmR/8aMzo
borDzvCtqD/0EO0zBTRhHE9Q4uZUMp4X/f3mwercys0gfiUjReproG/DkQ0+0jt3IlZKX2nuGAqP
rvy37Q7Z8uYwsYqMj7gZyIeQ91hnvbwgWJzmRh2IqzQuJdDOAUBS/cH1M7co4XiE74180IhrJg/F
Sv4clhjN3htefJ+I7WwaCYAiJ9q53wztsZUG1FzOxzIqpa1gJB1C5utG5gU8RV6ErjIGlcxRBmDC
klOTLWecvFnqae5w3tVK7Yz8/PWX5AWT67D8tlvQtCsyOBuAcwOPiDou9/tDCa/t/2c0LbCsatFP
Wio7AWMmOsdcmfbTTluFnL5azW1JzVKp4++UEnxv2Zc38j+fPqhuQoKrLaLZIEiCePryL5Bz3RdJ
ESXwvmA8uMhfN6SRZLNWp+A1AkKAxTPWxSPlJDIjaG8anwIE9hWIsfizayMNEGVtvLRLP3Uhzwcj
TtmL5dcERWBvAxQZwblCPweNPJTUkMAQJGtLj/lZN30SdVlQzwA9qgEiQklThlxGGWcCHMPukFuk
RlhC7qWUbguNKlYmZTkLH6ds4cG+f6n7fTEqCpkJZte9DFkKWs+fvimMLHQ5d2U0RqvT68ct+qaR
5oQS+HypujyGpC1Ys8PI0VCCY4dgu4HA0pfalpTo5zXTGScjoZvcRYTEvlXzhC608VUvJ/NcOtpV
kxO82CJnaNeSBI6w3FYlBp9ebJVX1fCMoSymX0w8l0ZwxsJv/HB669ZKo3weGzyesE8Q2m52DOgX
vbIu/kFzNHukzsq+GW8eOqAs3xf1oIgUW6oT0/oN3mZ6NLebUcj8SiqbTFdDFOvL+bOChPlAp9Q5
F8Ra6oWiZe3yIX4QvgQUdxWoOqydLzfEl9JsLh1bVVchoqd7Wrvm1+XO0r3UNYFxkGNY4qdMXHCp
HnvuIrsXLxa/hOO+bepcQv2fJAoWcm86T0sSOt6sf0maTzg4i/zb5JwxA0ws9F1RfjoYoUbQ0wAb
MdQQEvgYGmEIg5X8SQ5qRUl1GHkl24rEWxAO8alafXNZn08A4Beb5a6IB0OZ8ptiIzM3le74WN9y
IPXOy23FDBRgM9fQpW5S4Gnwi0F2p+DLD2DYZIB4rzZ+xkYoKEyUlZ2q8Ho17fGHUVdBTRR8BtvN
LPqll0TK61ii5LsR66PfCzBqQU4esD9EkiniqPpHmFBIegBiOfwOnd1id86db9sI/v3awhsTbG+Q
0VCXtEe0L9mr97FJnI6fx2CKVL6CVV51z+evfIV0vBHog+lsKeM+H3n1lF+1akvRI05yGiuHMI6z
9jAuiiEKfvE0TDPKZ8FyNKtvtFjqyCicA7FRcmolM1oT3+TsNL27/NPG/Z4A3PK7mWoXD5com8t+
pWLT1Rreaye+mKRyNnggt4poQc90txTqzFOYkicPzsLGa3WhH35DpRZgExmCMrpN85dIXDH/I9DW
u++mqDskOiyIeswrT+DxkBJqEvNOHARrHO6yHJgnQ+7ewpVtxJIubaKdA5pGJU3KZ+fI76zKoMFR
5wdQ/THrzvhLLoARfgvkzKEdOBAGFBnhZuYhh8l1xZfZNNKiLMmSGP+OyJE8lsVDys2/oLkVZ/ZT
ILgaFsF0/utyHJw0OMVxAgYTJhVH9ekstEF4XZGwGhemfONtjV51y+NeSKwdJL1jjQl4XhyfIyyy
oLx/UAUGiQBMJofyV22nJa5/ClwbCF4SSLuiGW8ZKSPC4x36jXN1bILEmwhSKvoxFLeZQU7DbhX2
tUh78gW/RBYeeuQi4Hw1GsPH0aPLA1pB4MnNSgIy8gEp21PhLViNCGa9/8iA4qZmDLyMggJy3cuE
pSVlzTHkns2/bdmR9Dg19xeGcN0u1vG5Ym846FIYrIfbyX9xZADvQYlsXt71RfUFjJKQ2Tpr6Bde
KmL5pq0yyFO1BH9JzGLVt0y/oopG3k9Zy3r/98FWuwKWKmiAu3fpxY2WefxDSMUGBhx9Vxub4Hpg
xRThtplBlRIWqlu5keu/DTlkHtqleANpDlqd59AcB1s5Ve+NYWfE/PdjH7D4pGW5LpGg0XWI7FFK
13RPw3aYsY8w0n/gPUS0f9fKfiFGPTxxy+VuIT9IMMVDkyz3syotpePmb1/1fh465qxl2UONE6HX
oHSAENWgmWiMpijC6wUblzOEOmd2NTltCGsJLr3XFB7TgOhHyOfuVQgxXkNQTxzMfk2XVd6f79K0
kOc4hb6qyUH59irf8OnBh/oYvt7d/hbgE1A4Ixo17D+Z7eqaWf2QiM3f+RDnUPKHg/pXHEKtJ8Bs
ipKaMBmFnmqL3cEvpqW59L1M13xei/GCkVbXrDcCS+Ujed9Yl8B4FYKclwWSFR/b16M2B+Ju3hcN
SBL3kUF/Lh2f2zjienTX4mk0pN5LmVh7XPhz8RJuUONTK5uR6tD+6LBgzShuM1QVlXERy/vh6LbW
TrlAuz5i+OKLmSc1Gh4sfEJixH6dYrL6R75sdbGsYFCoMW0yMlD/JxTd6enxKtJuX2/tAYvZQmfu
MIPn1e1CSvsEHWNIcg/id3XAD3mYhZ9Y2HCGnaj2jQG7ubjd41uwfPe1vjm7TWA0toDSmOo2h+vc
+M+9GH9Aan/W3IIm7605etyFLvj5Y4IaD6euFdHTSDTy6P/PZsALwNJmJ4b0Y5rTDODYbDAODEtV
OgbIt607K6oHzyRdWl1CIr9I5vUsb1VoVEI4/h6PJ5Am+caST9Eq/1hvqeFhR8lPd2oA7xgYMOCa
ERE5MOdigDmupc5IsjyJcldgWo62YtwshnSSpHS4yh8whvFLqvTQk6aQvPlwemz/GvRouwdVFCb0
gd/8yJwMyuhQhtqBqRJeOZrzJFgJL50ixZPg5dYIGvXxT3AY5hN0Qo7xB+BGLOrW8fThSPQL/okN
DmLByDzZJb55zeEnO0SFMPuas+NKcFrPl/Rllx2OeYyJSOSoUQiPHZdBjH7q8EXQxWNmKCxF4juW
E4iTqjED+CK0r5DveEzA8XnIiW+fiKqKJ7OUZXcqXxtv6ZYgxcgn1JJAr1EjGr4cDvcCkwEAC3kY
SevTBsQhKYU8EQ4Mf7qnEoIBKUpLCRAoDLGgD4tw7QNeDfF+/hv5CcbMaXgVtIKcxszPvSUioimx
dTWAYyaFYiNOdqcOuN2Ac2MhjFzkXRNhiNQOhBjIkcznn8bA+hEuWtpLb1kimHTzeEC2VsHId3KQ
WQWc7AfeL1jcHh1qJBfPJ1B3ugg5v6P0nMkiQHWsL5WuTy90AR1OhBeC/yEv6I74IzxrD60BdHzY
0t9YOS9v5BWgl4elDU8Y/tCi8rPkDZwZ2yAc/5G2sHmpAVkKBVa7nkAlrgmEikEy5dZNMzPLN+Ak
H6mdBFU31pAt4x9iExxKgk+RRT4rc09nfBN4GEd1AaQCBy2Sh3tEeFL7yrKdJVy+Hmgm/CZoIZjH
QMiaUQAO8nlSc8fkTNp+FBjbPhfVRzdZJbBqOfsbfHxGEGV6OlftYwJoeHj75BWtQ2A+7338t0aw
jWMVJVVHtV3HrexXEJJ1GgbeWwyFrtklbHQtgOPwmpq/R6ugaWXl/0oQ1vo5W5pdzL3w0uMHcS2Q
rx30FObcKJaYWQ241XAZdtZZtSiYZL7yypbYVttMeU2iwj589f7it+bPXS7CWw9dcIUjl90ewf0u
tB27iwqDax4LtPRzC13RbWrlkwP0rVGX08eGgL9yhwcWnVG3D1VXVH6WClyAysBZpxprDEE/HkW4
biXl0JRihp3wSBP1uBWldsilupYfEsZE1BWdeh85gDsrP3zkdJe3PG+BrnuTUjGiiNnUgfuWPvOA
fAnMx3MJtzpQXciPN0KB6OL6oZzQMFsmruJujKYgXFuOA7dUxNvOVddhye+LL9lFVZECe7il/kUt
2Rg0mQO8MvknVVpl282CebnCEeqZb1MIEUdEvKWn8DAosG946I+VPFLoPsvMRnYfy++x3NnkcmzT
app2aSA36mtWbN7/3T1vWlaz8IK9wV/SXTwOtUNE+Q/byrMIqEBez0oJ8z1BdxvTZ863axup81jb
7k8sK+xeA9xkvQEZL1f2RL04cWMBaTeRxPFWjtHzN5wgjdV4fhytLY8fAApXOXOE0Gj4pXvCh+x1
2ImxrpLUPOmw8xfmB1IlCwM2hth5pe+AldL4xLrDG03SX+Ex2/u7zUScY5b+cv1LLpp5GWkcTENp
Q2B8eaooQ7P1PL+TlruMKP8xSOd+24l/8cJYyOcwO7nLxbXfnsKrjpIN65YpASan52v1WNYVORsG
znRDJV5zohkmPxW6bxMzzZuH36sowClUCJYeWYgkemi1cFx0w126Z+ZYquEbUoXHELoG+QwGwSUK
2VEppSJAY+PGkJsTOMnsNONnXq98kwnEAt/HW7Fs3JgLs76LAXg7qUBv/G6zhS/GlHljyXw8Dk2m
1to1vr+oqzopRDTPUQpLb92swjkAIj9wEritV7CtHSYR2E+X/vDpaM5xJ+LfIXTH1I4zD8M/q2n9
Q97FCtIKNti9964VD0Jf1MVjE/X2nkIkouMpxWBY0VoaFGxi02dhKpsmOULeY90nG0/lADN3RrnM
Uc5rzSKfnrYJ8kt3fQ6YlLq9d4imPgVJ1dxFz1TSk6ARhdoUKC2kTWgCAX018UySn/klFXdcW6q9
GKBB0L3+xVNcTLshgeS/mKL3WO2qK7MQCqE7eYInruiGHMKzuJ/uFPNgXEGDkAl86Ce1B5BAUZHO
NFpkVYO3zw1t8XXASatHHUvN4RKBNF2v/ZHHOyuvnSTTNPn1/oPR/EEYVhXUcg5Zvq1zUSxPNo5j
0nFQIxpCXSIZaqutQPZPqYTrJ1xe2lSkor8v8x5Q18KzAuBtDpTr4Q7HwpnBaJYMz0iXClIeJUqB
yazXoivFA0p2tNvrqfV1Ss/S6+ge5mJWGWBqH6WLbDicOaGa0xn4oSGD7LlyXdzD/8h5tIE0t8eh
YaFEM3PkxAiajSzh7kEQ2/RFHAWrKQvtiLmI/sHlr69MF9o1GajHmTSrI9488hW9aXgYg7y9b6s/
W5E0HZOYqSNuM9zTByL/FqNQo4/nTu+9LCAKEuBrVjzXjz5LMRvH1R7NtXze80XfSgKuRZfFWy34
TTH1xJ1if8zWwA4Z7iHrAb2FBxbcfMi4dZuolTgyn1jONWqlWTWWXQiMBgEfSg2AaEgTlrMp3ftZ
ge2Oh+ea54pkpUwKtfed0yBKTMppWy5LD4GX7huB0VxpwOt7eTcHf/ckOv7NX8uBQa872QhMpqql
keuNWsc2sAHtrmlfPY64HrPHF4K2NedWJFKlM3FnWcOsQJH8LYecjX8F80KZ9QjwNl9ukW8lg+7V
FYMEz+dCxf7Z/huPkwe+R5qVg+Z034bPQOPqP1hallHcdX+R9XcOYzzac6yvlAKbLl4a5FwjPyXm
GlYQcWXvpP+OAyrx0QK6m9fo0aShIitPySP80LdDyKwDHgKS73XLkvtJQGC6gsA1+vwYgtMYCXqG
S2fhaEcjpns09bW3CND/jfR/SKgtFhIAH+axg+f2kJlc2ea5RbePlEZu7lARXEDIiYb6Ff5zjOIL
fCBurVAgtTXrbZQRqNeRgBioFgWRpj/b4A+yvhNs+Eg2psuw/n9rp/ELXPpecT9T7CTkl/GSv2Zb
KLnyDRvRlzF5zqIG5lflfYl1EtSHoiSQhjCgaHxNj+DRkXpHg8O66BtTNOHQR9TmECtX6UwdrFYt
f6kapsR3/T6WRkENtQRvmNJkd/CkiAVGIxPyOWrRI/NI/hO+UUfw10Nm0zRxP3AQgdtGMfv2YWen
GxMaiib1rH+RKzSh5GAcJUlwf6hNbdRa5072o55tuBdlLKrL+HDvxPzorfulLEsPZnSI4khW2qk+
hu08691CCV3mj/s4rWxwvQhwxcfqznxjkx++2oIs9nhhNoafzAwfd9tX8mrMjc8rGJZxud4ydBs4
AOydUrz1yiU6IfcrigJmeAJhZaZEItOgjHxA86XP6nQNy3aCiQScr7G+VtOy+4obf7KwanqprENk
kv56riG69dUtzJBXUrCBcCghNzlgddXGAeyVg9Dl+6GltwlhCw55uRyOslz+307By4QqgY0V33cE
Aw9bkTBU+GWkbycaoxRB1rF7eqM9pD/MUJ/AUE68yOwV1C0TYOv0sfQHTD2kSVFWVFKYF3hynZ+C
ft361RjLZUG8ffr5o/6MQz5q3denSF5RRUCZfkxs5IBYN1t6ijmkBgtNzE1lkyFANhOw2O1CH8H3
QZSK9Nmo+1ORQh4ov+Sxu0GJA3SMqlNBP6roe32zZ8OGNLlLFtDJO31E0XnIy2OGZyTA1v3KmJ+j
uX8dNnO2dmY4NKT0OvNNJgfi/K032aXn+SRuuzCoPeiMo4iu/RybsEIHNGOmAj1C7IYqyEq95jE9
vJayy9BYSEPPFPcS3uN9BBSOaBcndNNNNuPL1gWJzS6wbfkZytJXzuljegN6lyvcdu1NiMrzlq/3
mMtXxdqVZPlPOmD2pL9q7alQrPJHjiLhKvthHCPHJptkHYuCZ2Pul5YwH1fL9/p04WxZTYzXQtL7
/IBk6P1fgqOlQufodcJszQiKBIrttrnGY3OlNLlEHqpQFCyL6c3hM749YvfQ+8i8XJCbfCv89MxN
qr76SgL0OcrMNUbKYDil2YDDn00OKuaQAYQ34nQoTI3ej1V5u+DUsRoFPDc2zipinoBkiDxm5Lpl
2CWvX4y8WyUDSmzzWctQKRfRRnoGhLoe133yKfqGzyBqrUDc86fnJKcTvX9VgXQZBilXzweznX05
cH9Y2sy9BtXIL5kqgGDhGGzsdMCKMOM1yvp0KthLaHxUIPkkSAsj5yeCpxHmNlwlu+jm9L/Mqzky
DI1l037RIn2FGI+JoDi8M3CdahkrrLwnkqQr6xJTDXpACXNz/h8uSjJnV7XvSwdIelZnL11T/4yF
0cRktLqj0nvniYNd7SsmzUBGvjxe4egr9HD1sjAsBkLh3tBuE0Y7GTESzj92jsTodfweJ3OaUdFn
0vDOtPR0Dh9P9Rr9L9r8FRJR3t0z9OCWZzLRBFoFOR6jKilr759M2L9LlaHYBrKtoIa7oetEUkrx
En5mY3haHeqkKvGv0kpZpEZQ3FbgBvg2988fkEwOtVZIFeOfsgPL9EHUAGNNClsfhLtWU4AptCXo
ljbpjGdLH1aWQuOzZWSLi1t2SdEG1Jel2296ils9qruN910IELP6bR7oywQBhhDLrG+Jv8WLaZgj
8f/qVJpeldb6VIIgnb3NZeUubM6z2BPwZAryrKH9gXczRgtZodjQcsmmSf3QCdILiJkKMO9gGtQs
8YA597S8IIT4BiMAnw+Nm4z8eEBp5EtxAijpWsg5Ydh2mgv9s/awA5EI2pcyws5NEiv2k89Q+jYZ
kN81/YWYvS01io/1GyEwbWBtqRC+uaZnCYkc04OVWcXztNeVql18uK6dS/cJKDQz7RFfX4JtDnR9
6V5BRR04tVVVrT+huodzHtR9AddwJwHSpuxpQFKdDWZlf55RsuLqaGRQw3PRCxikOOA07F/LoMZt
aKu+OMD9ywaMhYhEhuKJG8nJ8a7sl3Q6QCYdL27pqNY1HVeZYIy6YA4RAz46yXC8aWBenCBSP+aZ
kxihg+CsVa7ZrFdlr799vvlV1WsYcPGKBZcohnThOyrloxbtlywqB93zktpUVBp60fLeoLRqeUlV
P55udd7d1Z8At2yeb6850oPzqwfD5QYzRY3abcE8kan0D4wk5Yx5mDPnjnXdBIz0Jpcz5yMnLaIr
/kJ52kZDsp9yVfPJfplP7cVPDJgjqWnZ5c9ntcUWpkzVcKrmN8lOLre9sATTxWASLhJc7yhBI6BB
pUOfq0UiuhMZCwnqSxvTv26Qq6D6nOgtDJYDWIdey9OQB1y/g6WRkQBrhkeaHyjx6c9zoYkjBywc
c8oX7j+aSp7Ddzwmjeru/wLPxC1diQ9HpgVSBvpegvWq4BmmXYe+wr1ZyKP1WAdO1+u3gmQSnkcq
yotu/wN82mIrax3jkRsu3aTXHlECcvmYE1PZio+YJ67wl4bZtRK2rU7TG/frBU+Zhto4702ywIar
09ATPb59fP7hNMnO/Y113GjSen/wDwbhSpKVllCNSTKcBnfucp6y4Gd58Cy5AKJixwcARTmaKD7t
eSB/kxRCoTJLMajiyy3u1qkHn2trD/worcA3SS6zUB41hA27ZflCf04iTOrH7bbjzZXoQT8hN2oO
JUGIUWmNFQl/3aKMf39+FN2Sw3klC+g+LH7M7KWUCUZnS7UABF1erZ6Wcv2C1ireF0xiYNt8yXOM
o4M4ZIxMRzu7fuhMyigH0iQdFEL351U+sl7mfvhE63OAeDxFC5lOXSAS0aYtmBae5Tm8zc8OcuQL
2Ijy5OJ/e6lcpjnwVQvtGjCNZTs2Rm0ryS6E+aJaYuvQPCU3ydXA12ruJrSdx07ST+U84uy6YkEX
BEZIrvm80aPgHTzVzuTk6b4qlbG4DEv1G7QJNXBBydxzJ2FowJF5tTQHOyzeb2zDIRwgYx7ecwQ4
8JZx60K7L3/aZFBlgSxpvijNsvGNTUv/x92Gr92akbJGDJj02Dv8hSylLj7zEOzQ3nOs3n3qL4xL
sEG07NdAfayE/qYN91fYw9qO2hekWu5dUmmq9edAKyDJvVJAzeBSLSzy3imcUVkDOgbGpA1DOzUg
XKIiYKXBR2+scIDo5hZFEei8WzLVynSr7k2Bo5Ug65yqiFAXY2V3TmKg5uAUxddqP0dUDxNZTFaT
j1dWak53cU1p6D9n1nHD5FGjh7rS6NcfgZWAhOiG9DMmZ/iqv+wSuBIWZg1bho2+gdOFMNPFzYgk
AkzpRH5eSqOs8977YfqwwiZVzhCT++hnw9tYCy8+32HSjqKyyM1yrz3K+hQ6/arxK7jxhdcr6rXT
8ALF5iDOdQ3lGDy6iG6IboQ5TcXFSXOhz7MgQslxgEVZlGdAYfXWkKe1y1W6dtcbvVAtXB6dZFrX
TS6cmeEc+pLA4HbFMC5xo1VW62zzGo7Hg2KqkWLlWEiDFDj2SFvIU24CEWr+CmGR7afeMKj7AEIQ
2nuBVM1oGIzd0OvMBoAZyzpJyjTnyG3PNTvsSXJ5RJNkvna2eeLf8sTNqsvDMtMEBIPD94EvhnLO
HdNjMCldr5JqMJcwrVPQf2ZEsdZE147a0EWXHnqe4kcivK1lZWuTiKP+gWwgNtQrmVSdk4GkJf+l
pU6i4w5qH6HjL1c21Xgs6mL9qhUgx7fG+lnGqvm1d52EWvO5VJoSz4XUMu81aXI+XZpmf6vgf18r
nyEXfE2rLE7kfVrS9kD4kN+PgWyzaqUeUqX7ystrnPmD5oE6vq4n4PWzJV/mf3b4OiCmZS+XNjxd
BmplYpDMZkjIsBT8s9VIjeBDnfTl8TkDnpZD3vZlzmndM5+CmZS8SBXfsb99U0D5vt1NRzXvHsO8
GkFLfeq9wL+jHleoRjIAgwZw1Crd782PjUKLp3GHctuVun437cs/pQNtQf4mccr63YqQe0aaMy5l
G6txNDWSpanEifMoNxiAcrVclnXLBlUiDV74phcOMLT1CaDEUqEUM/J0HwlRW/vpy9I/jzRh+pJv
t//j8GEFLqLEN4hG5fByM9M9nhMg/tyk58aLd1aAAp5aJ/AkxEmUlzUEMm1J0q80QFTWG2M39VKI
Ag38C1cAn4XBsegYuo2VgXhn/lPUA3vg6MDc7IlAk9jIW5Rqwht605Da1MTRCwM9TQLV/QxiOTzU
no6JyWFOJaFHjemuE59LuN0wC+7/c9Qw8euPjEzfIdlxML9IowXgfCX+oXCidt/uzAj+qvA+AA5Z
Q8CiJg9dk0tkh7TY/YB/76WS3cnSD5i1nGRVx821iF9aoj5Aj3CpR4z4gZu2xmtqYrivx9Go1f52
gqe0kVaWZjFj07rrRWqNLb1dgQh/C00kFjYS9RC4C7rTWs3pcxlVK5Kmhe2c/IXrxU+fDS9UxyrU
xFehFXdlP9wy13hXipLddETbjARceL9LPti7KSS1l0Q8YCk0QKl8McZKxyJgl+G6JmqcUIj/47fu
vWd35RcEr/aqKwM8AIJ0hMg3NeNB0Q8wZKXASHaiPR+UxfNhxLJuq24ZeUPNPJRgAIRxNr/UDxOf
V9KEbIQuMQO7NO+hSjPSXFzRF041euzQWfz0ESqVO/YC5XX/NKzs2HjonCN8KLm0TBR0JsQ6GW+M
IRB2HRsJ9ONePAa64TNUM6VBaUCVF1jzJeAOmhzEjq8wu1UGlVMB0agx+9ek6+WcsrnxUtwOpmXL
LCzvH0T7gklBsGgmoMWx1nRFKbCR8TfZusjAxgtwtE3DWNAHBxsPmVQRrl2lRlEZu/PIGqzX46yM
T4WJc/k7a30kCmxAaGF9leMnn3+5+dD86Fm818D7Rsj3GGdq0HKDwIk4xBCGKMRIFbqMGTYdIghI
fpCdfKe0xRycJ7tSlyMgFx80YhR4oAVli0jSlJB9ycml43mHTZTpV66N1/R7UL1dbvuqoU0/7BEv
Abdr3Nxb65BwEqLpDZ1CoYjG1V5UOBM7jvRlOLmnei6PjLxI3+JrOUiY00/Dhk30MicHdk2q3NAk
m75Xx4Yokb2Rt8G79undIF8UZz1PXrj0Amck57Q053cPpp6VMFrhyBMWRW1ArIrpWNtLtIY3EiWd
VkByYX4a2BT/WtxoMDvR7uoyWAhJise8WdrhhjbYw2huhOnoAptwI2PceDH/9zr3GkdHs9zSscoZ
PIFS+ErsDfRTE7AplyXRW3Vh82NyLInWtMB4oicEilp4UZVOLKbtI0zNl+WlrZ9590MyHWZFFSlT
GR4kkngsWMPi6p17OxbjMv+AKbSCBCfJVpegp48MJYkQUKWFva81vHoGl6Ou08ZpUG7pXGUKk/HW
GFxfX8nPspm1QFtMNozRTpuCUKvvLze5/yzZgVOJVViKp9VRRrI/TTMQOKWGMPczjRskYkyeG7iL
+ShP6n1dCaCrZGh/ZJiaK0k+D3bPykAsdxzNHcw47jZB4b2KxIAOtm3fFQEib85l/a0FtkQbGl3V
PiRNRE9Y7sacaJaRKA89ruIZ8H9LgofVkzv4wpSKXrMtN2O6sPk3Dl2/84PCv5yezAfK32s8fZbj
GG2XxJu+cbIUE2624Rkpcavpjjt/qGAsNA0xT6J5aMH55PqPi+sa5oQknXo+ngXYKQ9DnRosJuMS
U9iwICyCDQSqnwlWS0Z8C8VU8HwEHTTcnGelmvUo4wPh0es251RxfXdUf77CjPdUH/EzPOTGd3Z1
PwkRdHdkqq9O+GLfwOVEiizEBuPIsXTBHD0AmGcPSsoKU00Kdx/gYZZIAUX3LcYIRxfwx2Xfj1+c
dMQonvYJoAK0d84HmUD/tzEoK9lqbqi9laIK6AwbluyhxCYNm7Fh/r8LlzEvBKBrIHdw3dTiTr06
8sSKj0F2YdHJ+DWyw3hGvWmslxsvZSLdbMdCSJCn6iDMumCfyxaJGzW6V23qlPKnmVYCfXB1W+zQ
2Zll7SFuwxwi9VRhHNpvva3BwqDXocijsq2Bkv++H1PgGr8jfLUsp6nSKXwY4hUus1wTcsJQe6t/
OI4oxcfpeSTpXruvm8+aWzT7INoofnltGs/PGj/nNKdyj1JkcR2PGUiMd9PuF8LmmtqhcA+LHDUE
EVRNospB3LQ38ywYwpiPkzNm6pSK6j+EUaoVCYIZn0i8Fb2fxSHLNaRzeTagXvXwNDujHRcXN7sC
TiNWFi5Y97picraLG52djZ0O0ic16WYK8R2Evg66Tj56pYr6LOHxCn+/1hcHsapfCx2ypiUM2Rcs
ywe/RjnKPyDGtk8s21AqPtqcKqfRbk/yvTt6p7jfpvtYiv0oWsK+qXUtMKlt0+6vpeemAxQrTs84
zKWaxrxGq9cSfIcrzu4OsdX59dIwJCcgHkpNyREAmYSSdgSXfkwhJTqqbV0C7ipZ7BL/e+VaLT/8
D9LHZHc+bc2NpOOQMUfOcvinBQ0RKz8ShZOW97IW/rKRJxsG1FjthAIWiOQ0nKUEZ7kDb/zxzLPm
Jb9vuhm41bcwVevOCDPQsS1R4rHnZgMnwxdkznNwJCpjwoY6EY8bCqjZwq3VVRVdctJTQsfrlEmq
2PnLhkkQrO2pFEm42jTx9lXxPyaQ2zNfB/Kky1lVb2aAbxgDNZ53OEUNGDfI6VCFjBv2DQ4AcUnf
+Jd/AuUBFsqr7UzsotyUsSmQJCD5NZyxOihXsf6ootUoZfaht8NjDUnkIJsu6mk15bVMTcMBtTC/
NDyHuzkSLZa8c9wIApjgT4WUDpUCdy8Cxmn8827DQvX+O8FqFD1kMVvgo581rSHSnu0+TZiUk14E
TJRE7LROv8h9F59JcGilk4m1jC6YyVDkfTCjNYGke/gkvWzr5NZUd3PDLX35e/hH8ql5PBCXt8jb
Q2QH4eqQ7rZtdwhI1pmz2BNuGwlnZxz5qbPwxNwbyy3F6+I9xb5U6o45/U9uR1m1h6PCyWKlBSau
KrbKDy278R71bwXgz5SLm12GNKtdAhHrMNjazi8qB+tNeV3MgX7NiKDFe7IyLPfoyVr0gsNThu0r
x1elelWWrI5okKN3Us3LBhOdOxCxIMqFfuN6a4qD5FLRNFiJeLiZj6P5Waxenpk66VqRsfBFq0q+
L9zkrxpZnRS09qJan6RQV3uBWvoZGBlk8E/WKPHkffTY3H+E0bFcwCO42M1eyq+MGirWr3AH57AZ
GrIQbRJze8AkJeXG7Q56kE+88lHitcIwn8JtkE+IxhWrhMT9ysDQi4fEVTuU6dhkxYLZhYOiW6qh
NHudRe6n1ZkPPyGDHhDZi/P9EPVesFY984wDU4PH8hVo0py/GxNCTMy4h7ChadrnkPFV1O4MYZdx
ZbmvAfa/7kWvdCmyCqBgttWde4umn7cKSRN2BMZUI16Jl+80Ry6vcv4dUcDQuXXk7eJ7Iupky1sN
vcdMymoArbn6AGk8QMX4M60BOINObtHh0rRY8GQadwqaAx0KjijtZJXaauqiev4ngNerqcR3jMXF
FOM2Qk6xyFp76APw5IB8MvH2QMU5OCYGnH+YbEAa/eOqOPfI+uuyKwJsV7U5ZF54KANdzak/x0QV
QCyfDdNmZh3XrzYOw8R8qnonADqKV9YYad0bJ7oMYcGuZJc9LByDYKykg0tqGn708SA0OlsQVILY
ArKUiBkxp/kxf6Vwmt2EM1T+j3iGzsE7wGSkJtE5+6XObrTgWEnwZ2dTfv4riDdi0vU8ry89D4mJ
9gs3+2PBOIGwaC8sQPRzRSCIaT0dUUdGyNFcGCks7Ug/mT+Cvmn7XYbJLUW4wbXlZXtZHGhVLvgP
Ft/L1rCmewicyeKMdRaBqu7G1sXxutZb/ReyeW/HOB01qi0+dmUoxrXh8e0FuuMlcwibAhvr5AJW
9KZzo9Uk3V/iCMHvFXDAS78ORmSL2pIVb7Zn5TlxfW+8MSxDKV7vJ5ynKNKY5iP69wxM1YkNQY/u
huxggj5m1gNMjVq0xgh7etKjkQxn2cqQYhXzn3n7adh2ORJtqej1BSKKq8Jci8J8cNoysFpd0n1T
jTS5uVBAqP5FZo9DkCODONaKp90HuTISd/pdB2Z9uO6HhJpSEqXHJ0JhoFBbnMHxfbNU33Pd/CiN
OGNMRA/TNTkdV15djhTgDe6Xj2HpbNZGQtOBbfc2Lhwr+MTd6ZD+RmT0PDdTcJA0PCpQPdJO+MYO
DH89pT7HaIn6uyjDT15haMoaY1MpH1mwjkJYlKjA/jOnuRQS16OEee0Z2aJSpO+gcpAoCiTYPo88
q7XaXvRzuObEStsv/09xCvUhaH1ELrk0W1WISqtRHy3Ba9Z+NadtPUZp4vIjcXrNxBe6PMYnMXU3
4ue3+gENdcp2vjpAf51VZE0FYUWwRxGt6i9+U/qBirX/gcrhgKus3ovQ2SnLzfLeJAT/SnKoFs1J
6o1VyhM7qB3PT7EHPryCiyDHAHUEV6mYC2rgWOH+W8BBbjnvqBWjR0TvmNW5x2/fnUJMHbHDItl1
C6KFMMulJ46ygGyOzCQl5Iebh+1XfTG8RK42e11Yb4S0nyae4ZCRBKgrqb6OikrS5GFTSz80l/zt
W/rh1OUn5qUBc3tpSg6qIw4+nls7mCY/4CDEL1avmVkrTefKRdHS4oGEgUVVcFiV2f5Q5R+Uqbvh
AL541XX93P0Mh2i8C12GlpsTYsyoU360IZQGdw0LtOQZA1EEZTenJvd2iqfXz6n80vzKmE49pRBR
KKxH+nHrRnha5D6DAHzp+5c6KGlqgYwlJK6N3jpV+7+txbDIlvBaWrcA/brgp73dS1iGjtrETeLb
pIJcknbakqWL58dYlTWQ6KPhjyBZA3o6VgXTX00gsjx7HzSzqlkqhlj1+s0dzgTDhvYQqMtnIYw4
3jJeKXC8+9A7BFSQ3teHyTPOCp0s0NeGWU7u0kjJKYjsKg88EovC7eDRUKGjCfQnFWCYBYtdeo1h
e8X6Vw7A0iQhSupt4Bln25dVS5WhkdwLxVN/h9c+hVCc/+IED4Sew7X2YzvKDv7JdYbhiZCnf764
RPFK4+Kw7xJeUlL6otkFwYGaODNc0w4uObni8gf33cUga/UpMBAfpcDzIdH56zqAsVR9y3LDmGvS
KVRZYXGxzOxhsyqTL5PDoctvwR7N14ikAQU5sSEsOg4T3CmghcMZdtG4BpBtaZ8uIkfbX3cWZ1xp
xKECROnrt0A4+Y9Hk1bcFFb0O7U0GixPjKTstI/RcliJB/Aow0Dy+Qa6yvR0zz4VrI+6RobV39EM
biijdkZNF4LCEH0s+VnH6dxlIP575NDjq5hyZjwxatTSka2euaYN7BcUmIUqAMRU4hedQfbnr5H0
jbkFXOVxFG6xlSQ6bkE2i+OTw2PgrbDowp7cczEnummDoF+6A9sq9J2aT34yq6llb6Fl6rNKqYWj
Om7x7fIIMeTZOYFyhGAUYf61J25aILS2vfPePxeq+HcbmrNkCU8rTsWIjWtsDDlQwSFzCnUXZbBo
kkemGFwFSltXrChJ8L1sJ5sI8r2QTRqUqQmLnsQb6pej+hHKGmoaGomeripkNGUeAU6V9h8KQWDR
8S1KcK2Pk5JvSfqdsx/kNPKfGFiDx9xdd3ZOFHw/6afueg/t7AieWg8c8U6b+Bgq9bqR3HtbczYD
bAVzwdF8fpbx1cuheSnnbLR8kG4zIP+GA/d9fqtKEpbhndwBjTxxGVO3zE7uKhG2YAOREvP+dhwe
NuhvOJiyBh9zxOu7qmebIqtx1rrCOcfKaBdERhKOPnzu4ApCBjO0zsipIuLZdXzUR2E30aMoqxO1
24FpRdixL5W3MbuP1ADcU8HgWo0pq6uacYDTSts/OP3rfiVqd+QMMKVgcagDS5sUXQNNu9czaFGs
SpqxxENuerA0pHPQqOhqJN/nMeuWiDHRr0/Ntwara/gFyAGoYlX3zhDE8pTB6YMc6NEGoYsa6k+p
lfPtN0vSikHBP8NHa9mvknPjbg9oYj/3Ga9lIuLd/pVB0YKWV299sReNuJTDX2HQxBlHkRq6vLhK
8l896GSpUONxDx5B3h7Km+zRYVtIOgmS8WsTASvo6lCk3JqWvKiExl6AV+R4rc+5AKUPrfRr/PpU
Sr32wI52mNY/bXEvJAWtjf86ftmExIhf1VliNvWfSXXnS1pwMjAfLmc6/hPt4yrwMBTnR9Qvkw9a
aNUIsVJgWZCBHYUQZRw//xQ8X2rvfEevcHQ2zTQ1sbNB5VnVgSw76pdk+IdfecKBstsBBfGZDCxS
P3hnIECNgXqZzLQWevGrgAEsGXZuho5aChfTQ16GSQnMO4tw5NE3uUoFQz6AU/00O8FpE/cO/wCY
Xm3IHXyD/GbB2xbsjj1OpdkTwkwH38qtOLGQNW3+zF6EtnfWc7CKwl3NInrYWm3cQn99aZRp4Mga
GTBzTsn28hXKlrtiX7AWP5YUVWctSrHTAtZvEGrQpPvLzi6r7g6baIG1OCT+ykG2oh0M8kv55nLn
5xgz415oiHPUvdkaDmUAeYopsquBbDlc57Obhx+lJn9k7b4Sh+uIawukUnf4iQqIadouI2XF+qoi
eXM6ky/3gzHrarIvippyadaypvDTCxNHXlQHd1S7juZAg4p0kr09wR9xNhegebR0/0Myu0njTyD7
T/AwZhKojjqJFokrEHRuQLs7TidbpFIf4XsuHWfBqNhzkOrwCA123g3b8MdOtExs0UlpoTmkHDAa
UlRF7CQPd1akIw+jjbxL3CsFLfmfgQxHZEsjwb6wHUkF05W0bmYUvvkyA26PCNhiTsAjKoNEaLNh
+58sczDs2eYaOQYiPBTzF7GVD3vcMe8zKqWROA/kj/YB+74NZGn/3d0fDEZDCWQCTyqVD9FJyFuL
lytHaohMiFeRNCL8uJph0UbwryoUN008lVYCydsJ5Z3hbNjafuGcPT42ra587gghD4gP19Zd9cBo
CUXfYZ6+gevFLCbDDrygR5TsY7FQDzON6v1sL7dw0Q+4pOdbOZB9Ib0k7ZZPbRyVOPWkx81BWGy5
qX74cDAh+/AfLajGXezYYEtKNovXAhdHTmeC8nt8MFplgLs1DT7z9OufmKmPlbx30b55ZnIDXJyh
eDNPJ/158GEeGgGzWtEwHqIIIO1HknawDbIGX+ymzkzG5Ambvr+l3CzYl//y8Fwgq8KeSK0fB/ST
c3o0lER21T559vA9/OOeCW4aTSEq1IRWKIltrQol3rOhYSetPwCjyq1oi8xdTajUiHLwz/pwC2hL
a+APQU37+tXyPU6ZQj8NcnYI0v/XFlPZN9cEJGIsgnBDtHMvfQVz7xolZb8B0kHIkh3BwxJjRk02
1IFFy7gV3xvWZj7mGpvY/hTeLvQCYAz2uNFo2ISSN2ZXC8xGtr0F1uVAOF+u818jtmEYwMURvb9I
kED8+HL9YZH79trQo/ADS6gdzUPN+GRFm1HKwksf/y71btXgBtXKY0C/V0AIE684CHfQ0mWfxYLR
IsGzkuUYceA5oc3pL+Rlsl4mDl+BkkSBtxduJ+yLAJx7ePcoKlz3lXka0++Tk0dLeTGT3yZfRlmB
GHouBvCuR9gOdcJ41dTBj+JPdDJ4274R28kgMCzSY7iBljjvmrQzHYTkpvgFHbR8qTIzUmCT6B+l
QCdjEO43gOZe0bMV1ZwwOzCFpfFh6SXtXW2J35v1A7hvtEkfxBPmwKTQ0U16N4cl531sTOIUhEzt
IpUmPTvq4VLFsCDL4p5nXOFVTnLcydnpYwB9ZNW2/6btGdgtuGeqL2zy4+VBcmjTVLNjLusiB2sj
8dhSA5+yIhQnCcewBrWXFAmVnUpi7xniRpQ6Z9grCnEB1+m18tYyLOMiC4QyyjuB5ooStKFT7JgX
7kGEiYTxq3FVY89e9Oc7XVsdtdP+iuBijcnmi3kkVsge5ADDV+ubJZ3U/EhIYYkG6x5cWwl/c6LX
yhamw/RMqe+Y5MqpAH2k45jPu3mvl4D9E4LyHAOayc7s5mJSneF6SpLqNO8TvKkiCRp+LUufN5RG
q+n490dskWDu4MyiQGQRok1tMpnul30S1xKL3EFz7Nd+NX9uzG+rl4kbDjiv5dHkIVSnmbhtme7w
dRvWG5h+EQoeTbjZa7L20ktt5Ox3YDT/jvnRTD18briXB6Ry7bMy8JsajrCbxmylL39c0P0Y8IsZ
m57pogh6sVBHHNGbUfecFfcDGPXqqPqtNuNAtOhe9xWyw4qh9Gx82fLQ64LIf9N1WIty39dv9QLk
Ed96nfzA0w7cX+6Pc5Ope1TaO65A4QwEfGY3P4gTrFqXq50uSB51Z++61MSEmN16UgT+icVRqmTT
x521c40Td8j1kee5ksGIXPzwoohmkZZIMZfWZUGJvkglvRgrJUGDzTbgAha/1mzbQOEBsKwNDlFt
s54WVvx03j0JlhAC+bies8ixVZfnaUQnjnRSeph6eD3i6A6/83K6+WT1zTAE0tUEBngAZCrpVXBU
ytiyT7gqTWjJyQISFCKnYUb+R6pbHfHTUfihZMXmuqCx4jonFdO1dOW3RRVP/+apfwJBUnhwu5uQ
dUVnXTxoCjQ3JpHZ2o37NiZMGttGgM5Kj45AaXS0OjPp0D9ngyeT3845CAcfBQ0XqrrIFiQO+nrG
IK/Z14MqA1VJa9b8T77s0/ZhV0QtWhLaCjIc1PBLCHzGUpNVPtevgLjnUzOr3RzC0/9xkdyoHwpg
3N8/nXdqeAv5h+nHjgq3cq9hUOF9Fsh2IeYMfDgPVXt/5DPl+8BaMBDWmygBq5XaKWWYb0UfbJDi
KaQqXaImm+h5o2JhraU1SdmqSpnw2pathMTNfypY0T3XyRKjokaZZyE1uyUACqDhH2eFLi7MS4Sy
SH7qSoH76QN1DFwc1HPKVv2XZR1slMaEHQSsDORUOjZ18QJaONWNpfAyd5/VNzjls3XMT9IUYO16
bEl8m5db7sY8lj0qAZgRMZQhLJ+7ovMYIDl5/8hkPxQeVceHB3eLTC4Yz9LueeqrJ1EUkRNLVmKv
obN+GGDw4HuS7//1KTxjvWEVLrUYEPS3MUbVquSyh/K2wqMstWiPl2gsfoOvEtGezBtx3LD5Fo+j
aYIDiPIPlT/6MT23QBlLt5+0w0sM3QfZNJSTZU8vcA84NfL2kYkjU2+cWVdHPDsvr8pNIZCQMbVd
v3Ok/bFZuWpolfyunqyi/yXXASKScDzxCAROECBFQZerpXgTNmyfWzMbA5v4Duq7EcrWRRkzABeo
OpjHkKq3U5YP/OQ2ec4vZEYX+gD2McnUv+wSvuqx+eda1VUlVkSnK6G5InjAz2N9VLnPFmhJiAUM
mKakKjw9QN97JMIjuG+JYUx623ezrwHIbEDraqgob8Pd1zFTtBgamkBq5BsxWT68xIvtWH7D3tvD
9U+mB2mOc/PchpN4MPJ8n5vn5IsUCO8AWtQfN/HKokPKMSQ/3CsBCK+id2gK+3Sd0Miagr3kKhK4
RfcS/0Cl8KXA1K4TLy9kLRDwzYtHoMIPSrn1H6ett8vXdpIUtZ8gA0WiKf0rAmnnc8suoiA5R5ex
2ewdQAYajKBLIgUwycUXDxcwSx75auOoWHGugfk5SNBtXrg2WTsg6v33CN1nJPSXdoqedGlXw1HY
8EvaVc8UFU9rjMUxPKaZ04fNVRgBcxbrFW7kjAlqS5mOLkb9Z4hAEHE+praP42wO5Ussvj7p/WwO
0eAfGzprAKRFaUegh1mcEGlLTwOL9TLGn08JHJxoxQT8a7yh1cZ+eGUedJwgycC7rsRlnwJWjOxl
4wDLN7Ckc83pAR3kwAhztnqzSosuIY1+MMC75jVcAHP0wzWVePO+dwIbNuiTepdV2iEL193KZAye
Gvhl4kH++pJMTEDFXLu9z0ANeElLXnMR5ZZfIboqfy9+gCk4w+6zpZsq5fb5u/3ck0Vfp2t17Z+s
VGCC2o4LwhQjY0m7xr1yRaGsevNXkN4cYHoXvB8BW1LACkgAHHWBjv/snwqBg9DXxnl9jiB3MgF9
OBVugSB71L4wkbDyQiiRmaT6ku15mheZ8Hb4BnMlU2F1mL3jX38KDSxJhPPr7FMk1Yn6O9Nv3opz
7AuwwPNf2keO+d8KdhAL25oybww2dufIfEHyn4r7yxNyOjhgPBUend4VBqXIfOpJPkcxy1vl96pL
uzBhY9nE7U2OynlMYuRYdRQiIv2OgQsdKL0xht84M6++uHzTUGeS+E0ZL7UshVURs0eLxwnXga18
MI0vHgYeh1A28V1+Qn/1xJTfAdTMrsTXAzRSxQJXwlp1XuX3ujlzTCEVsfpEjp9hFy7VRr00k+L9
zHH6l0f4V1TkiRio2T4kVYoXvS0Er/7Grh1TJOfKkkIOfwOb+yInpSCSa7JyeKBu0BXQvXkwjwCd
Qna3F6AgOiTMeBg8mt2GgrZGkG50iQ/kT7aRyKD946+JCIMHaq1u1Nb505lpifQ9DmYMdnTpzTmc
QtA3ZlrvKltz0ygRM5WlIyamRbCiIXBR3TK9akEal63MR7p0MgbNUFcVyqGiJmYRys7whSRZHjhZ
KGqlUwZxLBNiZX7vN3DcBK8EABORA+31hB1l5qJ6FW4tPjq5GQFMZhxFmkI79fBDwNp/GXiHK6xu
a+57xKO3Sp86G49AvKrQiJVA9AgvIBSKjMEuW/gIjJCQ+a2xoYmY0fo1Lrb2auvYy6lDH+6+KPpK
IVzryisMxFbyJ+TjrrlJRVx61Z8vmvsJta7/6jFs5Y+FSBLynxAFPJybUkp1TQMF3++UZmqS7VZr
XKsuwL/uRRJmx+9kl9uPH165VkfguCvkYtT/b0ZYwAb9xYwiy2tXTh+G7nUnmwHZL6OB4HLdNJAY
7/c+ao/I4v06fbZfyyI12zhlQTITIHR8rwqazL8ef86WXccrLOYTK40AvhlsrE4qVTvJ3iWeAjvY
csPosd5wrXRdpm0SDyRTtCB2TGTNjMJohGHQa3jz55HraLOWxVj7mfOw8TYciV5rk29iS2KOdZ0y
8dsaWR+APyDAcix4s+LfEydlV60j4C0fSe5f+OJQfEnhyq8vc0gxikrzD+RDQr3p4pm71oIpX6pq
yn8HQj+67GWzWDfzO5/Wew24axxyWYnny+hION/aqYuI97NZC3xBeK2V6c911EoekbltM9S1w+9P
Cpt8debOANakzqeZRXHJunWJ4u63RT2LqUHTAsnZecVERgQ3VKZ1CvwcZDFd38EHsEDAXcW4+fr2
uvDbnCZGE2N6PD2mbx+vCaxRDqR4lYgAHrSRfDmIZsjDI26WU1zqm37AdsGl6x6L+/jHD54PHvwh
xLtha7HuaT7wW8Vfd8KzBUhoWga/ZkLhmxxYYeWU5RhPX1Bx2KrzE8tAf+BAKjWZDQRLv/XTouyo
iFy0+BEK/Bu+hD/t4JX5MxvXCl1wTVvKRMU220cvOg8z1+80GsnPe6+cPXCoiXDkw0qCywQVNrbW
gd53R2H0w9b/F6wqQeiV7BZgi/ocLKWwux+E1wpl0tvVJClHfhC3QAnVsHFMXYiqlMDP/y15b9zB
9qLxYDAJtN+51h97WmJvh/idXYUpvthfbSdvfRaGP/YvixE7EUWW0kYdFvkZKkeHVcm1UQR1kJpu
Z5IsYCG1TZ3WEp9jGtLPSIYfAH9yCkfDBcALzUE/TagU3ngkLBkc2FjOgxDfpDqIsQ2m0e4QTJFe
gyJaiA0HY3Ld6gc5SjmjQsx9VrW/Xa5/RCU6LY0ru2BB+LE82JcWMaz99G3BqJGLMRL4pvMEQCX0
efjVoBIIVoCGhg3BL/sJX6PiYd/6n8ndRYuf2lM4ZOrZlTj4JRp2G3jaHUsnUBnizacOHjlwCPi/
250mpJTwQ62eB6nScb2NUDrkQ4k1ed3wfbJLf/Q97e0e8m7WtEFsobjU1FmpcqSxp9M4tLcSwg27
zKClkP5qx9h5HmSTK+wc5K8ON2GvMgbl1SNdeM2MC89jh/8Jqamc9AsbMDz3USzJmX6nc27/RLff
D8xp/ZaZv98ktIH/ymPiJn0FcZaNDJj54xQyePVfsZXRNqIM/V33w7d02TNkuDqbajvidGvBrcLb
zmkUaJ0wZAhsvxKxONEPwgH9Pa98p2jYZ4C5LEosZRMpMN8/nvPWNwDdYtdcr8Q5FbMn6I0q7ajF
oCZEt79ajPOxMT+5RByH9wkjeB0u7m7WGL0oiNLx+V9v1UuJyHprqeng9dO40pyv8JBObkHAPAE5
su3ZepIdcgS0WSoEXGfBK3fIqUOqXIXGDCgLk9C17+XahW3jA014fkZByu0KsTDqsrDAKsy1hjXL
8ngcgmeTBk9Hl/MJrqEwOoLBZd9pfUdHNRx+3rQxcVPL547KgpAV5LDA/85+Plx0B2d54+4qwcgH
n6tum8buCPWkV8z52h82/EEP/6yHOPUCWvWccJUQhtZZzjQjfjbtF2T4qn71CN7xIC33TaW8Y2XK
OBQMNIehKR7YrHyxeIvGn43Y2C43MBsR6F7EbFs7ISpmRZ1EJvK2fRv0h6WaVXUbs5wrcT/zLuaY
7hsWNl8a1e2LuSbnsqkx054DGbDQvT8+6dO2bgZ7l83aD61H43noA72ECTcGSUzDlszR9jdp1KEA
kHKqxWxr9CaXTaj/5jix7Qjy9/kg0ahWAR5TB4j5yx2OAKamhDjwoTBlt6/dZDa5iYIGZAtL8iKI
jAmJXOQg+re+SMdmZoa/SzxJOJAH4sXpVIBkAIKWG6qcdWnm1DDF3KNQ9PaUUlKHXfjsvoL9KE58
rXztJgZCn3OtiJoxsohZ8sBHkTaSEuGiN0OKdqlh0XwAd8T+GzKRCaAfOWX5epe+sTcc03sj2uU0
0DUO3o9w6FWnbU/YipjBnjJvp07dygUXaQPTXMq09PQzx6K8c7qCekvupCpllHa4N3jNTsT2kEYn
mOAGc4mqaKi1CtN5yF1PfCvI8DC4Vx8HhDSpxiLHua73w5d/72uhiiE2cAMjBKa+yh4S6ERe/Y10
5jplZht+TT4+u2KXHeWCrfsrMqNhevlJEv2vZh8ZK5lVluVflM4xAgPPhYfIx5U8yaQeCDFqq/26
yr+A/3OxlQj0mmB0PR+tftaAPeReHv2ATsdKLbzHaxgQu8/bPy7ZKMuBflr+JFrQbq0KNxYn3Zkc
r4lX2a5/oHIlVL9lqnU6DJXTAjDSmP5RdfPR/87ApYkqcNMMX81K21y2ve4ZhpN1gN+nwhWDyyyp
ywYlHVBXV9qOIcdreBD23s9zMguSBnG8Aiz0KVyi2xqxEJbHO2xF4BYYHgKrWTCu8uJrpjczff+p
N6nE4yjj2mKzX4YwDBbE+0ou0+8HiIr+Yc15kGItC72QuYt0WBud33KS/fabAY5vwz2+jJj3o+UU
o/vqEc9JGA+bMQLa80M5OKDE/yA1JI9sGSmWsIySb0m9aX5MLQYsOxxuO3ht1GIeNFTl91ayJ7wL
uksKadLsbldZxHYnTelL2HguCjJR/4WHF3J6YMfBzrtS1suDPGw6xqFH1YFBN3ocKDQ894Ilcs6v
VVuWrEs83OYLbL2CyNk6BxvlGiTsIhHIJxn/prqRXr021h8W7whTqhERDhvYlMpWWNhRXXnzWX5z
BDbumuYRbFDSMsgawDVxtLlJwvzQA8Reu56pVslXoAEDweP7WAOrKZutJyabq2MRj9G+TX3gDbN0
T3Pgrc5KzBXGcEfWxnIGv3ViSOvYHlS+bE7Abmz5Yg5RPkbltV39Em8UJt4tPIr6e8YoEKda21Vc
5gzKCXjQV6GOlRIuqMroVetPcLKRW1m+g65kYBdxDn+kBWNx/uJ/JWQ3Yw3XTvJXL8Dq6Pgj5K3q
zw/0R5yFerMWKKhwbl+psA/w4CZMG+rDWLYsA3PFP2rPxqFwBvcPI+LaPCMsFf7YscUyJN9eWhv7
93+1dq8GHfwwrLoqsmlIacBpW4eLrsj2ZSskzZpKQ8dqMJq7SWboRUDrRlBZRXmLWcKRpqLM3Bgs
3XOeuz3dUacFakDZR33wMMfx8JgaEt8/+o6hUwt4a0mOmNAxAK3q9NCspN6rtWtZL4+RFjx1IxvK
ofxvk3C4TLd8oglk2rpucBiqwzLCvWl720gn4436L7aUFBVmRvquyeq5WXLV7g6K6SgE5iVqMDr4
NbCm5Es8gZGGfUcZ79F7GZ5vz1SJmlGIsURIL/O4w/OzbFEqqFZBElh51igbH7dtSKJFq7j0QXSi
VBCY/9EOHFvvhUP+Rf1jii/jm1U/CkVtoHK0yPHwa8jQX+7wLe+1lUkbkWWosLZAnUSVpBkmfkpw
+BBvklDHD/h9EqmmqbBl6BY6fmwqz0XgCGjWTe6cg6BcdZQm65304LC2rAJzf0T47DkXplGhCEDp
HVlpXhLW0TIfpL9IbyucSClq1ZaUKu6sAIOOaAN/5KPjo08HtHdx8Yh3P9UGiXvjbzT0H1c5JNhG
QmiWRsDsATtKizQDD37dWg/mx8660ZiQBC5XKLJF7jjRQVD5cRg06g/spWBgqtIVGJPZnakVKpy8
fh9atmg+AB2a9HBy7BkC3scZJWk0rTyaWcENDrhCqP+z8bY9U7n/IrmjXj453u/2YkE1rzaS6YWW
hLp6XRyAKMRz5HuY7jaKq/Z0CD6ZXQOUi5o0DYiWreN1KWWue5RQw6k2ZfSDNHwU76UQ7HqYfo8v
p0gEjz+aYaYQS4GbRhgEFEv4/4Vt/Q2lqfRrkhKQhsYA6PuIaD3arEVADh/s58Mi13MjSw5u7OFw
XEEhIIHE6hR+NkH5z8swrSIgVMY3mJLqJUzP052HLy/tuMLU3926eSL3kxTzevQtJXtaBPU/zKCX
CiwZ0A5JbpyBvcwj4GZDQW9eJGoHqkdOxj4A2Y34Gut0cjrfRp5noDK4trlLjX9oTrOxoN4Low4V
zjbCkpfBi9UwTEPxiScRiHRo1vaBAEPowKrI4FzGA7d2UZy00MW5UyQ7K78GyKPfJbKi+TuTntck
xskNzmYRAdiwdJVabePc3c9DCti8wXZiK2AkILYPOKdNKhPuqlRsWvswCd0dy9wlLbK2FaHo+VrC
sn1aIiC3kGR8FE3eaI5JQkK7NglvbzbCW7uTtbK+ENJhwRcciYmi35NzeLR8IbTWAHDDzMXJ7S//
KSI8MaAok1Rb83GVeysoqGQ5vp5etNvBwQy9wJ1bm6FdtMpBliNyuiC8WyIt4p82oATlOKIrb0S7
7QZVwh5RCoMpBARmivyjiiOm4fOZGOqt2BQ/XCpWE1VQB9Iu4HfUu/mheE8bV4rgDj9X4Xx8U+If
6XUk3WG/x4mUnpfEhgIr5Yl2P0H8J12g5Zzd87/zK9p/dT9uwf54UTwP0Xu0Ezte6BbqDCLUqDpi
3zN6gV8+XB7kv2LrGjSBBXsJzRyo5pqeCI402czrRW73qtLIdLEYpZeHMlT2EUwRgtVy6Qj8CBP4
q6qsr0IWq1VHfLPWdvoFRbrwr3PlU/hdhsxeRHqglYF7TWcpSZlWWDSrOQW6wTC5u3nQR3hm9NNw
bE55x0mRnsvnUscviehaFwUKw6GWtpgZnMm9lwiVS0qtrYpTVgBYkarwmXeTuH2oBVy5MjNq4ZWK
ZcaBQ9tF2Y77iJyZClmWK5j9ct+mJMbSX82jHoh0z8t8AdftaEUzDKyHet7L0dqs8WHr964iGWn2
pNvg+MxQzQ50MmXxA4wREwCnDOHJVZkALH95/FeVy+XM+G5ETsCSYiOQwodZMgLiePnUupCsACNf
iEsw64l8gPBFrvX9rWOaPP+nUtJ+0Efdkd+uGOXGMz11/96JIj/Fb0RMlCQTui+X7bPH9lkWR70x
wHfCpRnnrqXFU5LDobaKm04lxbmaQw249IzVbJ6VPbMnCQGPsZlzNRH3wSameayoA7tDoY06I5C7
M5RcQThP3UMjRnnApPdPEIp4mKzQF7MzMQ5dxCXDwnXMU7boqAIeWkI4A205uWpadvMeLqFeJad/
pUkozdJp2jRVaeyFG0P2XECfChk00wM5f46kWBmwOfU7snfduq6YoDR2ats2PvCd1l40jLGqQQ5p
S1QrYuZ0gcZ2xLY8aSYXJqauM0BrSs5r68r0NVHNL1ZtdfPIpr+rn4wKylRd+kvyI7LUI1LjzZGt
JO0ahbI5VDQZfXIvVw96751HgQvmQ7JijFE1SSntsRMhF7IdcnKKvpSCG8p1b4DlCJlbEYsnQ1xR
ottixRQC8ylEfszsDl4iPmTimdIsuMP6BNXM9p9KlSaXtoillwL8O0aj0HDDrqCkUKHEkVx0fBQC
xTFtdbUAntoFtr8dBvp+1GOS5TSuT43xX9Qybf1ILere2l2UD/i5p53i+nQjC5nyOrT80FZ3jkc/
3xAH4rY/ySSjsbhbVeFKcUHuNv538gCEDxAQF4ol2t9UeTcr10y8uRrMIjXTSC7UGbqRr+ThbgEL
IFbJam8tQwOSvYSodnetVQGYYhaKLNfDHZlsc3QCb9JAl40Ajg5+cYoW4efu6fSAoUbzWl/bQMEo
Q208gIovRQsR8xYIj7iuIB8n1C1JKqyPfeQtGf7NEj95F0xzUysEpfcyz/C9IM8vrbY8QISfhgE7
g+kOzFA7C/dx9OcjhFfU/qQl8ns82VSUK1Nc9q85UvRQ4EW32X/MO13ligEfhHNSh/FT/lebqgfr
Oxn5Zun/kWhUyjq0cimsDp6h7f/wj6Ox5GAP5n1qGz/AtqHxSqpK7NFcPfl8O/ZmrdSfXPM/jyhk
6hURYRySusDyGvN9xbcDGcuerm53yHlg7KDmSpvmYWYt6BnPy1RzbB/1ZjMeziA8+sQQqz10bgcu
c3jZTHbskaRW1OYzFK0ic4W0il/bpxG1Tvu+qJUfAl7YGlISFQdWmfL2X6TsTa3xfNKwbvFhTQNB
/HHd3CrXhDYwwdTFXbSsaXnq0RFf947SmFg7KZlkC1hvGJX337uLjZnhm8WlurcDPpGfqCMx+YU9
V80LUxHD9Xq1WggCQOwa9H4x4s2JLBUm9Gc8+Fp2JhMKmlAPe+DhLXQH8H4ZNPOmJLAHR0jsgwZ7
fiqR9Xgin7s/dRYTmi5r/hvkV23+wo8pyuSeyhZvkLRS7GqAczjeb91rSPRY6okRVMtnutyXyZ5o
+iVnD+fAvEKBOY91UFPxjxu1Qt6quREQ8JXnyiXYee8T8HoyGTJV7jT5tiSfO6Jf5Nd1z4xeOO5q
2I0tIibchkin2Y8Z2aldWUl+8VDp6RwErwepPaRIe/GUTWI3DUfvHSqYNNZImknaiPy9ulhM0O+Q
paj1KeClBx11KC5o92XnAOc0g4E/nt9vIjCAAGHf7D6K4eVWabCE58aWfCo0RjxH/1FPm9zm0vJH
0u9bpW0Kb9Bh6rccQByGd+Ndpb04w6DUdeUz6yllvdIw18aiJXqKpLaUuKQS1l+k8X/JedW9kSVq
u6EOFCEKvO6oJz98MN0dmxVmY/94pE82TPW9/UGFwKsh45hkFDDN4DJQO3sBdP0Afg1gIVFIO1Kf
2eWVwbO/A+kUSlYi7/Qiu08JsdA4XFXXbUmnDCoQUfVxA+sc68jz91A1PN+v4lP9WVKMngMKcwKl
9FnIp49vz37pqXWqPfYBOAfX+FrpUULy/CXcrcdxzIJCYimdwEfPngtDEx2xdrms2cYX2HnUayXV
fcrJyU5bPLtWGHf2mFAbzxd7LpeMzb184PUnWNiGeSzor3tC76UwlKc+EZRI/dHeqEXQC8icBAyT
6mhQ3T/Lt99agHgKpZwilXzWqGXl2vBkI6caE+EylEu7pSObwTmcJa/KoVPNW2DmrU8TgYY1m3js
pbSh6XXYtJl/wDih8v3M2bBwd3S8sg4Tl/O8NSjoSzs9lKYmgv7EzbFR4xgKm7e22jraem48j/th
p+3aQVe7fAZ+HuDseDY5/RYY6A2VwXulq0qy6EFnjvOpsyR7XpgvFPzI2aCG7bLuElN+QtNfVXng
WIavUy+Bqnfhjevpue48ABA/82mNaWghKenRyElPzvUgA7HIvU+4YGF9BaKiaocbOZ1FMGjpqNce
5poB8z5djnKdKd2pqjZY1MUWobD2lsC+zNAmjZmgHOo6dWaa1iGqBps3Qa8CGqiESNDc8gza402w
ubOwXbj19otSC4pKEs6GkiJieYOV8UfAuFFFLRZXw7AGqN1aneBXO3zZBl2cqTTm0WMvVH1g8Vb8
JFFRc3ufqfMBG5GeXNf8Ob7FrwjB2Z7SlnyDuY8F4uO49oqBqftk2FfQdFjYkkpuFmXT1ulB1VSm
CZnhata8NKXs1d5q6fXF2LVMuegJN+wO/6eaSWC++V2oup3xrEwbKbg9/v6Dr+52pH8wt2nTNjo8
5HyNlRrFtqFIZOlhdHKhHyYqo9PKGybeOaMnN0zeV9ojGT0PttEQQwICPrjgK5EApvjNggCPSdBA
f0Hga1NBwJFlN+69rGeRnmpDzLapzRgrIst+kyplZOcj2Ask/R3PspbxmJcojEo9HLkTqcwgRAMe
9Q6A+vR952s1lcYwiF3bUau1zwrfXbU9D9Xiq8bGD5WMA3GL/V2Vtge7wjOtirxvjrPi+IRY3Ebx
Cz8bl7gT6yFxdcAxP5xL43amlb/Idf9W3WqeqMnp5nNu4c00SctTMlNaNdK0SlLuKLPTkqSjDUPN
uFzjYIFYOBWuBu7EbwWBlm/xZjodcOd2i82H422nSeXxNJic9RdTKRoRwvCmjho5Qg6oDLQcwHE8
Eb9hJ1gY/N0PiDR7KqHKzRxbPcRB0v7sWqxAQEuFK2m3psIwo5Qj4EW2Eq+wcID0DOv82U/0G0Js
/vKQaLgERvr8ind69RvtUSxkYGjhMQOBVl+taNouRsx+CLw+dK+MYsdATwIE3PqWehW9DFvaXlez
vrOwDmAI6XCU8myJ+JciXBM9L5dWaogL8iWr4ZrU24dEINHB1VbWZckerKN0HkIZXspKVprgf14b
k0eXXuO0gIiwFU3McBFD+BfmubeIxEYjfrE0DOTM+KhavjPASvrFNBeVQ+daHpGYDVy1QF1IRO3H
bPgPsL0Lm+bmZYHt7bbUNL15esQFudbWWxRyWw8ABl8Xs1HmCU/N28WFPQycz+LyPFwE7U9bRR1n
0M96aVpHOP2NJ5E5Peqphj9GRjGcubZxDf1AGlIYbBn7aFpIGt72GaZsijJxmkMdhaGJKAOyYR1o
vXwUUinU0lGxt7QAOl+azIEnV5R+MHNPVd/QKwj7WlikStCg1bYWiDsAsNfkXirhPE+248/uiRQ0
n7gODc4acNOoQESuYArP1tND689UZkiPjIlCO9drNw9hHUqr5gF/JHEIzaMTzf9xU6hLDJPqb2GM
KhTUzBgZbNCGTuTR6vduDNPEZgt6uEIk1lqmudeACYDcNv4CHh5ODFEyZrV23uQQbP5uKRMRCCyK
ytzdSvGzhSetni/uTDNurBwRsjzKotcK6XfMwaH+7yIkkQxLC8s8lfz/CnUAOs2oJZEAmZhkPdhZ
g91kufge7yeZulSpfIwKHlhpkgCHY3mLkwM2xUH1kfYcvBrx5QJRRyvMD3zax+bZTmJeqv0BOlti
+rTn7jPa9wujpvXf6dkxZUmj+nhzgtym7Rr346vJ3GAmROVOyqS+kcYhNjDDY8iWojogVqnA6drB
uu6tpWIa+KPfEEqfGyzRSZ2t1yf+fxXi2WtDSU5vyFUAAYSxnx1urynZQZhD9khRUnU0l5pgj4zZ
1tmfsCkGz9TMClyELH+QXgyMPg5zoIDK8KXkxiqmUCfOEprEHp+Ws2hrWEAAr4r4b/f9RRrHnMCH
fcDYefDgMZjB7zAGlH2S7OTgb62xy3obWaN0b6kKEbZrrI0eyqZEoVOXRehRyxo+ACUUwrhccRpi
geE1W5xqpx+KHTmtrHELPWjPao5IvQCdiGSG1/W9YfuX998kFF/mOjJVKozJxawFNDMz13f1rHX+
UIoKMa2H0qzDfC0Yb5BAEfSum5BDDbWQ0qisU5hW3XdzOOtejuJSypdMAFDabZ391LX+CSBJ2OTd
keq1Br6qIdT5kFMreSRmcB6A9qxc8iGWn1Zjj82cKC81+ao0Rjnkke3rdkJTF3z0bTiMHbnfgNrV
UXhklbSjkkf2ndUbMXqqMvkqQM/zZk9nmLk8Vroqfgxe7isOMM85c9j8yovynO9WYRe0WvHNu31G
q1Slv3qz2umPPEKttr12l24g1Q7V3JLWAfzWIZMky4yBnR2HjGqFxbTBBY8r1cfWeCTlncHfJrcT
VBS11bnfwvXopq3SSSmKw6mhFkY5IFIIHnvhQqj8YOn21p9BcYzfq79s2/qELkE+WtHcSiKr4trv
Fxnb2LHve/y/FGEnP0oonF3tQWOvw4juck2wvtr/A5+lTlnIUFC9CFdvHaMyRnCXDiGQZTOubdaJ
tQaZNYGSv1vfrDQe5+MQ1KGtVOl8Wpz/9fRMEOGw68BmmpqK1W2jYP+7/RHftsFY3aMJu5rCXrd0
6B+MZ4Rjj2/Q32YDm3ZxQgBngLuGXR/UfVanIEht7N7M2bjssGv9u7jDHzXBCmnrpkcRad2biWNy
qrJLHM17V7eCGNoRymAQu0WCUeZ68xWH1Qj2hVRyueUKgHb5F4ESHXBqfUfXd9IXiTG5qcgxFZXr
elcAqMWJc+mYlPTyemJ760Rb6v4pLDo5gaD1xQCWuvL//DdkD7abOKtbDznkZNq95UO1x3jznZJv
eP6w8RgYew114UiXvzmIK0iUIKlsPNwI7GXQ0vJ/GFyEEP4fjXOnwfLWSteUrYZoLbfDXkOowtQM
p9oodvQIBccVtERY6b1H3obSUbTZfpnafaooEQOnRrjPdslkXKmBmAHUESqSbEsjWIuZlBj/GYkp
IwknZxMhapa4RmCKpb150hTJfbABsTGg1kesMbIAqwkffoMU9Y5LnJDg6kOfduxMHrsYCetkWzRQ
GRvI5JHO9gwHIo2/zNmRA4vFSGiH0pDz8UtfeXviwbtkzRtLw5DWIZxgSVPXFOWsvowFNbMGt3rI
2edQcU31XcByFctKeaqC3ALcFVseU7GtJ9jY8uXl1+fCB4I/9XJtF+uHw19+HdfK0hzUNxnr1PoW
WMy91FVTZ8sUBxy9iUDS0ra3dvxkP4E5GY2rxsjbGPx40WQUBtdwU0xhpyXp/SOPkirtMTny1+ty
0qpGMCnFGHGN/xPikhSeicr8s+sx7P4d3oHD9Z360e5XxD33oPhdG67VrvyHc87a7OgJAArbM8Ug
7jVcGmxfRCRfltXaOZcWIEoylQotZp3csKq6O7eub+oXRX/rom/NKZZVTDEezAiGka/skfCdPVq8
H20pToekGmhQfsIjYXNsA9DaNKm90Nm1BlbUEb04bu3T9djW/X5GPiG74QxKsUXe8MDJlwnA49Ut
4Ys1CNRzfHkS2/RQffFFbFbg7RFE+qF5fL/4Pot7iEJjErDtwwPZUxwXiukULoMnuMps29g0chlC
7VLjgVHuorg7FIzOmBUTIhlajkKdKlz5aMcELPeQ0WDzxXw/GIXhD8koBJzuGVivo8Ms4LroXc0q
xwaJ2bYu3UA3HgK3pHl9AWpyMUXS71EyFqIn9WwX4kciwGfMF6mmRvvRASdv6Ddylv8ew35jUEVM
NRrXcxbmI97IVRz4EGQdaIqnTmFz+M5bXxG/U8y+7qGVlpfrA2wGCz5ok2R4kEnhjMcCEQi/ZGZj
YQnHVCFqisnvQ7NCZvKkEXSrmWJ3rle6JQ/JgjLFBESZNbEf2+SXX5AAGPSp6b8I0+xF1uNQCqtE
6ooAiEXjA011lqisXUW+p/Sp7i0+QsGPRDVVFLTbVk+czWzZoD7TLEnDPfBsYO3CsdMrwmP0MKIg
dzvEWdmCAxyY7hig+fKWji8KpV/5pLCgltnPkfgNoA23nnMwjRYQV5TWghFO5m6A5nCtkEvLWjZ9
T0VYFDvziAVILU77WmyKETvwaEzmE4RN0rRj2UJfuyNRM4GYiTVApVay8uFNyies+HRRhes2uTZK
hYqMHpUnDbhAVCcI9E6vhiKzdUNRfQNJIAcFUc5HFBEC1A52pPHqJGAMAhGd98fimaJhCymaCQCz
8PZgXK/NmrE7CaAO6tvONKZONjFeFQiVJ0tSsFamMLzKTlLHIrcCBobbOpm/tpIVNvHlCzh0HVJ6
bPIcclsgFQc3ClmRtG2Yxm/Tk+fmyL2uZqGHl/jIt4WNVmWjDRnMJ6Pt+IDfDuFiaFMkSX1UUKO3
v6a8WPN+AHteJDhhMr331MrmEDH+dnykxp/vjGZZz7plfSxb8LFGISL/33ToR7GxUkED+NZbA7ZK
iRg2QK9L1ibbbYJutov+ERYLBMZLLNyBykWSEPZiq3sVHiSEBSB6Q0ri7iRSmlrxcxqrdQqw9jGT
gIjoVT4NTgs5EHpIYwT9wnptiwLQBMyyng95xJuTYojQZyF/AIOHvXO/thgmGFMM2gLgS7aYFInK
60j1G6eMSEzpGokemaFOs5oy0Tq7SKiQlPm7v1H0v74D1Zas5CVh1fs/RN4BgaxOPyyF8aHoqEd0
njjigEjE6UlQI7i0GcXnu+DI/INreTGdZ87FqdHgDXNU/4Z7kLx3LWt2wVZnhLBy8CnRbmNJcGvS
LTNO/YeH5J47eEN04Gof53XNYKc27X3nnhfzqFg0dljfsYwY89k4FdB1+nRgLqayM136fbqpI6HD
32ZH2NlSE+qDF7EwqVjoSPXxxa4Hdd059IRAlJRfYx4+0d25XuCjRvjWq6ftZbCH9LCFZPM2YmgW
Qq+cxojjLUvlGCO+ck7aZ7RWqNmvFXUStUROejflkVvIj/XiTz8+68RHFMSj8b6RMyiAyzGccrxx
g5BvfJR67gV/EuUjCF45N3VM8l6JywLN1Y2sk6cjObsmLA482OW3JaR5DXViq8kUf6Nwa5wAvgV4
1QFDyL0o2rCIItfiIlA55Gt4TScPoxs0aflf6aZgLlBYgk2GNOraKTJg4FLKsafWYrcJ0LVmvukM
DGauW5RU+CNBMvDSuVj6lBFypn4DAMkLI5IYZ4jn7Tt5EL55XM24sh2137tZ/Uko6xIcE9irmeiO
R8Kz0BwWW5rxQnsoN0qGc02ZDi8uBLSsjoCUYRMng3+/vaKbovpzWRR6KxwFLUCDFGVEGnvMw29y
lP5Rz0X4vbhkzJ1Yn4hmDPLHyThMDreSVpSElDwoo4TaxSCm4pyV2LkA6/7itIOxgykjjAEvLS8n
w6u8jnCrUhDFdlYzOYGfKkpo/zsB91qmNGGKORYPpx4wEvYqnm3XRahkbJliT9ga2GltTeMYjjqc
B1p0l0UbxRKwT/Ji4zuAuMz1YcL0TpQKaMxWAJVSPw15x6xjFbhg097Wq9gvqyhRzIiCSRxD++sY
MRpmIayDNhiCo8X41z+MDnusD9ytYn//rglUSmGqh9RUeZQarWPO3edn6tS00HPRaAsQavcvcdId
CSDaEPJyq9nR31LYTGxVzs+LBoMhjbXAx2qv7iMAGDjmecGTa2lOitL8FWOfx5SDgY/DVMhkAzV+
AN0uNvStH/i19hoY/k2wcdjHea21oeY1evp2AClZ9F2XB1PVGcOVdKTuE+JBha6J9ruyanTxVmtw
u7jSi/D2HoANQfRbYbDxyAFp1F6IHbEj8y/GtJaKUpjcxN+TXsRTNvRDm9rRet1EnxegHMQaeSvx
MzCkDqz9v6aVKjmEsSDEHduwjh11ZdwDSyRJBy4US6JwTOJmUxPoXmTIsyF3wPtTzlBm5nkybtwt
112k48SrXwAEBNLW4BuWAwGKcSDDAqG9QRcv4ExgjV1im8C9BhH/df7kGbzr2uyIIn8zRvyJMX4n
jP3x8mOCmXYTMoCtWcCVp8f0PYmyUaTqkZusIhIRovqilw9CJvw5gHaVcUhfDA0IqlPw5jFgVRfa
XC/AdRrm1QzuDwuBAHHo8AX5npxSZ/rKkiR+XhWXsfS9nfkVTPet65uyKSr3SvIEq8fLiA7Lgclv
YqoN+2G31qzNPX9VDZuSRLP3r9INcdTByYI3qxRvT2TBMXxcEB+uKRB43XhPOJXtM2RTVXKBkMbe
dVnszvtYDdTWIxxew0jyjTZ4pQggByHypRaMc2xyr3ZLUlBRWTqmt6lt6jzaK/hMY9sxfRjebqXe
xYPQmEsnfoZS2M7rPJZauhGVDag3Jzvepmt/5nv2EzVmf88K9rzGsLdyJ0I9y5CEPpDbU35MtnfL
NFJNBXV9jsU0CWa+wF2eH6RIx6zLYnnfAS2Rybl19wJesGxRY0xByaWV9UPA0MCz8Sz+28Oydp/F
qWN5FLMVvIoW1Ul1wkzObgTUOKh3GE7dqWHjzQxrGNUH8l1MHk3rYyXOwITEgpzpCKwC0XXhpZ5j
gAhtWP2mvjT6HWtFWu0CERC7Ff7bwzLnLWE8sO2+k0CDJWR42DX28ke/DQzKoFYEsUzFsOXEZCan
I91Ve6/RokgTHi8GNnfB6QVe3AqTeXoOueCUPQ8l4jjkUdMHeFIsk6zymQNgZ7bMED8iIu8Ne7cK
QVq9KIfwwX7KRbgwwk5PoChryZHjeZyw0SZtD+ihP6XyTtdZrLFpdJztrvzEltKfWQfM38HhGpzK
ZZ/cyIc8P/mtsE/G7lM+GRCEc7QEghQakOkn09QK/xZxYYDsQAuzOSHGir8ZcLxRJLLmwoLsnoyQ
V+yKhx7fC0kwXdRQXfz1E/VSCidGAU8rAkrP255dm1IdNDMwVPRt46xKHwbMu5s2/pV+A4MlRwYN
RVMNnMVyugzLmC53kTAgqJCOYwOCHrighb+rJfPENEOi9miVVulnQdKGpWE4R+N+k3/b+MGfOVIy
JnW4vH46TY7G/ZLZv8ha46j48Bs3QtUPohtsOuAib0rLyrOYIsa8+I0paexb/SNTYSPGMBa0iH6A
yVeXInH3LICsjWC113Z5cKWPQ9tQhBRszXnDgjwnUibinFCk/aIoOwFhEST4imaKHNkgmTobUYdD
Huk5ySPX8iW3KgyAx1r+b3e/WLbTGAOWmquq9B3UIRYElrPHrf0nXf/K0OeJ5HhS5s/ASEiI7OFN
uYmNN+63z0ibQPgfkzd2A++J/cis9N0jPvrqZKKGp6k0l8PLYt/GILI2b+fGounB7WkEGQLSTQB+
ihmzs78QHBGCCun+vQdOqZfkNbK0Nqv7xAgRxdXCn0EP3ptAQzZ9IhsdqqUBz20we2Jdsnj3hyXi
reUpuLzF4Fnee7txdPDxrq/xvLBOC5miMaEgeNFUests5jyNkgoOorY5sEOIVtdtlsV3qCqXZ/93
FO7cbJ7fxmGUDJED/z/hv6EXx6qDfBFBCM8yq3vgfpuiiHWoYDRn2JE7dvI5O/Vq65PuxIDgMDpf
dHw55mzGY5+3AAwXZ/NFba8gqoakTp/SK/i5dSi//LfiB96XowJ8qbeCA9MxUE2acWc+oC/Ajuc9
sOllP5Ux78Lhf6Sv/YGyNG24Nt6OwQyJFENWJ4qH96k9+lnaEDjKN789aLOl0bsNceAoYxKc7kbk
51iYoMAtuqK98KDwcLfB7uqzDvlk8Nji9eHEDKAXzZwAjbS+H5BfW5OoKn7fbzu4pQuL8N1dVPFN
cnaeLrd0i1Y71tRpKSNNnvH44EGDAF896uib2uXIReyRCOyWYdIVCz9WPVEkuyxyUGhd6lpl7AbG
Gc+ssCBw7Hd7jVcwG7kPp4w7lAR9sAw7xkjBgOhm2ThO9vx8u9J1CJmG/BC5F/36Ajyrw9PPOebL
ORphbhi2zlFB+oe9TcIGzmb0kBsBtn3iLEZy5avAsL6DSzFryGX76ZT7qYL9uyqa+09lYrHyTJ7P
BkMG66A0MbeBEdHxWU9CJO7mHPUtcDc4Q9W10pzLLueeoYjLhLZV0L+U4ifNRsMzp2sa8dyvU8X8
rXPNK4OkmRE/zkEJf3T+pDsiqwqWozim5zfINTWJX+IktoSg6+OiVYQbeTZW8baMD4cOqzdICrUg
535+cipfoOynFqBjPWOb1214yeIh75RhqOu7fM6IzkfVysn9F+yLNOnj3ybUVL1gTo5wFMn9uVya
ekughNAYOoJveXQZLWOarT57dFYT5LYwy+3+pqOMo10GPAZaXG7d/PWnZwwN5fnX7DvM+9Zl1N2D
dvoKlppVPdp9oY4uJVP+dnh48VHxiDAYkjK/K4IwUQGHV37iENGspacTI1ZVDKk6VNWjNcz2uUqk
4h6QhhlWsQvrqgPgxbxUyMrYYpJ0oFVdZbwpZ1RdtcYC0lYiaUaCgnv8cZmjOIq3s/W13y2lZUj9
50itu8xpvz/CI56o8ZsZjZkAufCZZimArxMYhd+jaNfrkxMLorCY/nLKiUeRK7qX8QLmWDSCMZy4
EwvcMOlNhepocDdKb8+v4SzmyU7EPnpRsiG+Y6mG1GGvHJEnQrdrevKqZ7ecHY+IQ6h4Q7xmY2hY
qL35s02qcfbgdshF+pLt6F+FbGMVP5USAXarHe+C3bW/eaBwC8T1NRYzNtv99rWhafheaUwNMQCm
TRsfH4zeySaPzFXIVGXTkMpTpOS7D/Mo4VTbWnFqJu6srWD7cLai1BUb5q7sxosPxGrNcVHShg7j
nMi2Lk2p26BRE6T/64uWX1lwLJM5HGAWX3lZScdaXPdK/unpUZmRGw9zQpsDftplOoa0Qcr99Fop
2bb4oT3EabgbRLW73FMQL1uzLdDyqLbsH15u9ZgBDUX6P+kbpD6ZsVu7OJWf4NucV6t9LMRSo3mV
JlPHmw4biungXZHLG+/q0x5IVBBU+EOGC4M/rOH7sRMiNYu0n8uy9gF7YYedxiiyysPZ2lFtGboA
lWWn9ppRgbYWKF5aIng/2DyZhFLeeB2/tA0M8R8GZWJ/Tr4OCrNpsLn4VNX0wSEBeZ+CafslbEI0
P2IzhlckyC/I1Mu81qfB+eXBQb02GQLBBOxEr9fWLRCS55CEkjxMXdPfSZamrnbVJbd9/Q7idizd
8BsZGU5eK7A4Kpr3qgvRY0KFtLIATYi0Lr203a9PloQLV5hUoeRz3d1fRUdLgTFBVYBRFm7l9pXH
kehRdrARU2zG2cGoCdDMsIg0F85yezVie46QjmtXbUwVJr7mUobR8Qhsv0ZQC9ukr9QFSbaVYOrN
8rJqZOAl4gljUmWAu2dhkffHujw2EsXs53g+bYx8cnf54NX+XT6MlbTq0sSO1+4aaufRt9r/XV70
8FotA52EgnjnvagSi1qNSsshw8/0E9ojjp4gHsVbOeHsJifo7D7kmAezdxwZyRDSjhEbpNzG+lRE
tjN25AZR/AF/uJCcFgHir8N6LcDWSbk/iMapAejdAVypCLX5rkdPHmayb40DEHmvvrlhWd3SUx2H
5stz/NAHqTha1iAYnaymQyaHySEJrHIBXu7gRlW2D4xDcpUZ3RjcpLC1885xF+A+5/R0nI06yNaf
2vOl59vSRgFrPIg2eVfyk+62CxWTcRiD6MoeZtIpiCXZY69Fji7x1JD3GA179T1ZXWB3pToHAa3q
gb7zMRjdtrdsh8O7knax2ol4rac0SABaY4nkKd2tZToJTrlNVAmt55CToB3gopzYQR562EOFG/k7
lMtRcuHC4EcZUCK1IgeSNv+siClhuKgLWbk0KrMEAWaRNiMskgahtP39HtO+4TbaBKXC+ZVTGipp
p+FoIB1tvACudJnTSZIJ38FhPxIaS71JIhce9Hn/xli4BwjrVDEdZvb/rdZyRpmYvFBmanBFSCRn
iImZnR1vAk2J7uQZUZ36TYDPTBj525E2yo/+8VSyGBSjIexjNKiCT3THA4odm1Ppwnpj+t89G3E5
1PMnjg4EzRatdrIuFk7qWy6aeAu+QpKWG7D4k5c6wf2hxaPWBa6v2WdTw7IgKrQG+3n0eVNwwcZr
VgRHciEjaeJCZLeBAyQCy1X0w6J3Z+efjpzwNHflSDAEPajQ/SDwG0kN5j5JjRBS7hkU55AOaa1H
Gosjt1+q33veIE8IazSM7zr5CMUQpW7ciH8zjjFs5qeA7G0frWZhj8Pz2UtIFRkFBv7d/qJaN1rI
RMGTJXsKM80wFiMUqor/pT/0pt08pHDfam4uvddiEbu0+AD2N5CILV1bDG8qYEBMYF6Hh38ofmE2
s+hc2jdfnOTWuCwn75IslRc/9VCM7kAtq0fidTmluFqI35DSI1J6CgwHec/xUAS3pN+BszSrpmGu
Ti0CH/fvlJxgkZwyHHaHDw5nakcViiBOAS9S+a6qJbg/HsXrntaiHgB7Xf2re/mV+XYNj3AoELfl
39bSJ4gV6SJdA07tTJ7XQysLTvMMXFyfpul4xKUlotuETkjQkUGofpNscb8H9h5bDinorRQaPVCn
4AgaNQkapHpi9Mu3fylMlc7Uv2E6+1Ldt/p23P8+ynkmooQWHrxl92L9WN4lJXMFbe4ccT01gUyr
fMPZWDRX0fA5kpgYTN9xx9xgoAm593ecQROf3aDfbew9NFLpFqAheuWxM/8GZO880mKyQlo/woK2
Jt2rGWiyLoZ4yv9SLn4vQipTQkK5uIGT3Mh59Lo1TGFXuECzGPy2LIvUsGb7a6FNfB+goohPe1vi
3nTWrWLHJERyjFU8zfdKGBo9/62vzF9g5X3yapJy4F9U9ebJjm4PBmYlas3+d99NG2f4tmSouv5W
FityfX22iQEMO+SRI0yzVOfaXyQOxgAD726QTrwOWoQpPJFKPJ0OZB/XNlAmLCxCVKbjWQvf4VJS
MtbC1QJKgLrIJ2zVUCuGsodgjaONyLX03qJUlLRHBIsuxQSZjXOjniUPwcoqRbBJr8o4A0HLvrOe
OnkEEcIuPcBVUvT5PTdrTd86BRbAT1IJHVtZW3vKIhXhM5ydl3R6m6mqYWA55I5WVa1X55CS0yKw
00V/lfIQEN9gdokG4f1CextPfQhTbCnQ4jhQmiFnfW6RgPYOSlJf3JjwXbues2wH11OOLhx3VOpA
/nuOvpsneEuuI2V6pkc9X+4sfHrqnyc3mUfP8rVlT/M63WdloYhQkUSYJf+vDM97ChI8SfhCepng
eztoD+5b5TSIQsFsWprIs64tu21ETnReqgTXTCsQNe8gY9g1Z4ynsyRJenkMqzl0st0NZyhiQ3HV
LFmtudjaFDxRdwaM9gaCMt4M+Z4o3BBBU3D3BCGmdmKUv8s7VICfGdDJ/IR5QPXia7TbcJe/K7qC
FbqcRxRUd/Brvo+fUTU4+BMJi3g1BRffyHai/Bv7ptSeQx+82VSq56geRAb/3JmGUredWKFQYyiP
34BEm2hIg/NigqUe82wq2vhGL+MXLF1TC0GNsY3VJmZ65HnewsaeMJYP0xu/aVxUHRX/PyJT9Otj
lUp3cOvqoV3pVrBd7S6AmkNR9+O8m+uvdMRL6efmjOpGO9GwgeIEBk8/5wHv+UornaZTD2RV2xuU
btTbPfdZnCHwVod1l6XHiHk3j7EMz/U8wP3T+yR/QTtMs3IAI0sNaX/VVMBWI8hFjrNt9ck2GVRE
gWecOafHmnW6TE+btVtsNfRdE6lfUdHT/2dxObHp+61tcm5CaZ4LXPc5mp7Nq4UwflnS6ZNs4/cr
C+9GDE44Rs8rbVtT6uOlKKK2PALekCVRK2nKdDNGtwaUmWz8BS4lT9N5/B8kl8QHReeFGOzAtHT2
zyDyqMHdXCD0nz5UjB7muTTa+JSkh6aaFpSm+fX/ax8wRR+Fn4DmTDw2PwfvE/7WRQ6Wf24y1sgi
j+OUIVlS4sZBRivtJGPdZcUZFjjUrFo5c3DMPHAooSU+DGfa7mFe2XnX+HW2NgolQrwfvMyoCII4
sGA+1Vijx2WX6cq5wGy3Ga1ox3Q3q0TrCwyBzbcy4lrdq5sn8bxPcusfWCgkkLA+Dy5Vax0qhZc0
hqBX4b5uMVZtWgMWOw3nJ+joYgopiAjKDpbdZCLlbtySWULT6YsCx/wmtlJD8JhCVnv7MvlPzI0Q
gTYFUQ9LRLGSrgjf4jyIFs1DlQyc498eD4uGJ/S4hbuMa4KaSaWAKYEF4d5nMBdHnHdlkNHR7v+1
2kRfx3UlMOHZqgzCI85f9voe3uLdnDlwC/eEuYukW/84KgM+yEC7shYfpDyMHCtQNAHwBm3z3di3
Yydmh7SpDELLB0U7RL++WarBEWZg1SCYhABFm1Ttx8+/XRAKH5bWORJsdj2JSBPfzLOBuZCV+fsh
YLoxHK5XL9LmhVqfFWIjcO/MINFE3OBDjHJ7/b9g4xOpNjY2dCDNa0NBoXwLrDbv9M7K6ouEsbUj
iKWlILG50qq0upKrKet21eoHGgYydxN+jCvqZUyANM2SiJJTrlhUFNtVm4Wxta3JyZzh29u29B22
jnuiz4Tcde7uiWQH7HMstZC/16tkJ1OYilOtgA0bOndQADx1AVYzhFkn6uOJbiz/lrnmL85Ae/uh
rmaL0zKtKvEsGjQUs3FmHaaaK6WL4ovvMEbsFCBe8N5lEZ7BclMbVhbEm4a5DifJr8dNCe7GatIt
1/ICCgTS7kWnPN3tpBJhSdxWrC3z8QM19FatUWeniPalFNBpGnr7LpwgvYzsDeBsUMi63C8JGXiD
27BzyjKyln1+MFDvikvMUlfq5RAp6oMMPYw3TXw/74lT06AJKEK9YWMH5h1yMh15nNtb2ByldQvO
obPr+uyMRrI5hOmAxnxhcIQQJelhBARq+IcOZnwrGe3jeq41QA/PoHQkluECxB+H0Y6UTbNft1Rs
4qEZPIyS0mmK2rC08/2chKN7j3xYth6ZNt00wB7HiHoZ17gbSePyc2H3GmZF8JxaxHXjsoLtSLup
3aDyz7PFmIUgqEpMuVyOmYUYhG0xv70ocNpcWdDgRuYQIZcI6qb1IOI/kiFAuBZcZqbIVI9KCpZc
y8sw6Wb1HG+iAczl83c+PQxigtg9aPPjVGWMuKd8aCgrtlD1lipAuTb37b7ZZjNfUzHku76Y+kUP
EvWtLXJzwyKw7luBIOwp4/lEousFVPfzr9i2F/e4L+XqrzejSyOuizJCO0WZOcW7i6ELMCTMJ559
Bfayw7BF9irqONPMJlbYeeidwqyzmA0hQZM4Ozee440rZlc3STH2zwhmSKtexkiYKysh9SW4Fq2z
LRzvCSLmmSkDQPXZRNGrOQ5/8tc0/TB6zWJyyWcGmvlCDfql7h3UgquGFrQROZIgerwwREuLxC/X
VbVt0GXWrS2ug0Psy8LlTeC8cbUvQ7S/vi4hdW0dKfOfr4dYvAOtp15oLwBSkW4jYUXeJQeqdhE5
NwCP5o9lYA4O7KIOmiHaI2EHktvENdGWkbtovV3akBCv93SQGrc3rt4PnnGE4H+kxvnNttqlBZfQ
J2kvkRBYIbGZ6aq+0DZpQ1DSaY4upy4/XxF7nWhkzMfCYOjVhff5mGmOhVkDy56nkYvCzofFzFIH
D7OElhRVByy7NbnXtKNrzXHlQ2FrCnb9N7ibQ1sCrDYamlXnQWqlk4VvvO3EHh3eXiKzS96APXZ3
9sDOd+4vJcFm/T3l9IzODr3YOVNWxYrAd6SrhU6/CLpX3qTJi2kc+22kttN9FbIfqtsPJ5g4DmwO
6lO5mVcNum9nfsPgLQyI5ClKt8JkFYrnzhLli8my64yB2gaGwggPuT6EoBjjbSTP5hICPAq54T/6
8Aj8/se7lJBM5uEOcwjSPvc1lh8bQO1PqE7KA0iv3H1W7u/5K32PLV4KOQo0goUOEXEF9NaTv2xT
9lau6PSWivmiVGu4XZ7qhl5OnijPpjuUsf/k0no/csdBjmyyFgnyprTPjebnzx+aTdMxJpolumCv
jre+BeVq91xcTv63U17FmlW0FwbtAYhnHpt8huipOcqthO0SxssqU5DxTu0DommNy9up992xv/x8
/RcdC3gKwGPYJeQZOpwu7vlpiZU2YHDH67/HPGyo2znetsJIc9n7fPdAF74dPhcl6pzfxGI9MKsh
gTb3mTyi4gCX/4g613tTC9Z5Fx0Ys1ghdLgT2CXpcUg1H0ZVDCrRrcQ6XQaj/VjcD8G73TssHExl
fXxyrVgIFMdiurl/RUtXsG66p56jOrNDqeyFlPADar6sZ5S9udb/fK8DP3LahOswDKkpR0X9OQRW
hTRIyIYTXKz4Dzc9L3vJF0kl7j7p2i8xywmAeLvd/fVHiJPd04i1A8G+ob5awTUL2tSqguQNwg44
W9Hu2IJ7zLo5nPagk9+W4e+BAXDH8ydV944FQomFvWga0A4o8veccJo2EZqugvCsk6FoB25jIaUH
hASfZG7XEhFGZSK9Trs8rN2LuSnWFmpsQTy5IpYOyqUOACRWM5fRdvMCP/P1KudYDh22yl+5BKPw
GtXvdKZynA8u3UiTXyBSAef/mUiQercsjY0llUv0+cvv9TpKZP76BkuR3FPrm43S653xUyYXbq2p
eaHeoxuld6XMlikmOgBxHO2nZldfExWDl8X69RalXsErRik6r+xSf2wW/urzOIerRh9kEQaX8vEl
PqiZOm3jQQiIESqfAN/JpstEVcsDl/4SJp8AII3Hz1pKX4Se2gJX5FBB9xVWWCvBxtLgUwzxCAG+
qyQEaerZM2Sgh5Upiz9rpP596qFMxGbf9YMj6k4qlPaVr+wEZ51B7jE2kUbxjxRdxlpeXcQ1EDXL
CBC+5JbHm7/0O4c68MPEF+SmZa50k3ZuQVuZpZd2tGJb9wueKrR64ZRMP74PVncC0L529lDKZmwJ
VqS5SygJi9S8YrKOYVik0YAi0FKYiMeIrfpJ5CiLNzI3rPhJkpE0z8VTTRcze+72sOWgq5iSusm1
s/jrqep2RUguCiB2W01a3weFaqs4XFs/borEpfllJeyeIL9NAp7fl7ed/iNhDC4SrqEbA/IgWAlW
IpjsSgGChsfZI/JDJ1ll2uiNcuQvByFkJj0fIIWJBpiH0eBWiPkj3WLdmbDBJOsMTzoLZBJXAiIY
s8+LJv/kggwxMw9pRH0ODhaY8o1Px7XMEKnFUfIrw8kaYQJIqqIWTZG3j7IpnbgnzWUNzuGUwlkZ
moHVGzHeY90Ixl2wR4rD+/Hr+hzirdbQUclsmaScrlVbHl9eBAHPn1NKC5MUdCQNs1SPIGdvi3yZ
qGXBP9gNnriSjAl3r3rp5HLCr73sYoCZHF6WStY91jCqc/SxJmdJRH0N/djLSUIH9zlO9kMOLkqX
eSVtJHYlAdrnDvEZQRA/co+lAGUdSwgLOP3wgA7dsfT7+Y8aRRx795R8QE0XLKqAq6RlZ2Xiqua6
2QskJK2gU9fCnTG3b6xauJYdlLbWQIHT7k+LdijJQz65aleHue68dvt0h7cJQyu9ulmcK/729Mvg
pMPuFvQNHVLH1bws5Aa2crV5n+E2o/zDO0rj7+EAXjdyBQS/M893ubXmcQwRAm896V4KOoVdfROV
crbopDHzzTWk50AsG2jD/m8gRb0Co2COfhtUopoXjlF4ZBPYjVjhyYXrMtquAIpC8IyY2Rdw4vWd
P18ooqdwuOsOe9TC5AYrouut+1npI2e7nlhY4U7ueVosR6SoyQ7eoYurxmZdIMd5g/SGrvPH4eru
/gfXJfsPN/oYmYD09lHAJYMA7YSgJc5PgS/V4CXvDLQz2SlXbcXqhInly3BdKij3x4ObEbDRQIq1
UglZ6astF20EY7+Z/5CzbxrI4Jifh68MInHMxa4RO/QRCtpa3KbUqfMfKcUZoqiDzj4TZvjma72Y
cn3idcpIDuEX2HRK3hKdc3eUpKs3s+X6MC9ZkVBXji/RWV0RXcsdYbXK0AoZ9di2eukvbiF6Nr+Y
5qrklNW6Qapvl7eXo4Hxgh6rd6tRpf43hOSsWL8+mR+eoUm5mff4v5rDBD92cR5b9O//pm2JmvA3
/vsW8q/CZeWPGaPUURqMFFQAcuexIfjOxftLh0g0I69CoQKhItWfIxxgkK/X2WyTHHd5Q+hQWx2J
X0z7aZn4LLf2Des0I0dHePfjGGGjbMG5ZVZnu/NDCONnAC9bRCjOYSIH372TxAecvk0uBqLKqNRk
78JblAmz136TWC7NNR4WaKXmZEewfRO4nok5AqxSndBHThzU+3+ivOtr2KnUrE2CcTXv9f1TVqo8
MQflenlkKcIoAWn5XKYuyI6oYkmzK6sd4In+CuWq90YMQ+PoT6rprYIPSbop8HjEKKP8sIKUgJ4m
hcXEJ8jnumZ1C9gJLh1uikH+sCyV0H+W+qtzjNSvXXowbeI3RiO/ODnHQz54jrNM/KBfjPpFNlkF
vDMqKZpqXTS72HB1rUTL7LGPB6ftEznwXO4tkGFAqn1TmYFSp6U7OknwhszHYdCq55ZfGWFOQ634
ETbQBxPti7s0pUEJZk7JIshHwkB1m+z9yRdGbbAgNPIMIPyPqsO/Hnt/39eFqktKM2yaXStaT3+/
WdkZxJeSen4TBJyKAVeW0yFVUTx5RXZVQjhdJsEbW6BCb24voqu+wsIIGUZoof210F/eV7Plgfyq
ZKgaT1hnfTZt35GZJ94TqxPRr8WIlovMxonGfHw9LcQpwCVPkwLhfgJ8sh58jxZIRqmmqvfiVjKF
mf+/6ViDK427KYreLFBIe15xRvZV6v1QB95RVNhH7ficHIVfTQdGKKc0JzPjP3LXYz7ewSwFBSWi
V5qTqAwUFPExNfaQnK0+uYdBv7fv0INbI6mu3YPkJBiTnA1o4Sf6iVujMYnNbKtlmi/ZvdFpsL5W
BrfSoeU9nDTPCO/Fdz06iQpr7qGGLDjgiSQTidE07Oyva0w6MhkSf/34YwySeputYpfDPMyaQhK9
Oo2Lr9bX/iZZ2rImiiu1VEoOGdRlseeqEkIkgH6Wka5ryuE67gGMK+rL38BUXFwLM31JrYvBGDQI
xNP4KiyEzEekUG80nMz8txD5AUq3OMJ+kO+E0k4Ud8Okd954EGKDVAHR8415Ch73pE7iXDhXVHWe
QLNXY+PI4rCzYaO2nnxG6EPr65uq2Ytr4lNIy5c3RGoqBokGYPL/nkqiuxHS9m5JjPXQR63a3kMU
s86Fby0OK17ypOlUfJJZ0W8/NimTlbQKnsuuEPbyCq3vxU8Q2dr1Chi+Gf6CmWANDTQKYpO346VG
o1woQwSXc3L4EvyQh/6FRd6ZgzogLNkb11k6DtJuBftStxQXoiPh7VaJ14vahVefsB3cPeyEpyZm
ZisLHStgqArlGxlMpQNeiYnnTyD0SH2UAAmZ1SFXB1le6s+H4kKanlM13bXbHsP9TWayPoLkKqj2
UVGcezZ+1S3j863XTHBatAevh5b/YTiPDqPEfhRD6t1ZkhohPu+9HPeoei6l3nTZd5XcIMhUN4I3
n6x3QLCBbvZegyo0P0QGkmwTcKrOYphE1x2+lK2LMozudqG4C7m6ZYWk9x2Tu2XS9kviCbn7B+Sy
z+1q9RdG/LNH9A9Jj7vGiqPnUZ0bNMj1sW2CXdUj7zOkjc8c4I6Ur1EHcTriLwsZBCSazQOyG8jk
v0lz/xJUQVCby3q9xfe8ZG0EZkY115L4GOtuoUEHwn2bo9H8IpTNNZL430oBkqQsIGegXl6TShkd
tC6GIDg2fosRcKJnkrePTTCXsN0paTa0E/Ea0R0mXr/D0OUxLAVcGbfG/zTtqJsrFWyGYN54uRno
cTZBt98FptMABe9hrFZHtSqRKdeKKD0e16mxeRHsJuCrNnTZxUm5yPHQC2QpXnJRrR4qn8P2ufwy
x+ZwDj5yy8VO/uhopMUIPO3pJQd/arxGakcJBddHakpS9knTSASzDk9ZnkPQPijtU3D1V1k2V9lo
w//8zF1udl1fDeUL8LqdcoEZfGlVT2Vd+3kqiH9FsileN51r3jKh3DxWm5nvRlrVzT6daRCseAjP
PBNjUdR9lUdXdp8zotpUmXVMVDEEdbs2jvI9h51jZnEmLQvAwgbTH5k8p3b+JO26ViKYxvVuyNQa
EitFC6ndVCki2SdJ2pTEXqujXAYcdNQmlA9zssSrEuyTwvOiKNl/jv+kznbqPovZcGR+c/Kvyt0E
AQ0E57JP5ZNvEehkzyquhc4Zy7gYG9LtY5ICzk9iTrJ5UZAiQNi/neaKoosNoif2odaqNRSkqO8t
LhnblYFbzluq9spuxZCxm9PUJmjHIoEWJctm5JMpdqlfexFmqEWDiAIDIILWzQ9hMut2esJpeKEo
290FEt5Q9b0uoVLwTqhRLry9XgLPOcZaFDuISgJWea1Wx0JOtCDsG0Z9edLxutArJE5eqlnE/nzp
ChQzTRZ6iMoceekuepqn52yd2JHAJ4yZg1KfjZFnB1MRUywwmn9mD0/VqJSf8zT/CWjzI69o+AKx
yRCQx0GJEx0EfgjZki0CmxI9TdOBH8xBniELUnh4VBTo1SQQePW2KuB4nDrc6fl2S6VxC0J6GMgE
mpgD2dqxCauJJvGDyGd3GrdAiEaRSk/uICR/4oGhpyHnzCIwtd0zKwJbxx0iUuwLUPLUpFsZ8Pud
k2JErKDNlj/UyypqBVo1npI9hUNXo6ZOLEvh0zYf+EP1ZaaoTn2QyYVKFLzr9HXMJrMUF86DmSAf
dg6YjvHJqrfgTDt4NI/sN3E3OrJP+5H24UYQvlWk3KEXDoIs2/GLJ99ucrScjDrJ0iZoNYLob6yW
0V47VF/X8RqzwqGvD5SISd71mUWmFAoz245BfAvKvLdSuuYpac5jHOmYLVn1gTvvHOcoAQjgGgfL
j/zNuxzLgQK0ffumV153hLFe40u+Nx/iMAMBM1FaPBuUmc29Ngz3TmgYGxSB6rbVSZ7BMsNxUXAq
wRGbM5AX/SC+4zPzxWla0zsWXfEpY5+O4EgxSXoA3qpU9Ar3+N1VJAn/UZK5M+v32gl9VQaxqszt
lm4l+FD+B3eprDoR9MUHDxhap5JbkxtcKaZW9Zn2Xz1hI+EbkhYQUjZREZ71Zddx4VJ2K4IO1CT9
mRye0kHPwXavJmDq0/BqJEeX15mJhS07nhj2Nx7VGkuHMnJB/BLG12PhtbKiSmWGAM4liEh3Nq+y
MVRFNV0AhOseSTSDSb9pAW50m6l2ThSwqvA3eHMW1oIQ7T20D6xEmShlXlWIFFBSk9LOMRTeqK5m
kw+x1Ahgad83pGBmLm7vlyxyl4U4QWMZBfqPkYYJCVmH8WfsBtWtdg/0DWqAbmawQ+AJaKOq0j6b
tV2TccefSX+fF6oi2Jg+NuX96PLPfL8+4onp7OJbhWw0mNKCWQk0lxqNDA1/3W6nl2betMufZdA3
LeZibQk7+sAKcYJTJe3lACMoHFvm1UEknrFW2xJKqHGmg8SXFAU9AQg2/kIz2/nnDNFhR+ewZS3x
tnMCREJF5RFw6VY6cSjL6KQPpI8Alo32g3Hnrw8yF+FJHnb3V89lGVEOBi3PEmz7CVfNNdJxCSlB
y6RR5lGutm0Wvkdz1scA9E2CJYfV6W9QQb73xCsR5x1a5djV5ToQMecKU1rDiCMKsbATucU9QCaw
GxLP1yM8Foqd9mm/1/USC97rODmywFPUJDTJpA3hH18NBwOhyQP4dacwD6zLJ1YAOI9lf481+N+u
Pgli/fQrHdUremSIZZ5+5fKVH1n1IN9CjuKVWIVH7/csZ/a7u74ZlcLAEpbxnr91SSlzss2Z93vt
sLFPiiqCbd9lqn9+9Nq1sru+rnRK37nxZyc8IWBO7ZpUrxBB4xSfEM333FgPQO9LRoTsL4sL6JjW
ijapz+N9i2iJSnt5PIQcLcjxxEAF9TnLNRYkB6B91ZvtWOnjc9mLSTmGWnb1zu1nJL5dmNQ1kQLL
/8rQJSTeOhGTvpLppkwY/XWLL2Z4yxgiG8/jnQQXix/QY2OgZ9jr8WzEBr88z+AAAlbbwe3P6TfW
Kw9QffeZgtyBrsOnbHw4Lw1jG66arhP2xU9QnYCocAPB4qgvIYkV+/IH61M89l4iLim2sy6WWaKP
MNBRtHQBiF0YlI984nEsGnLSjhMdDk5xNMwwBEDJmDFDLOUDFAEUK2OyMi8mG1fweyuua96fu4oK
CHx6my9CQE1gXfnGU4p9X8RGgQ2Py0KW9InH/AP6b2u9oD+c3o5ALg7vgWfCToIi9PrMm+TtTSDe
xdMIH5Vw/ea55e3cb/7FTl9UL5I9xoLn7Z16CXsO4RdaflhQyYNEdNoGN+g4WG6Y7oXvthc72EQI
7ZJ/E0jqw0Uli8vCnel9vTDAZeGKBrga1S3i9RKsjXEy6RTbMhGaC0yHYjwBpXOcKkZYEbh2hYGY
M9SSJJCedPFTjI+UFac1+oHGYGPQ8mj/MWvQhGaxKPZO633mCzRPsmRZIIHM5lVZvOE5401KTzlJ
5Z+kf3rpi2MYO9MrqPLISZAhYxKRj40llzHHjb9fExCjv3H9GnJcsJVzoYiYb/hQyAeq12ue0j1r
tl57NmQ6LUgegFugPL331resaeIc5ZPliEEs9yaQAiPY5kdMPGCIk1lKAEOOslZb1MT0UW04Twjb
Zvql/ItcCvV9mh5rHfJaFFIYwqyryU5klh/Rb2QcCAxcaF/QzaYvRbi+uE6BRDpdxroxl328I1BC
uPBKgvsIOSfhFk7lJEVUtTz9WG3DJoxMmMntKxA7wUZ+qcae4llzKFY55i7TBMjYX3BO/36jR//L
mDDI24pedusuAm5Uy+o9plbQmk20xN+YGN2zmgHTB+FJ8ir77jA4RIV7dtbzr+RS4LYuo+RhqXga
8QiJcIiteNE+QtvPl/UqY2YXd8lbI3VYHFinVPrPfMaja27BJTV/4tXiCxdsluMGqF26CnfNeu+C
HRgHCwEyf/OSmSvaUoXWMlMoFlMhHvuPkhWNe6qESMN+lCzH7xH+Liao00KLC3aTWzUMuMJX6t7Z
TVNtuSUYJM+0ttBgB6Ah6Rl3ph6Y5zQ64eMhVYPAc1Pm4OgGRV2CtNFum5IVKZOqxGRPy//KikmI
ZfCiUOn3ECMdIkf97ksegk0RsaLeUam0kD5Ha9r8OIYrpjOaJPZCkwDDIrF1DmaP9vEhwg97CluZ
IWRMDraszrkWF7sdM+To9J8z+WmrDSTJskn9zjoFJBXSpYeoYU+ARtQUjsWjHStjsz4rXycblCCY
6oZKKPONZh/OGvzgebvo6YJnekFnjuMPu9cX41Jz1GJ6AB8pqrR6fdfue/8fFNWUH9rPhbK94XkT
QVHoXsfV9TG80lOOm1tWJkiWgA5Ok9lo8SPsFa75Aw0DzxT0/IzUUu7aPo9HN107e3VbfQ67bgt+
+pB3bTciuNzFDL++7O72cjtL8/Ac8CitEiLyyvtTvHyi5yAa8EdJcXlTr78IV2gtokt+O6DyOp+G
YkCF9AijQn1yEIu0OdPKUhkY70yhfztG2dPXYv8QNa8TJ6n8/34cJYWZLKlRa4HbUpQHv+3Fd7nb
98rXoDDWALIPRqX4E9Jyic/n22MbSE3EHOLQiqPhCGSj2/nKoWwBVYEmGbYxOi3+Q4gqVZXyDQpJ
/Aj/icQgQC22C5GAMAY3/0SLxfxPFOERYU4soEGDGo4U1uj4zliTjIy8vVdowpnpeIk1baUt2gJL
s0tAy75MRD3UTGlKGbYKI1VIVw+VcLddJIptydUWtaIvdLFMDnToyy3QYLoT8lFmsbPDS4aBF9VK
Y8WreYX4zFWKn/FKGyoU1/ZwmorTcbBAUpzhTSOVqwgWeGUFVuULkH/zGRVTv9kZ8bioxW310Jbh
RSXlrCONz+REt7NdJArDO149Rveoef7iquzP2kicOi459FhX4GXwT8zjFK5JR7V7ilUZZRWbQQ8x
+GlEhbybVO/sps/PnNj5cIwD1Lf0YMxwXJe7YlKev7nUp8OYDv68szGq93hjgapfbtvl9l7jbvEw
X0stH8+yBrgyBa284EXFOCCgJXQ3pdlYxehqcqAbhN3qtDU9n0eVc63RvWaE8DMu6Wvyi66sHfxD
g2eKSl+1eT2HcVYwgeXFth665xHhI1KjVPD2Ty7CmY8TT/rY3up0KhA0oU1kspDDmF4PbxDbIQVL
89903P19777U/IwNmVqgzdaGzXyue6G6ILTbYUaQbn5WIV+Q2SASGeAgvkCQhyt6WvSDbQEuUf2j
7PfKlFZKo92eyP5+vGQhatc7LWx4cSTw9pwD4y0EFyl/U1D+2OB2Gize1ZnYUAruNyIMWU86QMWB
/AAnrv4bj+8Z4eKw8dkauERhbsXq9WveQnEdhO6TjzaNHXuWzvLPqL9IrMXOjsU85/fulc9CVIXm
XLCokMIDoIGw7B/X1jlx9rrqQFiZeMIKb+xvLjXJkDIEqa3i9JuCWYQJBAlvY1GHRuDfE1fWRUqB
ZsVit2+SxrH1pqmQvy2UkTCPfecEyc5Uv/XSaQ448eLwJ+GI40MaVHLoKoYtNdVzgFIbJ72vxM7U
6sugMo2ESTqivZ+TMn90I1To5JkrBKo1S3Rd9UVabtE1V/wBRSCJ8Wo3u5jv4IJqEfVZdSuSXeaD
hA0mOTWx064dR7otFQyQ1BxOgrrLxX7LX5Rht1WColrHLKISrjHU8bBzLbu3vo6NmtYuS86hHqYG
4hpXpKsX9XCpKD8MPJXuxvDyuUeFpE/5W51uZMCVtdzWu/bRDQ3ZJR9uaLYYIAFgVKhGRDJKIb+8
LgatrUdcDxajPD8iQl/g4pAW6Fnf3pDPcIoFqYO+QIKxGOcfIcGAsPbxXGA7nU6BVjtLkQ7PiDLV
TVh4z5Rj6g/i+8Q2sD1sTWB7ifWz3zZCSRIh3mfBFUlC0tyTkqeWRGdlgyRg7F6VsnH2sczyE+nh
4Vsoc4bQwJ+tNg1+3ArEJnFNPbXVN1Qjms0krQDQNazpFISgd6xttGq4ry87JPgAquR4H/PPqkcw
TKtVheF7ziyaBaluT0p4IzCKpR7LVppyTbPTxnAZmsYL7sV5vZkoF3Zkf+C9wop1/8aF5CH9/Xlc
vGKVDPDKBmuS20kkux7awqOCt0ZW8Nv6D6+4v6JIL2N5MhShZxUdtu3ZJgVJ6+WQgio/JC/m8OiA
K9cxlUjRVWAI9AcURhzMjYhAIOc6L5JyT7Xj5fG8MhlAapYwH1bjMWjaXsUHLhox2QxzM2R36vFA
u3Fukw2N1bp8dtG/lnOKjLlxKsaoXvYGldiKgdJOJBeAZ6bz7/Pe9lNfmre5t8n1SxUk80gbRZ0b
AV7Xi0L3KcfrIUnPXRYjrHZpufarH4o9ukasLQLFKdsZmx7jGQGEAnqkRYF/EOCHUqFxp3FGcwWc
HFzi0ETV211UFZIi/CvLAFb1w0qeopopbim7jJJC+62OfwbrCx8lg/6MACXTpowfcLIuZ1akk3Sn
O9Z3YtRAU8nnTgWO210Zw6AmnnCT/urOmR+hHVRszXow7R1Wr4kmwJ7FyIKxIIjuXIRDjG2dXONU
MHY7K0JU/8ABNmOTXsIRRqp86Foh56xb7JiLc+J01rlepDjrcJoVyKVWDkJkhOrbec58GpuCscrq
lEOOApXKf0LVM0RiQn3o6unTIOKsZWxKtDXsTlMjO9tLBCRkyYEEIgQUgGMl3zl9Y0EjE7HQyimh
sQfHE6IMKexuAZmpKBPgPY6AIFu9zJfNEuyoNtNWFidUs/ClyJtLa6gcCTCy1NEgH4E82XiyAOkx
BItlHkiDmwsKj7tQvcBGIOlDNCgNvCpnJf+btq4OJs04pypgxAO3F4QHW29+vQK+ADuiWDRZMmc2
HUNNXXY+EEGyfUIBRDw5SoBX0rPE5gcmxybCR/sJ//8m4GXvI3lcr8TkmfYp+emGummuwZs+vtmt
lRdTRN8JjBVu82PvNTjJmOXdKoS0sXBa0kSWztvBLld7XeZvWrcuL8LcCgkYD95iftcfx9zsfpuK
A4ZOk9cVEYDpE0F/6yCLnmeurEWOFEgbarmLzwalTEgSAGlXQMKLSlIgtoSfHwzAKnyck++Il1ug
KH+JN5X6YggGBqKE7+onoAlrwE/Duh476EhXDNGq3y4traO9rcGeSVaGGWG2HRwO1pn3mg2/XMLL
IqH0VrOxgwnkDoXcbKcmQbLFzsH1USFL+YdDueuRHLPGbDmL/+AWxKhWxeD1Ma3tIkZ7wguIF9xN
wiGGY9a7zTfTWTyhoPifkb/z7JudThVCA1AWp501Xmv2Wto9Xxpn9Kk+y9QxRQhyPk98K00FvLsC
aAsAzkvLJxunAOdNaiuIdyKwm4gRbJVMkMy1dDLFUJT0Iy0Kf/mWM4Oz7i7RNMx7WUw/IU6iyeuI
uLNaL5yuKHTYvzBHAgoYU7i1xHvlBatqTkhSMpD5S9YlUn4txl9JbXd/qaRa6alfHKVS5kb0paSm
mop3jSZlqIHFL8/BVcmkhSaRTH2BseXsoRJCdOVD/VEvAFDAaD/NgaMP9NgxxHzXC1u9Qk+yaXui
BJqcz18IiVNFY6LsBxssCAxqtJXRo/phHcsE7wXS4rgsAfzmrcnj9dXNXbLU67oFDUC+p3NDQ/BO
td7CNRpL7tZBiUeh1hoEPrqmRrX5bsMhqy8P6PL+vd0UMJBWwwtY5THzQ7sayyBEWAs9PgzbDEFE
I0mrwKz28QMUNBsJDZIkHUYjYruszYceGuerjovmC+hJ/0hqbwnDt7qiA86iVMvDDCDGO/8CPt8p
bUPNab6ICL+KWplG3hTmS41K+XmwWp0FjC+fwd81vqn64ik95V8uMqwBrHFxT3Q6nHVHbtv0r7dZ
sff86bV5DRwyXr4XYH4+AWpCzt9yUyZLlfaoGn/p4doTpkSPVbA4yRfMHrzg7A+Q8jyOv7e2KpC7
tQbRxWfA4t/1C4srdCDtSe66IuOxpvOMaCSayFXxrLAiqgIycoM3KqNwTMVIUeOi06qt2O2eKdE1
c+xu6YHNNkzyn1zvwN6pwwsUbpZo8Y4P0J7SWuGpow1/HUS5Zx1qos4StnngsWvVMjFhqUizJztY
rUKSK5UuPVGuqq5LDdQZb1x320Ubuvg+GEGEi/DetzBWdahqB2LInBg5V8Di7Cl0a3MZnjEfpyD6
nme4Xc3oWvWTCOBnqVQb/DpyFBTesch71Uq7Bjo/cwUoBd/KvThARiIl0MDHh2pDIiztlGCbA4WQ
uuEq3jXJT4XySGgD2iw80+5m8wc9PuYECWi/W9ITMAPljA6ZXk2pyXhTK4SOHNG8G83daiowROFl
r+lQiMluv+Fdmbv0CSzTQFeY9oGX1xynSMWjY2J0Kqaw/AydrrToBf1JLifBdHKORSQQYr86pLFd
RxZcT4moAvM6gk5QRcG6RSD+yfvyj/mNKzEpsHRzBL3ewgSsQi7xNEVJ9kSpH9tjS+/NID1NPhd8
3doY7/dnEJMhC2Wk7YM1As8pmr9Hf09VrOWyDkS+OcYPPW8sUHXhVWHoxxTKWOIOgQRB51BQmnQl
RUCZe9/1vDijTOVV/PmQllVVcku7Nly4gxVr7tj84b3Va20HLAwYjIk05tDcNngU2GPfGBA5/Kw/
OYzGFDwvAiteAeG/TL9T7qNckqCGuDAvOd322u+4SHdVKNOtNLYdSA3tgYfbCFfC57svhdnUmaE8
uPQ48YKhJjIa2asaFvxtTR3p5xJLnV49c5i36WQ9IFdNm9x7k5AY5Mg6bJ0WSHjJ3HpaUDz7S+Qd
fx2kxUSo1IdLZy4sl32JT6fVtJF2/eZwUvIAYidgzcP1IvDsSq40N7GYEFiDMDt+dMFIFd2GldBP
ySPOLvUAttvTRP/S6RB1NB1lcEa2fW6TZR92NnC5SE8hHlF5XDzUfGdngI3HlHTTdbPLgt44aDQp
OtXSMnHanM12kzljzmPpRLnpUK711KTAsMUH88GBX+QNjP/bK/pBZl4/rLS8sAHeJ3TcYBiBWxj2
rrIfe9ySkrUv/bqZmrYJEB3f2BCjcoPHXpLsZffxpbm9z/Et3R/sNN3GcWH1B39iblwCwjEPUQZR
PeC3XV+wu5RHshF7cNum1pP4RzEhdOuq78BbJIc23tlVRKkeIRwWbf72kxyDN164xDvtfTOd7f16
xsabHP1Hh6II9tai8goBVpucQlQIihpsNlnv/S0aLPwYubNW80LoLdO7wX+WZdXcsMocAh4xSbcf
wWvT2NBtpOpl0Ha2HEYZQxZcL+6eTX/cxfojd4kgC7HVOr8HrkZlL48OQM4AfgJ107Jz3Zh5Nfkj
fzZcVbFh5aHOor88HM+DD8pbRRJ/KBBykBmnHQJ0hVeOx/VFMDW7noyXaE+l5sNoos+B7k2KhPib
oQo68G0/rx478k1fPhlsFZ77C4OWWckxMPTLm19sxI7WSFxUsa5X1orSZd5ft4drY+yU97eiLPbj
QhXp6CnjnBVJ8owVo2zsxRLnIKWNNI/Xu9iHUXPQNeJeo5biSF+W2VVZ3IddLMlIPgZrG5x3q/+T
VZpABoKfltLSD5jY+hMxF8PGrfg/OEjxFxeQKdJ4i/3g+08mLFOpmPBHhj1To4XZysAjiwl+KtbU
s4eDo1DPlEKxaehFNsor9hRKBa17QlI45CiTKMUNcaVq0xAd+g/6jiTqYi/boiE3sUjIltwmRTGk
bDDMq405chfihsH4kIf3rvHEDfPD8IN5GCjlfhDR9aKZCRycpyrV92+/Q9ZYVagBMbz+HAdvOS//
PTPC5fqv0AlEimZMtrOEzrbdj7br2gMFs3zJDP4AsDnGkcOjAq2tITWdVhdn0EpITPTg4Yz75jvl
sgVvUf10vR/CK6cKaXNhJbCp6Q792EP8tx79uWhqrG11fyHr1aqwF1Nwwwjwr88UG1dvO3qadAOP
Dhy/Gd5cfQvluRzTqvEZsiNpVqOfOX4w/ePa20dcJH9ClzDMgPIp8CDQHkieRydv7q+4h+TuUULk
VW7NGUjVLpAZKPxiuDl5OLXU3Ye2iglCPLufUF1+CpnsXPCLpYUwgFSsdQUgaLKapxHy369Ozw5j
3kSUgYDVaWkaWNLWUK+J1Q0AwZ1oXcd92c5X1Fxpweu0E6VyEFQGb2buWriHlvKPUcPbNgArUIFO
sm4v4qbRLIfRJNn5Tno9x5RImK6zkfugWwsb8nEOgBWnG5poYuju/jGKfdg1QtWVqussmoY1B2pT
8li1rLm8t20L4EkyqwnXNN4qHsVK0knGkIMq+eYnoFFqG5bTH4L8NqyGVuCaTDaLXZUJx5eG++As
XAHmHTxhisiZ7ei6gce1ZOhYSLbwvpggOHu7g18QNZ6QrjuB+pOjobJGLXs5Zy0XXgPb/Efv+LrS
bSQXAeCPDrPJdhK0jJFPpsc6m9WI142J+iGmctpS0xZVGPKmbImUQtkUk/FJKAsFXwoGQSdvyVyT
NPXmjkns4qHio5qlLCSZUztYMsCiMPW++/PoKeeKKqFfr8yaIyNJhsm7SNtOz/jquBHL+JtHK4lx
59cG4dcQCZKzHBdSTX+boYd3hBUuP1r8oKa66CSSQ6yQ8hXtyHhAVpY1zgUXV+4w6zMn+HHXPZQ4
nmRxlZrln/QoZ5jNLJjeMZ43gRvgV/EvrfD2Fpodg98iQWIseJStRzkrXr+K+hp4J19Xvmubblup
X0VAKVLKfoWi95ezlESMlZbUtWMR5hfFkXTMu4NUrDnwFf6hBSGV8cyhsm1bmL2Yl8XTFWlj7PCd
oNxMtjsxJLEYvrzeE3iQStNIOOZeijC3rNIuO2xiQZv0mLBRH25l9qmj2/y/yc5Qo6eJbzLvOWnE
jaQcFWh/WEvaSvHL1aLR69APaTa6aGASFhInEGoM/xgh4QbcKbB8FRe8TSpJVheETFb4sSnGFFM0
zfmV5MrmKADSbj37zNofKs4ee5XYmVgY4rDVVMKmIQkvzeRG1V1qe0t6OJCD7Z8Pie1/SPAAkALb
YEgtLLzjBCJdfFEmyTfI0mneAAUvymQXwUqU/vHE4vIiuSJYPS1hURU8BeKZFkWMItW94kCQYnKk
zTxROCUc26AFwDWZOEniCSPUgajVa50r4JYv7uYvDG7X+PW90frwY4Cf9tlygQted2YzyiL23vh5
otJLspN9Y98ooaIpZh8LgCbT4t1TPmutqDYDIKxaM1HWbnOdz5Yq2J7b9ZfB8BKnxkYeqQQkSa+Z
dcHNDIH752WUem0qV4D6F6WREPoHeG8Ew99LfAYX/2oSWF4PQME2/0zYu1uVcrtePRGNm4LLSDcx
iFapos3//WCojlkA02K2Onk/sI+T2j6Xt8AZWqPHTy8IvWnO2mHm5NI2Ou3EPPINAzz2kCh3XwU0
aiXPtBolzEaPQ4gn1LKcPDBtfsMwGiXfo1JUUo2ZRBwCIo5wSJmokHw6OIk3LHPleaRJWdYYINQS
yPoW1hrt0aeOZciewxLbNCZtLJF5EDJg4H+R5RoO7zuKLBag4FOeM2Dg3tDTCjBgPyveEqo2DhDk
/kenEgdclp0a0tIFcKwkFxHt+gFU1ZBwezLtfPIlQAGDSziCI6uO3R6Rs6TODxxWFNx9iGTSIThS
epDXTLVmQ9CnN1ouZT4vf+/Zf38CnGgeH/Gm0U1bP1/7+oNZW0AFzxgxfke22e/Ks9NbxJqeq7go
JGNx5u3gntaio2+fQ+ygHU+Gl+ZDfLIUpHMwCCZvzGtd6ZloEs9+O6i00EA6WvqwGLqFfyOP+jf/
uItDoN4olDbsbsJ4HoDY6QCLmHXI3OUKkekyIBxUh9qin4hgzRYw7io4Fh2RYCWYNaQQ/wtcgyo3
moxyNFYQ6H7Ykq7x6LLN0dFunKgK0K8PtWqyj0Thhumy4CIne/vpwQe/ukop2rv46iW1SWUmmeoV
AXLrisTK76qwL1IcBdzjwSp6lUnx7xFmKqvNmyLx1xH3iF8oVTfM88wTFcGaov2gSGGhXSIFJTuF
j2SgBRX3WQXLl80PLDwcQAlLp4iKheBA4fCmwsjnjVR/gbbmdx61vIiJdFDEesc0CfEGRMSdORy0
pu4nl94qx0tdA5IHJXtgDS9c3fgO8I8TM3NT/fyVip300S/xoA7xrcEgSTCg4Nhqvud74VnJMfMa
4qMI5uqla/rrjRp6sdQEDJEIeYOuJeJzar8hUk+5QPrJwmmLULkor73R3qIoS+XPi/MLAPo5lMb7
tEUIEHokGLMJd0tYm03R3BnMDBKvGCUwknfFiZue9U7hMQc3Bk6au4JD+XHgght5TjuAbjXwnXML
wdffCLwf9Juoz06dhCIKd8aGuFtqH5cgp1QiL9CggABs8uSUqVQFtGFA503whiXSSx6vzEkLVf52
1d9xQik+tNWAa42BCAEBQz3GhNVX0+fb6yy8P1Vmh1zRRKeiCcrFGjQJxXKF924/79dcN6ZJdYt3
jz7rCArfmXkXo2uR4XpjsTuKs8oUtcLyrrbsoyk2HtaJ3U0dQOjl0CY0BqaLtShXKTEeefvmdVy4
IMZyRk0FB72PzOxc3AEYZIQLRwgqhw0eDyupgNtjeTqrwWXzt37xNnPXipCflaF3dTq4mXUgddvq
v3A9DyRxLY8xbhPp8za7dK2xoxpHI3JZsQaHCUMmNHhj25DLfr+3bxHUF74PpiH9big7WEVKiJ3a
HcT/o5gRpoeMDU4eV4AC8RXDpqj7bsX2UfMzuiO+SNY2kRBETdqj1lAplflCLSFXqDTkWwg9nOLQ
RyOTrwxujvDaOVwhwhOS2oNAwXQ2vCBXrHJJOyYUdQ1jK+wh2JbZxficGbi+VSEoAwjk88LY/+jA
ze/TJJp1olsW7spq2FUf3mcK2oVXMtd5KGMmU6v+nGjTJKgO863cJkMr4fFAXXC1/KJwOfD/mpvt
Lcz007G++tNaVI2WDopd8PFlLp+zPXcm5R93LPA9bsRf7zmyXsq4lAgjyHjUCSz4bq/BB2cgPJyW
INVRzivNMWUKHoL3MR/mIR+ZYSqGiSiMZw2FEBJFfFeGDmPKFlEwHh98dpKS1k/TBTacxxPzF08/
v3zjnDFYm32mDG5FnSOTdVIP384TFrE5wnNyBSGtYMnKDLRCKtgQMUKUK+pgwf+KXu+6hoi1+wIB
iKW9cw//LHF+Yn0wP1CCnlTBGAe5BOuUyvrlAeCz1YR+vO4MKt2sWjG8LB1e2PyEkAvBOmYDd+gd
Yx8u9X9xAgMKZoJ+QQ7c38yyPtaYmvo1U/z2fpco8RjXIqaQVdSR5j/ORY5REK+QG54BatAO2wYM
Cd1KW1hUUUqCx/BwoBoFjrdNqpVq8FKb28f/OHOSDRGy7cQkpxn0/S/A9RLvjaz8UHZRYz0UvlPX
yBw8p/zoGGbm3NAz2UnB9xVyag7y6bLrRtsRrenQbpCOJhGxkWuJw5q4cvWGgXa4y1xNUducad7b
PjVWtO9iuvGmxjG/rXZz8d/D03mwQPedQw1nbbPLNzbQjqjJVGvK/aD8DmELtXHnH3oaExjSCaPa
PGBepeFCA+gEGLDcN/xtGP1ePqOD7000qVbqlWvgfxHicMdbXtY4IF496j+PyYYbF/ZSmIjGsBg9
pZHuHNxMpk6DG2l38bJ95xanSt14HLJqtO1EkmxexCrK48y09c+PTmAsMZFzgGREKckDp8fdUbaV
61bTq4w2bHScO3gRMqkIKcZcXFLTo0LIfsLMGeBdWZyKMy5pfYBHKXqZE5L7Tk4VrhuHtnij8CIq
V4rjN6FZCdcC0TRLCvzO3VlV4axXeGRrgIm7jEDGhp7TwuCEXwsgz7XSBjwhhjSOf4ecOse3SEpU
MC998xmKsTJNyPXIhD9nlWWdi6aQ8imukY3zKi+AQQK1WXuVvzXh+MQoX726Rmwggats2sORjuxV
2m/kyUVylM5PxbG3z58tsdtNyag/zMKvhIhRqFzfetKwq4rvPW6sIhkVfvC3tBkgrSbBzO92FJOE
FQr0xrqFVsTdsaSqxGAg+S4z+HMwXvwnodweF1eMEZp5G8ax5gOFu5AYFFQBzfPPNAytI11GS/38
PJu3EM8K8gBe1+CIE4Yr9PCjMIR4W4Ydvpz8MHi9xFuQLsj7vTF/1v437CDeQWmE9J4roj+6iezO
VaKp+OkT7cIGChXD742Mo10360a4FNmtrpaRwJ0rzvuGnO/BupF2iKNStpHFJFrdmpBh9IXx4cuz
PJbRLerVsfmTIkgL9GX06FKJmyHAQ4LvHj8qMw5HSwLnobyQsPpPuKxyqF29UTbuhAFDimn/ymuN
ngtC22URTlQGbWLXpbfDmeOxxg2Vlc8rc1XvSK95XgbnTTTu6PQccNaCHWCoRFDfuQHpwtq3+sse
AYOaU5RkLSDbt6D/ZiHu/24MKBRWIjwXqefervRm3YIfodU0GGwbbziTdHIZauIxxfyRxpuHBpmz
8KQcBF8jWRwnWb9IfhH6TNzpdzh1Pszf8uLr6Qo+NQfM2QBghFDYKcZI9Sf/pANPqAiK0l5VEZj3
9t1tDnuWD+nG42FipikHjYw+hnTdMMcXH8V++jwnTjDgaH4xlRv9ShFn4rewbMTh6+AbpEN9pfg+
iiNTIhNzIlOO60JLhegdIDiC1Qqgi26Ln6SICARBClgJCblYG2YcQFN9zjCmW96mSs4SapgfzOg0
f1mxzg/RdlOdzUsk0Bw9HU/57UYRi7Kzrp/89h5H7MrcGR4TwlytZFcPyDxqachOLrY5IzMkWngc
BL0MoObrnpJUYCL6QvVwrjEMiPJAGMUpO5q5iTqA6iHmUPv9wKpFDGxsT8/FWouaXLEajI29I+Fh
dkPjNKSJGyJDWTkGZ41W4PZN4kAllxCLeP2/0P99CJ5uv8eTc5xxKaJwaFJBrv+WNVicZiZ6RLj5
MtnbcBq0wvixbye/7CvX8Z3oU67QSTg/Nf4UnOSgw+pUOprJKswduKH+u1NwZTDQIO72lLMN1pO2
Wk2uSTEXqWE7Zq+qwnwGJ9SE+2rkOE2k937eRecOZIQlwKsj25gTozBWvvJfKO4B/skANlnuL3s1
J4GITso8ZYfDyVN1eODWXrqeNyD9Dfr5omm/zFlU2iVbcncPJGkw3n9/cqqhxCPViarOKf8HWoEf
PTwyQC8c3Zq6uvY7uKWIUB7At9ruEk9cHFuEsE7M2cgLxZ3yLbyqdT7rCyh/G1JLUrGDhpHWyqQv
S5255JmGyqmJ/Dtit0vkLyM5DT6Kt5SeQukoaY/YeKcqfrNwtvfr9n+Te2bt3BqXgP36ajqHe+Gf
sT8NLetnseMbZ88lkkSOua9nUHM6fZBPhJ3zbkMTbibMOCl/uyJJfyVseuykxsprgDVGy/vB5uif
Ka3K3nNaxULrFPdf2ZJBbtUKwbp0/1deuIJTSMUmo4acT2xaLQnerqFUEPFgB8qxigeW9F14f4aC
JbrUhxkbpGaYieSdmC3/EXN6UdZmiVL5aTLFsLiA2GO+qGtwHh8GFkCHCMM/Yb+U/p0gZAeeod2M
lF1BVfstQ4ad7uWDa5MDFKQgkELZwsjv0zE0WV4k6oN2iINpYnHE4glCOAMZeplspXd3Q2Ehnjq1
abtbrJZKdkH/f93bTfscCDRqfoVP64DNx7LYrXvJ6+71CvFEDopui0i1Ga9ZY8BZAvvD6yumMh+t
EqTo0UkSi6+KstayTmWkULetHV1jdUIdDnNOVV/jVefwa4b01f5R6dnpHh4U52tsXyjSqf/b7uUV
usY8CH7P2lqei0QSHTX0dt8r0BUY4anqHCJq2vEa+57TWWNNooEBs3xmqRBa9uUbDbt6Gr+sbQEW
J57xWgNWChqrX/rg0aiGuIzBcGoiQILN2/KL5RWfQX3W1HCA14GkCrv3ui0Fwl7hMIm+Wu091s15
CDutPDUmkqoRSdfA4uNu59ys5Fp3staX5iNASF/qWHGjx/U70wQ4PImyeXRbwbEeO8FxxJWYxdPX
8bKVBB85ugsFuhb0Ah/c4Dek/qiQ9e58ZbXBMb+0k4l05HkXowVda08m4rjrsk+YR/0aaV6qnb2U
peLXGHY8viMPEF0U9ETwR8VOklAiUb4gldYloc96ST2EbwFpJAVOFO6ZkmNIcAahqCK0AsNveamo
j1NOtor+dTOt9LqkllkpEv/VGOiKWDjrQCY147SvpN312aScetXJvf4E5xhmpO8RZ0/tNgy7gjqQ
+AoJrBktvgawHU1eQLztEwBFDEUW30ybno+oQ58T7MaefzoN6+xiPSlUaORIGt2nFLNnnIXTfdM8
wzSC4XJbrOWW339YVav1TjXjlpTGO6BSiLxna1eGpaOK2aNQCXZWwjrz2Mjq7EMjSTL1hpVLGhmD
dqXFp8DoQCjXgTpOkMxR51ykeqedVU552h4BALWxCJH7yZogsOVYGGe6/y8d7Z2DWAvm0oMXdoIO
AUQgJhMIfYmmpfmUNrG+M120HreaNmKhI77QRqmesciaxApc2Il9n9/NNAbWLm/pMek1LRND8/Qi
1WzVFigE/dhQigPHw3x56KAjIap0CfkwDe4Fph+ANQLGfIj5izbK2UxLKpNKlNoLk8abDJfr/bxQ
lmnpITquxoHhXAIkAVbCgNP8wjaj9jWEtVbi8XiCexudz7UGD9duYEjC62kKQkenuMRPypmVGirT
Iad0NNv8qCBStnM3wElNIq/z8UWgX/lcO82vrl2LpVlMBpWIM8iMKkdu6jNtwJh24iPbTRo+PTx1
2tps74JuhPI2SYYWPP8O81RYmwwDVRm1i4d4dj5IG3JW1VZN72Ef0qWenUMwOBAB0Hh3elBXITBW
ustnqTyknkEPseuTLDTPtTV0JwY88ivqm1jX3wcG0YiNt8nRT26uSVMsgIQkDoHZ3ghk3xtkVkSI
QPlY9D6iQemmbZsGx+Q8GwcOEbTGlJ/EnhXj7sN/zkGfg2FZ8lwbxrs/4a4iN4ovsa/ySp39ENuz
8m9YYDWrcOsnn8lrHdOJHIHL90STaY5miwnQ5lxZxMiDjxfZRfJ3wkny2kcbXVfD4+mefWOi5lDw
5Di8Z/sYOcn1iqufxGpiFR3/9kPY17f4dz0Gap0VQVZ1zRtUXA1qMcOuvkS7T13E/+TnjBUiwQ/g
iHjZ+1K+nV9WsGCWqlVewe18lIsUrYgb2ineIWmh6gNliot2Jq0oix/AIHq2Bj+WImbDjTUBFhrr
v9FJviPUEKMkKeV+Xi+J+ixdJTHwTM28hpnp3FLGZmg1Hl6598VyMYCsgu2aQkLt2XNA5hMQ7kyO
mKGtPo8fS98lXVJhhRlZ3uDdVvOCK7t1WZmI2ahqehTYb9LZdftGZ8TOwLOsY5WzSu0+phxSpz3x
nmYGO0ld6pa5gjsLcPRKtrysosaNUX+zCE6b+56BVkpmVqoXIlgaPzluIwc9i4Ns/16YVkGLR3aT
s1BFL05uKVXJrpY/WozFIDqZ1G5Z2GcPbcAlVOsUhQjkOsXPq9BsFvxDXf5oz/sEjU23RF7jRGBD
Fx3h9avCanR2PTruQYlpNbEC14EtPzSx2+n8ImxWANVsgcmBZLK8GApI9zKjTx+dv8LJ2mgmTjG/
zSaR4pYSQjIlGqcQptmhUTURQT7XQzEGsRfkLmELKoe4KGnvMtc+9KVBGxMLJBL2B18is8jPJgG1
a4EdN/ANmIuyxvfVTeZDSD5reqNOFx5yKrnqwq2ttKpUGmAppkj1xABmTQz/DgM7obEljASrMfK3
Mtj12HvqDfvv/15u2DE11gto6vh75eB6OWFt9CpWcwv8yamvvNEfs4U+rOHFiUvEGHLSxnBDVNAS
GE4FfoK8zV9uf3DdqlSvIT0c1QK24320DCJx6C/atfKU75ek/WZ6VUIT5kxnbyj6Hq7YPRba6iOy
q4xFRUYlbKBXs8ev9ehe6bSkuu3eyD9B5CGy+35U3vQqY3IBg/RejgawAc5msZXo+Cmiu8f7HP1O
h28NTPV+PpbtHJg2iTmLSux+BmOVz4mKHdbyy0AEEDQLmrAKvL/xzlVO+to8KV0188ZAcqw118BA
d8w8DUjBcyMkJOM6N0yOxg9Us2olaR23V4Tg/Z9lokWGYQWZgXhs0M/N5AD/G6UbCL3GDdWc0tRz
ODWFygniZk2h+adZtD41Zqvz0T7lpveGKJ/YvKSNalAx647a2W7LHgQ+MatYhVlFM7hf3nyz+Je2
skCflYRNQ+2qYmMgUCMKhzED0YZKA/ofR84oL1fgu7pDxpbO7RvBlTaruZ1TUPGmsU+zLR5+9hFT
V/3uqufelW7/ZAPH//YGrzerFAyPJMuodEikM2Gm6Jt00SBB9YUxRnXkvRQoN/xh4G20+nkU468U
Tz/ijBFLPJjvdsXKnTI4+HxFGQ1Bu53c1UDXDw6IMiXS7VgX1zHyWu+uyVe5UyJoYFhtGCbPeOb2
u1CloqI8i4pkF7gnAsNMWc39U10Tv0VT+aENoZCTMwo6PwP6d9EkJbxwLO5cm/Y8pYbub7Kpere3
2t1vl/FQxB3jgF4C/DttsLjwgJOIqOsSOuS4wy5HKIxaM4Cf9QZJcmeEJ3A653Q5Tol3YvFhu4fK
kXlTsbCcal5t4rn+dvri+DHmPcdTTKXRwEZwvgkPFgEoG6JQcVjCJIkDiDUXoCbJsJN9/4RiAh8i
pnyiRls9Ww/ftd6T4nLv1W0APn/+BpZPKY0jQrfnmfHUO/qMjyx9+UyAqwdPqPKJd0fIjFJz078n
ohSVuARQAs0MxQO4EhWL0VAZ5gJJ5zqLIINj5N3ue0xZXr12cn5zFhe4mhJwQVCvwdGNIH2VGEV8
qRk4XpPee4YKhOUGliKkvfPJcgfu+g07d1cKEXLe1rP8ynAQB1Eo4zpSeoYHcJQHkwTyPu9LVq++
qmK0JdaUN7XNRynGFPgq2OUshDwZG1ZdcafKxQAu13nxsxp3UpPaC6G7PBjUU06fxYcWCbYpzPXO
o87DkaFpl4riy/dl9Mc4iCYWpLHO2QAljivSNiiX5k/wtEDymxSPkBJHKRJJwtlBWm2xHUFu5dq2
oQ8IsX9ScAzHBUoxWbgNg8gopJ5jGiu8uxPzsc/6v44i/b9sfUHckVnFqNLga0b1ifB5UcbNtQgG
XYf6QvVvpE4iaQJ0YA/3bhJk7fieDx9zpGiMkW7x5qeFW37MVdZBAJfGVvodd05wbgxnpy/BT+Qz
ilxqvMfOaI31xywrv49P71Y61D6NeK+XCmr/cauM/3bjq1526RapU59/xnymkG6ZM7ZOWpDHaOW0
OmdYNyCyxPWuAvZpSrXnc+wrS+4K9PNxT4rdWmMePy4NiNM8pmlQ2e5lEFhB69pRsr7WE6kwxahW
MOphOhvrrSnuOmIRVp0gQzbWB3Pg9WEbpJ8P2dIfmu+M36A43rsaD/IcDUuAE235F78oMyZg+/Ej
MlopcW1PQKrrsKF9Oz0klx0n9mTR1v9hcAv+Ks6r/x2j97naHxjvEY8R5TA0s2ZYC6gnBsTmr+FU
i/LLZz454bBmuiZNAghq4n+VnT0/yqV8ZPVZrS8QLQy52SpVbfyp5pVVxk+cfyvhOrG052nS8hUq
l5C+E6vgQT+6JEHis/803Bn8XnqE8cti3NBoOP5P1Hy1/J2ON5wogdnfsHY1ajhxwLToer5th7Ic
F946hmmUGaUio8cq79zkpmoXetnP0Rb/vkHVdqvr3QriUdCqYioiu645BPwTb9i7CbbkA54Ai3iW
XNCuJZ9oiBzEU1xh/76R27ZbF5dHzsaRk15blVkdjnDy1ahYwsAno6dFRY6EEljIM46XvbCZi3CP
3V5MxnXw1QrvoRytrO2GvMFJJedHeJv6KpiutN3EjjJiPdnoGrpZs5whfZqSc61KdzyKQznKZQTF
Cnnpfb9TZynAUYQsT8pZXyugO/GZQxFWtKyr0vi6nuFbrD17W4I+CkuvbXgoJ29wtyWUv6A4bAJ7
xp4h9WCj/wqDksch4yFzegPKXRk90prksYqtZi7RAzw03tRp6itf2Vpxd6/a4vl4aVMuzDHWEiKL
xxPO58ZOy24RcW0SVBO/d+qckiMaqek7BYdfkxHLLlSllDdg0TBXyXQKQ7MIEM3vS+gOcz7cZ1zf
J6092QS2LpM4w5q0IXEKDhXu+Zw/fywxrUjNF2brbRW8LoJjx5Lc3gdM29QVr6XOcVIu/rzXfDyD
zh177v74NMhm56TjtUtdGCB20BSsg6JOmtUv2xYMtOOrVwEtWzbKYyXsdpWZ2Q5qOgENHODEVhWZ
MQR3au2x6IfaRar+DajfCZBvCPQmJxDTZGxdv0Kcp/qWv4ctkV+NGdcKoBPzSWcBjlxdd7bKGsrI
fc++P9eGzIpTlme/hJD8KI/Esqz/J57lZ9swyBOQAA1COeEd2V1Kg+Y3UdhTiFclo4i/XRoPgckE
lC4dOrXBwVDqpGsly0HtgWPPy7zfQ69c3OnNvzaFGhH+j/GIP7cif8mtpd4nONSWS6ezDyI/Q0fP
dLv5fIoIypFUaXc5Mcq/s6U6F6n4dA+mZaNTWg3vk0A5kyZK0VS63Zn0RS59GGf9JrGIfA6Nn+v/
XEGl9WkEgkR6uPE1pJQNPNrjGWy0F4bBwNJOKdD+fkpKqDZCXwup0aFnjIx935nNDxeDOegK9hjx
sCpdeAC7MfwEkAUKEwLa/OWSm/dDZ8/b1jD3xJdey5C4Jw5djcKhSPqZ//qs887gDc5dsCV+utJl
V+iFvhBo6aV89vOeeut0x+5IJ6vc+4Rn8bORSwQ2CxdEr/Qbkow1Yx4aEFt62/k06paFjQYh67R+
4rN0FqAWRlFY7C1VNrYK1NPzCDzk3YErQeMG5XiLpM0b3tw3HasYh+rNIn597rQNsV3taGvU5LbG
vCnoNuDb7+S/ZQ6vJqib6FifRgIHkeP4ojz7uZLzRq/0uhYgOy1e4LBG4gPoWFBwq91eTfFGCUL0
35rryVFIAm2nvRIKs3wSNaB4gzivCHNEOZGhk1jIHocpdhAejbqQplgb/6FK1GrgAAN/BonMuNXf
sTsdqkPu1zwcxsmAAwfc8Z4VkjMcRxnG6QEyilcbAan51RY+tFkdR1EOqWLy+s1WreEJPoPYwVTu
dBT73vePo/o8QT7r6YG+nh1ZEjOxOSOwA9JulM2DvckblSyjlT5RorgpPf+8owrjRII0ttSZhm8C
CLR2UbOySqG7yqBM7EYEXWV+90UTQTqK2+vcA8bKq+y9AN31bczX3UJM3XoISjpCjK6Yhm1bpN3/
NenUyLrsmqj054ck+LzjaEI9+5yQPkTob6j5C2ZNEYsXcIomDyAYhlFDfj7ldNhTfF2PUwMSgQ/v
3Worq0eWe4/8XN33gmJfpLzKneZ1XMp9L1YzwYQ0hOwnIx9uZ6wPPmnfa4ZwfshlSegN+j00z6ir
jQWd6Ho7QcJ3rpKKkFvszdkcDWrbyis54R2KN/wqI4WEqLBPuIFf3dHlZ6/40YQFFlzqGXNIwMcq
bMw+3zmQov929Re6QOH2WwQAKQ/r3Hg9FVFLlF0LO7o6QxLTcXAjq3q/nWv5SE3yKVmuHYbv/vX1
FIuNH+jc0VJ+fP5Y9AKIGF9h/6Yoon9uRTFKd4dhFmLxoQbmbKApCX5k7J4jbNOZ46/2hV+nEHIV
Eikd4v3kGNTCW5QgB+epACIEHo/qY5MXp2PDjYwG80LX/7ZC3/SeX62jIAfGIQE4jBeNV0DlHTaK
lVXhyWPv+mnPAWoMUdz2pcef6AOW2t/1wBLOqBnh8d/KyYQHbqrkcbyYkl6hjMVKoJTeNUjV6M5r
/So8R7QAPPU2HXyv6+h/XZJE5Kqwq0wd6TRijtIapvz8E49H7r4o3CF86FRFjO5HBGMhWHa05qjV
NUqxKHrKbpQG0n9nIk8RqQ8MoORmqce5nwINXfi4jCyXwW5CNufu4pAhN1XNxulCD1+5x3NELYJf
FXZ8kLVFxzgatJ9iXQLqawXGeQ4FA21P6zXU12J8PYLC9t6Jitwc0So5LEe+PD+ab9weNuUNNNBL
JAp0xNCFTVBA6j9YbtE4EavXg3mWb2ssou3YRoEg9fbcAFuTvW4z5Ywpfnx6FW7NsiU++rO5rO3V
JCWFEAf4O667+BL5EYvqbW+l9j6YgKQHmCtSWnRVMf7c3f9GoBh2ZvJrulY8VfMvLLvY6wPiQ58x
CY33Gm2o6pZ6qitRpzx5aX7rH/T90A3HjfgPt58yx4labSPhUVcRjVFshzH/v55NonIOoh77xqg7
zcHuHQm5jeiZJ8ChwP10EVYwuXijSdeOOAVyf7jcg0IIakRvT6FpxigbOWI6RNo3kfvPSCwIiOKh
LZ0M5uym8bfT0yKZmMqHudcQRH1PY87nMmHqhiaV5bUfc9dPrVUYU71FuX8lIqUaISclAYUmDmku
qwq6urXZj4qQbvUPgjquKRNscavzo0PnBqUikBU4QBi2ogXwtseht+rzunkX+WCpCBVOmBEp5Spj
ndfNe7/1hucC2WgzdKM+BPNv1KN432j4pvpBRk1HwIraAGwpKwzbzvOuXGptrL1KIYJDK3M+sLuw
YaqHlpgzezifoFt1j9kg91IgNc/9Nzyu5JZyIBi5F0ZDH16/5GkRk+EOKCKeVWo33iXsEd/59qmh
2QrNZFl8wTXxkVCEk7DyeJX4hyqcksTY6Pj6Z4HZCYTKKbKpkM1nAZhEUUPVtI88aI3gqG+gqjik
H/XIg0jWvrE7LRI37YqDA2e75M3FTi1tfT8GvUO1/K3zgqglxwWRPA4UZu4xqXKZxssMEdjrhYog
uGByt2rjK5+fs4ZMW9q1cU+NtSfQoum2gbB9RdLZW1LrlHtgUOftIVBuDSFbJbfFrS91/2LApAUE
RyEIwqXC6vae2HvFhJErl5F1Odlgt59GUCiBwEXt/b+9uA+EBrYBGtRqlTh3/dyAICYgf36qhtd4
evclhz2Z2Dor4bBXAfzrbyDDiJYmEPWyrvnUQNHm8ZjLzALEmaf6lVjNl8vCuOrUXZZP7nfYRliG
KuGT/ZjiHqGCtsGvNb9gV9UVdbCjqvLpBW7drO8Wjoj3beGvFa4Kq0fBG+b25Uf9CC45Yfmt8G7J
i7hGRpyKQvFDWOZtIAmNhOu30yiU1HCRhzNUKMLLtk2NjTEfzyjyIRWmv0k6TxQs/ZATdBh1WqnD
vd6pQwecVgBj3AMFiD0Dg4irPE11mECHiazfk6+gKJGD8kJ4NuMAGwIBray0JhGxh1shiR2q5Nx5
RBSUAETUXy7a29Y2aWzoOeV2MUWQsJKSDObA77yRC6YFtZkjaN/JmAtGuIg3/kWZj+fquWLlhUmx
6oKLBJDrj57e6tcMMOyQbJBIjgb864tMboRGIx74PjcgWFRZBFk+1weARI5EY9exkUDzacxJ1Jn1
77Atgu2wp/Mh80GSbitFpkPZNvw9Zuli1DNnGiW6tDsAaSLWseJj7vEtvkSYwrY3EIIclluvqBsk
6Y81XTNgXLNp1CoFE9mpX7jvUu1zJErh7zPwwSdwFnhLCKQ+5sq8+LT6eTMK3BNuiHiywKWSsE2Q
qJUU7AJM3l5yadpSEh4y0Psj9kC7/lIk2t9enTjq9MB9zjFQwCdz74Qo5teQWlAQ6F8nwhuYNkjZ
/gXh9NgpvQ3CiqBophJVVQ5tnc41edch5UngNjahnSe3vhRbG+oqANjkQKQ9hCZdTXGTtUY6L4IV
ctiHNPGHhFN3p1owJRp4fZTrWFWNmu5aWF2VkqbGVi+3PRDRF/W9RiQGHZK7hRaO60Kawd3DeUS1
VYy42pdYFrUnCeySJK/F4Ckk/91YszH6q7cUALUw4H1X+mgtr0b1Q1sCH70Y8QoMLzTDSUpZf//0
ovJHU6CUcRsik44/g+pjGiPxcomBRhzlguG3UdXHNM/FAyeHbalaBbDA5MGAIMAvd1lRTZZ2ase+
8BB8XVpwOEbofeAf3rc7i/MhMao7UIPqCJduH2W/LDCllJg57kpHUdoNNkHo23Ik3vMXDNpVbhv4
DLBhiFRCv9lMw3sEoeOh9qBGrpV253hOksZwXVEwUHLUISygSBTDaJXLmxthibRWwecG4mqqQh7C
DnjVlAdrgym1CVTkdL2KJZDpwUuljB3QOODNyxbZ1hyUCfqoEibSgab9dcc3ejS17rC5k2xnbsfC
XbA147lL3EjVSG178aWBxy86iiufVEzVh8COsHujWEbg8YFjsKUTfSJ36AdO3+amGYGm03GhakbC
rzSQfii0jQ3+vUAKUVIlZ8Q89u6n5AVa9m5Vl2/jgNLUPVohMhYZ52tJHNOyq6Aep/3oFz9jHl6U
ODa3IRdg1LjTx8+M81Tx+Ng2XzEesOt9+fzH4Wdsvd3Udhz0QAq9CCiHtF82w8PmKUgRN0wMs359
IL3JzH8MPYxgdF8XNnHwAmyFlrAazh29HspnnOlOt/XHBNPZajv/ABJM4Rp/7U0QUetzSZV3WxXi
40XFaxT+JRvFFA9oeE5sBMik3dl7Cnrw1/FqeMCjvKLdKEcxrFqUURttgMJDHUG882W2npjY9X+z
/4Qoty/Tgxv8tOmrT1qU8D6osmyHLFgvjBlIRTAIu9TB5+g5mKE6zhZxnJAqh1LbfejchCfGKPCn
gJh3yBuvLT8kqZT6+hjg29zwJRQEzyAEzXfUv1ddIbSWmpsNVYMYcVgCm6mere/RMeR+iJm3JNMf
C03J0xGx1GU37O5VpH9LxjZP3GATgoGAXbxtsILMEiXyf09IaSb4zKkAznQ0437rzy218/zuFkR7
xDhByNCFRiDk81p1o1yrgKMRWlJ53vN/Z5UypXlmrgmgcGS3Cy9H++rHHM3g/Dkdd+WPSZuFeJtb
gCZqR0AFKTi0F6E+wjD3Da3oEiZd30dszrDCvuWx9CiS0mzEepQ8Iejs33dcOYFqs7UGVUGIYrGk
9ZVhkWqMZt63Ntf5hs8UGG7ALT9cyRMw4cpg9UDfGw8zgc9QDz+anrOf7DHnY1behkmPRfylD4ux
DVC4EERRVf0gCr3qbewhDRv3WLkPHpAVz4B3d2OBAR0gEg5uZFHy+wEE41OBi6CLj6gvsck6QWoB
+WAUjBwoc4YG4XGgsd0cbIX1pG5NwDqWRElVDCeqYw09hwVA95OwaUtak+XlJoX+paQ75luVM/hs
VenyhKwS/zdlWFWNStPrqVqF9uwyum1Ddkabc5OGMBl7ojd4NMNAg0wzKEwF/lwx5dgUPR5xIaGf
GtCnTX5BEa6ELZIXcHzE+lEZS84Jp0OQrZa8WXaxtsI85QcqFJJeQfHOpITLUL4W9WOiQg0Vme8G
DZif74x7HNZu+O/buHtxkrJfbzJDiNpCI/bPcrciuMMgdDDbjK2PTk83PK/5kNm0QlPlUJERsRNP
VR4/VSzKmlbrkeiLXdM2VkCIAvKCwzppbyuCgNr9GEPLwVlIbeFjKP137HAGXqmidarUQRJg1HM3
C8F1gxUdztmSPbcEeR0BH217HkNlHkJhkHB5b68etp0c/prW5f21IEsNIbiRwmq0A12MbpXOIFv6
IduIMj4YAX/JVc/LQmsIm8AP/hcQikZN/NUwUy9D4GZChBRwREZI56qsxNfXRUKineSvAryEEMXh
AxG7wVLbIV+auDWIFP/Vh9KmLzKUDpoSDkjfj7U5dlO6GEdycghFr5q78w39+9W3RsVMrSBT3E+O
BR0uCj5nIWNxThwJjx6KFia5/IyZ+q3Dm23qjRHiEVrFYWoRfD8k5xngjPSUVXlRgBUswwOp8CqR
0IqOs+Y9a7nFEHAVKRLUv6T1f4rGcxIBb7JB8OVNZZ1t4PBJkjXucUwdFNlHroPlAKWzQus0KmIC
qk7f3CBmfp2nrPtayNKzuTfCOswp/CATt6tPt4kFCFRcaF6omJS7naw1t5oDCGuvrEGpVXZJ2Ud5
ARIxJ3nzJP8gO40VT7TBPlTGslx+2fo6+be63sm5GlyNdLcAZ3msJZZK80YwSbEQ4cVPtEcWqtzR
p7S+BNixdu0NVtC6L73qnhGOnvfMrSem7e99u08arh0R7qHAaEirXxIOtCzBZcKUhKknwoxGYQRh
onR6YKSyf15RrsA/5OsavCQINlxQvEglkBcqcCOhMuBe1hWgfxNSJsKfY5GYnlLfqCiUOaK6KjE9
eQWiR3oJzdBPLb7dEGu308HGuxqr1bnRoe3HAOU/VEO8hDJFMwG12q3F1akD2khHYa5QyhXX2gch
Hw847Bk9C8Up7nr6BZEzMoT/xIE0ykwPQq4jxMV645FI7MISwntAw00haT9oCUwIhqQAiJpuvDjc
UvYsftRsaY2Wl4bDguamQwjbn9FrIiDtOhLeEpzJp4KLHWeh0WyDy09I+CSCsWbmMnVQm+jUYmbF
UBkt+Ph/mRLtPF3786sFc0H81Ny4G/3KVkcGYL05mhshFSA4Zo90Py5XClP+LwnOdHjK4nyFkkYr
3i7kWr+2wJLNZB2ePvvSAJiIoRXuSSBHr9igLtqwS7GDb7ylxxSYISdEcomfPKyhpDb3k90O+YBy
MiRTwnWeaFTLsUVEzcDhCiQnLm5oLmKE/f4/340kRRZlzYVIKF33izukUJEqWSEXWmFKm+3n6T0b
WkC77PtBOKdUxWW8IPQnVsP1zFM3LBa6REOPoxYqnkP6/YLNBILU/Y/riHY2WhjMHgsv3rtNFVBu
3S4vDeChBhPpB0NJ5NfzHphrZc09pPD9ihMzBOTyip8nfVWa7m6KmnCS29kr9RE7nQnn5D3A2PR5
B+ZdOZRF+rkgXvbYTsCbJN/RNnAaBvJ1lryrlUdO+dckxNG0mTT0g1LKSzDEt7UqyVPrP19GbWJj
pCC+4yS4RZYZHT4qJNjaqQBQqRR6aX7P8gK8pI7Nk4MHH+gyHAsEkqN5MQej95gJd4X7KsahXHh3
K3B7LnZJiiOMtZ3G2yzIZdym42eYio8/uC704Z6nrrKXm/Ji2XLOx7L8fWBRwwT6v+UekQ3PrHBN
IavB6rhJWPuDNMkSPVTFbWnA9kdwayp5S/wPpZnFJQ+viixJcgpFvS0yI4GVwWcz4O6A+N7lddgm
2Lb56DSA27JyPZ0zRdQmuy/uh0qyLBdKBU1qbauy47H34qHC2VlooeK6ilg4P1hB8yf9OLzYFs1f
swxDYZbN+rlT+XENEHLMl7BEjnm5veG2n8xYrwY9lmMaEFjpF5jaqT7p3cn+y1bfOoIy0OfI66Ir
oZ+mSltW16IK/LBndWvp6xSZfyVXHxIK0eo5Bi+EqoPsUzJnyDn8VC99nm7c7LKK/rM5gX1BA5vG
GQN9ugCRqkRlXuclGnhC/vXBC0YvdwIgPJEeOa5XVarhi3BBFEMcOzgUPRIUjVBSqJXkWwwwrCil
KFw5VzIFYaQRx14AWzKI+5GIr9c3yg/cHh+7VwNxtugOde0LKgj7oz/hN/VzS24ejxKc0XH/fC4Q
Pwmo6Zk4SVOuKAIjMyWg7k/SUStW3jKHiNq0hIWYaEnP8AoFiOcqZP9tk09/Dbcfy8aRmQEDJg7b
AvMSXpUa5SH0Fp6OsgDTLCHoqLDPWKHE13nGAzJVHD/h9z/0axqBESvx1HxQTn0XFbD1+AHIrSkB
mkfu+sJ0VvAocX2yMqpIrKYJqRGy8ZP7T1Uva+JfPCBdknAm2I1XtN9MemRVX/ZRCWEsv+eMOkY4
2iM/VK2RgECU+2tNbl08okLBgJQx9x5lAK5eCqbUHTCtjqnt+mvT3V1J40ql5AA1MV6I7AX1pIY4
do603DM7le9iCGOLleEw/mWTEDpvJ1MV5sDgThFf7UlpOZwr0MhOZshn9SONY7tvp1gQVe9RebDH
BtFWDgr7Ge8Owclp0Lvty0GmmZYOi0TGkEkCEejVJcLHsvwa16ny7cD79Zniho5dpZZxAgnm/j2U
lOyZTXScVq9ShzQ6t/KtKbt+noo6RpxP0WSGywToPEik25jgqOTQUvEoZ6+BdvREFsFeBWe1xDx6
mk8QzD6I2EDtnfLR1DcS0Db6muZMG6UoyuuWYZ/7cH1JxgblVCUv7znOq4uzTq6AEF9ChjANFU0x
A088CfXjXHwr412GE39nEolXoez5LthSKgsxVydPjtMurRVM84hFfBKq/BIAhWRjgIOOMNPOkIvZ
azzIfI4vCWMiYugiTwiXka1meDLVTdc2CC1IoGYw8cFzK/JfybG4Ax2ugLCIGTD1gF3O9mFqdfSR
DHTulhpDi8LdXfPCZ+b3b70OIA65X0GgOhEKzclvChLS0uzpYRDaZVYAz7FYVU3zgN1KlKMEknU3
0zdf0QcraXpDOk7vwzn0q2YzExxrkUt9QQNOit7bwM/Olo/7zxXj0mT0T1cgE6f00laP9HM9v/HM
Ew954JR9KPnNYRZP84/Tk136IbaICtmca4HHXPYlHbph/xRJiaHZCuiLGowgIPaPm6AChWg4DExV
cZOdy5YxcodQqSTizSmZqW13Z2s8WpIY6x2SqYlP2t1nyv34YGamH2L8g0pdijEa7aMeUjsXeTAn
uyulijxTYAmXIdJhPC5Hd1AvLiSCeyR3RpbKv9zXRJJi3M3866N2YvsVlFi9HdfyJrku4foJx0kx
HsgLJUg6TCaBzh7lcI0ZJjaDQhwSLGeoa7hcTas3BIy0D5+d1ZlpkcUjSyqJfzx374ONA5fvHf8l
7LCzVxLgfRVBwNUCkDj7uqYZsc6o1qox6iNoGISVW6YpjK2m1Y1EeKGeYhRitpBkY3Yok4d54/Dx
G4Qlmuqtm5OJjmKjDnsjwoK59pFDh3KpZyQlNKCuHhyM5vwdPBtrhbir2EhItuhYSpC13OUnrBZ2
NA7CVVWCheQQnVquRvRxhZLekVhHVmppJPHGZm6mLkVnEfwnqvchVQUh4fkItcdEKAe5e6orhnjI
2iJfSlu+aUq14G+zIjeVB7Vfk15b3VsrfZHtMuCO7AY7xs2STbOAeJ2/fYvXLNMAQqzse8HRejmP
9sRVHDEH+jYIUl0D0ufbdTpNrsfeIngm5kt7QxxbXIlsHqzfj0aNonIUFt1efXvp5VFJ/pXDiTBO
cHQ5abdNCsJ1VaWYXdNA9goaydCxq5wX1XJtr2bQbh5DmE+WnL87/6uxurJD/NhDCXzaOCKwbb/L
Fsrl6UMIQ4Fu+SSaEuX343IJLAOX747PRKhFQXBk4aQV5AVdmgRGH/zaaFmZWMqW71hMDDvsmxvO
wVGeKXYsJYVW6cYDMqmlKuuJ6LKbHkZyDyRfu0vClkECSrs8lG8ySsp5ttRDcgGUMGK+g0QkronF
5OyDoAlUGVq5HrzCXE8gNSOerycgICsL8pcjiInr9IdOH1np4qJZeKwAlOqXu9RmE3SrYvUoAWly
i/BcimwfXyQbfh8Pgr6m/7IwaChGdW8l6ZxfKnMuGqgb6LELxLNtAJY14A6tzNh5dN01kG8V30lN
O5mwKaTCyAPpDJ+/z6QERqTavUe5dPwue5KHtlcUZR919vXV1DtfijDlKOZQU6dZY/3Mi69C+ooK
ZdjiTgmRgaxY2MUsj16VnCP0Yrq4LbRrRYLrla4mSdA0NoLIinwSVTpywX+XheUbXH1ai/xboIpY
YW3Pgyhz9WcEd2eIIPFNxPI6Exp2+Uu5QwsZse6Q8nyk6EALxf5jVN5dRBSswg57KY2EqgbaJ5iO
uKGTBmYiHR6EfyF4/ME6S+rK/+EirnmmnoB6g6JuscKfGaD+sc6wuyzgcGWpCW41b1fsUDqjLL9i
URUlbh0U8TcORdd/IcQWSSrJRRQnJqk+TgGgL1KBXOQRn61zcQ4ABXzVkYub3o8+5uWk8tX0sByv
HGO4dzmvTsUcuwaRsjl8RXdYtnqmVUnIKsSKR4XVYrZ/Lbo6K2o9/UDjCKi8PoYvDeEm3qprD6qh
V2jOAkbphjuEnp4c7o/bbues2IkBYII+fF81q3cRR+a4BxjD9nTaeV9ksaXBeFrwuTFmJeyd15qK
xSGz/xixuVlx8i0bXp0Uj065pJdDVDD13dHt8WThStZ5s1cqB87I+A09oB7RD5zFs0zRxJk1ZON0
/+SpksWo/t8scVjRUkhf9EaUBOO11lTAvD/DgsEDeHVG0gkHkUXdaEKmb5A9agp6P2r3bEy5IzKG
fXnzsS2VSKiG1a5p4J1C4GNJQDadJXtyPkhS/yBiUbLltIPpdepJaEKDMRD7WYw7E5YudCLySXyJ
kafPEn7UT2zGevBR2QR2wNYvjuc57TcL0Z5a8N7ZfOqeoLRkEkZyLhvoUXKhwakubx3ytMdMLTnK
JW4F82Q6NpJxMTuuBQc7FdR+ncR/5yhDUjxeCuGGx6Sqg5hDHQiwkSF1yfj6gaAX0GNSZ00B7fHV
mT+dW/6F/tdxk243VY/6VnDT7XR6HFBNZcWPOdQ3ycFXGxN0EZXHCxWXYY6Q+fv5LPBVMFe08XF7
7asQn73pes1AUSxwUMY9qV0seEi1BmXYKSoJhPhZvrKwHNBCE4oCmM8PnBuy7/nTBk0mLTx1bvyv
aDOWiH1NcHgzaXSb8ZthHEOXwq5ywfo1J+3TFlwPrd6Bxdi/3D6k95jOjCshpZhWt2WyeolR62Sy
r3e3HXvae2y2AREMpP9LO9Ud0ImJC27EssY5mG5sTBguWfOwY2dnRtvxYmC/Lan6USPM/nMi08AR
ISLtGYmmOVgKCGGDbnQ9WLf4+RMMPwotXUbGF6b7ig6CZ2r9W77cMTBeImyr+pajVxktv31iigRU
UkUnHh2i4U3zCJT7w8zpGzY2ywG77XqQOB+K2JHjj22x3uhT/p2EcX4D+aOTMKOEC6qxi3U2sGyU
xEw4TlQ2SHs2fx9u3danTSDwHFvM1ftGKvOHhlO1BVwuMBnpTd8VLiDuNu9iAUjrucgmT5Rl2nUS
DzpoRsnGoraKnOJKQ7KZ+f8VBbbr/pQEbVFRegOYhfsekAY6mi6SMXGkIw5T7ojCk0/3AL1951kR
vmEaiJ512fQPb1b34wnt15YCDmBYrTvb3uDpe2I/w3gI2GJUJJ9XVyYUht/nLhSXZXPqfY2QDzwa
NjStky2LKFCXDxtSes8nByCA00Aw4xK8BGUJzt38QUhCF/9LAv6bSs6ib8lhpX3gF2CbEC6oPJfv
9FGKuThgE++L43U9s7TMF5WBODeknKRuUF8GRJTprvLDY0znB3jJEttwJ7ue+4h6lj6oCqNhnc/I
CqxRP7zxNUUHUmDspn+wPOsvD53BthORJ+2HwWGdSUEz8fW7qQvLcZze3an/IUfQUPGkdq5BapVo
M8V6GMoa1X70g0wwFrD0M99Y609UBQ8mDb/1ZRDhTjxQeXMJt3LjgWYbbWM83SgmBj7I8AkY0Aif
Eh0YYcjweeAjRn0s8SB95vpwH4vfkMn1v5L6tZQZwOfhDtCxAEeLz1wFY9abSrgdlxgdPF5jY7ix
DouMwk8Cs7Qt0OF+iHBtfXAWGPTTdVilHGPFpzDSf8vFPEJ/+b46fU5l5bMZwMjHyoeU8G8dlFNE
rghjwCo2MeqZ6wX9wfhd93iqFZMb6mFJvaZoX+nxinoXV+t2988yR06K9PTWLcFgDaFx6y/wqQOt
/QDTc8EWEc9e6mb8j/euNYBmpcW9uU9VnYXEJAPZI0Uj1Hjm7joL8M60kft/rcMQpKMYO5BKFT/w
nZs6JVoRm9Nz06TiX3U4egAh+YTMd+UnYNBzmB056iNpLMAoWgzyts7INC0s+pJ+hl1mEM/KwVac
SLhWsRt1/JzIZnfjN/3vqqyXhB5HEOstq5GVi+GOIx3kgSw+pUnaiqBLRnxmiz1rwkgdurhKih0b
KsE57ujLlaKi8nstzCskd00h6Zx3gvgwId/33NDV9KYfZg8jY/xBRBfNSNkd79jQX1H2ovv8bUjO
gJ6Uwch1dHhim3yMel323gbsYK/OH0EmoqXKNk6FngvjMRV86K8jHsChqqfns6NGli7khMAUd0/U
mTOG8f+0EuspzQvBEkWu4Pnob0wtwSQGVZ+XNkx6GHAXVgW8jshZt3QvpRNG+wP+/x7va1W5tBB1
Au5KzBCxKal+cWe5gcj41JzANEwhUNaBikuYXJUe9IXpUw50BGVdJqO3EM/a7BXjY0yMiP6boJAo
VFFdd5KG3tgIszYQ/zb8xTGVXUolEUFTpBqqL9EhuyaaX9W+oTiHltkBBzWY78DdA4yYv2wCoUco
hX2WL7RndXxdTIcVZTBCui75HLJlc6RSHnNuikEsQbUBDr9MuOB1wsRFj33sT//Rv9ORdFEHJLwW
K0mFIQPKUXS8PJNjUNFpA0gn4Tm638qS5su8Y78w1kz4XSYuB5OOWgFsjkzZTyOLDRyW2Ml9+yHw
LVEvCdwG/RwNBvZ+lCXUIqBiPx628AcqOnxHdAYS+x0JBswUnFHHWH4XTPGNmAFkBTi9WRWqL4Ul
+rrzJiPbZ5A0iA+RY+1oKU2njrJILLbD5CCXiFk1yoTEZ9tLQ8oRDTdJ/knANjEweYRTXESf+oUk
NpTA75uwSazV1X8488jQDh409lWPauoN1ipMzmRdfhdbPNK6gJEG07xedqBJwcma644ImOzqKL2k
fB4fuSYobR48Q7F+LJs00TqPG7FYVvDgGRD3NzPLAABnScROSMVAjU4FBrWeEWgCAiys4WT8WJ0C
VRA5Cc5MY2/Di+Hij95ieeJ0muovsoESEZvhVDQwhFJA6rQnVdXJkJdG65iqgDuCsqiHyhdarKN7
Rtt5QEFLcTy8K6LwXhXNMlvqFt/wsHMHltnMycQ2wJVAXT8K3ehthsfVCO/ra7wMoO733wjbcZA1
vR9/mKfNdDZiUJRbBeAIPa3xSsogpSpQB8saxH7V/LrMJPKUzeu5sKyod7gxYRru5Trh6GM1uy5W
sRuB+0D1cCCYpxwTYCo51uYEoaBEKe0ENexGkVZtt/zAA1DWjRlvLE18jewrG78qFGsQqO5bjGlH
5MYuz7P1zZ0xAS4M9cdKB1XckIBxa4Zfhq2zJrk/63KcXFpYqQxTd8E7mfrluh+bWmiBFQviNH/4
/7LICab3RaehLuXpW/toluQUwi9p4KRThqxw4oUo/ng9XKhkMOZVfbthMl4AAo+5ivhc+APOpXvh
ZxiPXccYzOqUWTKj/DNkZxoDHyZNFj2dRJ6dm+xbEdOF2RIvDrYb/rI4SShOrLhw2/uOEhBQl3We
CBlSw51EuBl1JhMqonR8S14EaxHA/3n5LJ2dmfZH0drARS512a9GAn5KVEYCf40KAUZoefQD31FR
Z9DlU5rxvYUWkvRn7Id/NkltGYoJ0txAJwMu7/L1vh9hhbWr8Hclk7TnkeuXT+qvvK3I2ZrXatl1
S4nJUOXdXLhUpIqDEFEfwf7iiG223rdvoWAgAjp9kKy3dx5Mqm9XrZ4dlyeXpz+ZpnY6rZ3KybOB
Qw+tU5mwwS7B+f8Hc+7Vh5vC5RgEO1gDMyxpdF9L6KG9Q2UCZc6dbqRgei+cdZjW4Odeq1qJ+grB
+GDAIn7TJCLzo7O9OutDMGcjfMlpsP3apbYAF6GTGKhWwp4xNdtHYNPg9dYrRi13xo0dCXz/uGwz
X2evZyum+mmPYa2UT2Fe3xOzkQ6rmEmv1zMlSFb9MNH0yy8iT+Bq73tJpP8fO64zjyr/XQwevfOY
j/JjvgxLBnvvcq5IZCLteATVI5bqF33QRztNt6gEv2PGvTYo7fbGpbaIOfYcxNbVTBgFrriOcbtS
6+wiQRs9istKrvb+H2WHvFN8Pf82mq6+xah1/Qf3W540bIMYXUOYAibnxaeDbXnMXfNcVH0zpdBc
zavz5JlcwQhFGT78ttBlmf+9qPPz+bP4/gGl3bWEZu2JSe4UakoZuzrB+pXt5ZwUPY5u1nAW9//F
oEvtGBdw5rfZV9j/baxPoC0x2ZaXz9D1usHUV7v85qxpXLdUWDFo9l0B2hZx0Jpb5Bo3Y9fyL6sD
28UiGYjinKRX0AHAdeq/zCv8iW1aWuE+j+26cQKILrctIW2bvZKh/zAfyABNgpE6gSyJ/HfKnl0O
XsoQJEOeFgSEdHhe/fyEHV/udHiJRxBZj5oq6U/BC4TN08mZ4mu6nkngQo3qTo+KUfa4/aUpdQYc
th6d4pDFuZDGy2CfleOox5VyFx+49EqTxIxIVq50vQX4Pc2DM1SSkq6wuzPmW+CGPphERHLVNNLa
Hc/2UFrQDbJDOoJ3MQTz8sLKALknr60xr7BN9szU5rIih60rbtY8qmyOUmvQG9W1OHdJ3//oB/UB
2C819tJIVh7Lp2sct+bQq65dumaotjTIBL00hnuLMPsNiS9267mjRem5d0cUhol0fAk6gPCKzKhd
YeprNbO0b21CVhPdDwfYG8cxLQ2YiQNMDz4NRUuVjinm3gIvBQ4+Jzdrbb2YFdamrBumXrlCDdRv
iWkXDHVPQwu5l9mSiUU01mgYNpDRv0zUnpRZ9ZoqHLvSPHu+5TB+eRjgTtGtU+qChERxRVYOXH1W
lpi/A2onEQwMYg4dF+hk71bPtuECGX0B6L/gkmZRTEK2/97Po9+u0RwNx5MkBTVaMOtYW8UAullC
qVmWPC5OldbIEcQihysvuzQwKLDX86rK2rP0f8eKgE/BGNdQkDvOVK40+4gQkuWdaEE/PPLibMwJ
hJBf2v1livCNCmuZ4z3wqV2l2jr7pgsmO5U1wQZZe26mX/fMLFkqqPTsjNFrZP6355ZIxCpUr6Rp
xG/INk012OQ4Kjw0ojfFzplBQ3A4IGFozzkCN+0renB+l5l46HfkljqRapAaeR5vSM2mrIAKETuG
Hmd1/ugC+LJal0nfceBoUFQ91WMZgBocloc7q9mVSL+mFVdouYCssrjSxTncD91cGGJyyljFTL3P
17H+vQy8yK9uXJEhkh+2JKmtRcz0oBE2FaErd9blluPMXsHf/T3IFurLW8rrJMbUoVkH5mo2xz0C
A9iI7Pub16M4kp8gX9eu1oqOIck7OWLh6R8HepdNWQIEu5uzPtLHOuEBdpqlIwJa9PvFN1YnjQ7F
hjecg/59+G7Fh+SYop0zQ+VMUchZkQW9fC5Daj6PhESGCdRS8w8kr8KiSPDCRA9OQFpGG4M4xFuO
qsNeTo/UZpkt0QTp723owaNaGQ7amTNleWqC61s6puidHIXvDqkv04wyg2q8m1YoD3ft7BlZhVT+
dVBO4fNMNZk/hD8FcdDS+VQzyRYYDo9gmf+Dj/NJqNUWfUR4cX5xp78vx+jyDt1IyFiMnXtlkh22
6gLzMG6nmAC2Ls5OCBbdsdBPmr4cJ/gFdWSV7OS8w+86y6I4XN3vqAz93GlvdxZXANGfRIRBJqVe
vsjZFS9PchxkCcqx1fcHuO8oiiHuptMWRj4yZfaoHUNgnRxS7DJmPn/KqN3mPdmMu3X6kRAoOnEx
9x7cKydcA/p4658srZ+waQxJsgerBnmprTlnacu8s1yADqDTKU3wsCNZT8kQXaC9Asrb52ng86iq
ya4jnwnSNFMZsEw3hgc2xrWqpw4pRJ43xoB7tgfmwDhQAdWiI0sVjjD4ltQ4m3KZ7/ttEAngUY+5
elfn0xeZXIFWT6zigx0/ETM12Eq6fvLPP58Uebl1179PtGCuOhRmNxf9VnlsiB5DuWrjeu+TVTdv
KYESL7d61jgUCBfeS2KnetHqn+wGJ5etCvC0VvpT+nWuayEbNvXwV5JLs0ydeRZkcUleHzF292gO
nwgiM5yz27xAh1uj5zpu7AdNIYkuNjPIkrm+jw01rzAp6vpoGrgMufkfUO85SwM+i4Q1hKHps6rl
C4jEvTRH1Ebdk9hxfF+TbEenA+M/0ySFzPRmMUNafPsn4U0O7eiWV/XXGtNkp+QYT4GW0chpIWI8
1JO1JgYw9Xbqg18WhQLeBEE/5nqREgSOxJ6yhcjJ9JX2djABMRWd7c93W1/sLKRuWsilOB+ioaXM
YwxcAeGa33XIg/N7XU9eW1uNEbnPpdMiy8zjDUC671MSOcVaXSv9EYO/0iWTijlxFK0siPUpOnE1
EvZL1z8QzPFeWTYdrDBcs0Myttt7P/gWBWsL+uijMvftJJFRMiKR2OCekUB1j9O9qG+v25+/b4Z8
4/X+NUa1pdv+HlMEu3raU938+DIGFichRZ1Df6JEKyb9o+4Mx+v7TBM5DzDdSZfw5I1bgK74taJs
10+5kgnIU/vceRt3R5Xxb+BBvIOTdQ9YIX2t46j6EcDx3BpQ3K3vlbgGFOG3/KdCt3LlOMi0AJxd
Iorz1E53GDBgN2dsTIYlS/GiqEbbXZqByb15/DFnZBtGqTsYn4ie/xjSDUnnH+wr8XgteRDsGY3B
521d/eY5Mqu9MtiRmr1K92slrhoYcoVX4LdigfjhIpVy4mP5/cnncLLxT46EbEftv+HkTquU5JZl
bDZvK+2Qvf9fpXCadfZ8PeTFk7g1QYviVDnnqtZ1oTJBW3N4MdZIQRce+EMGtRqglLSLJjEVyqhO
5MU94LxnqC8KOnaXQaAp0w2AQ6lBO0XJhozBZWXsmGQGwknbj0YEEFHcXO4v5N3FEC/0T8mQnSOX
nBsKVXUf/cfhFflwNjs0jvjKLVgusId8W86mUuj2k4hxCYJLbibCRj3+WLFUtcwUwpWoL4q+IqBp
VN3Rg781NPJjnvkgAzPqq6ymQiZfUZyGEgxKKAjCE/UBrq+KWl2SI/qeOMoRPJJFZqaIPakTnFxr
o/Lxwm9+iwS2LPEp7XLeriA80SIHHW/42+MAxhp6WaQJvMoiNGfoD5DrKUyewsdrKThfSiyublum
mN9jjPCMRyk0yDK0CiRR4hCOIT3jYuS6iTvxpz/sxuu24MReHag/yTq6Awpjw4agRY5IZupB7gDd
kQ4RarPdyYpJlKVe0G33pxbt7iw/35hmoXSvPsGRYTTInNnkEFXrRF0rPWHgfsAaaqsV2Lfv0Nli
NxAbdz3GdwoHBtcA2W0IZRVZ/qm5jtiV3aGNZxQxg35g+auPIbIfSGE2yUrXh6bVZV3hu+I82P6w
9KH+lDbc8fKGxd57KCkhidtU+6KYmtXrrWvhUHWBBxF71ssAaDnohdb5Zi8YISkH+F1Omww0JFQK
PUfj2PtwwNtzLfg2DiHj8I554nhP/bCoTutY16kDJCvluP0rgeNNut7wNXnnbwHjp+lWa3TmKXln
4dYZ0h9XEVjSLlcHQrIdJ53kDwD6ssVSAbSPTn4/l0s6OPZdvE+dec/WxjNXJuAomkxiqmH5V0Gg
ptN68fcJOpT99qmoQYQmcUGGE2KVz6una6UVIObPcgyFjWMbRrDkVkQdO2EtPaTQyTWGEKJDkXOc
HyDA+95IVWDeFRtbG4Pb8M1XPMMOe7v+HMQNI96gmXtREXlt8TXQ3cimlJmLkRGweOZcoWis9DoI
kUMPrUr/ZHtQFaR3FRQTqh+kj6ySaNkKof/tHj7gXwBFTM/Rkmz4RfrOQmFEAbnHqXPWH6xh3WkA
dKqaIUsiE9XVGjwH8Pvke1TJIgMxpElqzrAkPMoDVD2YqbMptEOEtTA3kXVDHn7C3xcVLW8urT8w
YskEYH5b4qt18WclfL5zxKih0S3nICqjqEI4NBVYe0v/gb4axvSDyebiGMptmZYZPvMKJ7Uei97o
dXsnoXagMOUvFP6YU3hWPyzwRwGifgZoNQYx76AFJ7Xftad31BYykBzCe3UdMLKY4qmgE4ppsSXi
2bO3xQTzFO9pAxlLIKGIE3zl5r2oXXbgvucsKYnr1JgMxrCSBQEvxVlImQNLseQ2Vv08ckYA4ogX
KjjoMOiHdKkKsuUpFPmjl/BhJhZfUYg7amswjg1eHtsGFtxB62skdy2QsoVXxG9+SSlM3WtSjJUy
fdXkbjSfv6a/DFjBIQhISDK1T5HRMPdijpDrs6QKKESvNHS8dy9U9VrvjaEaOrmUN7c/DPGNzP+i
fc8BnX4P5etcxEo9SMDpqaZOXdhPXxgKpD2fUIyYIGxCJUJ3Cpq+X0iVTMmPJHzvbdNpDLKbNNMb
5vVEkVSuwUVhGBUeJhoNkcr3i35tsWLM8S7jpBAmfmbZxKxFrSUbeUKdpODa1ZkDO62zbWwV/UGF
8TXp/hLp49yZU9dDFdn9toFIEZHsTHUI/JmmmskVHiGKTN9LIDkTGQDRcaP2ChkhtiTKmlCbbpnf
TgPmO79eiqT/FHHljTd183D7cOENTe0SZ2jtiCsf2D25BCugnCFuiGvNgc7rHsvnK+FzyBhafihg
thZkXhe4OksAYkhOGqmFLIvYouk9Xk7esK7TLsjy3s6vcuglAoG/FoBn5hBSZy5nXWbSO6emxmyT
QldrtxkNjpFfwKk+bf6nkWqAQi/jkPXJ3MI6QVPXYygcwSuWN4bTRHo763/DBue8qotGRL+7/bUu
AVzp2lE2dj1MiU0vZWXBENCLRnJSJCAZPY1A0r2jE/EwPkjY8xkj8K6R6KFyb0+c0Ttp+Y5D4gJc
iuvoQfciQYFdfjmxq+rMMlt2q1a74oipfvzwRk0BJIaJH2qui6/TB5iX6IhDQOQ6q8Y0Y+w/LAfE
z2fuNg2Dvxbe5ZI3DVFhRSCU9AUt4VDvb6LSZTuyh6C6UKgoi69sqtUGmwe+En97iTw5pHkxqpFJ
tmuQTOnJeUaFRUtwAdp4OEd6Xid6xqvvvJbsDsKKR6Il1J710zO03LjRX9XKwi9xZHAwtgS9gTS1
homE5+ZqlW+yVHUW9MHebiYg8/bh65Si6I08TB26bgaHGhJRO8woi8/iesUK2M6L+VVykc9Ff/p4
e+tOut6/QefObUot+mDKwFAdiU/ipPcA4RM0eltheW5M9SuFtz1NS9QfrTN/mwidF8SpNjNwKBmJ
wMagUpGuTBg30U/8Pru+AclIGPNH6PpvcfnuO+8fmPCdppgxImxWheDedIJKlJ7vAX8aZQeoFPBU
cIvB6DLsG/p69ZATWCEs0l6uqd/bYQBXWIuKuzhkPMLeNWVGXrQH9KcZ0lp5jgTHlx4Wk6Pe5/aG
/Fo7IkAj/BYi5haM7bFGdGJPSrDOE2JPKGeR46l8ubBBAwp20Fqj7V2X1wL9AepdLUM/qKvbBlVA
x60bty0rWhCMpX1r7gTG8k8Gly8qRnhSaXS1p8RGJWi1lsn+4ei0u3oA99taaRPr915uY7003SAw
UUVFMYlBtthQN+aLxwDdzxQwiBmKwNw+P2iTU+0f5e8GjfxyWnQJU4xdKI/gJbiB5rmhLUEnYnwn
OICr0VxAr4U2781+igwGcCcqNKd3u2kTSUtv2Ci1g0gpdi4H/C2g4/8NZgMp22fvZSKW7IqkW0yE
PUOmOqZDj990libBFMDb2d6HYTBHM3WzoSsoILLZBxHxojUWyna+KWjQ6K8b9jDijTHj6XuBdt35
JW8PmkS3iTB69XaApEgFy/xAJ5nuQ2TosEAJTwDRTkW7Cj+4DzxuxdR+IAFlr/QYhLdBTZ/0F+JW
EalZwFR45xQ6YAdZix1AVEXhDTIQfp4E7UMa0dqWLPnr7WQWmtKRJNtVb3yh79Plq+mQo69nkVjn
fPeAmVuCT8P4gVWHefrlG4X+gYMaExqjL2k+ebu61XhudAk4Mq92jqAFdmSOW65v2rLWQZKwlthC
c/vXAr/VJL2GYC3HoDPuP+KCB0hgbzUtSldSZap6ovqQl9hPcDpSoDY6wsrqEhUN/Byes5upXRRG
7TJFX3jeeFPWHMROTZ2Q+Dt9o9VBpZYMW5cer+bFD+tG8iqZhTHY5KhFlcVeNZKm11bD7Mb2S04K
OX2ixvOjk+PNyTwEp6T4Za8sT3sOyiVF5caXSwrEAGKmm62b3BXCW/afteZp03lpB5Kx1GGBJyzX
LYs4QQXqss54nyUlV+gMdStI7v46b/OnRTNnnNbzf7KmEvboSHtrk3FMKJDI49qMXyVsZtXBXXn9
DskTpse+Rh9HhzFADkP8UPzmwEUPAfEkCae7g7Ex4eTA70wwrBqzZQ3CfO4f9l9E1FUII6MIBBjI
9bjCLzSjHQrG+yHrMPkOOMB3xITqQ3X3Sdc+HxVq04I1/YXmsQZT8xs1+pU269TLZNfkRXZpmnp0
wOrZ7SQopZMdANUgCDrGdCkJBuQUp4/DExO6xQMasumX08EgO/Z03ZgbpU0I/uEVkuCQKnaoF8dp
UFAz78/5qt9UfzY5dzBKVC+8nAAcaX1P/g4H3h3s1SRRhv46ml4zxgu7L2W3C08xci3mwCcE8UoT
J5pgty0ctU/ijXTd+0bMauIbbm2Yf98h5AMD6s2oC1QQNTj7sokGlJxX56ulAKpHig8t3XkxtV7I
p7SKG1k48DEZ03cbC2u98CG+XUHIDuz8TekBT6V/Y9KH+vTyZfwIwQzwi8cPw9Pj4HnlEhE2IHud
w+r1x8+iRQwnmeDCCB+vZujAbwLoon/YJriOdSqzJm4YvKhhTLTODOUdsW3iJVtcejeagVgOiWWu
qCn85gD146s8drGmJebvfd2J3zCYvXMmdyQkUfli+UISpmX4zdUXA8QfEtVAMw/ak0EUORpkEOYu
KalFVOhmHZdqko83XLYHhgJiWBT30mycDFF/BWaJ/V7SwzVU87kz2aaIQF+B+K29v7fzzSxTHT6E
ohAiXYQbrxfPfAGGeE/MS5dv+n8EcN5fziPUlw3XD68M9Hmy97/PbFd3wGbeCouwjktFUezrFSre
jGjmn1FWv0ZRr2bv160Q3PW0a8CyqKnQ8+5Noruf97D72l9wkfysG8GQN5OTKFp2YZpgwo6Zd/fG
mL4e/L7t2UhEwckX+4rDysnJIvw0VjfGjZrcYsMSPDftp8RDuIglhAM5sv9JdEVxPEDNtyxD7vVc
H3GO6x35VA8ishkxxAqBCkh1luzYJcRKB0Yu6cmp6AvRDBgs5U5Cry/ZnAP3SKAD46w7hPjH/pIA
C47UTvteThmRxARvBMZEGFoAa5c9bLOKtcR3p7hUqqGRC/2M15R62f3e3ILB+qrN0sbcoSBcOKVp
aijh+69rC5UBhmH7hJpK82dAhTrD0w5IqGAssHw64x2Sb6SS1rYOf+iJimshwfaaoI0FANyfDzlZ
hKdOHVawUu+x8zcei0EvKgo3qNL6/NbVcBD8ZfcYxer1S3nhebKqs/mb/Mm5Rqs4zTkMxSQcMmqK
vxSXCw2x3qe669GsOGzHCSJmizY01oRHHhiax+c2fw0BksIbbTFVLngcFKwF5pQiRCRf9y00IUrY
ZnO+uer/W1Mrc1faphrPLQMo7adaSTeADK8kiVjMgDeAu8dFbCPhALK6bpjs2Shuzz6J7NFbWxCA
EUpds4s1WNAB7r52D8f2dh68pnX8ph6O5WwA5ZBTlKfcPKMTOLJp9/WPSYh9MRk3dYmryyNzVUv7
VcGMyuh+yXqJ60g1sTsoP2VQ5BAHDN+bhhDoq9/Ot5UGlfuG6ziPjsJ7D061USBZyFnFljEFGcNo
N/4iOnBMthTNtcpQo0XsOOHYRfs9YKG9h+EJ2v/dds3JAg+ecZDjOVdsc5Ktumw/IAf+pAmrEf2k
An8ubORngOtgDUh9eHTKAPjRqIOuydLAWwJvh5DR8T8g78Kx4ScVlDTRlCJBvFW0umY0JRN6H1oX
Qs0XoyYywuKdOlZcdJYzfMqpfSAJ4VoQYAciL18SheQqO5+pvI7wT3bQ6B9Or60LeNv4lViBddIe
pzVAIpfWMdf9BVPfhLLGsBcfwlL+E2jTlu61rEq4L3cAUge8sLsNQXAPPbaoX4C8r8Qe08t28iJK
tbt8vwtTtRA/ZLuV6f8BEndCkExy4KLwF4Ty3GKFqikmW1uWIWp19jUaaJimetDPxsBRGM08EOmq
R/BpnjDMFf5L0GyDwneg64t1yPsJmqJNcfDHrX58PXs7Ox5Atr6MSQDBFWb1jG8QL5ZdFTTwq61f
hsIGNxmSSWNZgjJp1ppwAykz9ImvPBwsct4FfyKCJ3vE/QUnKF0CNTYP/SgGZ0xn1oUGcoPd07ay
EJe8HuONrQGxAidra/YjTa/hsEj417oWcLGsnifcRec9pVq0CN3RKWG6mb/Ema840qDAmqdY4OXr
SK1BOZA+ZX0jYVxQM07g9aYiKrSy69lmyEbfoVXHr2ug8qq2En5oI0noiwAgmBe5vXcWENk3E9Fh
cX49By0tf1H5cpWxjBGzY9eMLduKBpsTSbvWIQHPb3vd+sAxLPTM6YXgj5OGeRZ8ZjYwxYXumZJg
LDx/WGCwNm4sWcDi6CndddKHBQlzVPcLPhY96tWY5+b6vutOkIQw81v1kIo7tdqKIBwH5y1aDqkd
brK6iSlmBcdcoYWHdEKguJklhMdFtZ5YUwSc8Kn3XR4aiP40483tAUpapA3fKQ9aDub8H7DJRNvx
hiE7t58+8Q8wIN5/eVP9sZEyYO6D8TWAzeILjH9j+QqA8Qr6b/h7VnzbMuL0t/lKDP38AWPqZ1vn
79BejWIMt+V/JZR5kKdB5917AqNm6KyKfngNlWDvVzbTw039XG6rzqFiURKSiGO6wKZfqM0v1dtF
TOL/Xd6FZcwysSc3daaAlUG76Ulbsco+NqLZ6AShXeBKh12gcbqTBfRAVSGlUjXmfPKCJZfKBQL7
YiCGd4Cld11WpU2KpsoDnmt/hmEApWFCr0CgjVzzl8xcBZQvyVKSz/SzJFQGZLPw7x1DYK1W7z+q
ZRC5qQKhBxF7p/Stl1QDzVcsnK5e0z2W15AIlzTyKChWZZX6D50qWZDgvjYvRSw2CesCmwBvrsex
Oce5MLTk+JUInQEE4B50n3MDLTpU+B80ykQBh69vA9dNQFQSJmlDUnL0TMLYfvZThoshn1JELrht
bOjgMFB95TlarGtnwL/jgeg9zY7jxnEur5A6ps3HQ4aAFWMGwaI5VNLM9v1Y/eyj3nHgn5i/s2kP
lT3t0NPLOk2I3iYkZa+Gp8zmhgGI8Cq7tac5sVKLrfkTE1cGh2j9G3H58KZcdleyLin4xvhkJK2M
dUVamb5+GLmxewg0VE6ObYXwY6fRPogbr09jk9Bk8SBreeWqLmkl2y2b4S15+HVwS+jMkzDXL3Hv
Ykph/1IdjQkTnP9OykECfrqtJ9BpBvK/HHs0XydN8kqnwyNJ5WnvWDNs8kZsE+ayUBLVWpy5OrJh
7/m7xXf2kFDpUFiUaovo8aAs0QLYKrOiezG0EjUl5oyexEz5JFDCOvl0+cJlNfkKhp2CAq0C2cWm
AtsTICO/B6gm1fJmSg+iyL85xkDDZ8oC3SDEAI1a64rVpBKvaHzOqTkJCImoyrfPCdFYsUIZxei2
Ov+s5HhzZbE6o5i1E92xYmyR5vwWHXSKuHb3GFJQ5jHqYjBW9VsFgH8IXoZYbeWGKKlm/iOyEMCJ
KE8Goc67N7XgosdzHdEVoXL4uRatWme6diwKagVmoc3sSc+VZZEVNqeXCHuC4g5rIjHNHG+An6JU
RYUoNyLabeNE5+ZVm+/lsfKFXLaOsY1Qb0zuQ687GxIdc2gHOdwI4Za7Mjb6vo2th7hPjl3b7f16
j/O1lwVYFmGKSfDVTDZCLBVO/OTOiHfj+asjYj7pbAYGoPac6QUIxLuYRyYr1Hz0GH7SxXJU/ApX
unAEZtqEV8Yza7nkOUsrW8hkY5EPMYjRcMnTraOr0f+cXC0R6cAcQoVwmqmjRXvHdRHejWBMadwF
D/n0HV7GWyy2cVMD28LHlgzQ8OWjJEwS9QLfXEvqz8LGsQCnIqNJfm5pstNbkceRahqP/y5mhWan
hyqo9u5G0wYt97yYRpPTMB84SRlvecxUsgaDVT0PUI0ACAigp7Vr6NzF/xgYV/x11NmiyFxNvIsB
z42sMtODTVG+XJ4p0KP8KiMxqbVolU3HObxefyjDz4JvdrPL8O9opstEJmq7zsMBTpxEbkV25g+N
WIvYrDtVpkRgtTbjrPrBfCvgF2qprHwdGDILokB8S0kJBP2Hr8ss72uCiAjOZuhh2PJhxgpuiYfL
JdrZwpzZ/KXb05EKKpbLQVsHa2cWUQ48d3A6jZoesroznJGwu3UQMUFdq7kRD2RFzW40u3yAqwX8
ujK8mtS3803auze3MW76LDrEX5bYW9NKdI4zWBtx2GQsQe5onkYQ4o9f6xFIcDGzIxovRUGu1P6p
QTQAhQA3av0BezRepyyWk5D1TnJHvY1o/YKy8jDrmtBdnudI7bKUt8Yyd7KBSwSaVKLsej0LiRMJ
7EeDkR0lh8XB4Qj82c5fIcTtc0ygqDpE6TH4EJCk8y/oe+ADEfdh/kNdRfQ7K1uUHLwEe0oQ06Uu
hbRoA3+3pdsZcgm0BmNOEnwfBp2ccZb1OmauDgq/9kgrl8c06418C6UtL7c5XfXeyOqlfEg0mEaC
feRYYfxAR2pn8bwODPbGytsdyJa/cF6awIK8mP6UR9OUuyPsl6sdWtCBGlgTV6VbWPa4fgGZxxs1
yfKhPVXyGWTNyQRYbCSRJKo5v/G7JiahrLoR5jCW0GJlZWcD+G1igpS8+liCoz7RHDWBjlX7ilm8
4QbkraAndyz7USlf8+cJOodC051RpgyVAASrEuHvUEhGWNBxSCE/mpXGcUNkgs3nIQjqv8QqPiNy
Eh3C/qD9Xztg9oOmEd0TE049tJaddGWmyq/Gcf3SAy2rMhhzyZYT3SGQBjs/zkK7FN6/BYJ6ki1S
7KzmI0BvEuKTOfKh+NlS9DC8C9xyugN/1AqQsW4yQ/4OkTZRDhA8WJhyb7W7d7wc4MqDapSnR9Hn
cS9PXWxmCZD5BCB+eIzmff8eJFGLgEzTviwnTmNq5X7aK+jDIOMJ41kz/XHF947reo4QBwU0Bz+F
+dPS3el0zIyWYXyhFG5WbWwPFTMPZ+5BN4lF0Xx4/cchEBhG5/+k90U7999/Q8U11mjEkz7VCaUA
uYz+TAaBLOcqTI3tr+6e8OjcQm+9im6FWxJvrq2RuiC1AfRGP0JkWMs9hoSw53wLmdNkF3CZ17l1
U6zWlH+wcAeXiQWwZR1CaU5YVrWf/QSNg6BAXoym2NFRgbKV3fablmreAMuY82bngfRx56C7cDbI
g/9dQjnIVg+k7NcNliM0iPH4l5aUaEB083pGs6hCsjMjwb+B5MOlbdJtmFtggk5ReYgAm5Nfk9ZF
f0Uv7GjPJxxxVLrVDT8p3JPEM92vlfMkzD/GEXk8RDV51gn9CMsrjYDNkahc/grI89REE3dyvpVJ
HHHtWc95+PSjCe/Ts15goe3K1rjV0SUcaq6axOWSTDwGF8+vbfSgKpHiHwKmGZuGGHaqEdRu+Sof
X+Vji1BlIhM4GIuJERszX0IhPO6m3p4eP3HUWC3mgJWFyS4eNqNS1OIZZPdt9mnqCCzr83OXDQ5i
5V/SmYBnOtpekENj1lpZAU84W8UEEdaOTE1ZUbyDCkQ/hf4yypNo673m+ejxPrFKwuiPm31iGpfu
PagHcVFAl0jLkb1qJNxTYc5fvreDxhSCwo3Fl09dhIMETYBRmAcYLdd2IPk2pTWV25gREfLw/M0x
RVNfdHhVfUB3Md8kfVdMe4+1Ci48JW9y/T+kK5oW/6Y8NSRTj4lSdqrb98eiOKmEoSz1+FSdqd81
28X5zUxGdeSPk5jAOYyMK+ZbmN2qURtMHMjL5gMtjxvXFK3Z5HfnEZUhdGDOhTYHBBocDUysUtfu
yXrXZvpk1sDhHcMKKF/dKp+dVWoHwsj9xv6oyjgD53xH8hV0ya7Xa18f9xU5klMOQruZqQT1pxjO
rifknp6PEke4qqV6sgKRX527MDqBeefXV4TrD6WrC1vNr/KP8wkJxPaUg8lQP6THXYKzUizZGpJz
DimdQmpPb+BOoCY0+iRIik29HtqkfVPtQ8gGXA3gQVZOR0b+T6fOzFZCnjorJzEZFlAJnht4YTzP
WSTzEafiVmx7JcLp4I+YRabvvEluFc9B9yPCwwOi9djHdQ9HI4RQul9ihXhfenaDHdOnO5zNbHTV
3PNSO/LeemlxXHQIYh65rBwf5GfuTDpqOmwBIXXZdQCNudmvNGI8sLCWP32vw2nlwk33dwCCHoAG
PQPAUKwdEgvVOK4UcZ2uYyyCq2rTsd4/SKxl3uvAAs4C11YYARCGGTQzk1o13MeG6Naxfj1EIKCc
jqexZYjfrslTw0pn1ymKVQ4iqCbeL9Da/vxHHXcgyM76ygz3JmDc0SpKhsqzTYdxadawOImb2f1T
TaizDRhV8XVZojr19Ym+6snJamPrNu6g+dtbBbHevjMPA4ttGH04S7FhLgI8k2sDAlKcAIkmAHov
5Y4NvEBnGjVb7TdwUj1iHHeCL1nW+kxQWK3XLAJ56po+GgUszD+kutn71h28lXEu1U9jn9V/z7LQ
D+XzKbQtPUCTwjVl+sXXJJkMbvWUeqt+sn4pzuq02RnSgVBlT3lDx4Sp5DLXhiThiiKTIfmU+Pin
qu07u2jQSSOVXB7mewNvWTBcoU9M22YdFZh5eI8WW+3pVamJwFCRyT7fZkmpZuHqDYgowbcM1b5q
OeFN7UFw3k1qmzhZrSQUNR4gv/8KMwM8AGMteXBT5pmrFuqOFniFpRFJKNomvddDiJ/d+v9MGwJU
hV00QLCXRV/dwxJrPnLJTwKNFY7isQc6j3APEtDxqL9TXlOpYDV8JUAFn+vboqxiYPM9YqBgzvhK
QzWIi7FOjgurBkwIexVe0d6dl0UiooMRROYyCadEk7mzJ76IBx6rqqK3vIp/pPGyZ5Y0oOdJNcEw
PWLRzglRqVvcHyJlkmigM5OWN9dg7GpP5Ffqh8yL6KxiD+c9FYpMiHCBa81FhuuUP0F9tgpOerZt
fSfuvAj8cN5PdHT1NsBecxYQV/CDf5AvPaPsHGJqp3Gbmnek9JiwA3zHSkC/iObA6UNKTtDetOqF
sCzWDznvf+i0YCy9hSrKoDMO4gZa19JTbhIvAToKrHf9KNgiVy7nbQrCSQoYKxrjRYLk9pFEhT4M
mCfH/BQFl6yykYsm4xKDLg9MPAs/2m+KqbRyqj3yu7p0X7s7eMiq5ZTUF8NT6/rn8fNhVczv47ze
/2MZ2PFn7rPrWAGWpbyqUZSzp4hf9CkE7u217gBu8JlpFxcVmKe5cSCWfma5oSWboXlS653zLDLD
ojn2qgmqeMq/MoDhoFsKYvwRm/FAKndBjGMLONGxD0ImpNMTVIcASNBKij09rSaGHChl8LzgE04C
Q+OgesPugTpLIbLZiFdXjBcLfzjUZZBKRTPdo7ULQHWaNyqfQKtac5azGd9FfVWtG7SF7142UsNE
FKPq47b5SJ/S4nhfi6pbxsQB8Aj0pd+FnIJ/DQsBVNdEUu3lHKViY/Ugd1RupdVHwXannyd9dGKE
xKjEU8JVmDbLnbcjdkK32vk2vy+DPJctpnjTckXv3ialJOQ2CY7FLMO58j3v7iAk8p2Twjp7As8b
+7bdsWJcAMx1yIMK+EsPxrnTB/WQrQpFPtDZMV5A8Bsa15zKmIVCwnO0IoVKNNLYcoz10oKaAhv8
ahIUJf1YdXjWa2isXVUznP/vy1PrKDGonkj5jyQWjQRpW3LHFwPZEOhSFzz1roJGYKfivAYVA5Z3
aD1YU0y1lM/y3nQF29zU7J/FeF2BlhvtVclBZ3ZYxyssGpkMRSWU2GlHaxbQGmtZ8ul3JeFkLdCL
kPGmNX9FyWIQCfoz07B1BgAqP9itTAwh+ZLGF0eSnkU2lX/iAl4wn3Z6S54GUhWTmna/MIHPNW+O
P8R8THUlRud6qrzeOEzwnBH67PnWnfbwquciHsYVwEdJHorJz+te8FUooioN1/GU52Pg0djjhyvW
5REyPK68kvD46kWENKzVmViq9X2aHRtdB4fXHnDMgMJ8s9Rx4+mTgudPOFchEHuf7TAjqCrK+AMP
ZHaqlqBgqkIkU/v3ZAnFzoRcLbUawNnuCUAwSZbDynGpSmEHjAGuU7UUXuTpxMh6bmCKLpUEyjkY
vVuIAAouLsL7tZCO73OiXQWfGkTnDauTdHaRVFO5cea4Mmq7OAGpwy9t80DqFymiEiMHq3MpQ7GO
OWIK6BMgKDFfK/n2ZahpVtdMD/DMUZWZooeYIRVlsbLwQX/rSr41upJScYEjmHcrGNS6Pq+j4EZ+
Y0lHC8KZtXTYgb+9CZl4WUCxc5B42A+jyMwPBnJIV312hnxKhNvwSHtseM3DugtfgZoHC5eOawQ3
vzqP+q6etak4KLH37j3K1MkCPqOrdFJR8UkoE2c9webh5AZb9EoXP6k6ESE6a32CX0BWqbYjGBVl
Fh1cSQPH+aFDITmQPjRQgHXcPJNIGGIOA70vT78HuMvYbW6SGg1zVKFG8RlzH5/xrIDi/OVl3OIo
l3S69nKxUWDZOZ5Zcz/kJr8gqo6lj5wMKl+cc1F5uKDWaJ52AqzX6fvqa+sOYiza0l6UrpL6cCpk
8C5jZI7kppbUmo1rWAto5rFnUyj4UCNke4h1w9cN2oaPlkf0rxOV74PTOoAEj5wcu2Fnh5nCvo4l
pRtBOnKVqepyS+G7u+VHu3sKrtzQtwAffCMSIsnpW7+oFuEAH4cgnKIZAWXGOuHfWMGmmKDzVzbk
eB95MyeINKatQCuNC3H062tQ23nl88YpbI2dqgibmuM8FhcTTOUAEz4rxQPqiuNRrpct5BsR9gGb
AiNRFSg69mgn80X00KT4PXagc9NcE4vF7O+ekojkrL0KlW46IAuhX4cnTb9uc2NuAtoF8tSaOASz
SD5cwJLrE2yTj7lCdRMoGamkm6n3OIt95mnDoQ2P1ZIJ0DPhA66lbLoVUVs7A/BZFKhSKcQSEuzK
u/O82dBakXvU+Ou6dio4tqdIOpjbuYAZ5IJES974oU0YWYb5rTg/l2rq2B2S2GxjQdaci2SAt0W8
DA62RbFy6vwfPG2qRvXyyK5wTAk2ncmnYSC4x/2UtPmweYe0vAzm38jRJKFuNlNmiKZ11APzMcwb
KszSeZwU2Ls0NdwTGxIEYlP+StJ3RugHSqxGfTzAO1RakQBPcx8sVqSuvXSXytAeGLqRRt22lPVK
TZX0gv3bT56grikTilnq3+HVVLkkCtYhHewHOWOXCRXOdodTFBbf0Zcr0JPzQqotJsgOWyq7AZY6
96AsgXFUreHtOPBBYcM9aGr44s/b5Hdn417NwW8gF2TF6LDrVXCoji3tWIeOUnwYNLZTG6zZo34C
KZN4QHpI4aGzHRetpxH3huS/sX2LtRvxUgQ2qr+71/P0NJOJbo1KXONgsrCW0QZr0WxVO4/0yMHZ
WEIAaZphVDRE+bCdAfRcc3iap5QAEHOq64sypOOiA0YqMYkUInU+1ALWALf0K6JJCiWdmOeb/Xwn
cX809z+fMPR8kHZ1zTM9v5PEWYvw+JGj3hmE3c1WJ+JjjlnvhpJEQPxowl1Pe2hHva2WcVs08uvI
M3W5tJVDIcXWpyH7xSTux44IZhtSDvnL2A95O38UZMmINUxo90VJTaJov+hJj4YR44Cmcsyod4Js
XlcA2GceOgGDBlZ8K5FU3LGyfgfkJKAZCK2hnkuHKt/RQfotMUf8zq1hvu7gRMb2+A7GYX1ENmdn
Cl1679L+X90JYU26Xkt2AnY2q3Jfaa6Vjfn4+uBonT5OZAFfrffVoahhcLSachMAcgu+37uFP8aX
11rjEB71U2dtl0ucpcyB/ZVjjqcBMs230NKTr23NN+ZJuX3EVh+yFsO0m8iH4xsXlBLKgHJa9DyJ
uPICiaD5TtcbOCKlrixkw+5Gxd0LDYeSPNig8Jo6Hvsq4s/OJvN2S8F1ckTxjdlhpQLYaDIEu9d7
7DtWF18W0gPsb81MvT82Ul73OeH93ICszP9RAwQdGglSveFhvRNN85gyP5vV09FRcY5V3GVrx9K8
KAwPxNoj0F7JZ/dmazZYm4Cg5V+NY5+9Ko6bcPlEM1x1LvCqMB589++Kjou0esCrqSVfjRt+Ov0m
GOP1q+cGAnPqHhI53jtmQEztnuoAijt0cy0pTBnM9COV7wcIybAbapLJMHLAGo1+PSfNNwjwctQT
5fqtpHa6zud1wM6ToVH3IyaJFNw/+OqA0LO14zm4tHscVOLID8UnIUkWlsMBCyug+ma1lRLEVgHH
J+FyZ8Ik5CqyZ7k6Herb/c96MP/kXxV8JSHeDy5Aj8P9zg+o5F5Db6kk+W//p/Shd1ciNZ3TV4wH
AjDX4XA9GYyobEOZ7Wp/gf9ISJum7TyrKJLQoTrJ6SF5+lc1BEUzf1iKAmo7JhjZZWWoKWNb9ZQ1
M+4ia5z1h9OepdJTcgY9YHHP8eeDvSHMrKuW9CNksgXyPq5rFcFKWIcNqTp1Zx7IAij7g0bneIVG
bwf/9RDkv4JMPh0wIrNMmPp7OFT06dOmi69XdE+TJ2k7Y7lKNKIC3PU8ZKOTHcYpe1KYwFvKjBSy
w/8nScNNbDO9rDA+Ux333SCB3rA2p1yKfoP+nkiPF4T/zfAkTx9KG4TzXN1rA7ixAQOYKDGnLlYv
Dg7C0THL1zElcsybZVwLbRCrpbStXuQRxcEQ9QIjBhUWoyo7YbiJgXoDxC63lKJ5EHB6HRwIZ8VD
hPTW+1ZrTpNyymCPHxe5TMS7eudLjisSvSodciGu1aJZEdXXv39VkfVFH4kq+rhEN0DuS4caAXqj
yJz4y2tyHnxAt7LemeR6JKsJ0T25inHiqbEINQAyDxHDeLN1sfxpiMe5ltCMHUclYKfouUjbCa4J
I7SetDI26oTnw61R5o8JFgtNLMrI02h1j09OUQj3f+pKpzsCfgtAKvmsb+E9qOaYj/I7jEfPxkhR
9zVBpqWlXnTXO+DBQF0XItbLO+Bir5Z7E9LCb/q3lZHYG9CHv6dpFJmaUGeIMJDpdxcWcbX5B6h0
Girk9nfzhndM75wCdkuxJqS+oAzB8yedj79vuJQnJ+dXJRodxFCp2/Jc+RBA0Lmz8gEQinm1MfCV
aANBojvkkM5qSOi4tM/y16Tt9bZ8bORn3EQWNtMiSEyfSYxoevHgvCXKbP+flJsT9gIpmmnWIofx
4XKxzTifunFg1Yq31thlgkP5hmRuGT3h1PMpibOtEBaPZHzmPor7T4W8EODqQcZuX0HmIk3txf2Y
kt7/sOPPHbP7tkQK91ZJAYwm57qjsfh6iB57U5B+Vsz0ecCDd/fX8gsnoTg6ZgLEhV/GizKNyHuw
YgwqYuhyFBfi3+28GEFKWQq0bSc6fIEfmA55nd7yVo2waZulOwKlk/t6frTrgK5wAu6LyrroVUff
cDSnvZ48j0GSm8IJ8kD4c8/gXL2IxIDrRAqFuJLjI4Yvk5iWdOGa0wdnIFd41R204JlDsN5hoImv
gh3gg8LSmcrnyV7VWjOrTMcUCuaskScQukxanpSCU6k8c5vUJ+kZc0AsuDlmNUWEKVgdQVYpTERZ
0kiadpyxE4L8Gy3n02Wh76QlR9wQmOrkP1uszZxFZCOgfC10mZhQIRvTxtcs1iWwByml0gASyHYU
7B7rdfWY2wQesMwpQEddySL1RNZ7xY24Sd1OsHBorsbpqDOqlYAT5pTq6cIntIq38CRWXWj6zZiK
GXRAu2v/x46KuSM3dBPb4ra8BmHIhCf6k8Tnm2aO0d7pvvK2mOTywRjpi1KyIhCtde0cFfeSDyZT
GWU9RiNqJrreXRmsE/JHUYDl1Z+mZmt1n7I4bk8BOGtTt3Cv792rtdO3zxKj+RQRzQXm0fxaXzAH
OH3uYQpgWRQpZXIDM+T/IMqRapVJmr1VkgnYl+J++u1sVh/S5+bVPZHOILvlGNKEnEy6GRihhucr
fDDiS8FmvCpC1NY7uRaLs+Ko//ALJi4fgaXUeMc7YIozOMNEktdYQSAM+Pp9KWpVQShMIdQ/zkWB
DOohl4VpbLaC1fS9ooIO2zmzKCzqklCR4NPss4NNFlIEScHuM6R/CkjXQrB0Drv2fABr6tKxBN+I
44sMkjPhiOzPKq8TGd0ppVrS/YTsvVHBeCbyGIsS4HZBRJFPgpo2gVQlcjS+/14lu1VRRiWh+8CU
QkBZXRbChR+1hhV8DCGiY8DNDqcM0VU51WROukldhXun9PviXJJlcUEWJkccndyGhMr/l10A8BqN
7oNSj7n66zl/d95VllACLwMjg7ocZK/+Xj3HihUxI8zB0MQ27/IPcBb4XcMcXRmly9pulS+bNHlM
JAK4hOErtjUmeLO1oJJvhO29iP1DcDUuS2HLVjAP6plZiwtALK1Xkb0hGOL8Ll4g4Bp24zvcS/sD
lNkO0QSOqVQIgKk+jdpy2VJpPAdMsxm5K+oiYIA1T49GOe+RoF0UWr5xr8JDaOQTXUHLZy9Ec7JH
ayWqCHV4Bp2pPLrTaWkjWRBTwsF/3/v2CLb13NNWZcwe4V7L+MpyAe/EYGSUYgswyIPgz4T/3Ibr
CNnFQk07lcPYDqkKb/X/IhxI3VhI5bbKytECuaJ46adqGlCcLqD8GI9weh+QKs6AlwbVPW7sjMPA
/QGoZhSSfNeXW6XOkj6xMC4YmB1gP8jHcXT8UASGQ3vJz1aJ3bijPPJxoQXX8Lfb6rmOOUu9vMLS
3aQkTaAqsiq5+TQFpVC6xdV63O1IUYYnsb6fJg7uRT6kLnm192nJ7FSgTzDq4jhQLRiGAsIlQfhe
KXqX4ODe/7cEM/Msoqj88HNcw/x9B+vxQdMSQ0MZj0K7KKvsdtP9INz5AnLUJkFFtYqH5kMh6581
OkavFXNo53lpvb1++wxSvlkXaI5KxpJcHVqFWFPmbU39KJx+r9t1mINhUuNe9CKCpET4kvgTQyfk
f6NBYXMBUNA6d0qPnAO9YxTdAh+J/uxgLX6W+aiw26rJg8gHeCpS9InTj0oRwP/il+5OfcwVxwLt
+cnVvdJFwAZ4whOD17oUy7b1KzXBDaPwbBjHkJERrYDWjnd48zXTPZaJKlwwg/cmURmV0RPzrP+G
n2U2blHZ/FvAZKZcqSj2v/V2P3yKFzmNYsU//2WEORUNRM53wTDzWWi2cmOrKxbKTXwqsWNgceNY
YGA6kU3SLgoz7QSEm+CdK7pkeew7bXsuOZX6s2xzmXDN3Jd4oOfHt6JmLpL8OfpXqGCR72iiLEx/
8q592VxDJeRy3MjPKCunSZAHmmTwmrgf8t9qAx7ok9+N3LEUFwCxclM9N9zeho4hP/NoXgAjGIiW
nIiW7yyUacN4HBbIMJfzZtH9crtRcTT5QcinjEh8GASzrEduMhBPijYhuhOenF9FXpW0+7BcZajn
zOYw3X5qML7WNDlx0FbunpcMM/dOm/aE/wGIT+Bb3o9wpguWgng8aZ6I3SPoba/J088zjdRSa4bu
37St/sE67R/LDsh+nRlCRIpTL8lUY69oH5g+DkxtdM5lXK3xg+r9SUeRRyWo1IA4SOOCAzbeuIOZ
mSNgP9lzGYIJXJJ9O8EZg+qs+TrH8iBuuKEIcVYI1J2D/lmfU+h2c/ajs/eSHNGhG0Cd3Si8KSSA
e2jtsMWwxFiEkfkPPLu+4URLhd7IuytoRQR3bZg1TAYCZyxEUEB2KwV6mqUtVHVDgF8gtin7new5
PNrp8Rx+UdsOWL6MYpbDF2MnsYhmw+WkvmX4M9kGWZYryNAM7N+BlZRQljRiLEsmnMLxsoaJYipH
XAc0xjvL/G0mJlPGJhFXA0IfrXiO6vXhhtweMK82mBslcPqc9DI3hnNcNalMx+QMVheTfVek3WwS
76ANIlPvnw72wekT4zbdW7uvujNW847ZY6hDE9MTm1rYDZOELZ2pAKhFZBsUZSmzS5f5ChaP9uGm
syvdk2AlZC/fgAQFkF9aJmpsUyQLM6Pf40bxudq1DVZI/+phbmkY1fIOhwbPEJlIuzecpF/PWcpu
ux+VPmw1Tkzp3L1m6Mo/0R+YhX9HhXDMQ5o2zN/6zLfVoFI1MrNozoqpPVsLtcPXacEQ7vioSXAI
ddV2VuyaBfQr522/XYZCw7Xcy3ayd9gAc2vhifFLVnQ7T/qYpA6D5VR7pcouJGxb360Pgd0nmrIe
y9f4ZPiuMsRE9avivAyA+cNoea2dSZv8YlqGDsz8eKZXqcxUnNVhuLTl1fChZNVkjCvDmJcz1pmg
n587K0VU5+oOhIdapF1LaqKRVXShSZiAG7MZMwG5D+5qDK52Iak0dg6blwGqG49iTHIegjaiGGN6
oexCC+aRl4dr2ileyQq7X7Y+hMJ9aN7BYHT04+ksJ92B+lwWyGDU30CaMlcBltGiMXiNzVWQ1F2A
7yY8UY8Sl+qCEMlAKjw2uZ/W0UAaIoFhwR3ZLrjZA+xC9R/qt/hLvRXbpIsa8H6vU51zl8mRwC+Z
nVpKrk6PfmKLmISWd44ghHVs8Vb8Dx2Qbe6o8u0Nxnt8dA1PR33TCiz+U7DFBTN7vQ1JU2EChxLo
nJVi2ziwDPzG0rBvBhPzfbd9ZhvOpqVi+xBsfgQd/14ffsZPRsO8xG2zBr+uitLf7wL5yaGS/XSS
6m+weWlz4AvfEmHdofBwZ9SMIfqZvnwUoRTrgqnuKm/q5UjpoGcHKqGiuAiIQ9joVdnQafJThbuW
iN1iN7Enkd52Rk8zwOuKukK9G3zt4O7TwQXkaE+pCjvufaBmv+8SGrYxduivmZGkoPa1DkVUi83k
FuYpm8e5Vc8l1x8L07wnk8l7H0AcGjmBDxVu69z0dOGkoNEVAiW1KcJkA2AClUbt1dHfnGDZO6YA
DmDtoMhzzH0n873XfW1eZfTEzOT94hxEG/Ozi+puEM9N38qoDOHUsUzbHHtYUX0kWgVL+dHOw/uC
gHg5TcBLBmSs0+wJ5KtGuK5lr1tyHbotmzEcpv/5EqSYtC/zNJEtFptjGMyiMSkkHeV5L50K6nlr
VDjFF9KPTRji15qmu7Hmhy5M1vhlneXgqVuZQEf1+A0WwvaNr8360dt0M4DLIMTDyuwqFAFhVbJE
CIJv5BSinmAUT5vVOz6smmDsMhkunc8Iavs2jg8COSjaenSSSqOhA4k//ubFitZTb+8Nf2dxE0EH
i7TVDNPwV4qQfrJlB6MU7OV2e53LLYNmIvGWQSwPH01UbY18YYtcz+N+UjRIfFkdlwCZr1tFGc3r
Q8eo6e7xXRZ0fjScbRc6ySD1sm1vhviP5VXY4hOv4oZJXKRMLhPs+1s3qvQKuOXevN4nASR/e+WR
TQ14BHno3YZrN4N+6QDPgHSoJox5c9bsrz53JLWnhm6qyBHBBOxnXIbJQ4jovQDko0GxEJJCNlha
hpZrq8aEhD3KJE2SxGF29VAAokkegQ1vedkzHfaujidjApRj8U5Uh/W8Z21ZE3xssXdW+BI1024z
eTUCA+S2F6I+SEV6bhcislaDlfz2FWPpd+/7jqM49NUEmFd9H8Ykq0zD4N5rvap+spB2boarJRQC
71EjH+kH4firxk+alNNFwpgOCfMQFAAWJ1xDTHBAVo7RjUZH51BgMljQHC6M4ihCBj0y+W0ZvIIR
Q8sRKe3c//jmnhef+1r35o2/1jpl+D1gnuMnnEKAX1VN9l2cRdftGAGSGFdSMoQ/OUJeqJcmYSx+
1fzU1dLsMVYTttyT6/5hud5VphnxCtvyBYzj9pA2LjbxRWTaVLdicKUCnHJbTDf+B5BOwV0v+2yu
4VXi63i6CeG24ij6t4vdli9LUZIqgtxUAYeFftwO+L9vVvSrMvZcIMXUSTxoll/DUTFV4pC2UslY
CMNmJuClNf6ioyxdk+CeUtVah0HbcscJSo9uyVh2D3kRmFZieG6vXQs89i0HPMQgza/OyZ27fBs0
+IxC2BpzvC4lwy4D0ktQm83PHH+40xETpcgyN5O8jfu4xb4bvopxjVRHlVL2cvMLCB5e4Fv5p+7M
VxTCNBNU1t8kqbwVqT0nG2XQhwO8+MXFyAyjSei6ZlbsnZmwff4JABsEfgKhlJTul2roRdSAPD6j
Jl+Pfj9ZZ/IJs1So/lUoM8h7uaQ0whq9NthAflIWf/pd/Eh/LJgWbhu4fCbs+tg+gLaORKkn+DYi
HSDyyM6lO7NBGuQS7byOMRmCmY8rFBQyAt0jwyV7/2NdaGhhFpTUG16aVwtNTJ5f9BxpqLW0GiGq
8L52ckT/OGO8jY7vP8ohbUMvxpjG7TdKcqsY8cNKiyHMSrCRNm3GhZfS0s6s6VxQ01BxWn8hN9sD
5NIE0YJWdK8+7dmmxJ9KX6elYK/OwfnQbGuiQRCPG50dY7PcKLU6rfLskmlz4nCw14dU+zhtQXpd
JsreLiwljiSVUaXBky/az+yvxvFPfBiV/jifJbBDxYjNrIpot14smbA6JOiSUizZ9hDIp5S2isd5
riAGwLLrBX5IgJsQX/8rkb19v3rtRoTA0stc+jJD+KyB/zsIS1NBNWn91hzLbkRVloOgVS7gu0ur
53Q+lOxjlSezAUlAcef2jMeuO7so4I7aK2JinxVeq7Z+WKhhXUkrvU+OhvNPuoza2POEn8zyaQSP
Nv+hMUTPeT1IvLMgxjcIa+RJ9tA3fUhsOe+WO8AlZ8y4tB9oumgABRCjQvnNHDJAqdGI1G9njx3y
Br5jorSSkEyW5sJd245jK13vuF8/d2cU5d/KWpG44c7Y42d9loaLNf2UCvC8IaznjdbOfG/gDnUx
7eGVP/3+wLEGTLDV5QEzCLvHTpemuNQcgKGkJyrNfIYvYsfERU4naN/vHltflxWroab6uOPuDKxp
OwolR/0YuLFJIeQYFZSIKN53oYH9vICV268nxReKpUdefPGn02PHLgNQ2xtdvWbjiXEUdPt8gO+d
PnAnpT8DCd4VTBp9FVnj8IpeJMW+67KrNiq9pcdjNlCixjDauloUo7IEaXatD7f9wVkWA2/EcQz1
Cp9WUYlQDgu5FMHysHjAynTi5BmarhB8/FxPx5U7MNz/b54+7c5btmTTUVHbmNtnpHRZd8ojt8KR
rBJGa3FqX3N9vxonskixTpPgAoVtgGuQw8RcLgQfOUCS34HgEK9yu2uPwQa5Vcn5laT8dNG0vYrQ
Frj9UwtGlSZO4wN3ZCgxccJbvsXKEVOMkiuGG6eqUzFGjA1xnjvEpxd41jw/l5H6yPM0gsAkKcCu
OA7e3ZOYOJfHq1kPdMdGAG8PysUnZFvGWX0E7BO0q7fkwosPiAzNuf1Tv14FuW/32+V0yOpEOf9t
H0y73+KCUAUHY+0JRs1WzjjVRFNoQUZrxRADAQChMWYfq+g8dEDpnY1Uj6XiTRTbVEmvmtRhJovF
xGzCgp9yJkI/UPsqFdIdVWx2+OTksIo9vmkc8g45fsQLczr1CQhFb0jS1aIufAUNddOoCFTNk769
8rIE543yhbMSs9aO3jL/B3lRcU99IEUCCysjtIFomoRgOcs0ylVNa/Y3UX3SsdS9Tjn7NFse00e1
o1QLrMzySIZDWCs87y8ktBcSWaSKKCSo9yW1Ni6s9sN+qBcvTCwS8eFUqguViNq361u4QCPMoxnH
Kpgd2nOLGyS1YIviGH8JORx8bVxjRVFcL8oeoH4eYAgXrRZdYh/JJ65a01FKVvcsxOkSAwDPDSvi
gkqX/bP/5vtNjXRUpS34spzPsAoOKazrXLOu4aoZfAdykoS+6Nc/X7+KLF0P28QFtxPXZpPIinBJ
GFq6iQxUDPemo9ipvljZsl7RKny0OhB9Dm0VoQ/FFKCEfxZ0vhSaWtVtM4P+wSY98f2iLxwkjUCn
zVMKvb3QK0BFaXclkjyQQKRoPlPrf3h5EqEx7wd0wTXO14i0eW92diXfyDzkyp3FxwybQ4E3msYK
P376Y7hlpdS3YP2Qh7j1ozU0AgoarQj/nAbW89QQiqRCOdlLz2UPUKMqzoaJf5mrrzlJCNcPlvDP
3Ph0bykyWhIuMkJE69F0kQ0TcxV0iC9MT1FFc0ZrP6L83k1K783IvcaY6/E/RLCc659fQ7AIJF/O
8EvFYjh2nZ2CvdPTs1wSrTfL7kWgrbPW9Tz7QM4JXY5qrln8iiEEp4u5ttOtUu2YuwZXsIPejkQD
zxydourEwzAxKa99HjjC8XPzsIYND/Brjy2rnSSQlJtlYG0Q5xY/Gu8ET6VplDS73QvIjsf1tVJS
N1eMGCeSK8GWeyTYHQAvtcPU41EYHKo+PJuo7gut/aIOVbNogsRyTVxPpEZigpJVwv8QFdnBKzXv
7rvnOraZUZ5gcX/afI4557XpYV65IhniV/a3VhjFk/Uy1Q23XK5BajvQ33yk5ckr8dYekEb5IDM/
Bh7kZ6a5YEEJuhcWH1aLAw0YekZDeQXYjaUU3vthFXKdecPPHKYAbVmzQZdy2Tgr1ozJwkVxPJAK
cggRpIl5ksNS5I3BsZAl978gYps647zLNtHLgh3p8FSnnW8nJhf8pZwd1murAyoxhBNGAoIWbDCs
KP73QesI8otG3gjKtBh8Oao/3gGvsw/z14+NNapS3TjXTMQ8ZvDBt8mKNdNPgZShXPWTIjn63+9l
x9ffe1y9OfcgUDGSErz2mdJsRFLs042lKndOSYqggBhcd07OeOgj10jmLfLXvrBmunjkaYRKOttN
Li1eBHcAFvpvsF8TGb4h8uLT/fDkRv1R4dxbQODRFvsP3iZevFoRCHAc/TG1nn7i+jsCPWsXpM7g
wr5dcnhJzQ8/tzX2tatme4vnlCApGJpve+wqyXcuUBSsXxUOwXAB/RdHtlRddbNBXz/Rp6cOBU3L
Q+yxZ2MxDIiLKxjZO1WyHcJuxsRK0iX5VjODn0nIBJx58L7NXqyYaYOFosyq7s7fxMmlkjIHmWr2
Kt0lDpsbiib6PQNbY8PQ0fh48Wjs6gKP1qSlATp9uMGSl5CllILvGJnlwUtkCtM2m0AJA2GaZzwG
HeCUxlAk7pzq/1Ge5I/H4tnG4WXGG6uJKG4J0Vvy6VM2uvELV5Y/DR23QTbz8beg+4IMvWBvN6Hm
8JQDV2apF2/qUGh7c/ESEzV63czsgYmRocerT47MFuOhWiHyQfkPUi9UV/zTuIFciQ4MiT8Nyys3
xHjorRr/bYZfNhxq5dJ9l+DEio/t5SOOu3zqEgUmk4WVEEIW31co0g4kyOBZmY0GME0Ljc7wuH8j
DCwnqct+/GnKeHeK+6SDSAMKzxKKr9RubDzXwJ8mQR5adMMoTCVokwtiDZKJFBY624z98vWGLKW9
ZAjFLmWwr5lojCh9TLeCOKQR92XWaourPNv3Q41MtXKaq6of0AZkIBbzYxEJ6oawCBQ6Z8U3T+0M
9rf63kv4ZCngXGm4ywTNx7akdwAet8M4iKNbDWarXZ6ySXr8l46YEcXDQwknMHKzCwflayiuaA4/
2951V2XHT5bB/F1OCsDPr1ehBV7CvtiAf3ep4OfpIXNjU7L9rE4qz+YoR2pGx6QFqqMoue2QfSQY
Bly7YdGo93bR4FTdYaB0uiJ9uTaAWH00LCyBaF0+RHk4ykPK44HzBmnykYeu6VQK8KNz7N8dK9+c
2cmobkAir2zMj0iyK5b2w01ZKpFk0x5O1nrteHDSjzcDSPxgQSEQYZhPfrtNohs0xwynCorHZZOD
7BGRIzb438/QSLWr34YDtml78SbkGMQPb2QtnNGrPUpL89M9uMxb+lHIxgy8wIQXa04itLQOhdLt
nIxdgVJrLwUutVMQOlUEpYVlhU7bXlNfj5JvKm/Y0Jly652dPRfmMi0HOH3CoypGi7pVUtYZkkMj
dD3eXnNkVO9o6tWmhLZ3gH2Hf2gMEWnxgXF+8E/kY2rCREPNIqIeIRB02K7xUco0apnQKAL/CFBW
JdrY+MZxldP/iJLKha9Cr7kv0nBBzc/8cxQvm3OoBKcDteF5t7dVOK/claCy8DHZi3OD7OdhvFr/
LbwSDh5GhWVlGvJwP3GLlixVzcukFqQvRDJawmJYZYEH9ons22fy/Xx3ibXzweznI274ZI1dbH48
9RS02o7jC/H98z32tnTJu8HKWCh2RnZC5gOmD9rCr+c6tusaNkBWg2ocktXxy2O2yaaoq2LlfO0Z
uO+2ELBVEPINjqTu8KFyCMDtK/fZsr0x2rHk8HMe3Bf7/3mDJbHoRW2Gedj2p93IL0RzmNpicEsa
egCO0n6fnxUUDo7wsOlCqJ0qJkehBmvELneWkql/pSCv1giOYMQVgCMVfQYJzfbDLcabEqqgFchb
hbgMlXa3hDbquFFfWCTSl6tnRTN0SgPRpT0qw1f71+dkUMen4dGttzyPjQ/A4tDFgvFRiKYl0+Or
Bx/RU97epmnPF8sWQfowzmwT/SlrvXQEny4gAksr69nyOwsMDwdVWmj4oWSHFzaP24g7JxElZZHt
+WrEwigYxGO0UmbU73guMxplydKxO852fJCme9jiMNwi4aL73aQvyh34RQXPTJonYlBqBMz8kgI1
5DCFHu/dZmOTeQX/CxqOuai44wtdivyXz6kyu6/mztFgGXd70+feY1lL2P9kKSOgHZC2Bq5yw/Cy
NhWssiHWYfRVyzF7pioObT02TMQVNoGFYaXARoDCKnRyisnLvTKVuT7ZZHZjF8BJzEujctXFDu4v
2hJYvu9t0QhWyVzegYPL4jpfrY5ykmg1PbbusGoqY8v4y5nI2foAdmdf4y+DM1YeXf0D0wfggHJg
SewjTPtQt8l/3gBmYS5lHBuef8e19K6/TFEmkSCeo8E/uEOv8cBkt6vR0hUYWPD0GGG/olof/f5f
4bkhuGSXHwVE6tb2qO+ozvEaTYRRdUt+eTt2hSz8+Zo0Incb4fdt426PRb2xPR36F4ebMXrMXbMx
ppBySq7obAlMDTJVzsxJoEsOJl5UTfHdyIQcpFumBNH2XhjbyZ8fUWFkVTcyJh0cJH73q+9pWpL0
YvR1HICqaxO5XfDxtux+rKKtI85bMkCBVeSB/Bu6GZ1z/4mn5hVOjcSUOyLHJz7cXjV1T4k6BFxz
TkOp1BbA8Qb6cMVac/yUoMz/hJKiDF38VWf/huYJibOk6xNbgzrRRCWo2YGQhhriSB+omPG64kns
Rw5EHBJ76adNL1lhMq3AGKulLHhha8a6rI7rENpDZlefRHd9WY4iGDH5ja1dllwwZyH/U+3acNgG
a26MNMsIjGDW2reuCjgwb9Qhn+MBMFFbRo3qA3v56yBzdqu46Tdx+i1iHskxTGH2jHA0Ri0+W5AU
QMFYs5r4YPOTezQhTHn6kOPIVSfwtfJ+QdSDFj4rXf6E3kIgcCn8bmAzFpD0IBa9caD04gJ4SL3n
7RfZ+FosHmFxcmf7RsPtg4ezZz37hidQHbkPG93Ju1N6dJ+FiSRIpwZrRi9uMnk8ohzYAkd5AEmy
vDum9ZDcyZjwSW1nJphjFVqndOKO/LnP39C2J8Bj5K/gld3LuDYQ/bEeKSky/M5CIDxGtF7W2fDW
plJPZkGa+m3oH34A9aAE/0PEO6BS7zf7xNwudXqCzWnkFB6TxkEg+w8cemvUQdJtljOH1f/LtsQ8
pCJTAOZSH521DgP3r8pPM9OKKtPQFFn6QPKQPK917qQBXdH73KY73sIYgMIXdThJ9OaTG4v/f97s
MMODU+YpDvl5ZUpMb6tmOYZ8bN5idIF5KFjQLlEcu1Rv8nY7eyDWZzlK8GdHZrckFYUQ8121sY65
RHlbVHZiw8L7U0ttip6mFIzJNaOQrb1I/HiP1SjlCmxdWVOVvFGIh8y6zl5SahpMPsbxc5oEbs11
MRPmllv4iKJcGf90sbd+hyk00pASzt1ZwiljLVfMdpBtzNTBycCVjfsh8wAr/ktMuCepbI5tNGcG
87iO6lRH/7Ou8soda5CKv9ESel7k/y4yL/IHh6FQW4qaAIdxZBu89nNDA6QrpEc6VWT2UP08sMOj
AFlBJ7uyF4VY0zysd8Am60BAnCYG7aDivc5s9hhdl2Gz8h08ScDY2fuuY61hx+vKG/nGRWdfo3KC
5/2dxsy5BjtmAajb9AbqArdnbv4K0hPtCmduv/pX694IhN2zVORpWIIFjLm77XZF3VB71tDuLr2k
CSZzImeBdPBNoj0MD2fpb+9V8j22A8FCuk5unn5O6hJjpAf4mkUUhPWeEzW2ZkPOlBXqxmUu6+4+
/Bzx6zDEgn4hvTaVSDD+eC5sO4X4U5QrNIzGJQ7oPhNUgXwl6Ls4rSRMUEHItF+X64qBo1Vlk+Wf
ok2zKq7A9aUjo6ZId9twd1SailZQxzer4SWeQy/fVfOU0PrSimLTMhFyhxqFqanZUs8Ml9BUKWSg
h6/OQEfI3pzCllmgJw/Di5QnQ1ekGu3Cc3DyI4lSnj4TvuPT5XAC1pQWpyoU8b6SL5AjuxNaBz2N
LUZzGuN9xFfKBso9vu42UwiORpDwMa8umNRl13VjiGSlriFgCY9eXocwVla8RWrWf5s0q3H2gdwy
eSoR8jVKxBBYE6qqKOH76mEF9lwz0y2fv6PRvaWQT5C3HJrX6Ouhmyf+OwxjV3b92FJTe2iD0gW5
RMRkv3PrD/3B6ndcsNLc9p1N4BQvDh1ooM5fOizu61cw/PDtMoJULBGjVRtED0MnH4D7inAGEEyy
jd02LF5Iki4QFrHt5QWcNKIQXByu8Yz73oZP2zipotZ7XZmL0rkUU21CTLTxXNX9ifQb4VSmwO85
2uoGgN2xgkQYAaIfVdwwcYnEedsufyEGwvAcNBpW6IL2gKoWqwsi061GheAegVl4mDkedNzUssN7
AWO2+x3mkRJszO23SIiD97+rSU29fJKQTWwAe/wFmTGje1xVnTmYUCU5C3Fvajinu+jrMNq9X5l2
u1euxdtmMKBJDqcumlTgsl6PySZfN1AxjeQRS9VfapMt0O7AvxkEeY33AnptNRp55WgpSjqn9aVq
wyxUnOMQo4Yn/m9FWtl+a4GTCCwKq4cvJGBsVlN3keBCo6ZljhDR2ks428HUfvc5wqsfSAxucS2L
3ztEw9wSykqAXm1XiQnaio4YjVIi+XlwwjAcK/P9ieYcOszCAY8HwUpVyPvm1d4kVk4KAEW2MYzJ
qLlbgFnCQ4gEbHFs97CDM4XB+U3CxVvHNZOaX4VXiYiii/EgPBG9Zp1RVA2Fi3UNZyu1nfzKOKhI
88vZxLX1I5l/jUQmzy/Aa2+H7jc68Xx0QquYDd5Iuq0p/EIAmrVUJmeZpSpjeiZiW6c2hdCsPwt4
UMExBS48oX1M/EdvLv/P7kb0wla6jW2IDz77rHtG/IYs+nPmMq1LItmROon4oR6/SpEHcyUX6R9x
dAaqd//Tbr8pOtBTNME24WCRrXUZQvAUsoC0a6W9RCbZMPLV+hf+01kRmQ8Se10BTe2q6F3lId/s
zv8tiYjKGyELVmTZcUd5knK1b0/PUcCaJeeVb61+lhMUK5xJ2rzX0RUDnfDN9SgOXfhu2eQtK/H2
9EUQD7gQPySzIUmGL3fq+v4GNPYy49L+kRDDXn4+hWZNMwq4tYF2rSz6F8DRR+Ln32khRffmwwlV
D5OVgYr7OhfhFkU7zyU4BRIk+mG923aiuVbXyi7zNZcY0H3mYOtDbnfLv1GapR/mOIDvlpV4bwaX
S10GfUfq6FaueFHm7GYgih3qXGhXvxn5LsEerZNpYZ9UlznEYaocfws1n2uJ3Jlzm7wAY4zx4kQI
bFUBwGkG8xNmp7giQ7KfYCyd0aFKcqimtRCINhCPIbX+Vym3kxks4S4SNVg9dNSlPmEOolRu5g2h
Fqjtxb3VmGmKSE4OrSc7nBBODWNtWVw3IrNTJ/HC7HgoR63GbGBAdcDVsDI81nOSVToc2XXKzV8F
HPLzW3EOjgZ23lgEV5Ohw/fxM9rUQ2UuUNnqaVgoxJQC+75IMhzJk8s9zLyjQvk51ymmd+5IQDDn
6l4z8Avc1fQNyz8Rl7JfMfRlLABwuucWWjI642Lws0KWA9oXdDsEjjdnl+kjXXmpFDoe8MQ3SN+R
UEGlaaAy7w3nothyMqul0wdDh1EbKEKlraNignUd3tMSSzfL3b/XxqGQyw+GCjGY8jPKzMGQWKay
l477gS+uKVQpzx9hjTtYedYWryI5mdxhOy9KoT6j5cC1Mwck75XTaQT9ZW+09dp8OfEi4Zqk67BZ
Bvd2kBli39pdQ+ut09uDkvkOlIzqPAEDA272jtehjpjMWIofczXMUUUubRHl2yU2rws5Woa9fY8J
cEC41KKeCCMwGtX158nvUSbiMzTkDTqsYHxu+sKZbs5KDqEca90NI9jsDVZtiHIDpbUfhXJgw8ZE
M5S9EmG+Ah7EKFc0u31w/JlxzRQd2u+NXAfFcLVspd6KTTPPa2Z7mnuyHe/Y18EMO/EyZ7+4+/3+
0ZgAKEJt0cE7nGcfqeaErIsACjajIyOqjCI2lk3r3kSRjxVErLq5dy6Y5johJ41wY02OAj8gJ/Qh
Bz3Wzw5e1LeRwFStt/2AZbR1N89QX96XnJ1bFoClQp5SmxxSd0YqHgk8v1OXKjaE/FwalNM3kuWA
nT2vIAG0ctyMjC4TfMMhQKchgNHhFAhGEWQvuX+/1zX38AN+UnWiwgdLktyYREdN9sjEbZLp6t/9
E1vsHShkANJ8vAH9t99gQ2eUHjhclsdnLUFzrEyy+VGyQ57tar7YW3PytFSUcUomq03KpBG7E+b6
jnjyERG/pftRTfh7rnE5IThKyC5wxXuGJr3vfsKLMGYpJeh8wDcQkXsdXmmpCMVig6V9k5TjxOBl
YoAs6d7a7rsZnf/+Anjo9qwLnFFRVrCef9UfO5y4FZ6y0LQyN1phrBJ7ly5WqvCjzRyqNJ82urOG
0KOPLHPcdprucuD+dhBJvtWSBB7X2nM0O6njmH/eMOgGtGjWvf3QlhE6aqmXxRNkGqAGoRAhhVT5
tdKTGzFsUZqa/v3AdThVeai5z4e0OgEkfRF7DYAq1DXwpi34RbMUtSPcE453VG7tN478Yd+YdvNP
Oi3duSb6Lx8HD1oBhwlfpcTj8zXY8uXRhsPw8KKKLNXWlMQU4OK4uhHZj4nbwt1cdwlhoTNI43U0
wZQA7aSyvkg39+ArpX+WtGZGlVGWNjsHlpADi6CozSymVA38X2IZjG5Um+xyUphofsLTf5DPMKzF
ESIH0Gnp4d8Pb/rMgIRSC3IkSYYz2TBnTw6TdOHPtfukcxI1wMyOtQRncnF/e//aJWymOECRbSn1
EYiJcKNyv6dcwnap4wG14/9oXGYdpwI/hK0Q6H1VquPtNi49mJhaMghY60YuMiWxWp+ZIwAmuKBB
mxaOPS4pp+W4lHpKlUNl2iWFHcJEYozaMobfoTNiqo6bXn1WJdA6TJImvql+ju9LhwNgbfhjZifh
+rh6FIuk6nfsV10JI1hC0B27Zmn07bvfRCbNnJl7rX+VkJQppNwcxMST5g8+efT106I+ecQd0EjG
ElYQqZX/tN54m9S0h6yNkkT0PPgdLlR8E9BZ2SaFikFQT7LmiNFcMNqG6/C/G96VERueOKlhe9yJ
+VwSnoEIQRotE/aJqHO5bJTMnFQxtL/wqaODMvAifXSvkGPm/89de2vzaMdE9WEySGmPoRD1nBur
bkt6xyae8ZnLsZDqsXN4dscJVbqtslVwvBvKcPDxPYSG66DHmQOCqpLuvLB6GjYfO1HRo8mJM6Ij
dWwHLnQUVoCG3i1iVuBaIhf0rH/r32H54lZH9Q5fnfftRsv4MgjyQr34NLqNIxvG0fwGSvuhJ8FX
3DNrQIexqNcFr0e4AnuyHvG3DGPC35UfxLkSFCMOaOx2NXKXlxfTL6Bk1ztbuNsGvjO/tMRQADla
5QMIFi4Ddhyjbe60GtdaLjzFs4Jxe2TZF2J7nA30ecWyuChNCVghuY1ytxvjt6rMFjEM/bSJwei2
ZzWipIbN9MhkQlnjnU9lBiKPMwOQVhAOXhVDTgylLLkPGfwTF0gBvcKW8OgXCX1J8XTCqZRkN/rx
m+gV6bDBYSuVrbYGGChvpN681Wfhen+5+N7S5qP1CgTjcsxgrBXJ1Sm86/DYXBKY7/f/GfeWL3io
m2q7qoXDeFmvC8B1eSRA0I3cI13zxcDWXai3nN2sGDRl+vT4HD0lZicTuMWIOMn/hiWGoH4HBEfC
7aw/ooHgoF9//eJXn0tM5H5qsqM9+p5hn9UzjYNuhfwEItWDxe5J7bcTwOfhOH1wI1QwMatQ6xpt
Co5bsOrrC4jzaY2xcNFtapy1hcR4OxOW3yHsk5Ufqq2bk/dZd8r/6qAFonuKH0txstr6yJnP/F8F
Mrl95LZ6RbIFxsGnrEbMXT6lM7GDYPfFiXzUBq+3Qw2c/3HXMOfOpdVn2BOnpaejzjgud+vbpOGr
PstM9Js5uEjLndPrZnyCThEjpvwZcgfjZhIrJtzlEJj24i4EOv6HZhQJvvISP25j+cBeMFnB2Hwy
m0mER6nwGfD0TZ5vpffUfQu4Y5F8mq209p4EV812VitdzNoX1SG5TDnuCnNq+YPg5mizzvOb9XHJ
XRzKcFTXIF1F0h1LKky3udzkuCHKmnZHz1yuujr+GQ8BRaJCzgIK9SxQuJSOiMi5uWoWuzcc76+y
bmtgOigKVOH1cgVXS/+2TbX4x1xkVoLc6ce75Sc94QZW4WAf8k/8XZPRGhjJ+Kd2GCy2iLVYHMUO
U8niUJbG7Jyqm1En/TfJfNRUJPXwTJq9CjQ9Aeg1TGfJZPzGmFVKrANveornD+bREvmNu4WFO+XM
uuY4gKyM6niS8iTtPnFRCPUlq7Y2oKdHh2Qa947VS/yXX8OGAFM3iqxNZXnzJ5Jrhdy73tgwxFxy
+U8aATBfXugvm7qojGX2Si7FFr4rNRcnifK17AguUjhYf2XVNQETY8PMlv1IvHlJDT0he4W7QY4u
ctOZLE+OVsiNpui84hpBkjOW2CzoxEnlg/XKcpnor0w++placfM1tvDgoupJkATAYmEdp2fX+5Fl
Cns+4lSB9oWypVFJ+P4yUVShIq6+Mvx2tjitnj9Bmu923RBZOTRS5K7dBdkN3/L8oP7jztZObOOs
HEt/OqBFhQSNXBWtrlIj9SFWZl2M0tmwCYISs+tYIok6BEee6RlgK4X/AEBRM4NSmlDWk7OGl4y/
1TbR2aVmOJaOrgF4xCG+QTFRjE1Rm2cPKMgv2sUq+bhKjyHCH0XrtGo/+6o1oGu5KHrqwHcYjlqY
5mfNCVUxaDp24vUKs3u9oRuypDBHdX8BS/oMNAL1oa0h8uQEXvyBaRjBiwqAKUpzSuObp7o+Tga5
AJHXqc5h2UCWgivXRjmBJvQKY0Dyc8DFcW3tboZSFYfFoSL74QgEBGHtXVcAxmjA8RhYUjtGzZ9n
FKLzdkgi17AkeWgk1bdZ1QIsmeOkgr6x377QSktMGGljpM6jxfeg7WJN/xhx0BKspKfgxtuBW9gs
1CjOX7nlZZmGuxuzWdcOFa+gXLB5YQy045HiLz1t68H/FRH9GiaZiraoa6sOOF32s9p7iUv6qyfL
wgpqGBqlu9XuOA/qGO2w4jKh7eDd6LLu59fs16ivT7yhpTZ86J8oQAif5jDbM165jGO/rDPsmE04
F0Egf8lx+QQzZ8sQ/gf1LN18AdsVHOGTT57naIADRJOcb4anLqncMdxAkYLjCAzsI+aqNxcB39HL
vrcMBwJxTz23lItYZgp9KboxWp8c4lFcgiGoXU3rrrWipsunQoD7UbUyIctkBW3VAL7Bvjs98ZBZ
sjYNSvRXa2B1/4lS8A1dpsso3DiTAGjDQteXtWdu0edQcdGIrEa5vLzVn5S+LOWeopybCGhT+ttj
nCJGcRKa2xWXpTx0B5H1lUKxX6k/UVtehMpD2+OmLo+slWP+32N4db0Yc93A0pvapIqDAS2MiUGu
qGaapuJDIBL85RFCmuFZ4L+2BsoEkqoqUfow8/JLCpfzWHb3RIPPnmSMHZ3OlbJsCIS52YUOdbfr
AQlKGG6JJdrF0Zeq1KmfniSoaLt4hTrRWvb/TFBBFvLztbL2ZLeZb0DpAWQeVN9PpZwzAEHnGp5d
bArV6BkrTRL4qZw0Y2jN+ZzD8wAfPuVaFgwdZRx7mhdP+fnu8BHYxp5WRj92WSlJay1g+cGAub63
U8vDTigUVg2XHXkgrc+KjXBdlGljz9L9DVrh5RBjBrhJOCQXF03pOqVn1SwCNPqIr6/tQ7WC1Zi4
jdeAqlZXbMdGLuZExQq1o3hTRD/7U37qj4XRLp9VZmUkSIA5QSdLRct8iq37hEFIBfwOTOKNSEBM
FLOT2+c3MoJr9idRG2+LSE59pRrCoTcds1rBPfVR64T83k7DnJwH6IJYj99y6LoaT+QQYaa87A1V
lm0iz6f0Xy97c7VPqxlCMWa4Dw0gvy6oYEO+U0YdMf1r76WiY32jgG0CtrKWi1c/36TysY2My6Mh
N6fafFzOdSeu+3Jymt7bOFJ5c7r6Us/YhLQEZRIpvkYYzk294+2/Jvm++TDScKXHjOOGO5qHWGo/
p4gpku8znDNaIxrTvCdVdAkQ25dvmmCaK08w8hMFvZAHl5CrX2bOC9RQ9VvDCObKPMAu8MJJ47w9
1gk9lZGidC4lG3bxJ7YHowjl3N/S6KOcGKFj7Ay7Ed3e+mygKc79sG4bE6XvmwclBAWoENNVLecG
R3LZkFt/J2XCL9HhbhbqhUluUw/QeTwR3nhVQs5zF7pyfBXJG+4LytRxf10LZ0COSVjOZHwydLJq
kCe1qOuGl1EQ7x73Wl8EfkR6ZtHOq7Om0zFwY8NpaJTkck+CPP/COnOP+EIPtbeKFh/54Y4qOx1t
Sg7KbZ66aX7DWDSEUDOtIMz5piTNTTzf1P0YCenKAEgAGn5InTVE7gVtzTQ9bq8WBJLExKB7euM5
N7vlJk08HjwU19Au+FVMixlob3m2UkTC8+8Ib3nsTlD7pmmdiIEDQMMy91AxFLtF9wL3o0vMiglF
FOcizG7KSlIzGhmSH0THUHZz5gEUeCQSRBfFLD2NRHxLrtr+AP16TnLjNsNE2ZJDQX26t3pEfdVf
uyamCywFfthiZqFE6qMWhyJDid9iHMse2R1VyEYs7h7zj5kwTi1SSUpMeUtpwwIusxj4/G9u28Hs
xNsOihEatrWFhuajv9nahWJlS3Sbu1nIx00Ys+WMKpCxdCZUvRSmmRwtcLeKycoBHsdel/FV6LaZ
5FbnVENC+7uomHyOSd+VrZkFh7h7BNrhR0cxVmNSBCscvUk5D8KG+Aw9ws/F6p70sXeFD/xxzts8
WQqfyHLXjrHIYEMQmj+uW2CAoT70ZMSiMGlAnBxSybgvA8ChvpWl/z6w4bnLJ233rlzFBFw+LNZd
Cym/mz87qzyM7o7kB+IdFXsdfLtVVTcUj4WHxWEX2887zpxZArFaMgDpciEcgA4UxPytIo0TpRo4
dJTD21q0NzWJeoIvf9mKWrM1Bk/kXMtbjItkxM6YpyFEqIY2a9c4XoA8WAW7comRNyL+jMy6D1++
XQQgwrswDyzlhuGZuKe9BWLqAb+Sd2FlxGzlHCN/1n8yQbGOr4SuATKr7CkRTbuJfnPWY9Z0u0pd
GvOljamXJy7ju7nqRbkYFQWyjfyKG/lQiFX71yYKgDN8qO879BKw3U+i9Qi1rsRZpRGHFbyoGYf7
VlUkj7Ti4eXmqtJG/ogryM04hl2Aafp1WKL3Xoic+7PaY4I+pvqVQfTbtVbchuchg4372yBz4s5a
qtzFIqF+CQ6LvL9nWuJf9l2LwoSgLgbb10bS1H/+yn8j0aa66H2FEU90VSFSFYXYQeF4YrKnK8he
ine62XzO0KUYQcnUaDe36SD+4QPzUhMrflwEbVMGVH8jYxPaFwBFQGvjTFO2zNv9JjmoCK/lAmkA
oz7MXlr3eJlSsalUxlhHuX4BRkaOLivUjxMB6dkY5DwEDyI9r+s2ZGv3RAYi0VqMEEOsFM+bwelb
cxM8WrDUfHeVGR9sJ9AvDjZ4SPbu0LNNi8WAt8Jxofp618T9i0nLD0EKZ36noQfppPjhsJz3Yl4F
QQN68FvUfeeUhf4H58zdxHgVPeNAVQc/7UJKFBzo1vURlbQIJXuewuLa8UuuFkSAieOoZXpXR0zT
ud+qPE4RFIc0B/4kEse1E43XyAMdVFc5MtIT0SMoKHAobhvDo1bHAArd9mZSpwncAzrwyXk0dfkU
6FQN+Io/pXpnhikPHUgoWt56XZ7KAqItVZEnbbGpdOYUWwD75WB/68riTxeR4eLLsjtpzPXmaZ4O
hlooLJH9FEs46LfruG0i++mgZ0AEk5UlO5OnI16Zt8r8d3/OL6ZCO+O9ne9e+iGC63I01H5+mKPD
V7lFxkdGobPGVHvi+C4sSKIPkiQ/9vOXGYfcLi09TG9aNdxyzM/RujSU3uS/aIjI7qUkbi5OWQM/
s3Zbj0UiYdvVA7QbTS+K7C7EeMV+FecKBJ0ZBs4VrpOscO2yu49TqRaM61Lv75chaSCwmA8GOT68
IbBGwNSvUjAVrDFgKGnAmBgQs7rCYNmIOrtbLswzVS/l839wxp4pje4MspLsWQ1UQvXYbPz2SnuC
NMDeKS6V2AWj5o0AU/Rl2z4nM9NHBWZeBkNxt15QZcmktSbJZZHvlwuEk2uwKCBI6VIYD8W7VtNy
jroZH+D4TOgNA8ybEjGQNhNSOkDK75lCh9KZ6wbc9Q+LnCwC13WA0r/kBfbLUhfN94UVQ4HINOaG
7aBheMCML9Jxk1OvRwqm07LToZiQbzLfX1OwjBYMMBOtXHZ0dWPnq9gp/LQTNg04jucr1CSHg9c2
gor0gjWYCsiMxSOIZK+hF8pS6k4oId5yWv2ZXlr0+ttNHXQseT10j3kALAep8QWumePQ+kxfIjWS
eu515PdBDvxLdaTbxSTtCc1QfacQjPNWF9LwQMLplF3fu4U32CTBLvdAj0v6jHAcK1ADpBu8CVh8
2L7F7eLGSn0/0wm3ghtUcL/kwJIh44G0NBjdDkpYEGpCuSXIzjnXPa+lL39znDOCX3yTz2whL4Qv
yB0efaoC+ob/VGjW3+HQoxxy4q9BAcVBQcZCbXnHglBkrJUo2UeJHOKK/Mn39QSHU+2fmeXUqMIY
vhNuFl+59eoxXbXB4Kd+ezUO2O15cGhfMJoXIPxYFI2Dat1Ow4LMgnCpch/rpesZyYGdoxw8xKTn
R21THZWeOH2YXVaGd/256uMJX5qp3gigqt+MGNonfmRaXWl3G1GKWrde7gXjE7AFLhYW/CJMFGR+
m7NJVO+CcbU6gyP/oGiKdWvUi+bgRZ1fs+tsFWLTz/ONXtIlZ1TkR3Eumrqx5QwNtmTRz4LRxpFs
RjGr4VCpozhILX9N6/vqW+CQ1LIknCWB01mStsO30oZjpdzvpiDsTq0A4hxxiQ2SRN8jW6iLQQS8
hyTScEbX5rffY982d2lZf8aO6rIXCn0uwaWut5i7cYX3Jrf0RF8u6IYEI69RvOoBwnano3PYHjqe
zIQMfaXiQ8Cx8z0uIFgb+RPrsITd8eGyEz9Kz86/XhbFvpp6+JtTaMSIklY936VAU9fllBxixMSR
+rqFo3yNrsiNhu4HppyZv56LFMdfs45dXdWls9ve4Xa1Kiqvu9KwOoyn3bAX7B1g1+jRpcqzpYc1
p6R7+xiRyfMo4spYg/6qSkLq7Ttb8SMjfB7nIpvFUDRpK4WWPi4TT2gf7xapjPTrc+uONL3RJs6F
3Nn2xXxCbEklHquPAyC8NsaqEMsw1qC6wXdaEHr2bR0dGwKWtI7I1gLuIyGo1DaeyFd2ieE3+/df
t04j4VI18YnolqW/Hc3doSCHM0zS8oBHM1VAx8B/SPMkqWr26AtJoMMn1wX+ZHNgbpL5CIbeTiyK
LA9rIEAUXZeWmg4mizZFq0rM7UsKR0ua2pYoXvkIpfqjiB9znf0A86bCLwJEvJIZk9AWnwS/e43H
ZJw22NM+fUOiHm1d6lZWV5NLy7qKe/7MIdTiRjReUb8fhgibl/06Y6rtDxtuqY7BXhH4cdhAWY2M
qFCxoB1oJeBpera4lIfXn00vHSnfm5algefT9S0PtTUk1deEABnQVnAzGYE1UgcJ6C9mufDHl0Ux
ebH287AaO3gIXhbHtSln3l2TJqhfv0DyDg/4jj1LcmgkCtvztqrNE5rJkmTp36r3PuPsl7B+ZtDw
xOIn9UesIVK3OxqpXDC5Hp+wfoMzAIm8XTC8RmZlqjGSFLP4rXRt/c4FS66j6rPK/u+HxdmkbGs8
avOB5yxhey1tGXfaUBoag3Zjei5nDTUJS7/4iw+ErZFdwtrklRkbKbZeCjvGia3uZWfMTtuWED4I
2O16h+FrKN2NBHPlI5dYdb64ugXTlU5CEG1ucfW8VdTGsUnzPItOfLzRgp0vR/R4eL7UFEHLGxX6
DGtt7vf9PSZ6BVEFdSO4mRPNTHTqk8c4XOoHw6kZgRugnyEP0rQHHub8OryUXtlyEaIlaxTMXNud
BKItV7N7zqhn0vCNc0vgPo8tgZVx3x7YWsQJZX4TLzxHXTk/xbWCjVJx6MXYIZ9Qr+XJwd6R6Coc
oSR5jjYIrbrULKGMgYLDvN53PUcm/tGBBpjVPONHO4gnpZDJbI0j3YNIyqWpkb+W2UrO8Dk5vroV
PA+XDnqPm68iepo2LfCyZbg9iy/ohOy0/MEd2i9zNDS0bckMCxEtEZgCXiQRgjazM63GfepwaFI9
/HhkW60bb4+MoCo837mS451gMV1aRxiqkN21oD1ZLQCAsASSF8XmBDkbtjZLTEVv1uy58EnKWGva
NnmsNAhrbEX8R7K4zWKQvi/VOcBbUKLi4LicSNe+BHnfMXAyB2SCaxRvekKE/qjcu0Uw1B+0X/nC
2yBdbHIb64EMvdj+5n5h4xD8AjhEsgDulSWRfaKXWitOCkD1jMgt29wF9t72wtQcI+pq0KjJvjDi
Nce8jaFPNsLNiDok7VBLEsWO86VKTmIMu4idv2Gvg4Ykh0rIpKXSwV1i7yKPANcV2wrjGOlmtl0D
ke10xOhuSb2G/Et/HzCpRIB4ApyJDd4UCdM+uYYWd9yYBjUFjU4+utMnTI7HEoYoSlQT8pOGSX2O
uUi3xzaey5geY4VX0NLv7DnKknHZ17nkcJguATiDTQcV1c3kTdZ+d4flsPGs5F3pSSZ5UJp5f/sr
zbYikEpxvr+PX2fHgGDuzHSSNZRqiGh8le9wYfpgvv+zyMbBqJIBmUX2ZWxEs5Ab8QxrwxHFvjs4
1NYonRJAw/rajWRctZKiwKeJ31ti/X4DN/FAkn8Otb+a2Yl5pZ70LPFD7i7lm2S3aoV9ba24NMt+
9P4OgecskkzFSS0XSHUHSHN+ptRKEHv1+u9oQa/BdDUkX5oGs03dav7KDQuXt0Syt2fyoGCf2dFg
CuGLNfprWUB68Yuqnqb34TKXZxe7Jw/aLXVawCJ8EOGaNNgE8Bu7QKyZbJMgJnMGI/J1DkIzn5pw
L5+e7TwiVrGy46z6BFemKnaYLwKLhGcis7i5dDFi1lkbIJzDCCLSajP0PrjgvVJHXZQNVmZOFR5T
DfAzb+UrXsSTnavrWEI1taL9pTGHbU/PRGVv8triKGPBvwlXHBcclbZmmg50FGpGJMpjAmIsnbGy
ocHFtbGUfbVCifzTK8eUdP0pfxiFiQtnbz3mR03cZJZCfGFQ+KbNV38CP1Prq5cC3xTfFw9Xs8rV
IZJRbCfPMLYijzdQ9wn8HPckScoTpEmxHRYsl/JmXeV98EnI1rurhoRkYlE+CXcGAu+ETIZTB1Vn
VXpncWA/oyqSHqjqF7nuxU7IeJLamO2C5poWxfT/0XwnofX2v4J5f8e5P3yovtt8BOKWLGtNkKdY
/mfqUKrPsBeajs5pDYvdMidSkygeCSwZBFSYaY/ruUjr6sM3WG0KpOubgt2mm0Wi9ISoTE+KJrSc
f2ysJ8AfKx6eZMi5Z8zMtoT7XdbUAcAIAV7I+fli22Yzb0AntkDF+XEa5eQwComtSOBwwsWNWU77
UdJDy3WKG2Nbd2oXZwiI76nRqMDHZ2VsalKAgzXUKGIhBacxLCUNCY4/u+BVxFN/Vkcdyky6emBZ
spd9WzjDBZBboP148zFQNxFRjPxbbn3bx0724gDDvNXrpO/NUiqFCPrwRoRkx+CZ08tseS25PkU0
PEXczpuvrAWTRW763mYiTOWuPxP41XjdKlxG+xbIVnMtrylSq8iVqqKkq9GoFGDSuJsNPsxoPw9M
ThfZI2tPqLtvNfxUpXWSCsAEIKiMOzjGd0nybsrD7dJvcWcW3Bl/GroS8AE6faEvOvD6NF+aOvva
prXn1yh8S1ccLdy5LaYPhWwFcdNsOqTg4TdLy985FYWMAzXIFoMeGDMe2aHomGUQtphO36WXqY9D
PdZB8PN80nLSw1qA9iItVt8WYrBmYiDLl9cm5E+PpsX0O0bRQ0TBho0KBMyc7e+pM2r0HQW3MklG
uIJJQxPdVLwU2gL9u77b+hJ0KjdgwowpUZ4cHkUvis3wAK9AW08ycBj4BqMGVxZ1XWgcEFqboQ3c
p6xGdH0C6wFzrBIYUZcA2XkpR4HM4gl5eDSTEjgNlQ56fLL7BdUf0ZSNtUd2L4vNYOyoGXES1YDF
qVMnQGpsohIwd5thYcFK82Fb5YJ3Ontb/a3nyBXbLgjCPRBN3fTYdhcKFnR0/tG+r/iprFBWn+f+
0/vzWmq0WYfaY0K5w7HVKwBZvxv855RclIgCHB/WDCqy4QrG77R2lJ/zgNuxPBGLJQbjZa22lDno
1uASHE9iLrwWdgslf8jX6/Dsnv3MQ3XQgVKTVDoJ084TM8IvFVuebtNJMhVql/DxaHWkN2QKoUkW
/qQLH8US0nryX2r/c2w8bnStPpTaNenyqEBC/vE7F/8oenbH8rnQ4eKkMqRbDyFdYCb3cpx7ml/A
9+Fyo+r6+XVTFzfF7x2Y+6ieHdNw2o++m92tVHd2pDZTgRrns1YG4coVzSFmtPzdJqWtcBV29OFL
1GC6BFio78MdhdnQdC0VFP45yOcBfrinQMNsqH/XuLnwWAxpHuownE3tR4NgweXB6Bie/JtJhIzi
EU5dlVhkuOTWWrVITOpaoI2zxn0D6KZjz2pdPXPWz1/iydRZesaz+M6JaqILZZKi5Tl0A4UWkBY7
abLnc0QjMmk0kXecVKHLT8NYucsaxzdr/ApHX2qDjCT8gC82XmKO6QrhwmvOU7DbxIVPtoNlmHjh
Jpc2o5sLg7Po3L/qwLJhlNSae4j/DZDlwU+IKVP5wxtizEQUnvl8Jt0StTc7VrLFJ9wBKzgwLv9N
4xBH4yyRQTLP6+GSq/BIIyzIfhe9LLSPottSo2ynYU00Oza7E5Ofw0abEzjQnqHBeyVXIV92LQEu
hKciywOpU3w9HVx7YQrKQ6WnE54glqwqcbGm3mKpgFcR9hdQeG1Q/D83SgzdhVDp+x6qs57lE/jC
rSeZPRuXD60q5G0Oyu4q7cYDyvwz0ezOpCct/tk866e7CkslJX/sTyJfSsS3osONxkx6FG5rU61l
vCZR2Jm8v7tRSqjNAzIlwgWzICXf1E43VP/suZ3y7Ft4kCC+AFv3o3bAYT0OXSF6SW94s/5vbGW6
XZevOWA2AWXg4TvViI86rpFo0Kaaxbzj6y1MUGLCTB9PO1bm82WG87uNM2kUzDs5Yc8ANjiznlu4
+dJ9SA8Jzd9pX+/lTIigAoeYIBdYsMp91hQwbKKGCaRNWH0+2qEh3LHxggOA9qgQZG3FUY1vnZYp
QKh9N1O/+kVTRAtKlat0GXbfQ480PBQrUAN7WUTG8oGDf2AKUUBuqVd1/gWq4fH8s7gn2oRJ9S0o
vMsY6ItUCYUlJ3S7CA5jMX5rRjrGyWxJkoMQi1dTZ40Sb7GMXaG0wj7xBW+HBxvOMqxydTQx6oq+
fL68zbuDfd2IrDZMSlFXk34Ew85feT6oprXOf7lyTsqeNoVElzenrfqVbTjrALh6VvnTa/pQH8mO
V+ZbGZ47Qia5fml/7PG8RrSM9ZZTqZv2WZVUQM8xJVUc+x+uevxQGfmSx7k4ERAlxT7CpCS1E7pn
PBDsXWPDEFZJTyLqpqbTRqhjV0uu4cA0m5gmTIgLerPGDtkAT5YX/8UFMK4lhZYlPjQIu7hBZECB
i5hq/Tz/PRAKOP1vOb5fVyu4LXKKU+EtnCudtW8eMbq0BlXnd9Pa7bre3GhPTNWzKFegRyX3ZEsd
C3LVOSWYJYPqHjbmyhdbAY5Dwfm/O0jH9JcuzgKLdrWm3rSoNlZ/uJI4dg2B3xkOzOC/cZw/h05g
nmAzeO5fkaxDFrk8WneG531U4bMkMuM2lydyE8tX9tEIYVNi35lzoxT4wjat0Qh7/S6HV2U24K4t
RuZGvDSL8ayYCiB0FnYzVCOuMCryEQL9W5Z4ZctOTyIZDhI79yk4YJ54zMTGglcoZT5dlDxWbhUi
YAGonmTTDptcRO0KaE6Mpob1xQQV6fC3DXNT1N+T4p1ESXEL0wnwKPlc9nAM1LDFhiEvirIY4F+l
kdxYMNuUlpptQk0KSNZPglfDBBL+2dM6TtbXLXzmRrG6myd/dFRRFy5CktiT4yXA5/CSMzcTnlrn
t1zbDI7pys2nR8VnRh/OmaEmkEsNnSfvgJo+0DZjrRcYRffdlhrXKyyzSjrxsmMkggkalV6PnrpV
YANwnZZMAJR/t+AiY/ArS26HaK/QK2KV5Qypke7J2tXb44wOLOI/V8siDChDLR+Gv+VlS/qbydfT
FUQCo37bHKFxx0Q8/jH2ru7mzlaSWilX8/+CiV276osPOHoyU6u+axGYk+eOA+/+kPJQ4/Jwd2id
FaWXemrkLZtUgkOdZ7o8zTru6iQclepXrda0rZG7n7A6bsgsaQeEzKjfLZ4toOXaS4suH4lQpiKN
0EfCE1MMkvHWkYeAoNBJHTSHRXWBBVXnfmxheiYafmb3U5mW2qIAh8i2OyKrZAkXG1VIVkuYmCjk
HUb9//vf045HXTssPwb+vmsi3p+LE7ZgFdFF1paOsOwSZAG6OdXiIU/ZIFjqBexaUfAi6aVNWwC2
fzZ9pbRA/1A6Wlz/ribx0J7FB6B6TN9rsKZji1gLMlx5nz2vHs1w1aI9qqJiZeJdhXVEsVmtEIyV
xDqKSGNMF7lHc+PqXAANYXZ4ULSgCXPVAnSx7HNcNH2xvPSj7F6D7PgALzyY9O7a/Gg9t/jflk2r
ZBro1HSq33dTVn8t3l8PtBqHF9xEOr2E2b/HQcDlZ+zetFQlIwGPwg7tOUztK68RrBdJAg/SWEsR
jHY52Xtfv8rxy316lkipcGKVY93yNxWDhrmy5VrfItfpiCh16/yHGCsZKhZoqyMix1KKxR8wVKvo
3q3Yl7hBN9EnNzzoomqWTOO/Ck4LocmMeLOVG3uPEcvc/yIEtACNJcxviFXuOYXh3UJGUQJRYzFI
tf8ghCOWJkaos9jCTzw3y+B3z/2FYUqpLc6+HgBoBkxhuQSNBr7YrGRX8HSAMXi7bCWxfFm6hVk+
1jatUd8ZA2C6WV52JXummzpk3YZPzcWZa1F+hWrTvSAE2l1S9I79ZdUfVzAw1334SkeQxWCxETKN
k2vItslr5viJe7eMb1kmmMSeslr0yMqWOq57iM0LMo8wLWohKJn1krt1ATuyHAzmx54GrTFGygqX
zr+eTIcVMQEpgaHywu9aBkNq47x+3glFjjUr1Q26mxWnTHTSS9hKqQX9oacbDqCn29eBw7NHESiC
E6vVvRcsLelsiXYAR/ye15ymcAaum1kW6UJ5a2g8wVO2DhciezXfto5O1PLR0f0t22UCD1xc/+k/
Q96Xy4XXbkp6k7J/Yy/Uuhmp70Noj9Z+qsROR+BhRtgsUiS6UtX7Uw9Yf+T86p2GTF/is8//IAC9
L7rEq3p1S8gSU/bAGH9o/v7YKT5YlMtNFoaIkPiA2jQEYGLkxpC4WiLgFxyiYreZTnBF5jYRYJNW
V4eAQP1IGAASEj4myoBB+nL19Ohe0IRlu1KbSXwZTyIRJZuW/fruCR+IGYxoYipeo2o6V64TAP8P
dT1fUR0QuaOYwFlZ43gUVB4/eOOkZ/RsLXEYN4S3LF/nFaSYtE/T9BUWBMWR0b7OhfqxuQkd1Vc2
eWgQzGBT6r5mbxKeVi+72RE9wB8054FT0otbE0YXTsO0C7/PlwcuL3KgL60zPPBsOApoc3JjlPTt
p4QMS4QO0lyMsPg/3n0/GX5Nmq8juFlz5fdHf1Y9vOTQrPyAP7sT3RdIIFvf/Wc3lmOyFbVdz2NS
8ekZvV8i/fFYFc8abmz+FAog9RVaapkAA5EoeEhnHwMcfhP1/U7ddJNweTZDGSGVXypPk2/9nwLC
rop1GSn5OMQVSUM0abLWupEscKW5ZGOt2bYrNHX81uZLoZan7c5eU2BU+HLHIl+gXR8GLnSbPlzo
o/k2e1aIwYh9M1u5+UUZ5vuzc+Im7G6niUNdmwB23XQlfyXdK54UV6M7KUW1tfs53LZSA9n84y4S
TLSVAAldO1AtYMeEGcFVTWnPCd6IEPKeXP3qZnDjhwBN5Ji0+76udEva9TKi2qIxIm1PmAxRgLn3
CDH6dgqHlYGK4c7/VaBDxc7r2eIBKXt0czFUoHZQY6FB7QIpNZJs5JUmDSo2pDvg0/NMRa9B8AqW
ZDohvokCJtRJ/db3ITwyT0b+4DdGEzFcjVuIodWhiG1zEMhO3LXvQDLJbA/cJWJ4y9Wfp+6lS2nn
l742LWxBWG3ZAK4zQWg4Qvgll4Xolonq7okj4cfieAlm/9Wz0at5I+oHh8o8tFcIevFEVXQ33eoh
jJLM13P7fTTIIRNpq6W4dNck6kVh44ioE/vCeDrAEtR7EMDKASgSvvpJeK/AKwPXl/SWPdm6By5i
R4pyhKTsjuNKn3df45v34S4O6D7W7Dv/PEDwhNd+4BYKwHAZoufhjHZJMVluDPHPgwHQPzhGzGoG
HxDcC4jLGnKwb6Ht7gyaHuI/vx6KPHpGT07JR3uHdehubmhsh/IiOBxmQJ6ecZGPw22VspolPZsd
0FcC2GxkSpQvbuxz4EnVGl3xh/PsgRHFVNvnwtpsBKFQLv43cyEykO879FPYeyjLNLjG33e/mlbr
yUWhFKAQpQwKAfukYpX4shOi1LfvVCVgYisXjgJDXYE5XRl3TlqSWoKp/rciuLaz1GHP/PWj2V9l
gSj+j7TLLwhCaqg//k9PTWxiEugzyeQISiDldkFwbljE4JqFA3r80yKvPawzEeeUGXiyWu9WucxN
buqUHDR7PYdVPp1GyPY9YCMOMNnY+64f64Hq0/Ycum8uWhyF1M3BkCkh9TN4GQwpUh0vjcvGlinr
zVe5QyedW5FnxP/LS7X8noYOoUsXNhdlYGiavImRCc9xW9hmIajZCWGXvk4IjEsePdcb67rMaf2W
EKayjAdR2K/6rEdgPwYaQL0oClxels/uJT1vVCJ7myATTWm1fed3r/NSUv9I0isCZl2yBny4GVSS
hkjn/FC44048lMr0MW6tSZXnvQlzgM9AGFvIedMOrWOBZXgNdf6R1785c9jQiBAoPHbLYW9Z9Y//
BtJRuiXsM6eiHqefeZ3vPVYF2sY0OpziClUtZfxiD/QkVevUC6/vh1XDEzUoMOBuiqXWk39SoL7N
5e6TWKoetdxwEzj54MN/WKPxOfWDpyJHXAudFN8VwMLDe5A492MrMHAVCe5NaFGmP4HLSHb6QA7P
nzl+bvZATrYVCDH7oujYzURFdo0lI/E4ENeC/slF+mo9phLzpaCk2G5UT6EXw19iHTwChd4VGxM0
JVaXqW6qHnipgHrcXxPBaZvukWF3PrBuMFYGREpVF8xoZ9C6LDdTuCQJP/FLSMoLsz+4iuFdFKc0
+3eHgvQ5vMayjwmVIPqO34d30pd4bp0bHROMEL9xAokUUycV8O59Hd/CiPoDJAXXnoQ9lVvpHAKp
Sj9BdAOIf/VDpzfcx9+Ff2QquH3KEt1raHQse9nKL+AN32CpVTaLLgRwMMKSZUG9bDTJB7Xz3/y6
pEABIROkKTMT5b5KLqONaPU1/vtev0PE5XzR99CblOkHj94YuekpK7LSiXB9fc4QfDBHm8o0yWcg
awVG8cjg2gEUFkY0OdTNpz0LQ0/8o8GBs1E/n+CSHt3YhTtfg6AS9mXNelHyuGTmPkSLNMTMBZKS
q2u86APiAjTLzu04TZQ4HBWztMrOGCghIGflDrl6CmaNrvmBPc8VZk420DrjJHSopvIDAuDjoCNe
UbfzKft7lFp9tJcUyOlHlSYrplUkISsRXwO0A5BT1CvsczVllb9OvO1XVhZFT06GWKSFFOZus5PT
oY3eLkhNR8yif3miyUoysYvw/fFxZ13SDnw28Y+VwNffvOOyQz/way/WfKj3ZevsrSZl/+UFf07U
4MkdeKbigorFN0y143r76aEW7+4Johr/Bn4VIssjaq4RdB+y2wBZdqIWMYB1ageASOljKSaqOsnc
unBssphqdTYj3NJxwQ9nOpt+AmBsm4HppHV4UuWHzxJc2bC6+yVoG0oU2HuEvTIKCekv/z80zeml
gdGOu0sV0LUhkahNvfGbe5RBjJCdwpH+yK/fhWxk0u1YJanUtRJajmVQUn5lxFCy4R3PzODpU5mv
vig7dYREed1vxogB2QjKPbFUgLCnjpBvOidbfPlZsjodNT3CyAVWsnCwONTF4l9djryp8tKFR7ih
+l6l9O03d2r5q9Shnln0a/5Gr4bCbKTtuGQgPwxFRtNryqWDYF+3Hu6tPw+RPDyN4ifWM5LTu44N
o483u4WA5x2VhyItqJ+UQFal8mhn3EhoknJn6jCYRMRB86dz/1cbKvdNDFbyjUxK88CuahWZTdBK
qTWztPxWbuyabhKDUmJtC+x3/HDEvJYCp7MkVkQMxafMJEJVhfuAPvoNx/ilPG8Fv3F0x5mQdVPt
BE5nIT1wNLrM4T5i58vK1UHw3diMFDD2ylk+VhrxlYI0reEqzuVoQpbqs+/kgJF3aFOTUOIbq3+c
2hLoZFVAfzWaLyEc/ib19bDPPBfFn/JP+Pw/kbcFPLrH64+l26z0ske8LeTdeDeeTXcercDHK9wS
zE9bRDo2zeSTfxRlNFBrD3BtrdzwlQKpaJJDQBmXEKgD0QYcfQPKkKcE7Dqzt5V2RuODGf2xs1TI
pWN72Tqo7U31KT4u4VbARObRNmneFxZBR4nf5FDot4q/9vAzM9kGch0XEQv/5Z96BxuzOjazICMZ
h6FJo4tCIzxxPmRS6zdAg5XILZaWO5CNG0kN7c2h33U11DYdmUxY8qSRpqNUW8Hc0oQpJLniHeeE
MmOojhg8CrHRN3O/FMOpQPtL3Iw3YcWZ29ePiZwfSptZsorb59IKCko6xeVP2ITCM606r92mBTjj
8IP5ddh42TGfYUoi78lMOO2Fml4nkM6zf89TKWjMgsqVN/tpTuxUB2brvtGEzN70iq/iHN+iiP+Q
M4CfZS4/1Pv0LNylHqGfGLgcFHxBWc+ifS3ElpeOQyqSzj3zebHWF80xkg7WQR9L44jVLiRts7Fg
xwBpccRHDtuLnZD6Gtnncpz3JWbJwHBb86U2LtKbt4R/q3ye9w2qJoi6CWENx5xjrbiGddtdm1y4
Tbnr8P19jmgbYvEXyZwF4WrV94htcL71CwokH6WJIN1XYHXht0tO0LT2YeVWVRdUT7Rc2scfQejL
AbpamcscsL9mHHmnzuIulBvjQls82VHbpxIG5o0CenzeTaliR7tanZ8rFuYABFL1Q6zGMjeOlFRO
72g2d6ujqW4hagyP1WlGcQ8SMhtALXMX7RdO1C8xxRtZ9sHu/hysZu4br/HLU+ge/IBLcArq1B/N
VPw5QlKIFTJqnG7fz1ztXdUWpURtCJvNeVEQFJAWC48x40xg4BdY+DB+UAF+rHQC66Q0tw1fp3eS
HP6FudfIlmVBsRf/c/DtUxnwALjBFcx7tEflTnjbeoL74rTWXVk9WuuyZVvCsdyK3lKr/6qRlIkq
HhHiGpbw5nzL70VehTj25H4JTjghUmqxPU5TXjGzvxPd8oXRkATZ9kPz+hOHmqN9hVRvqKp0R9vx
VbuhmUYdgP0pZVHdVRtv80+cIUrWxv/zFwPFKgoIPWt4oclP+h0IbgvSQyHNL0m27b7HokwOumy1
O3OKHuBF7c5ukkN+be/VT1iuKFIfD6PcAnQBHPhMuFmuZKks/m5Gd4CLtjmC7oy4g4nh9VOMOrm2
KlBwpaunGVJVNHaW2cM3My8Rj4jAo7cqXvA2RfwMh0rQ9F75c6SO/lkQxr2H2GftR82Lkz14OD1B
t7GvX74/6AGjOL3yqJhbJoZcj5ZYkY4p/MA9Q/rUtsoNKCJ0oYJfYQuGL3Tg+9GtSpNibEkYeROR
F8tzsUHp6FtQAS29CgpE6Zvc0tUd4PbZNuQvnBsLfTgxVQY7gskWjecFm0X+vg0JDAvDPMLV6ZMg
1rEe3xzt/YT7ulhQVBPyvm/gHCbAXmMufWhMOfqeIPba3mYi/oPy5zAvCVpo3zSkQWOm8uNEYBuw
PpWhJKL0loDva6MsrbBEKpEqYTOskKhnwgEFbiKOoYLFAa0D1hZxMx1Sz83wIHftubyAuqmG3zd7
8UIeLf5frxC4M2pE5wHWG+hWPINsdygMlIYge/r2naZO8hIbdrExd3WVMfyju9Wd6O3ls12xrd1I
sJlBU6omje2nci4FPVG7PvXuwWG8ike/c7FBFuKQDEvahMzmrzwbK15K21a6EieTfWl6bGkPfC8z
0arbqA+OpXJk+6agI14OvM6mTwPE6PDosFWMGm47z2zi1Ux0N4nf46NW30zTPegNUjOfTvH7D0ZR
iN06LT259oqDXDfS3w9Ln2Mj1+NBrPBxv5m5CN6t3SNoad/lFGUl1+1PoPCes5TfAqkvbeNSuh+6
7ohFNLh+9aMW5qmw19jEtbvKNCTLus0O1l/XNRTY/QqWLqvBj6L5nAykfuh8MbS1BCCZOlvzeyeV
+K/DSL14mkUiOb9D1rJRS1xgrCDQOd8+QblcQLK0GJUym4ltjrBrZ+0SprlQuMpGi1rx+BkmESJj
j67HnZJOQ2c7EnzHhT2Jcn74LNmRRLZByB3aVQ0dmW2bWUbqm61bPHdZkj/1+QRERY2s5Zr8oapq
UFXOPuYTSTI27yZHDR8DYhLG5GBDX906S/LSDqYe9xV9N+U0v374EoizAJfiJ4UxGRQ7gU/hb4Hh
Tq2GczIw2gSBQYNbWNqb/6x2TmvTPjzbqNlsOYRZwoEidkcS6U9Yc27T4ifnELSXBDJw5ECrY++e
bi9Jggv7RPfBhtg+h/DfKrAHSx7c1leL2Rem6OU4jsyabrQNbxcwvYIQ/rsD5co2eYaqM6yKs9Sr
DuqLstbvPaTirSvAGBFXiHtbV99SsBdSglr1vm6tjj7ylUiAdVjZxogoYVT8eex7U+ERrGC8TYmb
q4nyg6uyEqNMnnXdo35+apfCAa4NFLOngJCzZk7l9KfnqYsdly2u03zOARYixdEn32knK6/eZyCj
ex4H3ciFbIucl69J7/kh+sf5d9ZVFmKSVfdnujtBMa2Ckoyz/yqd9mgFjZ/rwEXILMcGMyPtnfLz
scGHkJFYHk8tg+OEnvcf3R8mGFuH8yBJ4U5B+xPtrJx4KhIt/PJPrIVkrbmgSOLIsXXg7cunBrQP
31k//x3eEeS8e9ELhF8hLnEU0qULEyPxbZ40GawwSPuI5jTpaXyDhIsvYxaYb4APByKqpaKmGQFY
TYJRfoNM67Tkv4zdzGZ9K08YUiaBUd4VeKyKwppaOElt5IIAYADvzDRSKV1/hRjvhr+YOuK3qKea
Iqgssphb4DrAU5bxI/+mVu6065A1VRNinCiqA1G83NLPDK3p3sqskL24ELrwpwVEzMkjaB/v90au
2yyHAWVEIdQsGWbvYHCPIbVVFYfWLHinKpIFz7ybTqqNz4I+5qJc2ytmGk9mSlDo0mTBnYNEi0Ix
GK1lUmu2zP2pRcs+x4E907VPLT92OmbtbcPnLMcm7lJNfqEBmRsFxsCf/ed5uir3Ny2amNALV11A
iompqeMGQ441iSsHAl8fPRMUANmv/h8DQlRTZZKFLl71PVj5Rcrze1HdqaskvCKNEhYqNV+RL2Gj
Mi1sVaCtf4dPVgYJf6gWjOYXQQTBuofgwXeyGbbrnOfJK8BfSWS4cD24euB7pOBSlOBtfeAPrHJu
DwQas5wh+InGdOuhwO/UI3LPGA7Px2BvhWuKxbqaj7WIpkprHSoeTCs+dF3grwr2nsfq3Jpore4L
Anc/SzTVlZRmNt8zDUMeKwogpOTtvRWH1ygYXTXOF3chp94yFumF4NyevvZvmFlwzIxsDrkFxfTd
MAAIM23olt/8jAKkflkNf8zXNCnic9pWVuiswxeXZyhNlif9urhcnHsr7hprZ5QT1/mO19Eue/EA
fiSr/7Ly3sU0M7zBXygU14BcEphDh1aIkPIrHRHXLrDIrNkbRDjK1smcRF5KK1e5RAfEfOQ08C8j
kNlUcrXcGfQaiGmhzYz8LXGY4qg/IGcvvi3JKwvBPVi2o94OYW9NT+XtI1dX6hf0gU5PcVO8bCew
O2PopTtHYcuVlHYchka5OILVy1blYYRQbMCsFUYKaSeJsBZSgHtvOuKyUUl49TsfzgSSgUfgkQ5R
oK02vwxb+9iKyFeqeDnEIath9Yz1hgA+dbUShduAoBMBcOz2XrwvwJNxa/Wgbc456Q5RmqBvGVzX
KMZEBQJFy3y+GTkl+D6Pq3s0seIwzZgViAQ6Q+AB5bUT44QLo/u7sYiq43rTlydGkFDNIewh7ToS
JAt5P4bqQzXnZ9phMmpDq7FEdH98e6dy6aX47KjlTkpeg1iE0KsAQbVTELDgO5XMXC9m6XV4aJI+
kEq+j9PsXRkkhjJSH1ZbOzU/nxgktSZT/CLw7BcT9Ew7AF8x5mq1OUn6ioFk8LwkrprmeeegjAmc
M+v2/gjaBt9MmD3fXq0DX2WC6UXfKKD8qM9mpd0rwF30U4YUWRCfMglPyS3kfYdXqUKXr3sCz2Z3
sOoEqZM1KalI5pR2+rGWeW5OwgoxjZuvzH86BxXMkUz198X8ye3h7Vb4g5kMQz2DVjLbZo+p+wLS
giGIrwWFtWdXtZR5zEoGpjImIUNwb4PPszUrEbZfeaWIE3NnmEkpP3GAqOpjRjuUiJymzgJ3gAJI
kmmIDyhKvjIuQ6m9kjDIZYmiVhP+12o2LW9c5y77CcANR3o1xKLIeOmpF0LulfAJRCJdyg5JH+Gt
aIUiS7/IMYyTsDQ25GAYTG1IMKDrCCm20+L/1ykgzKPE2WILryjd/KlCzikZEXIjtLAQsk1JQaID
TM02iJp+hv4+d3nL/n/lZJNy9twhExzlU9xQy3la6UAGDs/xpY+uV2iYMDN/xezyMq5VRRlkBzQY
XcXI0EULstNvVaIf70XoF7n4SnoTjfVap/3bNouwLyMcEmSaR2hQ2AZX9xoaOXIy9K6h7gURCwQ7
R1Abt47LPARShXWiTTZc57kHW8O9e0bZnzodyd01D9ddZWRkdeLX5G68g1TjTmWuP62v8DoWoev2
/xhnyWDBTpFL6A/+eTqJOHs+oS81ZOPVp56NSyDwuxXqyMCMAkpxGUHkBGPzJivQoglPxJsMq96y
d1uwHSHj2vh+34UHK9qZQe9Y8jXn3qofTJkZg0CVs8klkiobhOxoW36cr67h0b3pp85pvqu8tQ3M
ZclMxlCDqwzhLuW7rHwKPVxruCFgOa3AIyjJ/HRouHgH5HKcXmH2fxwViu0S/DL2b1A0YuxGMvng
I3MH+EQ0OQ0tfWffwtgzXaI80oJpmGz+mOU1JdS+tQrUfq2NoNeEzoIntNu1Kk7EABil3Yo3wv+f
8JmBpJOe7D+LxZzP27wD7Mirikz4b/H8eCAAVVmj4qFSJ+7k8NCzERAF/XudOazNoLpFn4QrPWKi
wgmY0ywy/nZ26QSGb3mVmIBWuJobiXLDmRp8FNLR0hbYR1Hk60idr8ozU/ISkKGqYFbRKGS3Lr3q
MBTt+r9AcPIGAAROfndfb7aqzFrrpnkST9jmBY9RrKe9K3l8ZuTmgimNTM8FLbRo4XObKuC854ax
hVNVGiGNDOJ8ovh9W82cQI3/KYHejjoGky8ND5izswkqb9YcXdxKh/ZZixdK0zV3FJhthVPvZV7r
fAjigY3MAE4YJQWLVOgp9b9koUEgTN9W9CQZTrjFKOyG2e/Yc9oKA8H3ScOU9SV2c+x5HU3yq6KN
dDMOC6wIDfahfqLUz6jUaeqE/p1XjfQinMTr0kQhQtfsd6NsQxtQ8loqvE0Y4W9+LQDLcxHYrYI8
lRGKWe3sPONmrrrvJ2R3aG0Q1caG9KXZxUexDF+KUEiNJqrdS+TzSyTm95tuPiu6csZZOPi3YGnN
eaHemGxGVASEeh5L83Pnl0cdhDa2nUTqQ4zAWXgjVRYIxgBURTB+eE72DJ6tUVF2i7+ULx5OKyrf
2yXI+mMCUQLqkWzd7qoC4TLoCXJ1+SbvpQZRQeoY0mR3dzVj3l385A6ElS4EsFVepDDLc1Y0CajD
CgCEm2AUhpREX0sITZ93WZYflhCwAZOaGSzIs8cHbYPbcVCKHBQdjYgYCTV/B2DrDTuHNXPYnl3U
v8e65s6rztWAA+APzrUkiZSuWKqPJBQvJJRg3qBxOUhSor5PbtTH7tNpzZFFd4VG94NsKwWNdOvk
ev0nqIrSYJQ6WRU0ufKsdVJzCDWMqjr59HIn7SuQRCx1uTo8NiyllHvB1XFK9/uhHby1oEc/E287
/SmHXGaS7Wg/MjW2lGw1hid4iMShTW0G4iyi27WfWlOFUUJBy0ra0ZejYQo9SrKO3QgHjwHmKmWv
GGaO+Ymh6cmDIoevftdsI8aRyNE+v7zYc2iq/Q4EXb/iqVajN92AfqHm/DBN3Sh12E5pnRbY5V89
tZCWmUjUoSjnGpnKlPbhcZ6AKhC3q5ST3GiKj2WjfYXbLI6X9rjEvlQNokCQmX0MK5n9lj6GTFrM
QkEHmcxpfKz8zbdC6GU8JbwfCfV8WnSRczjD1Mjo/g1mcAV6oIoRDu7dFDvG1juXL+K0iKWbENHo
82e8gBQCgpMMUe9B8BcsjfBhfvmSIV5ZKjxOhdCiYrlc9103DNlkIV+M5vKEaRrZPlV5O0odQNjq
FZ0waU+F79B/dzrEVQY3dNneOiL1OIUlqS7COMVbIe8E3WGxUYFyF8AW+jae2wMSOeAYGCT3Qvrg
vyV0fm+53esAYzIqRZqa5wRGw88GJd8peEzb+gzJPVlUe/aHacAnALNWBsMzrfzNidDJ2M1BQ5NN
jNUwwBzExdzQj/Dx7RdhyTP/gltMV+WULUhMCGDbr6WZXll9Lz4mFiFTp89WCpJLQpE+s7Od4RTn
Ve/h4nk7CZOwa6Hs1LrwA/aJnBT5ymb6WO64evhpHLJp86zvZGZIm6elAz3oEHVpbmpU1sSKcfWJ
adhw4gwzQBekocXskfkKnnuPv8WQ+j6vrrlua+R8LjPW0cr8YMIOO4cLWzafHX0Qh53YYzQgqvde
c2oWt4T2BLRP8XRrsuVA0eDFD4O+W5jpn/nzgu0k80lRV+DKYmy2IyMuqArUEEacSQzfeOp7C/aR
AVsayeyMJnUsY8Mke+jF5JKZipk2IXb3vGTqzcBZOkEo9fgcD37HKU0EtfUVUzcs9O7wPxYy/CFn
VN5qyr+LWR6UJ8V7/T8IsOQ1B08p6YgzKYH1RfECG/1PHy5QTTkUW1tlnN3d4Gqq/ENW+mSGnVAg
PQene4Rdd9wCRiAeZCJ4QfomgauAm9/AGdkK7h2+ae0yWQoIKGcgxiKOIah/ekh2V5wuKOvjRdod
CcV+bIS4+2f8ldXsicRPW+xuoUqYQbeaf++e74RzrMYK3DH7r+PdvFFFmWKvc9C9zJyspCJFIhrx
XlDe8uNsQqgcvTLRlQs3GdeuzJAH5Mbq7QJ9GboxUEypuSK75Stsjjqw8oCkkkNG4NhbNFtm31IL
1/8K3qJLHUcPr2EqSnYVl8ZndqcQ/2hYubkmVaBNp1Xiq0u2mi/qrhAuDy/14JxS4+fER+Xn2woR
vJVgNdorcyH/323O1zDpcOGrhk6vmiRzS8AJe6GG7gs6jjCECVvNgb1xLA0VliVJrvPnc87104LG
sXbmuCHlmLIAfSYgLOxa/dAPq0ECUlf4bVgPKUhuIuPq6SP+0kRhDotL6zgOSL8U5RegFM8Py7qA
hsiJoy4ijeOlNCOQ+T2Q3LUOASpGDZKQroU8oR3J0Q8nmHhTOnTAFozXlVo+EnDxDcIwJ95DU6KW
hqGfnVhL1s1Va/edCtnk7e864GICaxzRYdkaoVEFNJF9CGxsPFnM9NEzRUR09ge3ttA6QfzmNV/o
AiiEqbYttNEkor4yvjnlCPk4JRos/VLZIoWHiCYmCLwmK9HavOhrGVKrELdShMEHkLeugWOpHdfz
ShrcKiWL9G4IO7JstFdzdmyhSq/kt5V0xWVktxRhzMZh9azaI58Kj6PoEmI5RKyjKkB70O8D3NXY
jJFurKucPsJOdQZQWDqS0JYJh6p+ZTbwfPr7ygI3rC6Rmfknl97D45qELfh2pcFjUhwpeIWptvu5
p17LohbwYqG9qylroA6M9cGCSVtF+XmoJNrxaQI63Q1haKP4z32V3CmsbgxivG6OGta+XxbOHTwR
WV6GjewnvCqkfhPDpmQyC3J1YTkJktXCOU3sTOmi1a9jTNvgyrQVVYXFPK2IadHGL6tuEHpNR5Cv
7X54IgMfVZYT1GcOi5iueqJ/4HdK/hnNj4+SzmO+BuKlUrgncN4RcMN8XDUEi5FJtSUr0LHunk9B
A+fR7T/OahGRB/E8b1MUFPlL84Ha5IHRILTFNRC1W03XQ8MMJR1dB4vAkJ5XQTgyG1vEbF5rbYed
hIa+8d8wqVMhmyRFY90LEPyTtqOzkSVcyuA7T1rc9xTQIK1nYQ4RgtwDmHgYDFNj+CBFI5mqZW9c
twfOAqYdrQeKLqpDuc9Srl+vt4SQS3nh6S2EzQOknXISMa/+Z6Ryqz7uLJ6SCxt7QJMkjt5EqGRI
d3Z6UjJnyPiXmZtVEdnAhMUdVzpmY/w/+VaCdY2o+tKkqGhsrTgRbcUhYRE7BqvzRNup+o81qeZs
skOaSS5uFaToe1OdZ4xi2LEpjdnP3O4vL1fZ1odydjqfUM9i1uQAeOBaXhkGN82BTpiEjRkJzCg5
tYuZiHJbz1Cvz9SM74LAgbYYY3uNZi7neol0PvXzOc8PL4mpQx4M5/4vI+q237Wj4vbfN67A+9sH
WN2vOl0unqRTWqgoxmk4uppJLB2WMn+d6GmmMir18bgXWrPVrDdR/lnmNF/eIEQh9brflmDF9mTN
bSPV9koB1/Y6Wy+9SEgjuR4tsY6/yFn34PoJHOqnta3Zl/r7W9JmTXWZE0UDLz3SugNn6bBFN9Lv
a2WnFtII0mA0UDJws/L/z7aeXawOrtft7EcetKzAxNB00E2UPk4tw7NhN7kQT/kmN+lOQoTa609Z
awJN7HI0H1Cnse6EEfb96qm6Y4HclRwDGe1HbvgoevLcPADeTN6iiRk+UYbOs4tPmMOz7aG2Nh/m
vna57pLpvEmPggDJhC27ukUs7SPaj5K8rdZFnea/CfMR39OO+I5oFk6lCutZQMkP34elnvjw8EmH
g1simTtTQ/5KeKw+6QwqgT7QLMAlKXp6XgaFlRDukyAPDrwwo1NA+UyT+RjwapsDz/6tRfdG14v7
Q6aHbsuFB2jcndyYL2XLdn6OqfwlAlx0X0+dcl+Njk6dVeJLNt3DA5BCKhigaXu5jldNvfWr6gSU
Fo+NoHxFspI5IqbqqNwaXZK33dh2HoHVSAc1mrS0aZIUv8QkvUG1YsKkUwLYJpdnAMnfJHWhRun4
Z26LdxDXIVGy3T3Gl25J1+kKxd9u9zqR4946Rxg0rgpIS7YpWfHqNx8RvuAK+YZg26gLGFk5DThJ
gdsterO2GBxY6hULJjTrx/VL0IMmRoe6weCMEru05foZiNRFYh9K6LsmSroksnr99YNi84RwG2ZU
eMSAsDc139OUnyivmjH8E6t2efVBpK3DE34xhv9qFLxUyH3Fe6Z73081RhzQzAsGW2Au22qgv/Mf
etYl5oG1T78KgyJS6BKZo2pYalG4DcHSgPgAovdgv8xjvuKPCqt1WzkX/3j7CTJUDID7ilUni7J4
9OOyRAOfhpvOZeNyCbdqvUq4MEsDdTnbNpIzvkKHXhbz0Zl6Tsr8GVxhN3uijn+k+bfEQUuilNeF
vEuCGtFPVPIL+KacH+Ju0B9O5xZvlsh7TMqBDwq5NBlE6EMbteFkJ5zUbgH0QP2iuyahy4pEnBwe
sqgXSiDjTM1gNG5mfRmpTLBRkM7hCb085H5Kar9N1T5yq5vgXFWqI6OQLmu+Wm8hC4PXnD4n7C88
jAvRYGn22w4A66/TDF07e8XvlZucdeRDbIPrCHBAL3iS395MBK0HpoiO6mFmUpuC62jsCiCFImOz
lDpYjSIQkZR6qJwazq9UuW2LjsGNcU5URab/kzS3J/+4ihUaOLWFhb6XOMJOH380uYBJ53T+FBds
Es6JGbWSI713m48DRagDNszsitOW3v3GDuXkdo/T6QTNQq1URAb4NJzSBRqstfiCAIou4SDw5uGY
J5VGhvraMsn+juGR51FoSdbJGHhGT6saPALgITAm3RWKgBu/WeBdwP23BLCFgtwOmUVqHA/Z7mol
2nxhr2iYQ4Rqqi5n6gH01yneq9ar6lYahXWBMuHPJ5X0vIOhtmna3P/t0LsJRMZQm1GMR7wuSEE1
ZP8JekeMRa9tP5eQ1T97/h59N7Y2TH/3KbWsGlRNyqT9ekOrkEcJaO5ZltxWV5ukEO0D8+I638Ds
vohPo1OJsawac84p/XL+0+Irjkc/YEYgUKYYJP0yjcdxUPFunV+2KwwOKqLxToJ2qBg1kjuiQ6Lb
2GVZibiTWNf8RYc0fBVGIIv97jRkopu7OWrp/UhgfgfSa169k+Xs0XwAyjxzkZnnYQbr6meVxFTJ
Dh0HAa1eHJxB7GRsUyzFJNb6Co/LJp09x2+jJs9gJAk+WVwtJBePlHsHUTgwWJPsIinWC2cPkFXc
RYLhKVYMlSlmGpBjrmKcaL/+Z/rgUy5F45hXL3HFQ1PdjP/RtCpaZLuDt10XofkR2bIRuWJg+3QN
uMPzqplkroW5JnOZvvKSavAS2fEu2MTe8NopGULjKBC2FzyI/Xbp9xTWLDdW+7aNh35z32kQDaQR
/yAmkI/k3NgJTm9I50DmaJS4fygUVPREH0RNb/bwL0RR3YPT9EIDxO1YR2pZj/0/78rELcRREGYJ
refHdzI7wPtmGi6hjNGdjfRxMn/WVBshvP5BxsSdzNM6R0S4783ealGuvL+PtUYKDkJ4aHgL4r1x
3eGuUWQjIgsbV24FHO9iJwPt5iecPYTbGx1QBopF9KrHpmm8QqkKbqRKPlKCAI+IgPZTQkt5lppo
lgDixdv8EqxMSMljNolaQWev7abApmW6wIYhHkJUxaFECn98v4zFcbjKCrDVJ274LQbAQjEMS/mc
uPwLOFTi23GwvjLJVKsoPencrW+BrKvfw9oVZV5kPxZkrVYkA9+etABYgEbItLvfjnR+wmgugITj
4vEKk5zbO4J6RFj4lWyxK1OosvK9xsTEAyxPVncLHkHF6Z7QaxX0mVdN2KeKMu3Sp0ZdNK8DKEJv
w0jlAkfiJU3yyACnlL1tPT+Ryc1m9dDt2AKw/tWy+/PtgIIZKYD37slgnQ0Ot/C2MJwKrRYgO713
zt5GqT+0u9r5afxQKQ/NBOfIpyECgoORMc1zGZVTzcUFQ1lggNWjvwWUsnQ9aiNr0cch7Ush3eCs
F/oIi1WOOpSF0q0xLbLr+Y52NWIu1lwSH4v5lPvRqAn3qPUBuPpgXaGtRrLzXw7OlsVuUCRa99Kv
fY3X6aOdevJd646tHzSJRu7u4DnyxQ+mxhd7HbZ2qScUjQLGnQUzAEa9O+bly8Hf+tiwczHVnf0a
V+Yh8fy4b364TWi0lPAwthlb7kESvG6DD0S7YqfVi/sNqeKhUx+EQwBiTL4Ospr1ZuuaehrbIteW
BxiDQCDzaCrbPi2FhamqIY0nRglPV3BizCcsvslIK4CM49kkqvN4Ou9Q6K4WrxuKLFbMVCb/qBlo
7sSW/ph3+kIF3odKUYw2KASzwcANV1X7VlUpWysxD4hDqccAVT3GRV6ilXXzvme1h+hIFzQfsEPb
FF68KeaHY3ejH6SVQ7kjWwhhVe3m5wxBLwi2HKid7cR7GyL1urtpBM5HXJD3pteltaX4ceSXdZzP
ksI7ODFtlXcF9rAg+an6/CP6ZBQJmcyMQR9AmJLir71SE4nfQKS4h4Kbjgspl6PSlKndDEeAvnl7
JhB69a6i5NJevfx59EcKQyoBcLeXjIezeECEdoFIVXNdRpxfvL1LGb/Q7AmcFgbl6/TL/SrPEuZe
ZimcJNtDKi84ZM3TwH3cCboZL5x3KIUwE9OOc8rAUGMfT+ZUAJXps2FAIVa7tM6EtkLlap1GbDjH
M0rvLLmEDGFdBLjVyF4/vuNYzi3IiV2p6f5tw0l8x6nll7Zpj5yg5daGFUoytcbUhZ1L1ifZCgc2
caYy1/YBNq39J+hanv2uDm48GUMwLZXTyKKvQ+/JMGHpv7PBaSv+qzfNN5+pMlzdsU4wYQjjWVFr
Qhty90QtfkGn1czzen6WpJX+oh86jabqKiQoITFg24lI5gop4HX1WbWrno1ln4jhx9Z+/1NT/EX9
NJW140UKJBsbGdvychOA2qwG0pAWj2Kb1bEkl8LNYUhcYb+EtXEsrx8c++0Iu4STmEA8r4zmVZGs
iPJAJJ4tm6NYKUvjvdDS8B67JDzMYCVYvhC0WeEg6BadHB9uXYG6J891q0lh/3KW1HQtGKp3HHPG
NrCufzIs6PlxCftbVVKhrYMOq9RKbyzTirpnsG5kfCSOzW9QVS6Z8weXNXYwyOG6TLdT1M/VHNWq
yKcDI/Kzfg7+kYsoaz45vL4sEH9o/9z4Rap2u+b/DSkE1n4PngFZMs0JgaoS2mhLJyev/VXnERnX
51BLi/FYa0R8GvIhmVFP9fDGk5E2yR5yIPyqt+oIKnWwHoF3vSjBfryrJcyrsf9IEA/7nzjbr3/4
WHCBCrnTcXvqzgepK1eP6P8WFkYUtWzBoW7aVCe/IyB4JAX1RYm+/bXKJc/ad1Ic3Zqi2olnXHdc
iwCf1rZWTwEyqps/APtkg+50r04t2qBylcMIodQ944P4rVvIKlLPPeL9R0TpZdeoHBwuohyOxTbr
y6Twx+J37SzT4H/xuE685RpNtIiisB01Xh+cqlNEh+FqJd5hp5rmSyug3+fsOJZgNl0Ue+bhvG+4
XIxU4S5ixUz83/gEpxptqo1mxK6pEHpLRe131J+nYB6eyQCtxDELcxv3GnOfVa3oERtlwZ9vAmhl
ZXm2rw7e3tBaIEolbXL22n0iShAZ4NniMRXCbSV8WMm8hF/U+sDIJXnziv5HGasV8UdXt2Fr2X7A
wkWXxzelzeyyVl8Q17nK0se2qD4RhccQFcM3j5nwtzJRT4b451/wjq8Ydx6RhwFn9y1t5vW67k3q
wmERukxE297g/THvvXenHr4cT3eqpm4JgosClwMjKlHJskccdzNBf/ddrRjx+FtHvqtpW1bFnJOz
RDyrBUTpn3uO3+55XXYBWh3GKzAiHXmRJUf2yAZ8P0+m3M2AKQp+LGqaCYeone/G4EVZdtK8zJmi
IQh1+SaYyH3J27XomMY5bHUkDT21M5WGzhHk7OBfVNV7rOH8Te21JTXnnX4sNcr5xJKDkCHDI8+d
vFw7iiBqOuFee5NpsYxJWESw4zqgBsGWyveyITkGBqILYoOwkATzMdUuIrChknRNkNff2E0YDrOQ
f8jsCyeiWLe+UeAC78Dv9C9T37d4zoBD//VfzkDD1NZ6pXssBRDFJQsAqrXr3NqC02NxIfDrxie7
ERA04zMfG/fPe1sI5oYtFRnKDKg04RyJOildWoslNJcf2uSAeuYrp/5nr9P0l5C4mIu0qf3k/MuP
53FDElUgnM8QIOv3LXLYIAI8NP1X30nG2ROVTetR81pCqQKMwLq9k1qm5ehopT4Fhdxvmj9D/jGb
NVGJ1pOTtCvWd7ohIRkmmPApbe9uIxMsJb+dMmMtYthZAIBrgDMBxT0mY0Q6G86ABzHyTnhU0tOz
x+zl3CF1TGUL2T2g9ejCeUB6PLcl+fnJ7gnvBCev7JNkhKUApc+dpjsq3S93i5drJZQyNJE6+qrD
xBnlM/x5TH6eJYMdHvD7vlhATThHwTlvXbXHUn+SZjO6+nm3Jx9UNhbUEcUDtvW2byeV0dBCnsSo
X7P4vc4csraw39BeHC8LO5x9qrMzst7sAibwnXIk94Dy0zYNnaWwxuLo65ZpBoHUkRGNV266CUk5
LpRAjut3SRxvo/flGnqN3d2/emB1ETsdhyy8wQLsDtkCgdRYtZMpwnbvReW0nH53R8rPCHtr4rIZ
RR8kOTVdeSZq8fbCQNerVSxZcX6rKwy5j9S1ZBm2ipxB3fV1JV696Nqfx2R7xd/SxlphjNjBGGhh
4qTa1gxoQil8z1pk2+M8T6w6rCuTkSyoQzJjUANx/xzO8hOG11oNzKGzk8gFRHJMW8/aQQe0SWcE
rkWeIBYdFxdhT1zOaTZWTRB6fwqOueSu0/YAbcsiCBJLFO1Kh96u4WUXqAd8srDhLjFNW3jJHzcg
UUi/5eba1IAZYjFOghLZ8MPjJRhH+cb+2iHQQFe2Nw9hcnu9Kav7oi6IuO9Bs0XYhXkk7sBZehtR
e8Suv7NOv7tRAkXzZiiyVbnnCkLGdnb8GouBocO+HEDEhYQyden1PAph3+5Y074sDgfVz28kBOd8
VVVFW/OFuJT6BC5VtTKI7bclMc9TIZ49sd4R3e+n3wiw6e6WorKT+pIfw8WbydslarAt06NtqjmM
23XxyymE/aTgyfCkgJ+T8RVjvo0noxSbJOWJm91SGu5yUzuzxRWSWJaHqO6iBhFZjQ9C538eXReZ
zeep+YnRTbJD/K03sYeQUAPjMRRYFfhcZ5pA57cQlwiLGXjlP0U6HpECrrA5ytUFNUwggga1o5Xi
oK6tMNCu0P3E8mRfBpazAm7dAT1XYyz1nxk6PwSqrBSkybAsoBL8KLv5vpYpbPYdtdzZ6YjSZyn3
knGO+Dd3H7cxPk2VYwmEwgmkhJboZ4q9OOFjFW8MgxAEewXkM7mouQudpxDo9Ts8iF9K6xnPFbox
omUHQXV2nO5aWvCRMn4RDVZHduoXwgesTIaeAUnn6FMbXVYE6CUS0ECJkeW1weARZMPjj6GEFtD3
Tfugx8WgiYIVxtCVUjkuRBhOplhmOHoyhRt/VdE1w/IhwsE4onyF0CwxGVudh7TvrOd5mQLISXdX
eCtWs/jnGV1BqCltMtaxFFcUwVUc+CkKBDqpX8LRWEMOf2uJpQN0utfz27HfUK8FjnEFBWDl+Fqt
FfBLUWSroyOtm67G9Yp3wJABYUY0HRauh0lT6As0G1JimsASh3TrpqVobEDIVDYTRnAAFrF1m0t9
gwZ6uJSg8TtdImkay+h4oqmFdSFK/F9rez6rK0n5aOs3nQV5S87xekjnReNXR5KRckqxLAySIyf6
oOn1inDV2hxjBxLLfzvnWFpi2cNsEAHPuwp05Dr1+rfVSBM/NWjQWH55SdlI38kQSpUrTqCsQjCF
SUQgrDMu6e8wqnjm8bioKVtAfuseqB3akO6p5x42OGh9j+YGiLrIvE1+J7+K2PCkPq1u4p/1LICY
EMVsYA8+KWOBFgmlOGlxhTc1ZRUvW2jQBfYXfmcBEXQ+WMTV3MDT2oLY6DGHs36ca3PfUjRSW+WV
qUKYXoy1knGVvjz875fPR2qsKGRLhpsX1J5pvMokULxgkXj/9Wxb5twi7azwEnJPeymSOyaTlneK
9tsJwjWwy+RxqiKtN/OtHRdXDwFAOsPy2BxSqZx3t7WnE00f3QcXudh4yiR308bkweJitOujAfYC
45ZXtoipZAfdoQm+TmDCuiDKSfggfNQwImdtuUa+wR7X3yCJzrCS0Tm746HUfr9vJ/0kJxBoGdbG
mWm8mzY4yHBKx9AybxufgP6cGTL+eyXC5mwIE6njdEzSp5/c5g3IVj9h5TxbVy3e9jd+kw4v8JPD
XvYe8Hmo4PVnB8H5C8AdsVlYxCn7xbdewIcYTDdHRRCHyZgbbefJbipTBHxmHAHyFX0aa3TYJH3C
lh0oT9KKmqRqsYb6V7ZlzSoGE3wRiSaHYBGU4NALU9sC1BY42zApsCSDTlh+z9bdZ32eLR751HTx
D/7Yr3Qa6GOeoKn4C28gnXmoHEdjDvL+lQwLdlQwZVRFzoTYItknV3NAFpakfb9TmM+E8veVubFm
PCautjhrd35Ru2VJvvD0v0O8vZYRC9XqJev5Qd5r2KvINKzo6nRU4fvsc/IcHVFS9VtuWj3v67wm
YdWeYlvs+D51PK69jJgHfUi/hfRu77FqxIHtn+nD3XzmlHtjQK1ILvlCJFeQsqi2hv7r4tJylUdO
to34YbqWjcuXXXpOqRLNAyfTj+WYdam19fp28MKwQ/iXyDJHrzmWPRbKGusdWp9Xywm4iaqesXTs
keaYNgVs9wE/lRHBG46z772JJRmI6sObdrPp4ZcknWtnICD+fhjOfSbumeAEw49kUm4GP3UifU9L
a8J6PJen90FZE1ZiPd9X7M6ooGkuKvFuyDl82wcr9KxlO4Lu7A9XaIdEQk41Qb9yux9f3BIESpse
Aft1JxqKxL6YIij4XCvGCCvDLXfHE4fiLKBofAL7pRuH1v5jEpCljt17T8hmfH0t+TJKglNaZ6VC
e/f1ct/U/iQirc2lQKnCKNOCQkK2WcuSBNUY1GWfZB0+puwvpPoghEC+1yTDl5svAV9uAk9Re3c0
s/PvGvByYJSMJ4a0lxVQLDZJ/WRM2IrHdFe3lVNcHg3pzIOMrsjSTq5j5qugFI1t++uXXgtuIg6d
Von8q7dBT5RUB9aQ1Zv5CWPNBZIcxj28JqIqGdUFadCulYhVViX95u1tpiNAfF8cKZobw2ybh24a
9KqCyvlVh8NJMEuxHKtj9a4JhuVgig29IAYLbzHccx5UNgUp/S4eer7pexYJXXtIHGbbGEMHS6xt
TMuFIDQXCWiF5sqtJLa1OQioTDt0kmgR+skkXs8peV2fhDJXRJ1HZoyCfFwKFTDri7wfKs5pJ7uo
Auo3RiACwbn84eabe6fdjIRlljyRrGNlw1/Q/Rpk86vy8QOP7KqmPEzQcMJ8WYic7pxJINAOxYkS
ew+FA1rkxme/getqj51JsJsTFfO2f/TtFe5DG2iidhwI+7Sk+uGAOfNugOyy9uVm4OMf6fofkx2V
trcO8UzxhjydKjy9sqOK2zT2kmOqnRoW1H5S/7OcJCAhYU/3diqId/pp33y83+nNgrHqRlHVG9ld
m6yZ1TYYv7cAkpQRuPc2ecZ/zIDaSMrWaST9G4a6rJ4j9T3jozu3lybgRxds9qMLwywWt6J4MiHG
7DRuL5AD+E8Gft9WO7azGW+lM9XHDulAJzQjhSi68uvPysmJW+ysgeYby3DmPmpGGeeCmjZh1ECO
Cx6RwDxiXmfUq//uIkSFlxQluMVwXVNKJuBVhYvbbnGnQ8O08nP4jvy0i/LaS+znPWqN/DzJYgQL
Y7KYLQbPw8WQtjn4PjunRafuHGt4YyNDwugJGsuMnJXasIwFMHwSBfBG6rE9B4ShIFTY+tY1HGeC
mGf9qTIs+TyuTesc+/Nh1txgyHZGUd6/KTw3j87MKUZZSMCqDqhspLHeeT2pwMsi+fyV2sK9EPty
n7UhSJW1TEuBz2mojPYEY66vtKgIIibd2ezCsoka+c/dTBqIqcnO6RP0FubFyCXGwtbreaxsxijp
Fxg41JdqypO4DUNlaI/lt9pFDz6GCER+QFtgIuuXLNdHgqlI4IG7McA6n6Eydm/aKSt56yYzKn0C
kj+X14fxEGrPIx1nVYvnhPfYxaIOwWNxV65KhNRPbsbPiq0Uqo5M9687oYPHkC9v6SwrJ0Je1GKO
FWCSoC0oMQRubzpBHurNFC7Sn5m/afVU12+wRp1LoK2+5kvwC5CVn/idE0XhRqTXUOQkRrk/37k6
g4q/wVah+rLYR/EvDNw9chlMk9b2qLr9xu2KSn6MPImqkkiscNBngoHvSzyH7Li8Gvdt8bsKztjW
BPJudLydXrJPw3lzMzTYr+iKLPhWsMELb52+9kPo1kjy6Kxr1aRZm2c7v3DL2WGxWIjeQrX4jN6e
oeT1x3jENlZ4JymgfDRHG1e/JIsUpFVHlzZXvDbeW2//xD7L2vLQjEsL6iW6Hq70crvLqa4/HxPW
RECktSswBRYsFjqcVEfd5mFFQbAxqIq41OMYAT/9Y1RMXRIzSK/1a2JKodKnlFhiXz/3VO2zE13b
9kbQ81WrX5FVqWQg0KYu7pjriA8IB0awBj6iRQTpcjHJeYGomog4UBD798dTwbxzFMrIljJoeMbD
88/CCAyU5YB6O+zzLjBwaeyfY/cYmz3aQY25VIauU8rz5+66Z1rnULb8pYO+ayr18VO/fRWgQhRU
RNQTMmdxJbTKPZ1TCrexQqwtXf9Rp/pMO6GPVz+bjiRPJ9hPhjwnhe1MSCOUn/KLAOa+rbx+I+Mi
yEgP6HGBVT/c5nWsouICr6jep/LAkR3ugOnwr2A6rQYLjZv8pW67m/3vTTlnWIFqC51PjVCuAoW/
nJHOOabeG/RSyHsHQWUbT2BQMzOtPYIu5whiwCgOChiZgheN200DAMPUIfAhoqUlOJer81PBUmc9
Z8CeKpoVQb/jlkPyoB6wwnOGsTtD5gKxtNbwU6NjNui0yeUBUOuhj+g+o54xpojRVrNMWjQdzWVQ
e5zCS16PZlL8Gh88y2UntUcnfzYfsYFDnt8Q1vIMdcWBoblS8HmACya8ioHXdmsBI0BEyCIWbDhW
qpziiz8rdcBt4WGCP5lqKQhiIStCbqny5SOqolJ0bMaM15KCn7Jn7iKKpgE1ST9gQEjrO+BeGLKU
qbmkGC4jFqX8UPajLosWeVgeInn6vV3OC9tLwE/aKw6E+BAtbHSdtmr0x4PsAKzxSYdTiJ6+3fV2
VVOqE95CyuJKRsGeADLAbrMliVrMJk4kJ0Z141Or9cNQZyO8fMtbjMJkJTaEVLi4YPdG0Z8v8fRr
CI0F7Z7n5koUJanzLUd/Q1Hps2iqYFkF3XPTdG5YW5+SZdeLBYodQlHjt8B83ZsnpwE1Z5ikwXVt
tYa8dPJolVXFcL3HbUWN2O940Tx9CvCtN2L4CGtEe6JN0AEhuTyOYhfzeiXCDUQWJlRLX8XdIVKN
9yOlumzYNwquzh7vK+cZCcVr8ZF6nPbC/RQOR8yvBwpOIGiWOl7uh6WdGAuPgUxSzPvWEJHeQtS9
v3cPP7uP8kEIwqswWvoaMIrCv7/qWYRTCZt/HYzHqhBtLNLwG2vCOxW4GPZg7EwT/myJCYkExhjV
BH9+2Q7Zk+umSNaSgnC5sHg0yyZtlY60Lj9J99WXw0kMcZou+mYWAlSEIZsjMVjlqs85tfH6XAV0
LJt/95d2ANHO/OfH5rBP8MmzvGGT4D7Qll/SxuBTZp7woIsb9TJrX6nA95KeHBnTH2OCW4e/GJ1B
/8Z2KfPVcqiOQc66mKgRPCtMK5MqZb50JQOWJjusQ/3DXJO8C5aYeSC4yKZ3+JU6lkdtX8oBUzUP
01aX2PzZ9jKIlaRS/vkN794onsDKwBWU2Tcug2S5koVg0wFuiZlN6faIZSAQ/3wJEhhSWoEyzud1
ZAvB8cUw93SWIkI6ciyiePz5SlZpXhTmNLbZRLClvOr5Z0l1/zCFw+z0Zo3gi5PNd2YpXJr5Yr+t
0wTqWIiWnlZjPCHL8h75QsQnO84t6OInk1vrUsxiKdbNCc6R2UzS0NWtjTxCZrs3KHZBPzkO2KLK
fnk1qnpDU4G6xNAnFG1PW2L/EjZk1VN+6BGzT9ylJ17g7n5Ut0mzHH5bhojCsXnrDzghcE8Q8F9O
8OOa1/zZKYd0zrvcfojEUNXnb5oky6HhKLfV88bh+iHOtLb0MRdcnyWeIslA1WNLny5SNBTcQ6Nv
wJjjTz42cFvOLIjQ7VGMDi0R6NCbTfS16YkkVu9OIoDKYKDykoTNFuOpSA6n/h+XljjbPyWp5dkM
uQQbZvemntsvibbevRAm472ogZGdy44aq9RH8EWFi0KeHUyaw8WcINebaY24GmB+imWJSsaoJQlb
zfqPoWp9Y3F37RcMc8paw8C40/bY/LiyDC0aL9Tuff9OikNPe/I3sr0TLAHzm+gvWOdKo/18nByT
xj5oxndZSVRvv2JH61fK/9t1lD0yDIv2Z6eSMDSRje0LIqxoaM8Vj4yn/pUHqHOKe5D3IZ37Xpkj
htyfVsqDOVdwjiF+YaTfkm+QZ9aHzRVXdQfTLFIiOXts9qiD2dFFy+hyEy6nW82jbOXC9unUG4af
GvHWtMCkOk39uc+kGd85iqPnXZSZmy5nAI33xmCtr23aU7BhO3guttZHw2Ym1D2KCXarbKN3JE/U
okTTshNW5oK5mByVgZ+IYWY9pbRvD6I/yJ7U3m1jcyW5skuj2RVVWLmPnCeNyQ6RLPPGyH5gFHMz
CCoJI3ME8upKIvzxM7AJ6aLlOXuNxOCN6G2XT/8LZETkU7tcq3GvFXvHEFQzlY2V7lRyfE4MS9tm
hOACxR595NDxom3r+RGZMYtfad5fwJtzQr1RtBBAGntAXKdu+JX52a8bCNnjpqIvK4ITCG3iXGjD
gxOlLDQh9I0lPfgqFfLDQj5I3mV41AVMwCw0rxUALxMuDxH4B1D2RVzSz7ZHRt2fz0fNmowsk+MV
oc+OkYTP0CHaGd0PDUnl+lPebolTk2r0yrU68GKd5nGvfbkyFjjqZgRfOkItBjUudtslINaWX3HB
JAGVxtnhumg6lCkub8J0umQglCO4+dMueeLM2xi7xMcZCmZJPZBNU/GE5o4J0/kVLjWLSE31qMge
lTod4CphCQLNMv3Enz9jXfHEVCy2oALuxy3YIpsF/wCa/BRpG0h4SQcyzdJDCWMTpNtEFkih4gQx
TZhV/4IiuIGz+pbWzcc9Y/IPqtRXp5cnT/kptbBDQiTVjTH83qK3sEE17wqfDcwXB9Xv3T0qfV7w
jHt5NuV+HDemPPVTDtVKv/SpVaR/CD8rfqK50j38vkeMOZgZdJdmgr7Rs2IACcwHDQSObTetKiDL
O8jJoQX4HUxIWsiwIJHnq8WL+2tpopSn2rXrqh98VHOYHJdVWJDGXnVAR0p3rvzHtwqZd0Y5VmFR
hf3e0tB77aOJAJbkCu8LbZiCtt7bx1kjazVaIoLWKrjqOZuWOwcQUImYvvmEHfYHLeh7YYUTMgI9
5pjKzsMl3EXAnz8zFUH73jqncUt35PLIghEoOL40L729adzfCDI6QYryA8+n3AXDNijXf0HBwdas
FUxQwOVl8a69mS95CIueyNFurzh9420MLQgJC1yVqPgHaAwATFJnK9GmN0bCSDZQ+zOMlu2m13wD
EVYxKLi3HRh3cEZVZmhFM7pGPJU0booxxefhijuZm6HMQvdyCAQt4mDTje/5xwLgKAHyGW1g1j7e
Io3m3fdteZfKzDUEm+hNtAlF4OxVrs2K7wDrKFab51riyb19IVbhOu0mNc26bi4IJEwgseF1rr9Y
4nhUg5qyNHCSoAtnTZR6wqJsSdO+wDJMr5YKxzqGhNsKTdjgBeU+jd4UV8HiAxljaBWp6WLBDSGY
gmGm/cfreSpcQV49RFrW24e7IT7wjtNpUEale735gK7Nu/weOWx0GENbJvV/SvMmx/SccrnXcME2
J93y2nyYQELO0ikOSGjqzThbBPVSOpgfbWT85I/iiUUNcSttiuew6xluqK+DWp++lrJcIysNwuZN
bTMyNDUpWgdYp1Dj/DrTSk9anWb53jHVoQ9zHA+/IUJm0p1lE9p7VTP5VaiAW8fUkzGr/8MZr0I3
Y+8BciI1VinIzxSGcO/MRJymNOoGk0EmM2sp+C+Ui14GL2k9m4x+YiHAY6A8Kr9I6ND+L/sfrnas
wuG76dkxbtVbfTJ4LGZnTttLv7EqYEVfVWVIUZhWb9JrY1sQn84YlxGoqDPCJm6PVX8z3bOST31c
1urS5/yIaKh25YwrolHTUZDVTDY7b07AjlHgrVJWLPzsW3Law1niNtWO4oInDXXofORAtRJ8Yt+D
cEx3tJC97rw9ISHFPY7qjDyzAIc4zLVLfluTbboF0SpYe6kprswu5/ZgiduFS1fXupmtXJe6fpms
HaVn9nzysmbpNd2ZRqqxv6q1sJfpUFT37IgBGS88Pb4umFwOnVBy3PVWnbhvtVTBoAK9ksYf7VhF
z9yC+gMsXBWCn0+PrEL0LaharNIMu7l7Pmpytewlnod5h5qKbzhXdrUEAJp9WWEt1h0BWY43Smut
jv4m9gcLVwAA2yoUvaO9BYq7WECvjmnutSh69E9q5zdCWjTYe6NgIppeBft7N+6tnmeSGJTR8LSP
SIMuqazHjEND0Tb7dbVtg/ym5gT/PJmhpR/L6KRDDp5KvXn3/8E6SMBtQMMAShtVhoD6rqVnpcC1
1NDv1xRHpb02r9216vcgmN89kEQwX6W3PqfHay4kRPzvBDQ3nx3bIjQCPUg4jvxPJfXRaujSskb4
n2SsUDfoMj6neSEp90GMEVFCd89nIPbuLpRj1gxiUmmmozTqnWUzONjNXEkQ3h1cKk2Q3tecLMIF
6mHzWxEh3w6Fpvft4U8K0bh9qWewEL+2TUvxNlQ+/hy9vIMAlwcygZS1lEcTkO1AfZGKIpP4x10N
3rvpErNWb+xOznppivdaGa3hURsaB6XME/sGrgz0tjgSgJmlZvZ9UTBkvMfqlmng0qCPMTQz9LDH
1S8cFzCo2GHQudyhtyeu11YDZD3HDVI8sVju3ueiH/+OmV3YXT95bP6KruJgJra51tosXGc3yVD0
1YCykUkW1eKE1P6F74ZfMjVlFiLl2wlAV3ijTPCFOZeB5bOaqi1ITLMGKdxDU1f62KBcwovUil9F
RB612rU9uzn1dIwXSE0y18VQuIw3X6Qb65dCfH7czyb0gQzHJ54V4VwfbTVtgDMC9Sc+EHv5nVm2
+0odsRr1y+h7z20uppCKvLA85zkOmX+GCgitMyK7CyWgGhOFyeqJ4DYPqRnzFLDcCGVfyymykTO6
uPdBm1gcqwROPGULc5gz/l8ftdjsV2IhsidJgcVfEqzIvArqpzr0nj+KB4BufCs9TCLefTNAi7s3
DIV+LuHvUJ+uExYkOR+l2jpMdZD12Pz0y8aNdArFE4GKQCPiU6dLVaPmY6UN/lHk60TTr62wIuuO
lJJTmvDYB7yJw0PZ1vBmgcDKHaEQh+lvzTyiHU56HwFqXjpueFp9ibo9QfM46GCfurgP8J9NLXMP
EBl6b8OdrfSrfmzSYXxY698Eo0cywFB1Y1uFfCGcUZzAFt+W3bm9e4BD9AEEGASbj1XcgAuj21ol
DnGN7bMsUdP8K31xDSqY6Mx7xzLxnD5QTEvZC5BEBCshcTZSkKoIE9ET+giwivjD4+HdzQpg3TW0
F9OUsUVQT24mNpn3rPUqNkq4SNI7MLRRXCvmC1CJ6m1NrQOVgudz0J1a2PNX7psl5dAQ+6h1ALDv
LvDL9wJpIme08I0JHESXT82OZZwSZJy+57XRVOU7ZrV80QsgLL8bvp8xa8pulmnDo1YSnyTNiis8
waqTuNf7BHRZQ9HOznBRrGQlIxKTKPmMZXAo0cUY+hJcAh5G3NO/zBFYEqPNf0DTD+EPghDqVkx0
EGM/2GcsmbDSRH0vwS2ks8nmckNFxl06YnPxgCcxONY4JzRM9m480XZWUPmCblReGSFM71Fr/u3A
B29hMp8V1WfL+5xoUCOWWxuwkm+iFq1n51JvsM1nSxS70/S5x94rZVSDy8mlnnFJlIX7zdplybfg
lwiMShsBRKU4rENML8wR8xnhTzg/Adz3n6CV5UQVjRXdIqOoZ81xBVBIYlY705va9ZGGOCq+QA+F
IuUvNz0yhVA9Ar4zgM0a4dc3gwXp9haiM8xiyhsKfgaRTtmTuvj71sU68wzv2r1f1TU9XApfbf8W
SxAZmD5kJ+QjPDF4XtZUNKM9u2BuICuJrD5u7VCNitqvthAsm3XJlBMxU/FW0pYk9HRcCsI7yqoF
TEOlhXdWpfTgJbVBam4sQtrPGIYDtMIqKjFMjAIdHiocLJhmRy5xhHugu6ppvTLtE5lqnnWVICyq
CZhC6+MseKlI7x8rM8pcqDVGH/DRYbk9tLzUYw7b+F05qow/brK2P+5sB7//2LYScAwlZXa8/Vif
57OcjK1Sv1tKs1+Bf7TCLMh+UAJq1k/dpXRDGpxev0jyjbgMGxDIiE8zYs+VRXHcZbx+y0/aky9U
LovmiYGhnTTl2NWEqbSqEqJ8ePInzXy7i77Ze4ZTDTdeCFtvZeDdEqicdsLM+8y8X45DkaJvdoIn
JIlbcVEMEMPGbgXwE707ukn3OzmI0hgQoasRed1sy5A56nx88SrJnVFlUTwAttyRdjkGL6zI7EIO
99aiDJ7FwpyL3UaJsLl8aPQkbGTe4067PTK+1ccNc9nrRU5WcXsgFumXAKpl9XP4ivlDPTJT8tNQ
wqtZ9c7KSGgCgk6xKgrQxe/syHcwSXc0una/No6uNE1NL2+/oLLf03luy3/deCsKBVcLou6rMiAx
wAwUcbqRal5rEQjaSuCoo7KuTeYeTN+YvE8C88ITdBeaaFef6smUoQmf8/e91QLuklzIqKhiSF8t
f5G+aUO9jafTaVCBnSmEaCo5MAZkCSKzmiuhAFjjSx43WiXazgPphGI6zfV4/CBb5QRZ99ZcFCf1
VkgjBlquNwagofuLJ+wdX7YjQDvLzm/pXFaAA8sAWCgnvklzVq127Ft6uMWicBkp0f1MItESg8Oo
YPH89cJQC9mBb99nokZ71v6D7t/NXMTuuS1U0cqziLqb9EzODJO2BeXFZMN9k0G0Rx4/Wq0Fal9t
vXhuS0s37MV/4h24NajhqTtCSD2We+YoReKYhCJ03c7M1yhOkjofFnWJ7DoJfRxx4DxGFoOJumJv
E85+lLQPfIjUO0SFSYGRLiN3iHobRSYqaJeyPQc80MLBHaSH8TbNlSVplbR2EdJpPKVDycDxFwAZ
J2XSFV/64wD2rYnI5kot03TzaGk96L3e74wbmip2DAi5dlNkCBpuOKHSQnAE6e0MiRAn/hDSTuAu
cs66No9f/2Qvnn9nc5fQe0dLz0je1Mj+/3OPWycMk+KsDNF5Fzo8TZUZXfEjbysplju4cMYOCtHB
DD92sYYBNShrVfd5QfAU8i37a1rNHtR50hYtvVYElMHMDaMkMrJ92DLWC1YENGw1s63TMa5hg2bx
MKZaC70U4WF61REqOgkj+bsEnkMelIYYrQbgFZsj8py+GZ6z+vkSw+Hin5t1qeeRlP6qGyHEnAab
v744tvPIY2IXLUor8j1Lw+sTFYfCvBRhIroWsRjWmDt5lipQxEMVb396bu1lylA6vMaH1jAjsSDM
Wm3TDUvwt0oEomHccs1uh85kcANNzphE5vkj5mH+E8QoZwVfbhWm+d2X9uGFkcFP43iVN661OOWW
TcVx320v/rHGaLhJHW9sdb/uY0Nkqu1mgiPC7VwlVt9MM/6A691TsZFopZeh5C8lqLLJKul3A4DR
XMHkUb78bgOyyt45KVrzv85wIbYdY123h9UqchNHfGNC9FKTnbR5K9cwdtcYNtePhNz2re5kz5y1
VgYCFBgZv4lPBq4Cy+Ubek7VGHWf7fA12fHd5etaz1B40Ti81yPxTRwoT9f4cBmvq7vHPdcQqwCw
RCxwq8pXtwE1uEColEqnuXBbhbuuf1yCxOto2JpmPfCUN2sXwhLlva8koF6wcLZ467K3KkNbenY2
Bm6a4Dn0IVN/a/edX0OYWtqOyQm+IMEQRP7lxcWTBPGXBbxrJmeZ3U/jbSrJTnC6h8a7bqb8wdfW
FLf81a03ZVOz3URuNXSwNIJx1wWDynSnxcU404L6mItRLyh8K6aQzzaMhdNkds7IJODWQQDFf1O9
EBIh+W+ZMNLglGKuJERE9Vs4mD6c6iAofhWWkF9Qe6NLUG+t+SXXOIX2KxnximCSq3fqI/YQS5yS
ZpksrMNQJb+o8lLmK4LeFvZc3Hbg3NXhN1cbXfM9ZEkWnaOGnemDpfsxjNZ+DgzsECLnZUQBzq8h
icjvYsBrNzwZu5Xd0/xFPyURzRaSIJX8or+9DPqckQkMzQbz71A81ayHLpkgp1bIjwuUybIvllMG
0hHg2i5EEMHLcBN/V8fERnzBBjzFb1ZjBEVYYa4LRl1rKexMbirSRnVX1wZlhUf6EVcLp2bbsAg2
ScZ1TKQPupqEJXNMpVYiLh8SAG2+L/zFHJaju38QzCxZmlhQuwt9rhKYJcppMWPMp3dpui5li1hB
aMzVoCSzBpP8P4xBe7TgAAgSGo7PXUstqiPuf848c4si11cMRMfWV6M09LxlqaL4kHSTzRZz3PAa
zTJPRg5TU75rqFIWvas62tLGRVOKq13gqx0KWKRLPRB6mMfpUOD6sscdUu08P75XxF13LvPtnT0P
G9TvW6aGHZE5nULmnja1ekyC34l5k4N3Kyzpmzbu869u70LeNP0qA5GIASyL1KeNnbiC7qnAeZN3
zl4M1cIWxfVG2/mjydz4TmzYPGIusIM5zr97K86RFXLK4uj/7GV70n78dznRxHakjJuXH8Kz2hFN
oVRIB7aY9q3CEoI4MSHB/IYAQMj1qFfoaoxaurheSv/61HCtaNN3EcRYXaFd/ATWcawu1kP16g4T
bvf08oES3on2j0LH0laLlgjC6SUzlOzSDyDQoaRV4RV7R2wSU4SIeVm8LIOviLpdSadMfd2420vz
2PPInC0+w8e9fkNLk+KMc39LAriP7s1Q4rkRLahjuFHxPh3bkpTPbYOaReggbLBR+bOuB9smDNSU
E7SKTJtwyPg3JBztzwgL+7eghR6xgicGLriu9HzMoC0SQxxk24yVHNBW+tYfhL25vbx6r3ikPj7J
FcT4FPFLyWav+1szJ2BoXrChwhroqOSXgtyb8Ad/fpDwbYo7vM2+tmeAzyhgAc8y/4i1jcv/hsH/
sHKFhRpMIDu+7iqZhcgcEASA1Qc1r1Y/TxB2pGipCPiXZSyqkV1mGjOTyQW2CJkWSSqrdwFASmlj
cf5OYv2we7dkoq3+mUisocnbGZtQNsx9PQcM+v6uTH5Lie5HLj7BHCBRJT4i1csilPIy0MN2/b6F
G76Zw9gxCqdOmihVJaw7sXuSqv6CHxaQwgFVIIiexW4d7x0mp180n+54LrNCHV5Ob2ZzHOXu63pV
Kz6/YC83yApA5oYyLntfBxUIg4HglrgSXrEkhk9MOFJz5xcZUj7DM8syZvMewc3eYk6pjm5PRAaI
LHtTrPd/E32bkAOoupYug1WBW/KF/lDgU1kbIJkp9QAtRy2sUXZBDfmXjL4ih4dssRLbZ3kxMmsR
aHu3pMpS6ZcfNe76wuScx5S+1jn64Z57N2Wd2hlS5jvG21rak2T8O9N6a+6bWLdeapLo+WJltMmp
BpiyfDZ3VkCXqah7WTKtbpErD2ixXbvf97ntuHrl9XcN0huaXsoYRg8eJEQR2ocwGmkWj9Epf5qw
+UqJIcwCvUeDqVltyC/NK5Twdyndxa1lDjKdapZuwdWuXJHUkRAkUKKcrRp5ZqGn9wC/n7H1UJtM
GqsX6E9Qgomod7f37MNvWFs8pgeXU/ufbrCZIalP7Z+AKok7G/UdhOmN32Lw3nZWByZRUw1wRSoq
4TrfjYh4wMGPiDS2U0gscaSXAkmkfOPMC4jnOE1EJbMfJ3ISKKVaovv0u6ZeJuuwEUay3I9JDPRF
Bt8LRmIo9cpJWz8s+WuHHKOyao/x4RTEsdqLKogqcOGZuWWVM0dI818KWFBuKaAyN80vpqK7yys2
rvVTGyObSpebU/g8T9ISCQoeoPCkw4e+PSwSSLsdIW+q8dOUsfeg/faQQ491aytrcX0nvk8nYsHE
stuaw/6x4hPTyCiBiPTn2R2668GCbnM8gKXhg+K2ZBYNh4RGGZnHgW52L16VX1HdX3v0kaIBXUZd
w8h7KS15FRILj/Z8irwL0iz3JlF0PzFkUVAg2zeAEP4vDBidhYWO9wkE7RNvATR3AuvlmOKRO9El
t4if/njNb9JjU+tge28GZ9blQXtnWMJyNiw52A0TLATrRqY8Ox5oPD8koW5L5mMs95bg8tmjYmLg
a1HydvwGjVGtWDUX/QxOY3RnlUfYA/ImF9+AIWDp3cvtOygGpwiODlfIsZl8bwQRnQI/s86NEUWY
mCnV3f5mUBTpnMvwNoKKbckLa0C0dfaaJ59rCm3HC3cxX2BZbDf5Lg8TUlpyhQTxj+5hFyNG4nnV
DAFjriXlMhypfZNrhQ5K7RGbl2p4+ZkuMN/aXZDV56Wz66Cp0qqkgoxbjTjwihIS6/IrB6VlF9/i
9IhikraP4k+2/6Kd9H7SELKLjBVSqnIDVr4Qjh6W7BVXmMiQoHINE/S/0V3pyFX/hBmEOmSqaO9v
+ydJICnSyTsy7p3Ru7xOjKho9iKq0hLY8dcXDvwhUGh0THnXc8b0Vf1HSLjfO4B/hJnSjxOe9q4P
G0WaSp/O4y93W8g25LBWtn9vuD0bwlZDQ3Yvv5fv/Z/5MYCZnS7MMmUKuqZNOjIbjF7n4QLThonZ
Fe574N35iEXSdfcdYm5ccf2/gM306f2VluSu2b5Z37pmJh55DD7keIHY+7FfOkcIZdwuV9l2zBwi
eo8tvekuuHEuBo0XXzMeiAI2HFatE4dKdQGlTitQEaNU9o+5W5Kcn8NoIsyiS4sadKrCsK1+/PpU
a6xa0Ra5pDT2eFBQPSp/3RJf8mpa2r9KKBpg8oYG1XWSRh2lsArRQ8HU09wuw9onyxLoxH08Ubh0
88eVRsNBXiOZ25ltM5H0Gcm1GKMjL1TZdsdXOow5CcvLDcVe23BZHqiESUpAzulYVUlHImUxAQTr
Iqh6NcbufROQ9ZxhHma1fF/OcLM8gS9W/6uyi4DVEQQD1SrkPxcvRieN/JNhXbVgAIIa7IvJAJhq
zYQ2SImIp+2R2N6nTHNoch1n4Erpg26icd4L62M2Vch8CyLLHoJTIwOq7z1MxK+HMyQyYn0VC0cV
EFLL/xQiXKFh2pHw+c0PAT7PJbuuqpyl39IS28PB3mhg/203m/qOpCZEt5hReS0EI4QjfN5mBD9/
XA6IYgBybsjC5hQD6fhqaX9MtjcSQ3crcwj8CX3HS870v6k3eRQwX/UQEFo5TNnN/aMmAhIY3ch7
LWYVASlkMZrzzOhDDy+U1q4Fo6+INxLmXHUs7wPbDWX6AN5o8t+/MGWHyGiCwBcpMgOzvpstl0d6
ItVOKKGOkMkytaFSLrCPpeWeG7povJfy0IH3d3x/NKrl5Cp4EoazCbLV2SqDa7kBSkfdksVA0SvX
hyZwshCjNU9evJ7zoGYb0Q91KEsHyf0o7BKIpKBYoNRULz2/fKlTBoBDYNRT+otR0am86QJ1z8jK
1Rz+80N6L8xYptVt5l5jiQ2Qs8DU7yya5jYNWYGqqzWQQQVQVoj+x3tSdCwRDQcVL369zhmgwt0u
Vk2byiqel1KUhndmHBT1NxneG45J//8fiUXPD9Qydr/3irab0EvOCGNgV0F+SJkCfYEBhbym/nKC
GimePpl3CSiLWzfCO+nl1Ro0AisZfqtHzCdKHeRVnh3mf7sWO7iz2Dogpu+5wPelsFM6zWPSpdD8
x9DRHJY9hvx3mYtvHvGS1bJof961Cn1anm8hbnXAvouAcgskSpANFXx7ArHUVepQOy2rOsqcqAD4
LyDgNcH0iEVCsO4UOwLbiRijxyhG96bZUm1CoFknNp5WVJ/3Px3gZKZKpmXB3xbDlrgEVK7RCLRH
Nsx/045AH8lJgBIL5szxTduLAVfCMN5bqMcH8j2zSC0Ns+r8OTU8y+p1ALGeY0jW4mcSXGsg69cL
XOfTQij6lLhhHngoktgDSdLlwlFvwUfJqHE16URP8nLb4GbwDoKl1RsBH+3sFi176XmNu7XvJFWq
/0xh2Y9UYIKljzXQKrFuDuUjZM5BKgXPpQekBOCIvvqIYprKernkrFai8DMy+3iU6XGaFRBTXtFX
Xj0nl3JaAla6WiP5+iP3BlF7aVoLJE8Ma1qSkQlqfizQo7fjsbjhBGAw4ti7SQrxa4phJuLDObsI
KI2JBSu7nIYm+PBzS5TZY6Fj2/7XpFspQwCJGQ0/FXST/xhu8PV2r0hHNW0styucwLnx3fZp7sOa
nN/eRnQ8xRxurf7korOdqzNiSotT/uFkPaDTRE2og6vvSG83TuUi+m4l7nis7saA6ENmAB4FG6wR
FEIdNXAkuCLZ8BIzkGOc9XIN4p2ZEDs0KPz5tnnQVGi6JqPgHl+nh5Nmwh1P2n40JK4OQOJKaPjk
LSwXhhYBPME2n24zGqX8DUvBZwNAjYnH1aZnrWvLRnleGwMo4Nh26xW29ZzvuKxCeEr+EsOEhDt0
fRJWU+6XJ18Ds6as2BFC+LZCMGg5oY788WGSGoLvbWOgmCnFgCIH2/RWSBjdL6R5XZxBvTDD8/yL
zrxMYifY6+mQCkurgV9xo2e0Xq/3Sqi5QG1J7j3pxgHBrpZ5swpTJmxCr9efkL2MppPN7d3WSxbJ
SXNbTGnHdXSij+Ybo4aNxOEDbz+VK7B1we3g1jHNK1duzR1xJnYx+x9y9MqJoW885crYwy3YFL0b
PJUkRQSBvvwN0fO37TK6LyEG5P0kMR+/czIxh4PJLQE7N62ciG/YfxbLpU2wXLxJ7XehOGYHL4al
SpwWN95drmSBdOjpLfLXe/MdaTKaMMdJLPBKx7+dLgueHOWEdi8FXbAKYMFzANNz392DPOTLD6mq
aO5/8g3ENZv2yahKBL7OjxuDw9XBPjwSCN4nrtP28z8GB4YDwABrq3vEkhi+SlriEJjB8vR0GVzr
nuQsIZ+kPNVOutNjJiZs5+6c8j6b+p9JaESf5ZfhI9Y5dVzQTdhzRnDn969Ksa7rT6qk3r3W5HJS
/4gKwYe1hwRCSazaas/YBGKmWvlFq03juOIUWN+rvAQ9E+yX3fEKho61m39LiwpIYFd+n4FvgS+0
2+EosrdnjdSc2fIroqH+JQYSp55+7oZfu4yl6BykVJTAmNAM9Je2Xfi07hJ1oTrssjjaQUmblF/g
KCY3T7haxWKwCKK9FNc/ErRNqk2QzhvsZyWHJeOgVbeMHk9spV5uYr367fx3wrOIdB56RuEkMVgY
ljYMAExJeRTU667fl36BpJaD9NejVbSEIz3N5QqB37u6940qbu1EtXZfjFMgSA7MAavfeiW5Yz8A
Haovjcd1jyBBjJ0uuoQbyG2XnKOdeEi3WcZV/ph7ElXB0ImXnttZW05tgP9yPU+h9m2FfwWjfJ/L
o5/IGL6SxpuGCEVlLNnFCyBUJ8o+8AusBWLizGpwT+Lpru99AJocNAmLn+xKDlY3AbGeDhGOfwG6
d8iYx5jz4L75k7a1VKdi0Gwe3KjLErsF9QSrP2az8PMZAtXBQcnSUmLzNl3ogyf0LZFwq+kB7+D1
9Ff6bpdz4KKzwycFdgCKHsaoTwBIneFqmWMw0CbeP1dzNWgVd9x2zYDEFR8CtccrapkzugkcTwXI
7ApcDOSLSobaLUFyrb+3xrN69c9mVIqJ1ZgBNDVjfJUUJmKyyN7W84jP3+J1Tt5WZT1v/zNZl1W/
0Xa7VnVhssvRxlo/QsW4Q2v/ShCY0cdcBRNrxuknN6F1xehx32KNb3zOvE0W1yD/kQuyUQVzLV+Q
A3f/TYkjpzBaTc5IQOtvHECnE2QnBwNd9aJhTSAtka+F0T3ShsqbmfQVDtXH/JfruoY1nTbMhTXj
0GOJB36KHYzsv14kcH5h12FOxXKsf/RoUuZ9OhP5y8w2obf323pErByXWGME7aSbqigbEu/oHU8G
wznqY+RmJqm3iJMErNUuJg2faHddNLVW2GWWok/kVruOuPiqA9SyCL7Hfu2lCCXB7G0bZXaQ7PAN
wIdgQ+ymHdM+/2poAtcPT+ruV9KwTnJ1SMX1I9bqdbzW0Kmy+kL8jNiT8wzD8emebHnb9t+cYj3w
W7Run5y7pYG2AKJmQXyNfHyAYdB8g4O4IIAVu371PlnT8FAtJifmryQKKwbV4m8pfXJLll1I/v7G
3OZ5CerSx8vGLUiKxHAtmIuKKeEx/cKFJzmQJG5+IcHRZZjpk2pIM13gPjaW8RW2DDomid9VtUol
B57/h66Z6y5m1ICuTnuv7ZhwmRAu5UiA8iS7uUrv+YIRM47doX3yOsF28pI7VaP/nxA7yn49amge
uPTO+GY7t4Ooq6FiRXLMI4DZbS8YzxwINnBcatI8D5jM+u2OP0mCO3UQ2ZfWWERoic5abpIO8CHh
l0dBf6EKPlWkykqlUVyEHW9LSsZBw1Gl788K6t5E4cOlaPywRRK2vSKoMkpZrXgyIWDOyBTdIzNU
xSiBT5nAi2lEMmcHA+4YOEXgdgDd46aDz7AiWDRZV+/bsbUszbCSQG6fdX2ajUxhHf60+8VWcvFs
WAX3PDDqFwuPQq6ve9WGEKO79aIXD3P8+RaFrwnnzkooK0RY+LW4PGE12a/2AgxQS4PHtGbdjImx
U6xZ7bLkSpPY8WfkhbnfZTclTDSQMeOF4KNkBGal8eww2xJxQbQAnnM4DkzriJXZ9m7cDcEiY3Cs
OHx3de3ayuLb9nSxCNiImqtXIbdgNdE85iWR0D+4qmNXJstekAgVwkgzSh/DBhnZY2RHR8Ngl6Xh
xuw3fxq+3/OdVCO5wSJ6daBFktXDimI0Vds+rX8Bn9GwLtcysfj3otrFoiHZoayN2WL9CvxgxhFl
P/rhunfspqpGFd7Ksc+OuGYp3fgMpLrIOyIiAPEEpMgva3LuwyOGT2+bj/lF/MgGx2s5PZ2lCGhI
acZNUdZ2nuQQlgFRaxJ0mM2xbxryC8ALOJGDQ9V9hVZ8+Z9yp2fz5JpMEApSD8o4UqbfMo/BpiJG
5826Nzpruy5IEtRMonk7yJUDm2PtFbaBeBAsjsYvj1zNifxFCdBFHnTr2gwcBc3Op923G4GaB0aM
pASX01hU+11xJjvRGjvBO8XBqk67BVnrgAw3JtOcWiBubKzx99m0j8TJAu7HVXMjHTc8A8+V6H0P
FsrFGD5YCwS+ym9VTzFXr6wB/iG08cCPmiUaJimAJOJdCxXKJIc5pf9yPzwkUmdKZqTomYdbjexV
/vUScK1Q4lXW7k1WwTjI+FQmA/lFCROPH6BoitGWMK5vbaHTh6mSVGohDgKdU/aXqgCgSd7ZPKjs
djtSjiZhj6OifhCyqWB7+YH68gNBWJ7MMNx8F/n7SjkPqgGLsdpycg7wyQJSjAYI6tgJF4vW1d9B
dsiV0u2nVvYZ1rItIdZi0aWF9QIkY3J7wUskoiO0MWo0PVdVCuySNT6IRCez36kfnSQ6b56aCCF9
IDRgJbNgwrmvLfjAjWt1R/fK3WCKyymxDnB4oEI6Jshad51oGL/PMJqm5XEq09jqszDFclEAwXsT
xhezzBj4q0rqNFzSU784NVVo7BbajYsmt8okVnp3jDi85IkSuw35f+S7imljHWNACmjhP2kQFVEl
HT1mX+loCwFMldBqPkGZo6eSIIViFKBP9rHWj6Q20EgmVgRTuk00Oh32ICFDp3lV/gsg4Jbyw4oQ
lWtJeuRDnCvUTmYVDSGXyR6BEb/Waz6NPjNmTe0cL7/9GNKIpflk/6oGOh+p49yCVj0au9bZe9Y2
nVI9y1La9LTFdhf1x42dn4NAZ58xlIeNJbLuxTBhiO9j3/lAztH4fZ7KU77hCRVs0gvZNjaHpHj9
xPlHvMU7/vMhJhq5H6uTGtK2ih+crBm65w4lwaUoYZ6v41SHqobcgLjLO2A55KijUrS4vn4wOlMt
1ivjhd7dBoPvka5Czj/G8FYR+zFoHxcSswuCHStNeer9KxtiR6dSZCxvGRIaLKAZL9cDUNbXxGVY
VSc80WiiS+r9pXZQdWDifTFz9ZTrQexlD5Kb9Dp+kb3ygzmAC2jf0cJ3qx0pJIoSUkd04x2BB8K7
uBjGI6sWDkX+wTFFBH+ilMXoQDD8o81U684gRv0B8lBp40wVJGM39QmWP14om4UqGLZJP+JHYFET
rEusaJWsK4MOrHtU7guTP1J/pOdQNPOMxfE4qWq9HlAZ7lEuqxGMu7+DHHPgOW9BOMOB1DxnJZDr
kNjC95N1h+Z//qnrL5WvuBOGDXw6oQxrsgtQ6f9w58EoEaf4y2d2MUgRxeBW5T6A7ayl/SzvAdgu
HX1HNjMbvHXKfd2VOQqXEZITkaRLi16TLrKCAFCD9uJA33YH/R4t2n27nOtWv7QFq9pkTpJyn5SQ
QUtyfkdP7yH7ymxD+BzpYrKuXjWmS1jQjr5wsaUCZ13+pMHh6mRnLHUwsx4ZrNf7n/nCL4GZXr09
oVubBffgCLI2cxOS+H/AAQXyN/MmxyDUuAgonAdB3UL8BPKdr2P6n3tzDV+o35dT/LWkcWKPx2W5
C5YF/INqRIwb6KbfmEuuaIA2gvDQeaiO6uwVwOCCaWd5rbne2nhWXZfOSusLx9NdBl/doAVS/ruT
0RsIcWlTMhCtjcSLN7GvneYqiF85jWSo7KE7v1FJXO2LFYQjGyAHPqzTWAeRrROSJwBVmYYdgLlu
2POafAmIf5e81b63SUSECtu7fxdx1ZHd4H90H9ibV3sLcOa0BKS1lKMFN7OnjDPcatDo6fPCZkpK
S4weCS+fv0yMuGnt9K/f6qs04mIoYBXlhH5S77MCiSeStu1QrzV3j7SLqKNXRX2NPpO+/ZmcKFOw
PHJ/N0GbzuwApbsbeKp+ORX4HchLLOG9KkOl1t8N+L4lq8HBnkQGUw3Z5iFXxlCV5s4edfAmOBU9
wyoKk95ey8wIHljPFdTWbwX6u4VmMBXKeER9wxdEItoMRm4wKg75ITmt/J7vaTyK2ALDs4Z1vvef
H/GKWm5ng/FS8v5kHxJKHSPAZ7IRfcpcEn7GMGgqlUyMsbpQJjDwOd2WOf4gQvt7VwfgMsycF4nS
Tz4Ek8mLwO5OIsdMnoh0IOpgT9yHXEMuqJTwbQpdFZ03bIV0kbb2udvWRm7wGrIHF0v8SHuuecpD
QGGcwx0wBtGVDzyE8MxO/L3nw9EeQ7E6zcYeLbxxllpxf3vSNr9yz6tE7yXuJng2o4Rd0Gu/6mQS
YcWXw/b3J2W3HBHcNkdfJ3kS3xTi7o0SFnYMGebbolriwmoqLF1Amzd4PXw6mDQs62IC4gPreL8j
T8YMprHYyKzl9xSqx+yRuH3FnGIwe8ExxSfCwvWR/8ta8iNgJjRDGM7IuG/FHpWAkqWStZHDEm6V
eUkrV/gxt+Dntw5EuUTVZhHErYzEbma9cDleGr6SMoYefIV4KeQKbGg9aeRIZIGJvXw13NSRBUwW
+aAFQfn0t5KrCzrDgK/ns4F3OW3I9fDcx35mioBc64qxrPvu8LFE0czFh3sED9PrWm3L4yTcePEZ
OeparzHvLXQnsY3wxTF/aVO+sioiLXzea7FYc285MLaSgExEE823FxcqaGMG4n6Wede/x+TGOSBF
+0bTHhLNnGqjEzGVgikR3EffOjBdqBDtGX+wjvsTXz5jdoltWtImV/yVmbhjqJunCFOB6AOGEYmj
ooPdP7SRsi7XVHPrLixs1i7Kn1Oiq8iOhqUq6CoFELYy9LJt+MYFv0KEnfZT4RVXcvJVQ1uAuLhj
Ta6KMMI3A9yxYl2v2iWltAfnkDu0OJfzpafm2PaplAf/Vnr0Y3HNoKhhltCEGQ5b3zjE81Se9wcV
dOkf2wVQToV1vrz4T0HnMdT2E7krwRQN6I6oS0lQsndC8rdlrm0SyIE4myh302NjZsq7fTpfYKoe
1GsANGmXPEdn/ymRyX5tjFPjXifsrWl++cCkhuewxVYh2HESk7NCInBAiTNeuyLbNCicVsMTkTo1
KXTpC+l/xGFbeUsaAL0YOw7EaiSu+DOUFRx8tjC/icPp5zIHknaCHYMGjhE5Q0CLRvZOKXa4KfKJ
5q8FwUzKvFZEY4VV0znDEe3adATRNv5Gm7f+HSJbUl1OhvM6zR7XugamRJO4WRB+8pvLHE4B9v1d
j2FAioLYF3V+HBFnWYpN2T+CPFmxDaTxc77yXokQkUnsXRNBdzSO6n9bSFEw+7TLl/QTbOwK6Cn9
DiTK1zy3B1ehcHvaNZifu+vbPTkcwe4eFNm9VPFEg+Axsd3lGq56GDbYaiZOSna20dnKeOm9smGf
plrLy4Jo59yZPNkxdlzZtqdjY+dKRRv8xHNgGRDOfU+xmnHrVCfsRUVKrbwI3b53H0wyf54x8W8/
rNAQvTdpjQDXSFVyJQrlsUfI40cLVWHqbaqT4p95rfGKZ7Z523HxSuxL6P3TRSUlWRLY/7XaxuSZ
wiUE3pb1b/obNFDk4gI6YQLkqgyduil4aOKaDTpWDN5vi3d8A5odH7WtdtCvxl2wMQ2DDzr0dUdF
oYB08VNpvVxY03Ylzi1fE1/zrSJgwJriCIQSPZOOO4zU9qW/6as2QZFADE73jGJdlutPt9QsctiR
eJIgq/6XUQmt10NiBExHtXuj8fyWoll6djG+OBcW7fzRE/X8pi90ePmX+9Y30QZtaFF5k2fzyC7M
265XtH6OZ8+Pw4r8aYBOsTWHZ0HGhO/UGFFnLPszwPdU2qTvllmkBt9N6yDrY2mN2lSUPUoOwNh0
JwznMlncF6g9n/HVI4mi+sC51flUN9BTyMwcgp1CF9sYkn2DJTA+CAkN2RJw4TxJew3i1DASYYUx
C7A2RrAJnKSiAJ92ASgN1MML5LySrW47im1vCTJ3isaVnKnSPDgdArVWHcIlxdc5sSgiyTpWVkLJ
s9LaWHcpuf5zsLEkkSVjPuxvvovFrUzkiPEed8qLEKPJ39XbpvcuUDgVgak4fXHCTGZoQ9WWIf6P
ZvP4vZhZPvO1wIv5ytJXQ7dLZwyQF/us36CAHa5cBlWLmHT2+BY6wFt1+lWaiWBnyWXS3+VwXOew
2YgEd0PMRDoqIqk36e1oSp1l/NgH+Pab4ulx6VFqWHKFcXn1OPDK913aj+LhRjGwdV3dLRK7rk+D
e1P1EvM2n0f9k4J0BaWRFugpqP/s0m1IKL1b+MK+QJfQnJqqZjydx4DjZ++ZsJbH6ir8K7zEDaND
s7pakOthJIHQYUPqJEUgJTaHoJIEoohTYfmb9x1WyG2Lm/Ix8S9n03PonbkoyDa54PvqwQcvaSDW
mVKZ79qlrYLjwBCRBJpr/Tn+Upirk22k+G5naqrJTZTycCkcQgqEXsY/pqD7DdY0MfBnolkSKQku
awMUW8FriOy+4WIWCuIuva9F5KoGqtaAJTMZkLx/HXp2sMDXdjEMi0xePy9lM0lxuzma4TIuHnih
ZlJDaKvVvkJRNSTx2obUcNLMW6yq97dATRPK5qHrumiOSoz9jVfLhRgfLZD2Zq+fv34y+PKSezrT
gBw/PWQc3NuYQefsxoan6RpMKAbPbTAWWByjVw2VY5P4/IS0yd31L04jQR0A6xHwRlM0R0m3BQAr
aBG/DnpSLMAEhFKPHPXUZErfWTiTlx6ujPJYPs8hK1BMewFoE8LfsuosbNzWqRsTlJz05RQcuxSg
6o7+NZwH0o37YE+GIS5rgJZCgeAvdR3n71d/YixbWiQ9NQ5WjBZ6Ic9iW5IUrPl2ENDKq62RpRb9
1AH2M26B2NgBIa/7eR9rvflP4k5IyznyUMLsGR+vhlkLXw8k7WPUpa7s9meN6d57h3xWlrf4j8T7
WG7fha/Diwv0eGyqmbfevBq3QtoE7xogXBWZ6lbJymlE35nmQ3IPYlLFQUAfncPYuyGJR+dC98OI
2U/AgZ5AecWg4nSKY79wA5mBOxC2Z/B/lgAl64/xGT83yq+0Sr4PhaRlY1VnrHOxDPBT4OwvlV7d
Yp0XUJpJyfblTHAovrPzRrsZ9tlI1C3WZULgzbLMoRYWPhnPRobVlHaT6pfxFPObJyS07T1JP/9V
zd00cZqgbYs6zYzzpt0fwz1peca+EfsJvVj3gPYE6e+8SCsSeh5ioLmoZQiuWYj0gM6gFHCogLU0
CZOOaYd3W6LSY1rbdrJT7F3FWGH6meUSeYCkSjn+gcFx3Uo9ANtK5llwBIFrBrj9IUbO67ow+OHs
aHG7f1EtD66WuWfqsg98yuBO8Frt/Y99vPc6dmwzrl9EMUUDZMJ1nf9BrcstMp0pmPrOgKiJ8P+l
30snXyvVKZwCVLEvXGO7sonawtMYytWvwRbaXwU8Lew+MsJ2Ri6OrMWqidCl4FlvHwCHQ9M0Yo+N
686dRoitoVXil7ryHiNF+VWLu1DUpSJ41iCAXFZ0yidhUmNwvDlT+DSIixs1Edrd8xRBzOeayyFe
Ztj5EgJrklixeo7n6SHqzyX8jkc3xBwuT65TSDJlKFXB3ahV3yfmLIPVpMaxMzA9nlVJwdVgZ+6S
7piTLywO0P7wyjL4zdXKAZKomCSaSNlWsTyIpDjKZXSx0M3lGoU9WBaNyY47JSC2jdRKNKSXEh5O
T86lta9KHkYFdBYGulrwFehSIqGCDak0emNUYnQ8rcJruLwM1gtI2Hw2P2amklq8FI1GX2JCLd9C
f39RUy6lxKXuEQJ6YhrYEtvqgGbHwxmENuEBY7jL7N5zjtRSTnT7e+jQGlZQJJDaLUVS7bWzeoyk
HsCQOvdC52qigoElLC71grVE4x++Gm+I4jGvB7n/d0eK8/xkHInAMEmvmDTEtdsEZATauB3WcHYb
hBNCYTM4bvoXMl8ka8S1yJgxpKsrkscSgh1gN/pP0Ycnkm3idcEZjQBY9ni214rKNo8ukzAK+kVT
/YlzgCZ5PQ4gm2EA8W+8G+FSvMymefDaKs8TMHb8/EqsXC+qOQof6mtI2Eo1HceSWWgwLsOcseIM
FvAQVKXuGj0khMOiVnmD0rcSpKMzHe2JY8chEUlqhQpKpC7CmF5H/WEUyTEBO1jR7RbBjAEmcJIM
d7mqrh4kPCnTwwkSb4AqguyMh8LvMcQ4oIgCOwfwuUZ06sK0AOIVCuPtZ9QrTmZFai5/1wJiOFeU
tr14CZCKRJpFW//RRrIR46LJq0EP5EWpR3fUR2jhddB+WtgOKzXZ1D3KCc4ulpZQaF/He2o+ANU9
Y35cuR3BIE2TJi3MMgn+Pd5FfrerehhZJi/kCqgKOLvytkE4woWaiF/GVCqENgtfEnAyLazQfeKj
AI2exs3j/SuCgt5fOldKclPwNm9YcY2zlcsY+UgN7IzQRIcQBsREPlRGHeB8o25f5lG7tBM7UKQG
nDDrq28cybmwQMhREEEh3fLwN75snw4z18X76vwFopmRoNjOuGtG/HlmZWpFXaKBGPX6hqT4rXp7
NDx0iJb9Mlch00tazf3ssYfiTmN3w9n3AS6FkSULDRSXX1sH6FMqRmBl5//A5KW3kwJ7PoUchzoJ
kZ2LU4SEu8iEKVFCXllmL22EgufsLo5Lh0DKRe606XBGzcEHNy3h5NbtP4PZmaQr8IHLhnW9KIlH
Xvf1mqgREPfu1/ILxiQ5C6XipdUuIYGCfZui779Mz4tXs9HDx8umcWUs+XaNuIeTbZ3DYyf0NPHR
uhxOM48ljT6t7pokUfJDowQfKG2pYTIXd1WVPe7QbVcBgJjh6DO832Wz+LzRri9fAs9MNtvpc/Bg
1d6LShsegtTWTHsZThXOS1e2DgTfcGswiotV7VQloa6tcc4XHHa2DUTh5+mcbIY4JOxP9c6ogfu5
mE3sV4X3eil7GMqXo0nfzz/nOxmqptgY0TjaiMAKRWgHcyCZiWp7BjNOEPn5pp2/03GH+vhctk6N
DpCSCg/eJtDs9uTITtJkAHV0yO2BF+LrKF2iRaDxJmlAKh3pyAPqT6xA9Pe3UlyCqJYB6F385VrK
T3+ooZPqYHt17zsM92uFwqpNxIE5/Khnhe6m+Hro2dlvevPq2c5A1zNOHLP5FWdGcxCPMDbGqEdf
nBcnQsQyPoUqDi9CGgTKPT/Yg8ld6s5s3bO7VIQBERn7CMqEcjASvQdtZaujtzaI4Q+lrfzzHxeL
ZSQ9XZUZuADWhmMzaIMeMj1NIQIXDku1Cn+Pps+mKfG0rIyxdswDivPNy7hIEPX1ocEqcCKh6sWO
ESV9fok8MhxQxgZP/Du6BAtJ9cClGVi8tM26PdVAalBrasF35DKl32Domg6kHsxoJ0FBRUzGnUYz
yyfQnzfs1aeKGNw2EmofJrOWjQ66kHsucqL6eLdcbAeaIDhg5Vvne/bWrKISAhLmGvE26VjOruB6
Tc6ZJCNeklnKIdk7fN6EQ5G80NOmz3oqZPqL9bYAAMxFfe6ZWUEPqaCalKPfHeK/Jg+sbzCPQfJ9
bGke8g8Cx7yJJ1S4vCUTDOKI1QoGnR1o/C+I+Gx1n5YvVGZ9J5QkEwymfBb+W9ZgALPWc+ZD+zT9
FUZ+T2uXH3cEFe9xVz+4VFYx0HG3hHj/+fR4oANLd61QJY9kXmkxOsw7dreIpDYPK31zR7CTaVbI
AfW48lUHiKgwZqvpWMXgvWF7G7ssrIr1VN7HL2Vc7UY9fzcCi2M3m85tK7ROacZIdhWKhlR8oW6p
uQJRWVCThpuwa5Ycxfdp1jcu2ncNys4GHj4Ne2rNvZj0xC2vLYMqLkeMFOmqvtGyBgoLoaptNRkj
Pss+i6HtIGGmFkMzP2M7L6HEvwVDOE/yqnnSHyh/vapsaY/sLMbebLJ+TcFn0E+mKSBxYT4wzZJt
o7e5tW8oGVh/caOg1JQ7wpZ0heyoe92UGtYLmGg4Tkx+rPbwi1BKqg3u2g5lHeUczJTS72SzQN7J
sKR8G80tIzbAWET1phdm/C7fM3fJYu4XlhheJSHjHbiGxUZ3opsYWYkAL1F1kZ8l5KH6OkG3drw4
khHdoHR+yMLot/NyRFpogonwP51dljNP4Wf986hudyUQ2WXcrBNm/CqoxOR2PCjza9JmuTqzpCOI
uWF0VUdDl10z8JUqAMhjp2mg04soPrNauGVkLNmYC1VRRYVRqNwProUNBQYRmGLoZhbNCVLUGhx9
cO0dsNq5pvIOVjtZxjya4ZMgtqhpCDaGIWDQalXzvvtbZKcPL8besnAFZw2Dl8dSpbZIJz8UHnbJ
yI0Lcta4Jpn9hSDxrNPqmT12HDIVGiJxy0vjEXTwyiFLO0XP6ywYUcnU5XqInhWEqvRJdvTT2YXE
uD7NE6RL32kk2vmOimCM3GhtKaLwAvZrPLY5h1D5yCCHyI0I4DDCkHjdHExcfua+tphVo2CiMaER
CGIy7X5d+hEZaicsJ8kuQRElg5SsVpVc1qV+/q53t317TkpX0H+5HNI//xnRgPuN9f+G/5nH+Qcd
nKUr0oAn1UjEGayHD3CLCTueRwGivX0hMJXUBU6PTSD0m9udCIiUar29bJEseus0Wjx9RGuCZiDn
jtRiU9BdpurbDgGG+rdRu8N62SP/2nZ02eKSHqqeOV4v+EEU0DtFoSbHu1h6x6OMTb19MZTpWvUJ
FCurACzrq3b1EDRz/wTeP+DgufytITbfj6M0Gx+Eibj6nZ1h8Gz56awrfcHYSorIN054OBBIW+bW
yue+uz6VhhsMVEKOMU8W1wDBJJLkYOjIVTGH6XTWRDG6RdR5K5kv7IPHSt2tAeqUI72UB8Bhb1Tj
sygIV6/7RsXPdU3i8SlS+IzBHTkukZE2tDj9DY83QoAcg4uBmOGyse5JV6WIMIjL+liz0tmXxjAt
OVFm8140b7cArj5hvWDJL4igr3yl9iXncK0WDARF9VJdAHMwLnH8e2clRvViqXg4y2KfAYPo6yf4
NbLXkKIYFO7a3O3mxvEpFb8BLvpgqk3IY6P6+0ii+akbml4xyGoSOKbuv0miEAk4/lHVUvLWKhUr
qXm7f8/iHFZjpTeKMLtatXKr2lGzLHSIitfJQUgONq72EE0ARe9VWX03a6TozRb6XXyh10xQ9bkt
PIefxXQmpkp+WnySOEhlve2QG9UyJKrbwhusEeD7xu6AHRvKoQbATQqyDbTQLBVaRg4z2fYQgj1E
yt/YlJEWY7NRxcykfpuYld3QWAhaGfIv4gACuVDt9ODzZvzvAgl3RrJzY3WmacmG9yXmW15g6sAT
UC9wdK0Gc6vq2dwR3JAWqHIs+0L1/aC8OgBBMnrNGuUmmhszSO6WZTOHODeI4zdkDHmmgyMMSRrR
gjuLyNPovcyvYI/JYgaml3kK6FUTCre4dw7tFY8Qv6L0o3i6ScFZGeK8H3mGJ3PLoixBnaHSPf95
Vg9QJ0eshfDr6Cea4vGujGYrkLk56Et5WiDA1a9WgpByVwwkBlK1llV1uCalZSWIyabuLMYBhdYd
uf+xYy9IbzZra8BUW5uc3L8nl5nmc19KevJs2wPdgE6C1WXbRpqTbL9u4j8gRbJj+hvZzREwbvtt
V0buBcHC+pYxDrnRJ2PDWO/p0zyw0HclFMxWOqUczq/a4i8ML5f91g7HJS5XsZ2Fr/YmTTdXLxFh
9cAFPpBbiLts8oPaFCnXXILLvVpNy9XBMskRpx/AOR3gSefzp8Q83k0ffoBLqd2FSlZ7aKlV3Cj1
VQrSRvJD3eJI8MkFghxbMiXdzCSZbbkXGsa0MjRlJMRDLNmtzijAuANvLKEVe8IpLShQr58LzdxN
sXl47h7vAwkuXH0HIj5BiL4xqQAX629mqgRAg8w3itYfm7VV7Qxvv2W9zDXTWt8rvrXlTWcf6W5d
Qbi1EC3Uk11VTXEUGIlMwwru0Pgsh5s7CQ4AgcQx8244qjfjdO1pxhJUCz+ge/cRa+QJ/DkPCzG+
XMuxbzUhrHGRFZjslx1LDmtogS6Qk7ZZx/4KFlRHfzTiYWM/4VoRYBE5YcQ7pj9hIPoaT1rNG2vZ
XCPH0UDBAK+p8/gjH2nbS7ecNzWHueqn0hi7ix2SD97BolvWaFcXKoI+xBgTeDsPuDYTQzoFuIX8
w+XrMsYvt9Hcv7WGmomVg3PEmKvA7W65Ux9CgsGkMEXOaiV0nwm0SB6yKNgX0mvw6+qxjTvG2jPP
IrKLsXN+ivnSRfcRyTl0BMKYCtJbqaZHMLgn2jRngL8SlVwzQ5dBQyTi8u/aCFSzxx/5Ve9wgjO7
CeeBdaa/wWXzq3bNyK7n8ip7bN9xgYksDZtxyC6YaiN1DwZL4FMLkTyAZwUCFINr7xKax5JfOn3N
AyJE+sI/aPSDkeouZvKZE9tyixo0YNuFZSfIkixH8jhV/m+S4Rr1Bo5/vaLr0/JNnE30hjLDjjT2
l6W/3g56NQmikqQJ4n5rGybfKBVqc9fVWBla0Fg06zlzL9ulrvrWF8ZbeXgBV1gim07VXEtPDA8l
fdEf/2crnazNngf+fivid8S2eOD7cL/TI/SKWPbbo1KZqdC4juGNRqas/0XcLSXQgHUQznlf6WWU
2lHwFd/5L1dZcV4ixsvqtfXREBg1k7yIVZnBRpqTUxOTm7CV966hryPSYt/HCwU3c1LF48ZpN6IH
cKCkW4XCKKNz34s/nVjSx8nQxlqY5RXj3IL/j9VXYE+bKSDbo9Acy8cypb6fv5X55aas7ImncqbQ
zlbUxylzfne8TAlN1+aBas0e0nzQddGZWpDpgCOo4V7SAJqIRcSGZdmLiLgGbWmyk0L06hBUMfOb
ketVe5ak6+euim5AeOgWltCngAOy3VLx9DTyARglyNQvGw6pFlUesH6UJzK6xIfYLPmeBGxObj6r
B95rwh9hWSIIiIaWFs8CpdlcBN6zAiuThe1WetJ7KO0ODRFYMDe/JtYLEpfVHudpUZnKjK4ubE5K
tbExUn2aKE/nKKdAAdi7TvQLmBXS3DfaLqba5UWrhnLeWucrO9LQbp7wRb7MryH0D+b30WI5qXzu
sfBe2nhAeMpDZPEyidx8wiS4scXxjv0SLPGADa5lUCG8/J5GpKfyUqPtxia+xW4yY3l0IDcrmIvv
SaxEXYblhwVp+VU3uXXqUJ0XGz7v0o2JbudarlIm4ut90aFkGmYuyDejVye4Ra0m7/DfROXtDYuK
MnQoWh1qc4GrY7vWBM1uIaH93ax5CZ3wQIZlWocdYsij7YXfOWn9cjU25cVDRQ11Q+srEjNObNOv
g/tsZpnUoAvBQeQKExdnayIy+zDfnJTJt7OmQUqTVNPEUuekYB7PxoWQV63937CtvmO2Vas09hDS
+TkBWhM1b4kQntxXVg0wWTdgjAqH4AIbxuOZvCEGDWg0cmQAFdwnrjXVfQR7X/r1poVEJqE8OHrF
tO7gAm3b+x3xq4YhIWRgQgCCV26K6w1eyyYNTlUS2wk+PocLREKpndmDDH0wQExXyi73lg9HewFY
yc6OLybxRayCLtC67MIcXVpxwMeoNgiqCcRz9PB1NsTzfrXpwQaqLt9sD5TQoX0SNAziHex7xkQD
iiFgyHl+NAjVXWO/vg2/bDajvCcSYd2AyPaKOBlDpPEJxPIHBlzLzVvwyXDUT7Xh7wxp1eD6rysa
bmYlUIezzowrMK44CZOb/BELPdUpfcy1VqTwrl4+mTjPnyO0Hx9APid6BrJ0lJOejpULtAxUW82L
ZYqEHOkn2sba5mDq4Nn54Dk8W5BJkzx/T2h+C/SSrV1NpUVcHiKgQmvQDdwJ0IaZB0RYgY66sr5P
BqG1VklhUAh+U4dD1vKShDxTSwfoiIS94PPjDT/cV21qphmgknm81o5LuJus0hrDwsy29dNDNpEx
PSrxCpG241vF+Roa0svrynqp+TL81oN0xIWnObY/4WYYIsIPY8ipeDxKzSGrFG2VylrXbBG8PW5Y
JYfPUlSFpCjX/lCd/ucz4BVkhEjgD/+hAfVDla0qhwJdErVWPKbOcPyifltnMyBDZpZ5d2h9zXA7
z7EAjeugm2ch4ThxggtGpPpiK9KT9wtHgEAj7u/+owaNBqjGzvUylZiK9F68O4NmtjLyt1iOOYty
Zw8zfBYW5LAJeIozd9mBYwMYjnQ6MF2BDvBKu+GNNX1hFu9DuZurLSKiy0/WsHnzU1E8aK6QTWxF
QqLE0bKsuTSeA91BGSNI6DsQuqQS+az7un8xSwSbmkPipywzBlaqsoux1CzY5svsm0POvYuK+5Wo
gSiFUwGdfAwWiWL8byZETFW3Nksvi+7j/euOLO4VUncAyjzX/ZySYMnvWfjLWkuBgy4Uj21EKM2g
9C/DVBGjFfNy5kxe63eWtSwYLKTOm8oK++qPx5yyIRcA9bNTMYam6djeDAJYDzsahkucW3B/bQZO
qgY9WG8h2lAadl/IGA3D0Sz09rPMST1aWr2LEuaDuvupztqu9Ui+p/QbvLpg49zkmSJDviw8xDTF
/BIpreSQd4+tnR9bh8c8lHzARgE/cbE+jzP3gXEncBxCxKmLiY7is8jkuGF82euwzgWB+IkM54+3
eiaWhyKGMJjncDDHBBRRSQigGUGEWhjI5oBbUWx+BJPjEUADMb98KFtbUdCwP070Tf9Q+SeAP8AR
SEHpGRslxuagJi/QjZY+X9lHdw1lrJROrb//Abc+i1O9wO2nbfoJioswjpKd6fLoiRWTeu5c+WFO
ildyEhQ1lJK1gqo+HbyiHk/VrnIVuWiabQ/OHCpzq+m1jmCq14+8ZHIaApvQJ2aF7a4ygQ+zOsGn
PBzYtYS1TxBgZyKD2UHK0e48LHGQ4ILXYZUnVqcp5v6z2XVlTqVk6PxpIvsn34u5nQ7XojH5wGxz
4Eb3e2xKI9dYT7Cu8oYWSm9eZ3McJbjf8Ouz0Pn+ySWFnMFs/atO4KJL1FWWbmoSX61yo0OWpfBo
e6T2U1Gz0gn6xw/93Zjpb6S4d2dUyWpWWlt0jOdEraJ7DEC/nIrlwaKxiPRcU77yrgQCAJQZ//+D
VtMaILavGdYVoF+9Mrk/EDpl8vZD0V9eqEvTtXMbTbcFO2Lba0o5nJt53veaErwwl0xoRhyuJhSC
QeL0cG7/Q2zVq2QxZCpqNJvjMNjMWMh46Eg+m1vKwwxG0NSASwO3d2+NliH0JhFrFdf90xbdm5Xd
VmjrqPMJ+IMx/qk+cd2Gj+ZI86+doWPwSkkMHsFbaaXVPf/nUpQ8LJ4tYBZSgnhO/+u/oEFRhAJr
ZBp5xwdQS61x0jNVlCScUbnb5TY19O7rd2RckB3CIWHlj3+kECfr896i4UMT0vstPs54FWPETlpq
Y7MF5VNlVsXcm0j5RLKUIAz0B8dxhMzCEpWbAzeLFNaGIbYaEBz1hcZjR7MGlv6DfEJ6LuGgRne4
RA/2Eulea45FXB93R5yuvqDdPI4C2U5SsjwCLPp8H6pr0gB/0WiU1mc2/yte1/2yr/XZaz5Lu1gf
mAp5stdtv76QXKHlmWGleAdVEKqN1NuCMHauUetSa52Ldky/xL6dJslo2LWkuxChS1eQ6EY+i4rI
n+9x+wniJVi2m5LOMiUuTCujcRXOtiem3kcn7PrHwKmDtZKHzHfKjl3Je7PD8fj2XZSaNVlTovPQ
eCg2+HP4WQupU5cmXipF5FdH4lPdmnufV9N9xxFM08MqzKo+2hldBdb68CVA51hhUUQEqnM0NM60
frRK8swdGwN939WvBPt/MyMmV2zB84j6uXaQRTi2hE0KWDG12Kf8WxnFw91a33Vkrz0bNoRN3lLs
sgG8wbuWt9ZikwvY4Q1bpRyw7b37iHQEFUAFtfXrgTJpQEXx0nzKERIbC+eM+32fLWlPcqGxzUXg
wNYnDYKHsg28Dn8G4sHDzl1uSUMwt1zQz64Ge9xyyVBaukVGkUby7H4O2T7kqwn14fo/6ZMxIEn8
8X/EJqMKTn1wAUR3wRjFNqdb+gwM8YT2sQjO171u0isZal1HFLiZid09M5OohLPFWn0oiSfVy13C
oe+UfujT6i9cz2F3DsE6thPAHYlwtiqf0SUxRrqXV0SNKyf8IxSETIBFudajQ4wp9Ny7Gb0B/t5d
lfEgmO2KO4Buhout6C0/WSo5Jv3Tp3/6nZ9plIlD+XR7bBJlqWN6SMzGTEQaw/xQMGQRnCa6qqRg
j1c8Vd+5Ue+rBvCUyfZ6OYBXkIiMsi1pD+/eoNtdTT8VtNT2SDmr7jdDZlsu/uOm7p1S971gp9vq
heA0Gd8Q7CgCWM/0gsqHEIfsH33zx3nbYTVQ2POx441rKzv+FPn3BhJvFhZeHs7CfGkJ/GCJ1/yV
2MfVQ2inu30n6XoGpRoEddduIvDfOhCf6rtBOfiabu65d2lVw0Il4twLOxDdF9iPwolfi7fsbnso
WbFEIQssumgjExBz9TWGBN5keS6YCmcByz6rqvPWXwhAsOV3Q18a58rnPFmyp0q2DQEgkFFiAZ5J
hde3UV7i9YTW026E0xCJEVot29GfvSoPX3swa+wQa1HehC9QGK34X2MxaDj6qMbzSybaFh2myQyb
JnyIbHg2sCjgIZKRvj5BmTC5XXWNUWlm2sYbuDgKp0F7CXAY88x4noLZ1MJrT+9RKWoYBhkJ+sWp
keCQ+ocoNkoY5Kqk0uXy553nGEtz7/r8cBRPYUBW4h+ZPTrI+l+0g1Bu+nLT2n+q8jQGXE6o7OU4
r241xzQf1T2gZ7/6wn9m1schmcIK66WX89AbwQiZAMN6hgXZTJJ3osjy0gno6glmDz3SNvSgE+ak
0yTUHmXKsdXwNg6BtHI+HOPkF5XxGvqy6et459mbkQFbqNF/uppRO5b6S2fH9sD78lGB2rSFZ7KI
uBFSsaZTN0ElvE/L7P7ksJ7xxLcPhzbdtJR2gAPRLa3I4urPt0VIIguoadoFNcragvSok0xUivod
t9MipT3oCh6K2EqQ+AhVS/wbW8Hoeez8zNnwpIgkkxnCBNzSU0B36lGh/88qXBbpzrnArGkyXA2s
R7zSNZ7OYxBg8o/5DyHW8OpkpAHM2zidug2ztP4P0x1bS9zCPyTeBX93jNiQkSxlrYrE/E2r9HAK
39sykwBOBs7+JMz1dxHCSnhunF+N8dRA3IIcFlizIGmfbM8Akrl1GY2c1ndpwZCjdHHwY89ueQwV
BIvFegoPpTC6lOri0KW3U+HzsJrCjEKEiNRKaooCebFG8V6qe1lKGE66kc3C/fPgiGixZ50fBEc6
jRZXCIXr4n1tqLr8esFWPvxhj/ICxc5YmdKjPP0B6AZyIbtx6WytqOAmQjEFB7Y5JXRmf71jz0he
89B0mSMe2Dmm2LcUeiNCxtDjvIJwk/3F9+WjrD+Kpu/wkw715vGjRyZdieZFOV+uwvOn2JfjaTvG
Sc3DRYTuIpQL7Ch6Rcn3Di6K1oSR2b4rUMccfcN6Et0Lddd8B/N5G7YH9XjlpaMBFvDwleOD5Guh
OljEjB5ZNxca/hFvMo7mHkyDudfUfeu5OwYr3ssuWOF2I5JvKJmsE/AiRpgFPTdxYMVrWRt6hD6K
gR1pMl/U5zh/4qgkTI/9gEvuFLwe3gm7YFAaHQpiBdBgLdirjeIvXVaOpJoA56UO0D+KftVSxel3
stOyeTocN81J4aqfac3aVq754LBWVCADUr+Om+ST18LgH1E+weNZxPjdo7kIjOgcXb180K1KLA+t
nSqjpncVdWnEi2B+h/i+A+GI0oJZahdzxocaTOAInfja/CjFxD5c5nZq9Hx7URzRRAoCM5b8n81l
t+LW3GYaKtFwdbhw/PuARAbOfYug6govJYp0Y55RfVIZgmDzgdZ7wyho18RFVN+MasXlPMqIiTKy
JjWv+O7vxQ1G4iVWUX+Qd8wy8WjHFFMHCrABbNeb8nvs4o9Qmuot4SWqfQYYjvwNsg5xP7dcSnx1
LUcb+C+uNNHOAWQndKuCNIC9PuAUgpGmq5pFu63BQSMKhjrbwCuXFSmUCwNp7s4S7r3UeYXOVgvY
OYcLB/m6Upc5DpqCOiyV73/p5mvCSSHkahkmAGn1rSAmoaYwL75WnLGeIx9Mbh/px0efBUYwMpoW
m4QvmQt4blK7ZrYGnFlpQ0nLInjW594+DUnptbqoBjJR3Tqu+diSvfhLB9W1tx8bbp+w+ZGEBWiT
LPvaSspV9+TfFDT2EGJMwLr5Ql/oqQEtnOTFJA/m5udPf5UP11Juvyphqt+a2pGdRDzru9d71rQ2
XHVUKASUwmm5cuLjyeeULRec6BvfEkYuPlTZK2UAECBBWPpBpgF13qBbplIZJSF8FKbAGFA9ASTf
FvWz4BiLMGTatmdSVNwdWn66ky+m2kMafdPiuZHUT5ypF+aTu4cIIfdoneVIwKSKSq2Tc74CvUmD
RfNanSmCQcl4cwHE3qmpIaQaqca5EuK0Qlqd6gSaQUbyZtL49ypSwFuOTm3utsCb707CUdwB12R+
YrFd/SkCwfRWX3CtotFlx1FKUrY0a4VFyjiXc4bWt/f93tSJ8B6dbh2OB+h3nQ9HbxSKEJLB0y+w
jxzBM+eh1kWNQjKGcN8OkIQrT0srqKElqC+04BVFfl4dYRQjBRR2N+GaHxUIsQUQB8Aei2z04QF4
FkqUA8Xb/uvljJdJtIa2FwwMtjZP7f3cMffJChMibAVhffxHuI4VCgwhCmbIYbhXfNyCCK2zKaQS
1Q1R4Q6NxztngiDX9srht2nGXyltkRz/h4RwJ/sGJXpOpzz+KgTjLly0Xie6FfaWYVjZuJKXqBER
urgV2IFEuESWhmSPd3zBktpjVl2da8vxcmV5JBTqUa6+uxJl1b0swnqXOKMVgvPwmyfY4zlv+/e+
fDBJf8/pRovmpYGbs1Sbng1EXghYE1ScgesZGBgSQl6FFBTNhbKGqe921XS5LrMBBClFmqch5Qk2
988ONOk1ez93vKy97ITi1fGZ6bP5gTzeb24aWufv30mYmHquuJOzq4+laHiNZvbJIK0j0v1X9ELb
hCpDM/oFsirOtLicRTq+NmxmXduYe4QlATES5tUzyv8eDRcP4mQyeUcqqLAP1IuVxkO9o4hjhNBA
TbfiZ/ieO69wTZpQjF6thWdC2ZcpZx5sHwYYHZV/8vvcKA/yLaDs277CDXnVuD1hywckDHnXosIh
/Fg330k5UCcBl+m+YM87PL5p8Z04XwjhZ9z/qNHLl/VkzTN3RQpV0JnIr8utJkfrV3rPNGCbKolB
Sh78fHnHMX1/RBaO93dcjeOzS1d5RAZd3rTjgJgWxcw8FJaS0/HwOiXKpsTFBixTHKwek3gELpK5
jYuCgcMSVk5Rbv9yTtRPOGu0v72btPx/hrUb6It6nshS/U6C8q1M5jN04QRK/f+4YEicnnPpdRbk
8ux0NvtRqz1VVkNvnod6lD5y55wGPbiHIKUx+v100xBVO8Wuxft68VXGnDXfNjO+jAgSHWR1PCo6
/RGL1GMF68/Zo5GbOPX0x7i0JCci1+01osBui9Tqsh6DekVuF/QXjjdcuTgi1U8pwNHGc11Rv6po
Gfo05Sp6jtKoja3rPJ0HiHV3d6mM/hyXJJWrXKl2MwIUy8WzseQKpMJaXlE8FuaCrhMZ14VDzNrU
xDr5P5sxkZGAGyAq1J0ZKv9tQ+OSCOnOT2ioK58Ao1B2QykojKuS4hX+0IkrFHJ8RqEAsWIwTMa6
Fo2uAAGg3KVbSozU0qUA4pjNL92iKayrCrrnhDZ5s4uNLMNxVp5piORnsDvTDA3pUk4IdMXHpgMw
sUQT+VA+W2XmMGUSmt3D5ZbX9yi4DLRng0/OaUU7Xiuhrx0BSuzwUmfhTliHbDRFXXMBJWcaziX+
V7CqZc1hCXcFf+cOi5n42qbf39p70SVIkChhs2UGv22fBrNDR1uxir2/xszou3MnBrLk/zigh/oS
fRRjXfVvfDAfb403Oa9iXPGgTH/vSVZeNmp/YIIcVaktS1w0dNpenpICrtGMxPPYG8C5s/tJtROG
guOFVndg+Q11RpVl0m5aLQle/zHo5X0/UBCog19zexzllHV0lue4uGfSA+0t48gs0ivvr91FtxZs
hPE3sJgj4/AIX3p6iwZCWXFvyHM65L+ELdPUe89GTiP9Lt2ZqI9+VT9qPrMeyis72dXgjGbm0EcK
YQFYmxrVNLDjnUPbCYrtO5lbJS1M+TrwgaCIgetPX2bivkn28r28TPcKpeBxOtPBNzAAU4spMywf
pcaqVqWYXje8CxYJ5xyUnhdh9kyy2bB7LVBvUZQ3/ZOG5qwBZxF+e+9HyHSIBdI/iKEhpmpyJzA3
dJY6lJxgrQdgJTzBG4rqIvL7U330acnCWjwxgCTDrBls4PXJd/NDwCTEzbJAfpD71PhGiDEWvujc
sxycFVz4WpcZ3cWPeHzdsMHbXbevQFTLafnW5x9+K9U609DxEMaTq3zI8m++p+cbUWd4iTgNytgy
QwlhjfO8el8NGRE4GU+1cCOGvF7hjIT7y/AohtAzcg86Y16zidUL21skGBM7ep25J1kvtMeFvADd
GONYPSMQ+abDRyDLEDEWDWLfRu23atM1hxwTGQPCWbMs5EEm9RknHSxvPsHZQ6Q+8bKEHhS7133n
/2Ugf+bH82kTuSegNl2nSx94MXtZotAcmWuSCMF6hatxyZkLFWN0lw6iWv3IgEV9GiKoFoXXQo7R
oCXr0SBpsOlojvc8YLZmIE7119pdj1A5KmtBHL7z5f+ZOZYpSYKoHspGn3V3h1on4LAYzjOH81Dh
m+qu70fPDowhoMJmirHu79uAdTezqd/yBiPL8spemtLmlPqMi98IEjIeXJiy0FKdKMGrA9/NrQ9C
UJm6/tB7/4kDClu4GN+ON5x9PIcVpHzZAhdHtnVz7VDSFcyP3JxMAK2Zfrg+v0VYRdRmK1cygbYE
6pwbNKv28dE+eqGZ6lON7YCrIhgmWS+QDil2H48VLx+8UsAv2nfuazSOsNEzBkizRUS+CMQNg7E9
hbWdvz2lgeVSBuS0roxZbVrjIpHnR/wOQeKtsQDak7ThD3KTutXPzLinDDjyHRvd6mHOlS4scdSD
XgzEQPpYpuaVvnzSyLLWFLJYwkbbi0j0o37rDKcQw4MCZQ+fXEUICOfzLrlYtb8M9TQR65gyWPid
V+SzB7vPwme8pG/dgmtIMqxzC2cAAoxqyExEbkME3Wl6SGm+hUcGMpqFgWbDP37T+b1NMXBQKlRT
WQpqJ549CXIaFzDlf1EVOn2c9tj7zfIkRbB3UCGN9x+C76xv5bfu5YJzcf+WXKfgW81t7CiE0j+D
A8wftxWQp2MFH3NyVz9G6fGaIigiQM6PX1bufHixVjxVNOU5QzjH9OcZZqJUvy7Vs98BKdM6Zt5W
+kplMnw3lBr00NNWwnA0Geus66zFWLwn6wVZpHk0OLyLPFizCUWz4wI4KEDcuRJ0+Z01VFvGn8O1
/HwrV6knHZxXzSuFHoX8bgEEokQ4yOMIkVH1MPrX9DnldXPo6hZszNf25V5taxaHWUguvPF0sKZD
rOBLHZYsbqkvpyJsCbLLlGW9Jgt9JGNTn5Zj17ZxNtNfSACFJEXGjRM130htydAtR8dpUstVQc9c
aZRCee9rSqvul/QT+bozKoPKbr0bK+3qJ50FcDkY4bzECBmUmfZwZqSE2oTZ0TgT+o7tUnugqX1D
/EkwBSmk4AcaszEaKxaaCQeMKzRJZ2PNdrIJT33s0gxLOzwLiVy66lROqzhRL/r8+jgtt02+NPTf
6eUvcaGk/jS98rx04wA3s9CamypzWVLjGAVmB818NQOxz9IJTSRpcLOt2+W7jk3rq4+8LnD4UhLk
2B28Eibk32WqNB2lX+FfMhpb1D3W4UWTeyxhFUiueom+EsOo8Tlbsqh1AnjwXWiM+2jKPzgB5Nxb
buZVhCBIcK1fP6+pwgoZzq1kpnxkUEXCrn6JJul5lVUgqIfdE8cdmFqssl2jO+T6b1zuG2aoBJEg
0nqt7yD0TMuxHIMcZWwMu9sMjUYtYcFXqUR9mtZyHHNXQ0/xU84oABSR/m7BVcAxZRCx/yg2KRwS
/3DGBDHNLFn9Ui12fKWfmstUxoLg3WCZcdsRSPYTb49fxvKuMv4a++qLyTicuAC1cJpepHSxv7yE
/LwtmyrTqLeFNL2T+JLJ/kiW3iqboQjCK/n7NymYyFDqcDNuXAeMr4wXGTlvOb8/xWj6S4JFQd9i
bVUF0lFQOq3Gn/MzkhKX45sbz+/+9Ch2YgYS+2J7M7jID5fcLhAkXQwvK4y2ErZFUWnpWxMp4ICl
Cm3E00EnOGuEaITFiiiXeByoEvvPJli1XOwBwaohgUPQySkfimjF0z0TFbdoqByP+V4v0HIapqo+
YMUt1lc2a4zSfNnXHEJElVbQjeKeMjriaFY14nUWo7gC0SEX0SahCU94KQZXgBAjEjvSv4JLS2z4
fy7UNBw/xzoF1wHIE+iQ6seDgBBr8eZJLebwaqj3OINZGgcQvOFI7AM2gtvz41ECFUX82YwppTFf
TjQ4s2+J0KhRGG3BxLydy66niD6h1iILTKUYZjpnYJ+JbPlxI6gH2lGRstUoM5vBKN0QnylRVyQ/
slGIApUwORhwCZGBdz3iubZAosB41JskXLeWllUMHGjoHet0o3AzbIS0HXUOr92SFSji0UjjU0OA
xSPELJJOWC/wmS8f4lC5wCyKbJ1WBoLf3nBiLmFyMi39KEZjgTTlcdYvDUIF2fcAxjhisLHoJCRi
nPw2N5YHtipr3lU/1k8oZdSJtCFZZbaD4x5Fs14L4s8FJH6i/1bvPwca7OEUr5Omou5tjTgvwrhd
CsH4qv3Y9IN+SiI6hLZN57rEOXHoVFUK0mhq9NWIHaGz1LcrHJ8sfDb0aEbNNRtBQR92y56cEolP
UXKXua0wHvPcv58UpAcPjScufV21ZUd1hL0X2Jfp8oGYrsLkqNafXgs/XKhSxOS1GqbkbifGPc4e
33Yu+2p/PmDi2JOZCJ/8K6H3VPSjPuQgsQ+oz+/0YSTUeF5pB4tLglTMiK2y5s36sCJeYV1qL4rH
UbEMmIwuYwvTm78MM66STOwkibf2XmGP9vKlj8XCBgiqKAKq/PqY42ljWH7B6rTvA/i/PzAGP7zf
PhjLiHv3T8/6B5K93VgkAlFAtaSzFJuf8Of7AcUgsPWmOdelzf38zA4w4e/CpvSN0kgnzMZzprWG
b9sMQuWrnO5bFBEqt4eYqWB7DzwHPohALaJhj7Swvv0HydaJvrLYmSRRM8ZSq5AHgsL8WdnDDJz1
AuLvJZt0677WBOtGBfTgmZviFSMqjRVt4kZuJIl+geyTBANEGZk0jWcSE5yN4qhAbKkrUwQXqmCM
kODMuH/pjy60g/dbbCYkW2LXk5Gpco2RyfqM92dAGtmaIk5456cRXc0AgOpnkJuOQabB+1vb/QVv
6RBobUgcaBzPFA6MoDtvIBKm+B3YrqDOZ3Ph7UPb5ZmwpA41z9npzhAln/lJoLvfX+PqWNFneIho
0jMT253cxAIhxQP/PV2w9cP03rzmDqmGBR7ebKCgdgquBGpzQh41TGgfKIoAn8zaEoEgSO/r9zTB
Ds/eTpyiqCgyA5LD5bjTvFKeqKih5iENDSkeIWKaFpJzxGPKUAxc/KdWWeb8oEPEMECdVStBFpmL
hraLVNmjc1D2rpAQ1y9BtXoZB21qXuMB+kKfQkKIK3pj2P4uLyRE9m5vr5qKWeZ/xIJIx3iFe2TZ
lfdcoOmHj5Z+KJyBNQLyyCxaoGIJ9wMLYSuvesuwlQ//5qUGWtTsX8vZtyFxNvqsc24Tk/lj44AH
at+pytgLgazNekb0t7jHytjpyKH+QGd60LWFPQdw8e/CC1ACWU1u3bOqIlY1jJBfLswGRJtCz0IW
M/NCufJMFAxLqSl1qbb6acEvul+llqZqnNziGOsKtVKD9bm2l/u6qTkIiJNd9czrTBlmXVaykrXh
3fpSqiib9p2OYvAafa3/1VkQoN1OBJBdeFmmu+F6IGDc0JJb2wK3Y/hCcBrv+iYmyAgGmq/SOUuI
HdTZCgEu78W1LlLAwaymVZHCe6kOLUbaozadshAtzpqmDwXIPIYO3Sq1CRDpllESPRNb/PpgBMVs
mARld1Tt0MgElnsmihNFHcJfcCOu6+f0nH7U3mHjvAB88dsUlhFDJu8E36DKC7D/MJ2m4cLEuYuu
OiSt8dHgrYiTU7Wjhb0FPJzNAFoNfnI0rXIvSjoh1sNGCf1+HNHINLRPenGrYAacF1rByfZX8Fil
zVnEePq6qSypLJKtTJzTuF6UWWaO90oK2hndtdkoWlhzvPYS5dD7lhbpWzElIMuQnmeCbS3EoRkZ
o3/v/kzTRI5yHcC1xyaltJVD4tK92XmLKh3kixTadvy/tlBIjmqm3nJdXDhYMbL1hvDxfcuexxi5
Zpli2GYn41CEPNsFlGJw7mMfib/wJbImR5EmidstKZoi+kCb0muliFdbXH3ztmlp9ZXuvgvBNKX3
jJjdmFFCK4F+FbC7FYnDmb/Rd9zwkn136GzjopbeXeqs2tfkoGilNpt8LodRUSiEdJSjIyQHwY0B
FbyFmNasU190usw6wTPaADEe4pQd3eMPZEgezbPxPM2uMhj4zih8HiTDO2m5a9pjsVPmoKH1PVw4
cn9MsAoTO4XW9J3AZHbncx37gN51o7sWb5cPXQWnbP0NH7GXGgwC0jV1wJ6hM3PdIdC0puY+OEvi
bZ1AwltzDsSMTdX/AkpabKk7hyr58t4nhocYUESGHDfBIQZHyGZckuRjGGP2UJmA0hacE4Ly9b/A
gRlhgRgbapsdxMEzFIfhesy51ZfZaV53hfPvYnoj9zonrK+KFjn1/BkrHEqTlTn+/z1RuccwMY8Q
NAoqSo94tx1f6O6V1mvkjfNzqpX40etrbZ6REy2I0u1kH7P5rAIIwLys48RvhE1YOFT4+bzcd24s
uNZJQSC0qPZJrUlZP/VfY67+fvRo9rQ63aC02oOkPgUP1cGtFR47JG+yEs5Q18pR3FUtsehiDBoH
+Nv1qhQSxJcXd24x9L18LV/os4CQR91mE+6u5+1PsKgJCOXQlPwIEy/qcdQ1En/JIa1k5MlNl3ah
fIOsXPP+pr8cTCTc17Xl5WgN31KdKLXwk1iFrfaemCC9HfZa4+aqHwEgKPq6AbLlLR6urTd3K6gg
0XCJHzYW2M3NPKCnVxoxiZV88m8bZ4CEuTuVMs0S4dRLIVseqRtxH1grng8ir3NjEa33eGE4i9MZ
BqOvYLrVUINyo4rqUf2auQi10BHjFFpi6cUOtmIYPtVrbH25sDkV6NbqAt0ehtp6aTXDob8ES2kf
rTxYPLGztU1hZjKALdLirzGGLHRo1cu9F/F4hebhHnIvw1OnkEjuFSEeNu2uLFtBSuZZE33pI93M
R67DAIQmuZgM3TPldNaWUEKx6gNUprMplGHLGpFl8Y/70t6TAqX5F9KWmxvzoyasgwU8Yc+IUqJb
jR+m0lgJz6dCr9be/sTD9aOoSDzM/++giHkNkWsMzOoOQUPw+FfEhVCGvfR5ZNbJ0a0es4ugz+AE
oc3di7U/yh7MMcQQStpw3Zu9G22d+FI8Q64iyUihEyXK4b+TB2BwxpooqrQh8DGnQBvM8uheP8RU
CcMj/uDx6mbFpy77JGX7wTT0fSmzsWzgmGSnS5iFsMrygNCluDvDegDBeUCiRgCvLAMZCCAvm9MJ
vl3PtcEGCP27tjKxLrzdFRYWykzxiwZvU0+g6O+eFVzV1WbkbnW0qp+NDrdB63eXlBHMUep0wDBr
6LjPZ8tFKYHjyHTbSn1cD29nPDDFng0+iLGJlsCMAcYMVfbUjgXbE0Hz1+JGoCLs4R8/s4cvraNl
u12GeBnSU53L+FZER/ea+alWFdrtS1rDu08Qusg6XqiVE87glj8fK8hZndvnoe+3c6D+5mj0sOzG
/cNl3AhMyFme/FrKUbgpfvamr5+8MHnK8vOQuWtTGWRTMiBSjqutlejY/5t1uupzdiu1p1NcSK5Q
R6vxU3NM2fzN13UINMEcQbrdq15HcUZEAJSKK2JIQz6OZP98ZtRqg0gUh/5Y13XHF28gR2vuTjgL
OOkLeswqkIAjORWnmWsX7W8WjlN5e3GnFyXmA+1m7Vn2frZzggn2bnAKzaO6H10omAj7dXQ1KcKj
Tt44NhLQQHs+bKZ9rfd7DGDiHaUjFVCOBdmIPWxdLsgEIJ78vN/D4HLUyQKjKskS8Ny0fuodR8Wa
Yyzhl8w4VzIKagl+5zhAZRXGTK187ci8czIzzF1EzIS0qzkj2BgXGIQqGdmanwBmsWV9VdwYS90l
fUD4rrZ+6Zqq0l73p8LqkAtFt6X6+QD5vj9OhklAX9LGnz6q2A5qpN0xBBozCqKFOTPqkZv7OX4J
1rzPPmzO5I8N8YBwa5ULelqeBJqGSV6K3QpBfP2LX8SM752sKqn2VqBlMipdZqqK//g9tZRWaopb
yuy3cl9SqDIOKgqBepPiFhPRvUVWLU4Maki2WFmrMwekm/GUccLlEzMFNo28zQmv0/jwroxYcEVA
VAOTGYDNaa+b94rYvVDLsVkLckvYwEoagJGtA/XTyBWyL82mdVGxBA2x5weSHpP0ljtw2WtZNtos
SlogBp5ScUW9bi35zQSfjMk1Wao5g6rtti7P8vjRSVWFUowN2NqHAVyFNTsqCzmQLkzQTvlxEhLE
h26gS4JwN9h3y7Q605+SsshSJhLCLBhqYhO/+lD6uNPwMmnEPuUtlXRz0Su7MKga5cCmRdZg0QSw
zDj5+oTgmJK/5vtRNkgU3mGqZXJApy28ZOY/0vgpMvm6nKV/LTyoDsONO+b6CExpnoLU5s88fnGr
ya/6cnTNrCosV2JwUIBLvbKfutdBuy/2sAnN1RVUuzUUeS6fny+KzLRPVBy/zG76DfSUIaHi91qf
WErJ3WZHaUbWcoR5Ww853EC0I8FEzYmcpCVPFCZnMt1+WeM2NnrqGcTLo9ufKJssq9vcfio3W0fB
g8HltQybYFfQqqgK2o8aX/fX4v5r6Aqte4eKGTL8+uWeS5FUhprZYvhRk9sCP3zP5sLMlJv+xl1b
Qsu5lFwf0If5ulBsAQnv8Sh+gF8fRJIhHGEk6xj+3kgZ8tcJukdAd6ht0/ihBayRR+/XpcTZSJn/
6rludZr1pDP6S6KbnNOX93z4sirV+cw23oVLzg97SUYbgZIroYlZcQMoCTvNyphsTxizEVVd91am
lCr1K5QnIF/pN/6Q2IcFHYPEnEFkjwSbt34vGAcnkyD7S+KHuAMg7Y3+esNCKZ6FMidh3ts5Wm9V
q/n6/i6iK9VErjHjvMMbsNMedrQZJ9AtJd/iNXeOyDUjmMbGSYxUdPWfbUEPARtWXuZhj1TxQhzG
swu4f3CbDQYhvnGjFkg7a04PykXpJfu90APociuTa3WYr1Sj7wJQU6uQSkKbJgjnU0v30tI9sKkc
zd7ao5v4AaweHWoQVnlZRCXU7PAHDND/SAj2kRJ0s9ASXkRNvfGXefUgilGbgxhJZ3c5CEN96YF7
l9LBlTimVVNHsdEt7rC8/p3maBE8RVKmgV7i0GB5wmj1qdQCQZugHsYRfyC7qYyYNQbnxob3SGv4
MwpM9ZpwdoZ3+maV3oo/7AXDiyjGzzhiYPv/VfKT0+1FGUbTD+vuaoIO1H0tf6ILs5NnilgokBDX
FrhDm8M5euwssr54+95i9BfUQ5egGN84w9UDIzEF+stS4AiFd5jthgHOKCKyNQvO7hCx4MEC4Sfe
3QWJ36Kkjaw6y+tcGG/dqrnwPuS7nh4m9z9NMsYC48wfpzgHuo3TOkIzC9p126oxAKWlMUnHfpTG
IWBGJsaujjjMdj6Y1x6AVsXHrXbt2kATd4meaCIChO8IqQq7zUZ6G8yCkUXEQfKsC7nhW0lKdg9Z
FAUGRzzMOW7EsxvV9XC5Ck/IbQ2GOKA1a6iUtNrViHVeMx1fmAfDELUZUlOQ60GDnkQN5sWvRzkk
v+Dg8OJ4LNMzP5G/THwbZLICYTtEcC/DaPhXK7/T9Gcghl1QF5BQzUg7xVESSCHKAHW3hQLxGHb+
LqPxXIeU39dfrN6W8BouaekakHhhREdURO2cQ/fb9UtH8XIAr7WF0O0WOLTwqq35SSGXJdbyK29T
bsvEuL/tRW0M3UjfyLAMzrx/YQmH3M7JtV7IFMD+jRfVFTlmWG5W2axCMW54qIulOan6c0UqdPsz
8LUl1P7DoqgsZYO+QkD3TkAvjOYmEcvlz+wb3oD8cGIk3FHKLfECCvfxfr8weyTHq/wzJpgsrUlJ
gEY3dUcscGnW489+j0dqn02Ec4aaMw3Y2EEeB4/1YXoZj5eGjsMSfAhbvLS+bNW+NoxEO7zPN7S8
8yX/g3/hHWe5CEe392nkpXDtPYECKi81KShaoBFlmxb0+e9x9fChW1qXQjR9OEg08s5MozMtWOCx
OatB/hfdozACMHrIrl4DfedzdJR0bPlBR0C7Hi1FWfNWLdHxvAHnUInQn9rPMilZgupN5oq+Nbo6
GU0sETR7TV2SA/S219QVtpsbC8ky6Il00gefNur2T7QVLQNvHLyP70MjYn8wKUSarSrvJSfBYUg5
0VyVQySG2YVYOykyevMpbVH2TzlZ+y0ryI6xxytwjMM2ePTbjwqGzy55GYbH7NvEIF6GogvdPSse
FuSETyrrx5IVy/HXBbCeEa880PnEIzRzYq4lpgWxrXVpB+7lneEyyrPAaXTRhs33NLtmayT5/qox
6vVp52eN4I64aKIL7vl4frJWHnClel4pq/Y1X+VvVN2qPNBg9GpUAK0f88dnQfvJY7/zBfL28iuk
etlrstuHcNq4RFokTMPLZ+HOGVJ+HLvW1nywQ6TJs/oXRrjV5va7pW7wquY2TVaRc2e2O9r49Svf
6HH29D9qsY1fVvrUDCztA4yZjfDYfVDrevkETFUwB3H81xVohL/rIQD6ck2oQLOTvv5aGT0L5sGS
OJZdQ5LYiESBKejrjUunmOixeNYLat5DdMaztSNP29JAzxWWg1wLYT1HoLh6IMzUR5F5LEt1b39O
23Bs/ZeOfY3zxXGMC/kEgoAFwPCmNcZhhjCkWd4pEY4soT8pJPsT3+hppmmBTWl1NhneDjQf7z32
0Q3t/Myjvvw1lcs++m/CJahoqjpbaQlbeurBYzRvQDgGd33aDQ1+E+xYUVKLYoa/mvQIYhdMpuw5
VwHjdxb9d4asW3jYeVJ5r83+QmNNvCnXKs/TcnFZqPnj+UJCcKIB6PpPA69ht5wwLAKJQ58we9Wr
AY0GFAqyYhqwHDdi2ZNLEEybE5o5gxhRMJktdl8PL1po2g/eZiDWwGJ1vTYZX7JPUlCIUFc8pOCQ
lmuSVdSRlwq6DTb2wCpgmLVHNHXHmLNEVHu7waPT2ZwojUT5EJ+5eaAdGOC+fjZZwtQC97gaWnSi
qJw+wrn8kHfUeHagG15eGc2wMyq2rW/xwP6YNavZ19dcYb6LkmZ71rXgyHBcwUSjBqCcw6j9LWym
3ARO9+uTLyREiUQLAQxSDSxWkQxbGXmejEFuuOx2hwkAWrCa8mIzZ/MzJwNfechnO7G18MF0PoYK
eFaL2wer5Hrfp8mMEbeLURNU4LG5JIYPsQr7jp0X3yOSHzdT6fGbCJFQZyYLJrs9fuv0tM3mheer
3imge45Ui+koH2BHbt7NbHaBvcDyYpJ5aSCGP6rtc6ecgfJ2Z7CFu5ONBJ9SK1Ozoj6uLpq0I2MV
IB0y4BmcYEjFkT8DCjWYdfq/wnJ3/TFOh73EI6dKWxAIt8DiqEGFao2LSqtmVEqKd/qEFs9w0+jM
yNKUyZzAphDvbQd7pDrSFPgYxP0Kgkh4t5Xz36Ucvsh+P7Xi9cClrIFrAc6nepZfudOGBL4S4rFw
Do7rHM8T71WSJO5DvxwEmYzGH6fyxGzds3DXU5TiFDwO6s1VAOO3sOhZquvNTcw03BweRqZtXgMh
qDhYA7lmSfE22EKih5SPviMrWd10f7Ah2P3tiosWHwsOTY7BxxRwyqhylDhG2Rzs4K6uSmy76HI1
ZboPtpLXWB/5UJGpxv+HV9VXAC+U4YLMbgLxPhHnrPuaTV741KfZBsHQrpwFM0v9l5XPf3+sOYgL
4i1kKlm1oD4ZDvgQoP8TXoaEzCqozEbjedkDGXCboH+lqnBvvbcYUmIPzqvpfE36dhj/avnMXMyL
MDEq9f5v6dd7K21/JPfyqQmhJqSoAqtTmRuF/kdi9yA1HIf6LxNeT4RIKHB/TS2Aup23+IyjIe9o
Ou3pbleogwQqda2JGFEdJA4KNzF6PT4X/2fvKxJxxbtCKLp9E5hZvDqxG9vAWNdtTAtM2ItaxK8F
TN1YmxiueuyFJIDJKjJCUL6ERWWf6bvKTVopHcvZ+RaYfIN9/IEwxa+K0EUnOSEwO/TtiSZ/Vq9N
zu1DzcAtDSCbmsDt34ic6iWa9ZuwxAC33dy1puYjGoH8sbqhlI1KM3KRpurBupmdPGJCk9veAHRo
wmu5txq88hMYPIsUhsQ4fUk0eMZvbmt+bMCByded+m/DDegKsGG7HGKkGTzkGfXiZWeQcERGbNsl
WGvFSSPjGHkFSO6+dK+rEc0LpgCyhVjOdCiwQlfi2IHECUJAh0Y3cY1qrEFbo6AgKy9iytMKhjeu
f/PKp5N+8CC2+YrLnH7JQ7V1odcfIGGPGbot7VcYOyOWWCgAP7C0lwOwBSUWoT5ZCgDdE8VAzUpa
TqZPevXC43CMAx1bESMTI5YmM2Y+hZvqwpo+rW+P5FnNq9zX+pvFh6kcIz1G5J7SG7kcAsg0pTUN
hzPCsjE0aUzNVRZpLGntZl2UaKXR+m7Gbjegt4FnmO3Sn231DR38Fzbxk+wG+hGRpYmbxCKg0qtx
rd3cHGUD/6aOuwLfdOdQQ7Veww45T1VkN4z5yA4r9FBMqHnlPb5hEyOU6p8zcW0QtElYlRz1NWsG
kXlgfOlIvNoErwGJNmvfVhGBFTyzX1S612cLAaUZxDn8IVJqy5trSzCjqwnTatIsYpKI0EUoNqV6
G/udSDhRlHrIRuUsa4snPNUXtDdKqAYUh8hpPAY2ol85rWtfnYn95LsNahsGj8GuyPmd3nSbNtGu
ux0Xkj7ukhl49/ujo4LUbfB6rUDUhUFMAiblfv1qFLbQNKlRMBHUXL8/5HO3zUBG/5udJS0G0BEz
861LzkjMvn8Kmde/czU9WnjQYFwpDyOcwfUjeoUwvX/iB9I1f/W860+wXazFrUgrzJJ6+rtIgUyM
ZaZHcTro2GPovxRxaVCwldE7x0QNZkBhvRp8X068TvWCkGS+jh8UohYwSa0lRSrPV4E+Um23TBx2
woWAW6Y51S6blPp22rxfqdzc71Gch7j80S1cttjV4sC4n+2yEU7xFjCxLdWkvZkCLvMX8Kx0NKKh
7yn+Ywr2sMNyeHEQPqRKYvR1tU6pDUpQooaQVZULe99a39wsHRs3LQ7gTGzxDHcyw2/t2DQLnt8m
o8m7DGR1G/N44SUDqHiFHN1t17GPwKz6MFUUgEYYM90WQPgmvXQeIXBtYnB+28q8qgeV6lgblZKd
gGN5NovCzytXY+ki5V7GmsnOl0PbnqM9pxXE1keEgq93pufb/3qGIBV1e0miV86+GVNiT9CQXJmQ
CLJsRM0Z7e9RXrMjKuexX7G8srL0oW2MaXOT130NjMSLcPx9Un8Mycr8heqGIiB+JI4T7GXw2mDu
pGjFZ7TwdtF94bn7Ocy0PE/cBsdx+Nh9rvDl3PxC8LpPgbHJIcfAWl6vqjsbA6vZxdfMmnmNDyF3
gEJlKMRoyPE1wD3aSvCeijqr4DO9UxSlG4mlsR4nr6Ux44kyAy3KjkxtrIj0eim7jZr3cDApuO9S
f3XKoqcV/Vmtq6GxnaQCiuk0iDKOVmnGEoGHwyZg7MtF3BCcZ17Lhd98feDVwaho2PIuMCMZ0MGc
vHFs7HNqOSI5S+Qc+JWR/ZknGgFIjUlpgPBXOqItfCiG1DL7AbUym9eltTfFG4CWz8cQhSqn2z6T
BYs/AvsQa1zaQDx9wTkvU1BrjKzlbeXz7fvMzcRRLeccYF5WTrwxGUB0ktuCuUIM7wmH8f6q8Axa
/f6qkxoUOxdSAAupqJHopG9jZXoWTLTp8QwUOSzVaUFUdbV+Nk/taB8F0QHRZ5ZzbY6JlxWlFAg+
x5O5fi0rLh8P4yH6BC654TupyiPNuAy0NGzt44oamCgSk7C+RClJnlvSjYi50gbzdYuZfkSfyom4
bH2F4hAQKZPZoGuwnJin0FIJkcGOvXCM9RqqYSdoxibhRr4HQKAG+pCJjAIbvItvqky7uULliMP8
d5OOaCpVzI7yZ55teryRIE5WwAwUqhZ5Ch9V2phCZLTF+qcE+a6sKtBQKs8y+kgbylFza284brjx
mNyWxBJcKq4OaMvFabsZCuk66HodG7q08p1U46zHToGEAEQX2hSQYwWCgqDyMjp/nqXx1IVn7LvF
LL58B8R6nd1F+Xy3kDA2jUkjJrTX9oobFC2uUmOzMMwEgtQ40GpkYHfDtunMDxQfgiOvuB5yc5s7
xJGoZmiG2Ls5VPVI9TQOo7SkkzJhxHRrgNfmkGI8Z7GRJUwtupFgXT2/jgdoQAuzdQwV8xQ4bUyE
bI9NXIUT9ZgdOGbHdxF/LelbnHad+sNROYofQMw7xyddR0eWZ6oqXjk1+/47OGtNviwD+rmgHzSC
LwV2+T3lVFZzqqsIlLAT3L5reKrstxAjZ6MLZfhZlhGjipfSWY0/c63i/xYb88qK1k7CeuSyylqX
aeHuXm/IIJItm4DQHNeXGmuvbebRnm93MDN5g1M04bklhbKtf0OsrSOP2CR2qOrvujtD7peHNARf
P0WSCSWxmeyj+pLQHMAMG8fqleQj24dy3fEaU/sm05451VrFu/gSZGwJ4O37AZweg3CtLUTD9DLQ
zFHBva5HNnIp1rPK9EuE2LTsKzp3ZohrGv9202c3zLLUFZAZ8IbCpq8FadRDH2REA5oQpEV67abN
fXKAHdRurlHObOrrJxhQKHrhRrDmbB63Yn8DjHG5WTCUxotN6ZyGn+0l3f+NSoL5DNMjKJQe2Eww
WxmvQ0WzEmnV2KMguK7HJ48/Va3eiuHEh5uD9uUb5a/loEiV4FEJ1WLtReCKloBi00as4s+PtrnI
0KuC7Z6xjEHL4HSVUpAdXV3HK1oSWzMI3walitFje8EmMKQRcECH+X/SicoZ8YkO6zBqajBAqnqJ
I/bIsUgRrJpJyv7TEi+29SSss5jaktEZeTN4CpF08aZNL8018rkZ0Li2/uJpSTVLIQhYuBd3uir3
NdOusxXqUwvyCtzSJPx8ZEFdxHhHcFnX03yRgZY2PMZbZTeDh1UNDfF41QWs/gosERSbAoa5YQ6S
7iGWK2Roecaz9Es63QrDlkeRcbHgEL2G9cMdJxwhqz4jklEV453OeTeYCvVuJa2RTYGwj4AkFoIN
fxXt13OJVx4KVPM16ygw6Jgt0+5nA0A8fsVVHPB1NIQ8xxDCYDe/34NwhAY2fgG+k9l7FRfJwKdd
9qRKtewPxVeTIgY6gqXbB6Bm5VizQySbeuTxjeMoDdmcys9Z1AHEHuR97jeujgJ2kx2QcPbMcfII
vbzsGv23UoC6RuhHx9J4ZS2KFt57HVrmLsEKcQ+5QUaOb6lTYSGvYwkMvUUFbssx0HOdI7DFW1Xd
ReBdgOo3roPy+F4QknHPcod/zxce0wcxjWw6elh4QMjxGxqkatu8DnW+QgQVO1viobzwTv4zhKAL
ZDJglUhjW6qT7ldCJ/Sc+d2hgqlx97DXlwthj4NzbsHEMrwtO1odhGEBB6+g9DoOIC25+BmNtdNg
kDMKLlFNQR0d2S93xaXBacfh3N9EEw/EblL6hW0Qvwh2RTYfNm6QcGYs5fc5lxq1oMuMgmZ4BRGB
8w6J750sZboTxj5CRZSFAVH2Z4FhiNe0Z74aNPpWIlTZ+FSFp/QJ97+s7blY6RPVnV+8JTzrh5sK
i92ffLq2+c9/e5Ih001N9HIYVkNIffeAarhoP/vqfrNHU5EKxMfSWkwDUKmA7+POdTkYBIsftBAd
SsvHiW/083LLwGd5xfqi+uL5OvYvQZbFls0I8l/dt/o3qPvPTORn0DzzzHjVsqImRZqWGVrhhIxk
TRvaTCQDUxBO9OBzluU7Nx3SXAlKB2ERKAWxKOleacURKebVoLgsXYw/BWuU0J5k+8nUMPHsV+HF
fH7yUOWCToqtUiyvi190ySJERCSvJJ2nR67ItI+z0uxr+lFGGqToTBrM8xPa9iz4r0zCQz/y+AZN
Ewb3RffOGcnCvyt+BdCQSs5WMlQRNLSBIGMHGI6f6DPIhbblkM06lFlG/vWHnfPoiE3OS1Zn5JsO
e9VFBywplHY9Cm35ULKmmdKf0UHUiFW3HyL0RByD6mESovc8XOF9voyg7rKMJAV9bwpH0I+Phcy9
reowUNpWWgMwzClZmE05v2Mgp/zwuI/xPoL9UXz+z/jF3NIfIRft7IG+jG1KRRuMjNPkvbD59ku2
8cXoAoS737s/ooyKGD1X6HEAy3XTl5+QGreCCZ0XOD7+KmI+PNpSZh4jlAtpEDP5jHM2ooDJm56G
hA3AEeNtC6uMbVZKKzq90DVY13s+z/spPF+yCNRiQoBW2PbTTjj7YZTCLb7capuIX4SD/gLPgcPq
wzBC5Yc0S1FX362BtMLNFvdbcEWY2PdgBpGR83JfNjLRi17NLgAkMfEpWKZuwEXb948n2MXrAwoJ
UtpGuv+4iQ3tjo1Es6+LBkNAww4z2CNeVWYCRHSuDAKU60hGQ00qz1EGGgm+pfVxYS3MSEsAKixK
0YgSiOVcKtxUFo4k2bNBfAxCFekybElZCpFNwHkgRrenfFKgd3hkStbfFKFFfi2PlbD8vyJ7pNj+
C1han2cyKAnK92pukhct/5aGXN0TyZOnEhzJJxkQNi4fEQ76VVYiA7fE4H443RFnfCl7f3037FXd
bgV+up7x987GJ7nq8odPPMt3/dwH0bc0Y+9N14QNt73VeM+wUVVywEBD20vndMgajr3QQb4t9Rn6
naXlkn67cG8SE++4b3rnVKwnGSrAVlJ6gx4vYMpXc/0dEDPuWTBwxrna07Jph492INc28zvbDXfO
3FrMD9wMGSciHpHA8R4CdhnmXxP2oz5Mmxz07kWBcCac930goEY6UCKj+YJO0E/LrfjBJVYjDOCN
bUj/f2XYGzmfYxjzMNKtX8A+mUczv4qpMwa1WDM/7K3vYQRxyRMSK3W2eawh84qd0GLCCYspSBr3
6yiULwz1j0+ey4aJgwIB92NZJZW4XyqQj6mVR1SPaXrWmlgIYpS5RGirR/fpi9RfXltPkdhAfTop
dFSYOxAhrdfv0HgCC+LL4c2TWP5wNhV9Sl0fQyDrmQsmREO8T3lZBoVmwFjuZr31ZtZhd9kdAFns
pmXEX7pWCQWLvtr1mRunMLtDqgOq8BNayVPchm1jPQJHS/t3hZUJorWt4WZoWaXgtKPSyrTFjGyL
zuNcckPqVt3tC35nBxrQoem4xoT9Yx/QpRbcXr5SVOddkoswlhYkzJL+Qo2rd3MApEjbzw8W68KZ
jExSOEYH0yrlW0iTNu5pIeYrcceDsiGHiL3+pAgOtxzExuLR7rHtoDc8yIdi3n5kOtQ8kzOl/SgD
jy+RsGm6cngrHCigFJrIjluqZT+c+1jpgxMscQHwGSl17sDhwI0cKxSrE9tkhB7nuabdMyRQc+k0
d0zHVRk8OFE9rQKRnJ32Q9OpQm6IbAkX4h41k2nIwplZwdJ3jMmUZ1LZnpe3nfJyGfE0G1lWwzNN
K7/zTuSe40ruQVlNzewxklj0M4Px69R8QwOald0HJIUDNkMtTDzL08uUp3abdmit777ha7fVJB2R
z1F5vmkbO5dV0s9ikmuUXAl2QaRgLanOaHhtxJUG1c5GwoI+G/hXdZzKUsQvdEHsK69CJsIxD6xV
GMYrx+PcmHpv4CTzCd2f7Gkj1ngdsIYSnC5jpNL+jJemTgAeju3aZPMKTpiBoOp9TT/VBnsT3k95
W+wH0P/rFdBvDrT+rmqdceed9c5nuNMfdOZgOuBUUn/COHjn3JfZ4lKAZcjBlQHT164KeCUUi8Z1
/hhc4T8t6iO9pltE/FTc+w30+5s2pl6VG9oEeyRQ+LgAr0n1EKtbAFRKLkVdtQzeE0WHzmjdajTH
5HQGU5d9DQI0IYIPBVx7HVwXXzkyMQFh7G3j8wg4U75Z9oGNchzA3xlcHdC4Km5EQoI2SM/qQczo
E5kigDG4E49VLEskpel8gXbqTlce5gGFbSdZgJAF5l6weM3XKtbat4DcaFNXXMsdrsMj+cPSrXxQ
sQ7CEnoqNXTQltj8sEWbegFMUyFLoPRC3537OGXLG1zhCs8FbHdwmze35ld1XhWznDGmXq9vimMc
wHRuulKK9fOr1CivTB0KvBm1wIEFQ7qqiF+OGt6WD7TJWH/x1k/vKr8uwBVJvV1w7k1JnTBuPv+/
Dx2X3TJCtyNAYobIxN+zdxPdgO4zCT4raOSEgYDerDUq1MzWSq3qLen5YaNjQCHSYIjw5b4Tvwrw
57am1eQAj2OGWmEdTweYWzO0imjfKdGB1xVd78zKTtPm85ZDTbrAVcmNI3uZW9if0/yMmjaGQg8R
LNWupqjykKi4hYyWYu2gh2aufJ549h5kWtGSLPOkG/5bDg3bLY2cZuFk+Q0rcrrL/PYxGvw9wtFV
9mhaw+19d/E57sb0SgOQi2F9vGCYPWE5fWJB+4Y81nGGUaEKBxG7sMJmVKgh9Tv5y+R5hJOpYXeD
oss2WO6mC2RF1cN/DHGLkSVMJdmA2Dzo9Yv1lnzuCBCuWZIz9/cK6pJ2FjUjfLSYMxnEsdFk+2D9
wzY0fp4/zdz8hiFgTFOQZMUXUewtoZ5e1H7MHgoimv/V5SQVhzKc9GUYP90JzGntRPy92QQuC+Z3
Lwe1bWQl8Ft+OfdomwjRBp/XKwH11O/eRWXPUtXVbpfp/uYCgH1M507C8zcwru6MGfp7M96BeR2I
oN0v4NUk2S+Ovrv1ZQrGAOSjDk6G6j5+C0G5C+1WsBd1RR2U3YVt2DJQ2cxYis7QRnPjjHLwBjV1
QXjKUVxExS8aPMkyl5PgbAobP/8uFphlgV0313gd+HC83D9+B3LTIWMql/S+bWvthPUlFVLtAlQr
ZzmPJdayg1nwjPkRT1h8BCO4u9xZ1I7/NTTNVPBw1WpO6gDvMmqfeRB5gPROpWcFq5Pb58yJbCuX
bXamyhrx+TmjkJGzE47Q5PcnRybseKPzjiRevKBYlA7LS9U6NcHkymGbEhGp4nFZ8yuCbXhxc/d1
RMNn3Yi4j4NJYte84b+fr7UUa8uVatCfHBakA1PCNdkDxCiACg5PIPZ4aT5u9wPwAHkmc31Yt2/m
H+kqvBiihd9AhvvOI5zGyKT1SdqPbX/wUJO/qLd92+NCkVShAK9Usov+Pk16AoxHTUlwxnMEJeVT
khmnWl4v9g28ENt5+jhiMOgiFxqh/WGyr2fHzcmlOU8j941bAzMgyn8s8GmOsWHE9jzS7srGZhCE
47fqg1FN7Auj4G7S0e0TZwFP3zQjXv/BMEgZw4u1bsQv1v/9SPDtBRmndedu6eJHem315E63rVzT
as/8KSsBAq+eFenVPm9iWCzjiMivdmZiJZ/Z3Wnt5RsUnqyo0RxrA8Ai17BrNvQn5+bU+lC5UoMs
80a868/CAF26BUGBwJg1PlTYzVPodWTaqLfyV9/Yl5/6JHuWg16NqhZtT5NUs4hMWxRsuFO4WhUX
pBtYBsmlPaQbV9dhmU28RiDmJ/Je3b5lSodmG/8E5lG2j8Lh9KBHoNza3uobyO51AP9yL2BFBAC3
vGkob+4jFnw1jlofjZKh9advBfGAff/d0sm0cDMdmPv1TpZ1aXOERw/qLBtZbbOpVNGEihVaQkAR
o/dvBbRwOxc9AyK3zpBJKXB8UmZqzlR8nt5xbU5Zn7Ui7po/uY/9gqJE9+VbnirNtk4yYm2xvLI/
nrZTgw4a0Y7rdjWAKrACD4GhuHywobj/N1mI0JbASdiDQJD2+hZsORf5Un0JUkTlDF9RWUJN1In/
MXc1JpZ5rBPvxx66ZpRjaXK7Ouo7I12PGXB1911Fa4RL/Nreu3tPMZjiwyiDqJlOxruxWnlXsp2I
pKajSjdw5HjNJ7FEmbqB1sLWhNM49HksXtkgn0BHgmXboNsSuS7VRE3ZpSd71hPi5WLHahKmnHhn
5wnXzUMOI1Z0WrHIkt0AA9u2ER4KmoX/DaId8Bm8Z6OOw2e9GRuoL16bntaKXTnUbY0JoNE75VMf
euBgw4o7Gpwh79GkXNxa6npc7fu+gLY8ZT0sfuCcm2Wq3tJmZqo8IhEUYyYodna151k2eoD9ZD4H
RpJJvzPjl2QpoPMmn3+Y6jyRcNtNuuCzga9LTeOKpad4yaEuox5fNlfcppwC0eJDDTiyfC6YdI8D
R9svKxrQdiaoJtGu/XG4ajpsFfzhyGHzc50ePLUe0ml6gE2/JuwzEzDVypnU0HWvtVXI1E+Iiquo
5y4ZCsiqQJX3IVc+FdwRiHxNN2j7vncfG3EpOGRCsGuSzy8A0okw/9282lj8ssfGPj6X4wDN6vS9
XY9lkBw8Q18P91lTmU8Gc0bDlvEV7gyy7DzFPt6bKYFFQLvbpB6Mlf6FBUoFdoqmG+EhLCP3vFHD
+9lpyCMlZWk11TNzu3pFFgmlE1ODqB11RQ0PMuID++iUK1UuP8kNkg5zwwr/x6o24cZwawa5KeoC
vD06PPBXaXbt8cbtnqpGXDabcWQDVLS9lKX+4J7/3qr5qS9vEmaIj5wUXq6YYa/44e3T0+Fcm9iX
S2Hwh/tUL/TKzuSLfB4RCQJZmW5WcLxGj6eRx3g9oNbmauWxhezuHyn2SPm5hGQI26jy5GseJOaE
59Ft1vKKscnCzWYM9N9Uf7sSzysFWYn/JS8xA6BArcZ7OlCkrChRsvA/g7v5EysWoLIK1406U1Ma
f/l7GHxpNHgmKa4UmBBp5yjF1T0cXzyfUFB7QdN6TkLCgs4PaxlpVKRzJ7Yp5+eT3f+Uk1+DOlrG
Hp7DwjtUrVmgn5f3dYRAhuBisY9RvGiRCqoXCywOV+04Fes7/WE8dGP/5YemuarpG9LcYns/Ig5q
bbaiNG9j5taiBZNPYDQe1+AXbABS+NjyNr2yMBT8bpscYN8OsckHaKACOa0Dsl5Qbpsne7r1/6q/
hCR3icZa3qiEoGYu3vxvfM5uqI3znm7FDh/jpeeeQ6t/EqS4TVamifmq5kUHgpdLhiIO5A5JKkg5
B14bFQO8C6d6Pn2AHhp3mec5v/2h2zOxUsCR5rjwNulcPYsM1PWSSbGOHC+5OmsNDbgfPnHhP5wW
Qy50QaR7d5T0Lkv0n4yAC1KsvIjkDYHTYLlf4i1yCeaPeU3rgbiOBIqMXdrlakVm1Jsz8ppYaCwY
WnWr1Mnle3YJ9tTjyA2W6BEthcvJenF2NWWJnz15/8A0b4+sBsFg8XUEc3/HOssc0vz3vMnwYsyH
VdRDO+9n5kbYjK1rvQswoqeDg3Eg/23iwturSVAvvNTJcBB4U7l/YSlOn9WkR/3CxLqjAYgg/5yJ
uf1jQfNlg3Q/hJ9ucMmyAdIdYGAYA55dklTNXBAb9tZay4ePfZTKk6c9eDscGQss/1TJO76ANULH
DXlTq0ArcXu6PNU29nSsiOyZjBvfKPTGCy3/HDzhZBT4pKrVQ5nPihGK68MZ3Y4HCjBTh3l3e60d
C6t9ZK6VMHIT9HnOxse8wBKIllqdEoQiink/JL6US+1eDytcfigklySIGVJzXH5GHK1bOH4jwnWd
316iIXnoKAvzd3IsOFhZrLMkgkCPY7TAgSjbA5EcFPj7+jVBNUrtaLBCAy5x8zHgszHQqCTRxQ9C
rGIWAphpKGmfmJLc6TzU8VZuJCMdXiWrl0e9cbEGWm1Ic2KdsNHmUMGnwdJgkM/Gk58aNTg/CzEZ
oRUCyDSqPa4WO9joFl/wJ1g6RgHGzuDZ0ymLSBEuiincENnxLOmVhaRX32MBUssBKdN3DxztbY1z
6V3YFq0B00Exbz8tBlnTc4Od6dCikSvNE/gvirKWfot1tUgi2dOMFPgVPHc5HaiMFlZSq55pN2pu
oIPFPQ4zFnz37dhLSP07Ywt7VPJ+OorE9b/lvW3/Q/QGZ1qqsza03HeoRdlkFF6bbtnYrdfrDiX6
px4drj+rVfKjYWWaGVfdRmQZTXWuPdyt4lVvmorlavMVJlj2b4fcb0wrrbdvXcJSk2hVQUNIMix3
qsFpiQeYQ+x66h0qFpIfoHMFUHUAIg0i28b53EN4Z10zed4pzcqrhr/QHco3yyimHyZTz3iRCmka
jTHPY2vq/RUvnrgDLaAXbaYsPCl7Jch6aul/xl90G/46TrWg8JNiSUF1KnB6vJeTGiSJjmQM9vZd
2OSSR4I4tceTOk66dk2rVl2I+DrwONuOjNR47TRYFyK4mqi0zv2Qgf9x7/rqH3Ib+5/C7jME1Zrq
2FSZLe+ZhazOa1cWXlrSilNo8AYgsCWcZcQEqmxq/NhujH+sTZs2j1NwHLn0fYF+WPDHoyLoliOh
qFsml9roT/fyMI8cEAc+np0ODIwlfviEu/k01eKh9768m2Ca76fvDAVxKlAy1f550oTNMc7q8TwS
AMCM8FUb6hDSw47MwIaOvXE52i4xnddaKXletNBTyA3g3fYZOfM1tetgbCOJnAmwGwnutRHJMMyS
vZR7Zbhcw3xT8Mrd1NW8u4yq4GpnsD8p6KxhViydgLcdRBatuNUHa6RRXkM238I3ZlT4EVPvMws6
Ldrrf1Bfmp5VlfU6QwfoRNe8N032MS4FrHsw6R1qcAIsYcSj+MagWiWbcVAI8uDsXBOKG2Fd3GJD
tQGS2jzfFSIb4a5GPCpM6ipXzHF8dvL24fRn5rC2p9J9fLkilx++BXg8gL7jgYVyn37wwUv9MyEE
KZi7IjQjPSkjkRSErW4zaLfDRjRmtcB/2b57+t992ywM+uAmoY4QY+LDGDy59hfTMyepMPB3/hF8
Wu8tjxfHFbmDcsZ0QZhY9gH6BH8K9VfrYZ/3oUEAgAgKw0eHBtzQq7WGHokAgB2VwkW83jojDkLd
JBgJlXcOqyMZmcC2pB01SaUYP9HLEhdZ9fI4zOUOnLRyCwVc4Fw+t/ANRqbBgXzQt4ycU0CPZ1Hy
f0EHECwc6qcxl2q3lsw5TJHFe8Ajmwdsnp03wq8ywLrn+KM7V+D4cyxwaMGXlgTRFmCV/rHncHVW
JWYlL1dY6LVCBdsEATF7uwrYPGNCVa6YxdYuU7s7k7GJ5y3Q4AHe4it0DhFCLLs3NeUJcykxgMYi
Vtv53ZK+WAiA98MW3X+HbWHhMkugEWbl1XxtRAk8qQwpGjvdfOt+McXCUQWXA6xS4Dl3KgZYXhtt
vEA411d8cO8hQRiQA0RUYIUaaxS4SGpcjSSxaDCgwhk0UaZIYC1T1yQ/PERICkn38AXEyL9Pb8zl
6HS6ryPCDgbBnW268oZ0obv5PpvK6MKUtT2KJsgyJ3urX4p7+SisL+Ndg1iB+CA2nBumwCpOp6gh
aKstqFEERpXGJqvCYx+Ag1wF57Dgik6l2UslRaELf+MBsa7R/ibJkMD1FpAFWXo9R5IYcGd5Apew
JsSNL95NWwaCG4QOdZUy/uCXFV5Zt81SApkIRO1rvsrjGqBhVKBfJ82TPW5yHOBitKSL1LWaYR2N
lAoHOLoNsdaoUE2F3KTc3xRLcYH21ZHRdWsaN+spgRmUZQvdCSd2HKiHN6A+hkGWWxEtqRO/ZxkJ
spIbtZ5xJ8rpaRBJb7UFAFc3eQDejZ3vageNSfdk4zmv4sEQV9SACw2ncGl0ubXB/Z0ohqQ8Hm07
lsgIwKrYbL71imGYfg00zZD5Kp0pqDwFHOcoBfWf/W7DBBJ2meDfN15ilwS4XxASSk6VUoB82WF+
7cdx8Pn+UEtz2aCv7l4g+VDakCwIo0/X1pzd6fU4oLzrPW4rBDvj7m6xJ91PJHrFSziZcxeoF92/
NKKjp+cEeNyj/e8MMXxKfUo1sqQXGmVblU2gyKxYPcIJXFGP999HkTzYqa//ehB3zVaETYUrC1cD
ozNJJGWZBothw23OPxS5D5n2SKzsGFv5xcxJMMWYH0EywnA2t9K3wo6NbJhjs0yh7dV383EmC1Ah
QgcwQkJSs1iPFhvO6YirOsdzejpVfeb2D85ckb+9s5plwqCOl65nqTFRCTPFREdhRIHnBZhknrYf
p3X5zLhB7/bu7ujMWaNwhrakNiYuOJBsc8tFHuk7tLbmz1VS8owCDe3zbjotXX9QWnIcVmzh8pV5
3c9A7/ZazrIfy6FEUtsQtIV2Hz694ltOdscm+MM74nfSQTrFxqIZ3vOTiP2vsgpMpPcNdU11a2MS
yYj5cP1pzD0k79AVVGuSFV6bC/XiybTeV4LHbY+Z+6JJx9DmfuS9OwOTgdkGAL38nMsvGXh1snpW
4K5i8YHvBp6fxS3TJCeS0SMFE+55abZw+xaU3UfcpozeDnDT84Rx2Tpg3A0Ihxv4fXrAOzKPAN7+
41TKnAwVHqOsN3QKRyAI4SJTfJyZDSdHC/yN2mxqvFk2feIGujSeW/gDUGw11dUwMnpZSP+gvYws
FfSUurvM9x3CVzyw7AZR6VqO/ceHG41r0bFx7irw4qAA1oOINrKDZCLqLmxz83gCvXS+qHHr6lPo
qW/prn4E2We74+lniS0pGAvfTbmwy85mbznh1GZQMoh+DECiG58+HmncDhZZ4RGmTEVeCYwTrXcg
dWuQRsGSFvEDha26Nhea8NrVAFuFv2XNuc9e9qtH59xng1FbzTO3jkDWP5KYg2m3wgimHRBfY3Cz
07UTLQj7bEa7XstLAD/90VwlmQDLcnz307Qf8pB3+U/JUJLZdF8m/yIi8uHkEPczvu5leDhGjDY9
fOPw9Owf3mzhq/+Zy+XkfaRWVI87bgaw/gx7SJT1kUKNxw6Cmp0xs942KSjWqwKa/L7WLVFXxzPH
7rDFhViae0Hov6D71SHy9O5z4ccPMgVm+7bEqbuLFRJM5gdpM6i2/ClPoq/vfHGQ9DEzYZb2c4zU
3pT0PBKy09ku9S5q0z28aN+vAA5WCJefoZZzlcYwDXPi1mzEYxneW9ZAqjM/bg9ldGljs0Myf9ye
gWS73cr9OYVihcH04gqwqJtM2ynXvPbcPTX4gyfNfe4ECTVr9N8irWqrHDYoErmuvcuE8fmibxqn
gWs6khGKzqhzit/saRo7HZ+TwoHWnJRUEsHqPwmzkUYuG4s8REiT6BKZ+myMsUOU6Oi/ivBS08M8
/NXS2uqD0DJDRndOTxzfDHl97UK4AZl0GfcH+uAw9jl6pfelxHOmLJb5QHeuKMjsmF6aybbh1aHj
byDsRXlxVvHHFkz0yaXuwdBYVS+UgkAfv4bbx9ds6DutfYpByF6b6M9TIyapkejnFOcjqmucrtZi
JE1bfqlctiEYPXwla2Zp7ds9ezjZjyOXMLe07btFpqhqS+A8qaOdvheoSJjVxGyhOFtjgL/0o5QI
5JbH/M9DBb9hoX3KLFnH3MyqlKk6YWlfL7bZGV+Q6dlfVMZ5lxl9H4OfatXbImUy4mhhXJkngr8r
vUJoGjBQsy2uwIGpkHaU7Cd9dpK3wwT6SRI/ZxS+ccb6InZu+WeKjJ8c2P+/jQwyG4PCKyJEMVew
w0xoqbCx4LrQKP67QdM1Yo+VPEVimJPJ/NZsQfp1/Fjhgg9xLQ7+tIbeVsA/uRtZdlKhBfbyLFEN
fkuD61NV+KGlXgBUkr1iKwb4k0JJWsuJbdilSLBnaG4xFN+/7xZuHntnVnjuHRs/XJyFGEHWo912
hElDA3Wfv+sogzbSjw0d6Ae5xNnRgzmAgQScuzfqthKbNP5bBobHNmzyk0NAyDPSpjmP9kOSGpTM
A63UFqlmwitcxokxxssfEGLpyF+gaCUc27f/hTxUXO6yN8Ib8k/JBNrRT6CxRGHa4GwWGD9NFklh
kOTK3b5C8YW1BOx0qRtXYxHmmYK2CDCr+iwKvU95aRTx2F9FQoizpBXKaTw30+xAkVjWya1r1zYT
AreWvcXbeyEB5dDC7MbBBsd5g8ReOduaxIYAe2Xf97I9ZOZb9uu2GrI0NEN/Yrs8DRUu6ryUvmF+
hhnrGvLyYZaaAf+9s126LkcRHLnFHKScczzoYq2NXK678i3RTkxO7J72fMYtqpzxzb4/1t1VtR+B
2c7QURY4+G6EWw5UMlKouLh/s7hHozjoUFJpglkvGhLnyJixVWNt2GYcOLz9/2KU3v+rYtwHeUdO
kyp2ptVdUEEzzdDV9x+Zx2arBu6bwUgTH50AVGQDXTM1nYAyYWXg8v2VG2TuZ2JImqp+cd1d576+
DATTTZJxwEjJVhjCcKYR7dSAqVEfaJ/NdQu6MyO9aLKrzgh3n8yTu/gyozU/UfULZaljP9HS5MaA
Nq2Xrghea7TQaeJjbCLN9KOVwr7CuXsQw+vPjBC5gvJwKfA2lIG9d94bzQAOMeUd8UhTC3YqCtt+
YCV2FyqCQQl/ZHPXyb2F6hIb84kzO2ifpMaV1B5wL9s8TxpBLNrGfE+V0gDuPo0IM2t2BwQEcALq
PR4qpCODgSdqAL6cQfXMCXh1wZ57Rx6xG+KyKF/F5B8yQ8ZUK7qENfXslk8cPcM8vw1MuN0vHMYd
yUqc25HfrhiCmDyu52W0daIz+ZJR+9ukj6L2IlfmdvyJWna4TnhnFfGw03PgbtJXs8mKC6u1I6xG
2t0IHtgRjkVv9lwCRn7TDaWNPVNf2/AS/Cr3uAIq/bgDJPRxGyhr7yhq4FZS/+jYaxUCsOuFnXWg
sDcZf42E+MbI6W/oicg6YYPGx/tf/gujUiKRWRNkt/a1T3ueOrPuZk3oVaDxK+glKmLTfsOABw3M
zIF4XX8pXtfO9Z4fOgrPzjJmyOyqLMdgNfvQscruyJPkT8biU0BAZyUHTsbtfwf6ldKCfV/iSoCZ
vR9HwGgQ15xmhBQseI56ABSh+hZHb69TzQ8L3df2tb/qV+GnUutNPJW7Udd9rVddFX9Tv7EdCZQj
NqU/Fd54GIQQ2/ka+QUVjHhXqK2V+JUw6y0jXQ+hQr3Jqw/3v+u1zH3eGgMs54WxCNmt96pOhtXn
fQ/mqhwgqbjdqhPcgvCZkGFHuK2yvkp1MTCHaI/QrBefUDVuRxlfSdA7NOQok+w7ZFtQru8Bidu0
8aJqIJEv18RnfYlo9IAy+4X36hTreerz7xEYDAW/YXk2CYyVi/sR9vDQM1d5SR5U9lakjgyN6vxa
9LCDlRIQA9P3jMWeKEYKBRBL4brRWhM/6Pmd0VKrtp/wAmVQFmF/KMNgxEER+1HYgwJn6n7BLvOd
SHTc1iucy1IObL7PHPwZ67McD/qEVbR+Oi7SakkkYJ8ZLmrtiL7G7ajBzmzCv2pFIB0wsjWKJS56
7HCB6QEqbHDK2WcFkYp+0+8K7fOk6ejU42IAKWWq/O9vRQKJdFMNz+DeJ9YXdmEzDEDkhvoT2h/o
ONW5yMO5nhiZ9XTHltQRrqNAlwsh6KYzxzsr58EILPEhDote4ztLH6n1ty6z6NvLUoxXZaaQQM+I
zUzt0HNHBP07jUSDk6TKpG2XlHjnhXhWAug/U3HQDiDhVmag3nuB/s+8zmLU3TWQZPGqDxOU+vof
WVB2XpPfNN/DvLlAFXbKaYYlwJKCyLnmKcGGNnJxAR6LTcCBwU3yuMsZSNTxHYRZt0WSBzKvxXkq
3Z/Wodn+bIbJ7Eh/A3PI49BBThtVbDvmmmExxG4YnMnUP2QnXI7/X/I4neSPjCtOGTqDDhaUy9nl
CYhiem6wThlw5qtUfB+YFNCDj+gi+SgGU2RFPJ4kXFu+ebMu3r6Z3HHw36BuFJ500ZsXYcwLqkNR
F4h3yUIDF2PS4KBAv3JhPrId0l20ifK64kCTH9bJmDIcoqbHUv/Uo1YjNh9Y81WwNnvNi0EAxR1r
08fWnfrZq8zo09qVi0oM3+Qm3AE8UdR2XNGS7r5CYeAXr83ZaIP1JEKx1vCcKn3F9iZdqJqO66Yh
xaU/v/pzqjouefr3RLTgHGaiL5+dhBytmAEg/3BC2W/001dSo5nN4TRj68vzOi8xnG2dJL97g57W
by8cdZ2yGIPDUnZvopxqMqq5UcSZlX+R98mgJL+VRZSJ6iDf/4UP4HrdabPTBxlB7I7O1+CLrTAJ
laEdc60QYGygDRDxrdAPYLxpm3JNLD6NYTeFQdWimVShrem2w79y6HmoK19gbV6sbsBGzQE8XZxO
XMyohQR3A3FBu3MtMEQJU3hoAxYYv0BwmQwWIDC3vyiSfdLL9CrvuIwJUc+Cu1HPQHUL1kI6ysfY
WuUwM59mpOjjqF1KVZsbvwxgu3F1rpNKguX3s99W21lsdMq9Q+uqFrSC1ywi7e5jrL9F6gbcI084
YrbOmaTyTwemjRleYHcul40mj5XtFEBr8iPtXjGlKOsAQHuL6B8l4PpPPi0VKvHctyBN2+KmRnBj
KrdigbIuWUzXCR5ML0GHw/lpY1t1MFq62P+CNT09tFmv2Ll0KjHuEtStY/e/cQoYJGIWBHiSEj/I
Om7XRrhm5BFPWz3sFfgHZZqjTFNNlisivhDR+ZX1VhahxJ0mRNFFQZxODCIEbesQX4wBnXvf2csY
vIEH3Zk3eT9ybHTaF6KtYtONsJR0Rj4928gA7ycj/mqtYUPomRP7SyhSoxTYt909YaIgnIuYE3GO
RJUi/2ZdDmaal1xs60oiloGuy5wxpMKOwVvVckTYIHqucaV61Yfr3N3Isq+pgec+sOUAXw7GgV++
3i6rH4XlQVnbOniWcS9IRhH1031GAUE1cKt0icI+tAQcYZjUvtfvJ8onjAd48R8TDroYcBPJUadQ
Jitwq812coRPAIskezYC2LGbvNo6lVSL7Shm2XtLWHmPN4KBL9hdXV8vvXMWDy8rbJxXOEoibiZ/
GFZoZ+EMsIljmWoee+Ad+CovozGoS2qhJzzaEjqMGa1T6hOZzhQbLyiFmxCdem52M/bHyWf+mra0
RgVW2hOLNs/9Sedh358cc2Veur5xBAY4pxiInr+uOAOCwelUcj06K/7+fMKYB/HKc4b1def8k+56
eJgNdGG6HioD9Q5dvCRc0ZhweJLLSYRxDRMSKB50vhb04D6HIl11RkA9O2ScC/rHoedxLZPTvZnD
H1wmH30VMuUCpmLU32dNPCWuPyiugreXrVTZa5+RpNJeJ8c6l+wRH8vRFZjjHTqy/GDqJm9iWrQD
RiFR/CkzQ7z0Y9JXOGLl8sDpQhnzHFEj0998R6a6OolODCaG6CS8QJcrNpRD1uIKi/ueFgUYdxDZ
kcpvQhpOpDDEyys6vb6y1KbN+tBBWXFpjc2TrPSHkJC1eCpyvbffPoUJvNzxJ/V1xaFI7xwGQcrP
HGbBOsVfzERshN6tbz/efAinhjrJWkQYMzM6h6D1KQzLXnXf/0G54ZmQgin693b0ukWFQX9dliIF
8hvONoqYtBX3LSWqBUI6RW3QaTTYexGBbzZaUbgAh+zEOWdltvrBC4yHVF+vdxsS2M5JT41ygzlb
MUAacXrFkQWe3VJOUIMd8AbWFri6648MblWYJUznkG2jJZDnABL9OT8c4iX9k4dnItQDwGZjxI+L
pYKMwN/IsyYqVasbJTTZqG8qKhKoehPT93eQueHGRaN5mzhDI0fzRBK/BD2QbCR+tB7964sCi7kK
Q0FHUcKJ9IVScOtPgCDTMDQCpBfD8IMT3Uls2q15r7bpVj/EjZVdw2AKF5Dv4ChVpqrC/Kw1ZYsd
Qg8sFVLYcU3w7aBAc73XuAUiGtsyNBhjjiOaYIpqOpxPeedTjvaxOZdjwscx1rlLZdODUcPcqtOA
NeLCBi8YbaRnbFsEcyuMhWYsC3Cc6M5EM+MK3gFoxBrAUb9O4pwZrVpbG7kTGkmA9t+GhRlC+Vh4
Z3ciDdgcLRmnOwy1/TuXjVAS52UhfhlSzMhhvH9bmca0ehfJMlzIsNoGZdGo7s/ePXWBHAAwA7WQ
jBnYymADGhEoYNKJllHDqrXuezK+97FH7Q2xOMTAXS/EWgD71r4hUHCENsXGcEuJ0jz2XX7x1pMx
vYJH3mblYZgaZUG/useva675RYm8Ju2jvF1mY4xoFRe2k9a0rY8ILNnmp/dsKuJxTy2wBMuRRqBC
V2oInifcRzB7MGDVlMSvbYzvMJZHgpe8EcQIwAUZJNFNonkFfyNqHeNDKG/4P9XzxVcHDZ6Aj0pF
FXRTamwTb4kFcJ5RCGrjM7ma6sqrXXsS5MMDV5+j+a5aeGgC3LTgFTf0pPfd5ru+2LO1G2YQMBDn
aJpm83MOqbA8/mqiZBu1qwdYavu1TyclbCNMVd2p9Xy2r6V2vaez5cyECn0qAfH4Nu7pbHf1x9yA
lB5QwYM3tQipFb2OVeZ/UAM2gMkgT8+JK4Xhe6qdND+i8ODW6oLikaXukBWLvePKjQbaQq8pmD7q
HczujdLUOsILeiu+4cc5dIZDldLrCF2Xv9R/0VHC5x+sfzmZbIOlQdu8Qe+Tugev8QhNA5efr4SR
J0MtSQTKOhR0KOPY4G++XHn3FPKUEJo5qkNEFWvPVi+lR5bEYypRahWWCu/w3Z4kdYdLMdfBWsX+
SqHrm4wCbrlbDWkSqB1zrXbYjpi3FUkouCablHuJnyWfELoL/IutItgvaV+6i7z+sJ0QVhMDcEdE
Q3UGX0qe6MnnAyLFEy9S2qCF7OTdmW3CZTIzPmt30VdGsYIPKuJvHvBqMFK8gBaaTbkJl+G1O160
JvpKva5shk/EKFILyOVGfLIktPCkIpL8bgyYTul7aJKW7sQ02V17SrxuBeJZvx5WVIjmeiB+vZEd
Wn2BRWorKpmBSs+uks5/+2d6IevDPJ+qcjuYi3lzp4LwIbTLQhgQkcOdvdUatt+P9Pfjf64ZTWpl
BDjC/RgxcGCRO1SCxOqhNfTVa8LQRAvS1QMknUn9eoDLBiBxc4ehhlzeFHgd0mUDrbDj7JE3CUl6
7XYzfsx0RxDQICk1HcKsMLcDTGDZNxAjgMVRsdFgozHf57hkY7VOJ9tImdFqHz1KThjCaeE5ASh0
qwIaGrYU0U2c9da8hxl8I+J4e7qVAL9Tvp1CJyaSO7XTtxgJ/Bq1uA/5kiVBklcVcABD+QNn3CbQ
zOD+Pk/DqLtfg2mpxMC2ZM/1chedcWhbRrIfRvPR5HjqNPR0mBV2m5FEdPMsjhuXfmB4wboYxbXD
uXDuT82FHGBTR1rw27SXdMLtNvrkYBRJ8esvsNDIr5gee9lnoXlsB9LwertQxy1P1FOFXD4tNyUn
MNLIuOpntq+6tjowtI6oHYrZD03VEDzaRbU+hpm8fxu7T9rphkqdggN+Ag4d2XVvKkjR+OS++Xd9
xBYpqHM3crKcRXsH6VyMcHoNB3F6aCXuIO1EKjaT7OcWknF4wyTlA8LReXYJQ/CiQzGL7mimIXlU
LaR+9dBYJs/tVFbRLhxdEsHNsOPa3LZC0UZDMS5PH7MgTkgttoaHmfG7IT4x+lpuFr6OlG34IASX
bM2QetxI0g/YLiV0Vu6FWQA5VHScCiB35lGNpPSG2hcIA/dZUwDzkPJ4WH+a73PlDwt2XME2LHCH
x23z59dnkrLnUPO9XlypUa0q6or9G3IkY2Ya7cRSEXlbPHxSeakwjDygyQGIVpg178tmWHZcQKVv
hGfoUSTuk/pCFrUr7rgHqdGV4UJXgq0HiRsv5VmRAh8G2/EJlRQ67TaGq+4I+3xBNq/ZUj3ojWKO
yhNbSAmx5Szu1xip28X/nj4C1POj0vEOc6OnjuCmv1FbZkhqHtvv+5iis3yGmQnTcEZJR8mIHY6A
NVPzTMpv3h719VjB/gd67gsAZoO42V1ivMr4zVtE+cYjvCJM0TKlPlw4siNuGCPzDXUx2/tQlyRg
jO6Rt0VK1umbi10T0aBxVi0OBySb6g/xR6jX2cSZXSFNu0AvZl98wSmgz6tzdK+pH6qidTydCe7g
RGVXNuAf3cuN8Nb5NUc53s4NqY6ywyWJqHQgo8jPj8xIyVY9bUkIHx6c9KEDG0Z8VKtjUD2AjxRI
Wxl411zcqat3rvU7wdSlwpjYu46h6pvp+KCLl/DbAeGQqeg3JGYnxF0aWPXto81OAdAhnpfoRnJM
68a1nuCuueLupTiOJ1a/LSnDW06NXGAwczIKAtyUUs6XeKkXjXF+bMMbAL0ppfOgm10PP3Yr7Myd
m2cX4ns3BB5WxLU3/V4Ky/Town/A0Md2dCH9n4KWvMTtRBojA4y0MsEiT/4O5hKrMhLT+x5PaOtp
ro1Rft7Rw2li9LUDwaFp9maqzOnvYsSk8yF9/wqCVPozylXEJLcDk53tCeu++qEn9SKD+MBK25Wt
lqdjEg3I1PrjGayePO0AGrUC6+PPogFyd6StuSRNmPbzZYnkImbAZuAiQWMFQ1OX3nu8WWqbtZ+3
TB7vyttws9pmm8HQX4doOmjw2JYgHDdUwTRp/vsajc+fEJsCei2YO1/NcwbKFjKeD1sCtHK3lSTI
LckP9UFdZn0n0YFA0U0QjE5dZKWFZwAMnAlskmxEywGjNaSDIdlBasNLUNgDGu2ElidukxEJTB/k
M5Klw4GSyoaauP/XR33xldfbB2y3zI9ew7p75P4QbABEPoHlNOjqsLzE/wGThnnmF/YaukHONMFf
oCYc0QQd5SjXhuTo+BRX1yFdI7+N/6W1pLHz1iFIgyRCggjA9sr0P75ggNGO6BKnC5ZW+wxtF7sz
XExSzRKWku6z/dpCUFu9anVaCwygVkxTTszD3aGeQYhXSewWsb/PPqQbb5Nxwp2rd7nyOO8Q3vdq
kmgRA4ibMwQzLro4H4xoLYd/vgAEE50voty0rm2zplO5s8yihzgEtvqbxnG+MQn/Tfy4jtBL83WG
TfQSBlgdTo1t071yUCo7CqTxBKPnjrVqW9QNvtuv87A8ZwerffI95QiSpSOK+fsSNR7l9eIOnVZ3
u308Hy4ve2f+R/k+DZ8hiPB4AmQrVaRJD1hoO2p7ugrFzm3AFUEN/j7rpJFLQ6NSidZKxTp8+Qrq
hs5Fj/QqsKYPHjLgLdNaHrgM4BYlvNhNhE+ZXek8pD0b9l7A2L5EROgYf4miFMGImBBaamNjd2cO
Q9+zzN5gyJYtFBQ+Q37q+jb9sDvzfd0I1myIWFrpfG08QkAfhs57cl14H/8ljXnJcqi87+sY+oZ+
LXpbyzFlz8dZx/qAt2NDicqpd27Bw6wj4tec4M/eWJJ9qB5l0FfNJuxaaOA/fht+sHac2GhciRNq
xQNKqVaNc5dMSllDBgdGaO+0GkLZq1hE2W6j/qcjPwLV/zB+LNIr7UCAicA1klSka7c0R+9ODk01
R8iDjDELT8c32BNXiqUJysWBQ+9q4KuL6wqw500/Rgw6GwQdZRMiSGaRmua9CHCF1iFT/i1uHvz1
K4tRHgQbjhBit1rpGzNSWVNt8jfc9olPn+G14sDJeLbHgENZy8/0ci5qbhAWZY832DfKUXZrwmrw
zoNx8X244VEasPeNkxjwLU094D8Upn3DqWVu9LvnhLTjq9bQCi/2ZkSOqkqS1+jtZQLGJaAT9yYw
NXQhcpm/5QTiV+iL+FWUhl2LM7tB/S/TNf+rsOX+rfrA9LJeRkZxTmMsXA8jMyPOz32TuQwsAXAy
8fqaoN9z/M6V63d87DIXAnWtwgzhiePpMUQ4s9JNfuP9gUPnGAkPQ11gJoQvMGwKLwOGmKHKXbWs
XkV6rrbsQOhs8XuH4JRCOVTy/zH9AcBfSD+Qe2vcPCK3mvC813vw2UXTI3Y2audGpqGLPoh+gw0A
mazvRr4xWWcDvpvXGGCEQYoATP5btdSn0DTnC1IdmSHUVl4fSpWw8ZB3wxf70lMCGAW52Bif44Jn
hPHUYssmbC/bNX0pzcyjUpEmHXXDOtk/AlApg9PQ6DQwAl5+RkWb8N2Wj8XT6wJvBoY0C2M9QnBW
AQkJczoJdTKCbIpkSUGt1RUWgpLTBj3gkRTVEW/IthnqOILnlf5mwOY0GqgMKVDz6/Gyj50fBY1w
s/A+MiBIYMVP2tymtsuUVysD5gJ3xARuLweuyWSWjDOc+JciDZKfo40j9DN6JSWpZzpkwDvjc5GD
cGGc8jvhedRL18CTv4+TZzaJoSj/HUB26y6/qzZueKXj9WavDqSAXhQifKObff6k2JbBgr1j4H8F
S+8X+yNs4WdDFNhZCYHnl4TYFx6PG7f2+cFWlfhJ3w8e60PxqPLkkUM+SlEgeXM+uZ1ftCzJSVDE
SautDROgUcs32b7GfF7TSdz2kCVSZvDklGt6RTiXY+ysxbBBYzf2AEIC/l5Qf40qnWh7EVXOKMxY
TsC7taVDvyYTDUqR+WW62tgcS3AOV3jPlbXMB6BdlO40sRUrM9xf1fuyckbcWD4UoWAL9iikvoZ5
aREu3/+4fMngZbvhnmDJydlLRZmSpRmY47yQV2IWvdmsgI+QPB1Sa6WOtQyLHt85dfoK3VICGoQv
4DgGtNhVrdtW6TfAqghFQ14tGPgx4kZzO52aFqdQrONz1Jwf5ACNG66ToG8h0gZ4Q+3bZ1sVVGQP
gpg0AMQkx64HUUnY4u6/ivj5bW3iYM3Q/UWhwGpxIL1HZI4JFzi4T6pMy5QG03aS9Z8HzEMAREsP
VkY0sQ7JGKSi9cYCqlQPuTwspv0nal7bsmxt/kWoOrQ4hOAWKPu8m5CNeVG2V+seNc1rkkdrdpJl
uFmhDXgiyWvF45OHvYnv5XF/jnu2h+60HPrS0jmIyCVAhBOwIOx38J2wYqUn9Pc7lSkpWTuanHOD
4WvyetSGyLpPeFUK7sdczEX8O2nMLeKJ82ZVyz9duxZD5u4N94w7sTvXGJFZc4V8UuiNzLxRLqck
RRGf+qLIguF1x8ta0g6OuMhy7iYrMsascC0NwZso8iHwXs8VUWuoLkDkOumS/gKMoXXE5XCavHXG
D09IKWin1/4JIFiHcY5o0fuetZId8nA83Bsb8ZlzgyS8+xpblFJyA6vEGWbdDUYd9mEWM6nCXUaM
K8t8EAnx1WZ4v3n3EWvPwEwd6zAJ7mAK5EVQQLXzAaduj7sUTpN7HblACEQdsnG2JhsK0scp3nfS
DyS92IJ/LqD5rSCWN09tTV4w6ZvBXaRryGfFjMxxbuBD5H9HdZAtP71lDM71zit1LRLM41RgqILY
avAEMwSCGZk86sYKckyRYNUSzSMEdt6FNEDMYThumHWs9Jc45Rj+o6j+vDNO8kIMb/3aoeK9/JJN
HzBT1eFPterD+Kvq18xu//u8HW9kn9Hj2E8FnomH/CvSt7K+baJCaW/lNBAV75XP6eYPCqnTQ1kK
SYjy1fQgJLubkIcsaWDsxMqRtzzYlcVsNQ4f4mgzFfGvyB1xNPQ+D/CQNN3L+H5LLRMht2RCLov2
JB/Cg3Km6Jg+O/4/Rs3TvFSTJYaf+6bNBVEmpihsS9W0Gr9EihCbpm9QgXtbwnnpDMsiI84hRPRZ
6eoEJqySWaWKobSsHF9fCnhcmjoUTt10dsvkdkE8RzbXQkk46M9u2PbHWY+dMffZyub/8l450QIY
AcOWcoZ4liNZIcP0Ph9dVflC/zVgAP20j3VJEQuNyfnJKpcMt+xDUDFqP7/9tUWMkhwCdC8iNg12
xFWW9pWbIEhVJ/+Kg8k+FV6p178M/ziwu39o9e1snLga3ljnlVr1yoIDNXgYkEJYZDc8RpU9xtLN
be+s535T20658vvkXb0uTrbo2roSC0Zien93MpVTwYigD7rvz+NG1s9ngeFr/Zc8eFtsZS5rEu7P
9/ETucYKlXsT7xA2B+ruaJpu2fetDx5N9EQI0ySG8YuTPDLztOa4eImRZpNDiKKDrGM/xF5x64T8
ck1Uq0SO1mWRhcIb418yxGRggpaDjZI8uedUOOXscq7gm3DOYBiXGkH3KhKUsaqWKO6y8cq1BUb8
Vymz4iBdu6+ZUmZ2l6etl3KZg/LZvUDr5kukpWO+0NxFPTWwN+bTWeZtGwScy9scxFyS4yPPCTMr
dRYEKQ3boh7LQi2PTZBJ71fKTJDx3b9X4Fp7J4L0kgJvdYwHWsAcXqBT61qZi8kLbaX20fZzdTow
JTjMFAhnpdlwT96QzxYM2Nos33yeHD5JvghTBuAmfFoHGZoPgQZ7/6sz4irFsXOl0bTnCBryJuJ4
13q3NSL3A3wtIKlsg78JdPgibPxS+zC/Mt2AgB7KG3n6hXwY6d88WZ2zdX5MtSphZzXzEUXZjgr5
ceildNNRv5EHwq4nQ1yyScKsfglRm5fl1fh1LpSu0+KvdtBLtzLsOdLPAZwMMvL06cq277Jq1kb/
IGyyK4eDET1/t/ON+wGHKcDH6S9v5KphiYMSbp3e7jJQc8dpxyiYE6mb3vTtL0VKOeHIpPPXrylY
GYu3afr6j+b9TBMsDdz1H+1YrYXJkHJg7tLj4Gm4+sO5eVhfnDHnvxEBL9DZozFMvO9VJ8zwGz3e
rWkOezQ+/JV+AydZrKj38B6KnYVdPFHbO5y8emlIHUFu2cl0l98XqQhMdyRhR9+bC0s1qQVmT3iq
a+XILOV2LYTrKxmT5Bh2941fgubkP34hOAKOeg/rOlE9YbmIXH13V4SsBb4RsvTuXnWSLS3HwORl
+f1M1wOI1dvG540rzFChTJDe21ayTVHlQ7tnOZ636d0EAOn3ytXq1xvlYbX81IcF2F3yddB74J6G
nmRl/GJkGwQyD2RccLe4ZGVNOGMy3EhAI0iRAziPoM/sQji8ATeBCmalc7YelBVdizeSn+2Aa3mU
tcekam6PrOdlc34xqQG+J3Ygs5SE9fAgTmknX72eD625o7w3EB0LJ/XeJp87418GjRfEevvbvWF9
YIq5eHOKguFqkUTFTPxvtw9V8KQp9hPdiBgWcpz0VD9xjTI0eawOQMfigqt0oJI5eDHrrhvpNH/U
D2HWAzSjIQMVdx2rYl3DM7Rm3WgkfXggyac5o/ckQeQyfKI89Eyi1WaIZoNvWMDJ/gZOuopOjxpI
TxESNbOZTCUtfZNxczaOFzUe+tBi3VJjItIjlwcXLhxMIOJhmflr/WY/Ke9djBl2HDCPosq0LyzD
207qllXKxGc24yD9aLnqSNQdaZ+vDinVo3byE6uGaIPsphSMy3E6vKeoDMXXC3FCamUDVThbKuHc
NSEDU9aHQdt7ae/SYkGIB9K46dPS4We8nMxpsWzf27+Wc0FB41X5H4f15wtuNejLb9oGVLOLQgvM
iOrs58/cZjPDGmnyUfL26qA7xwkGeLhBJbz/ubITFtQ5cn6aCDh6MeIxZ5XfwBSR6KAqszZJ+MRr
oXO1knIFvTFN580Q4uorjdifzRIBp0NAAYxhxBAC5ziscIG0crLjZ+T2B1OTUubUSnc+LRNzRPgS
1a2uKQAhHPn5cIxshP+0CmEyq2WcBaM7JUw46rAWCfdY8359hI1yxRYCcci1WuotH99EfqFPeBoy
xbp/PUwR3EMMYFC1PNpbcR/TsaeAaCktrDoZfoEhj/PoARe9lIuINdQeQCyli+/T1H9OiCX+UxT2
CzuWLziK2vhnaE1cTWr8WdDlGR2bP0WnS4WHRR6boYLxCJvITKFrytRjVuAsFm8CJHXRiMFJ1/wO
DYu+IGxFqQHfl0aegNR3MYNqEyEjmrNqkO6tuwpAT8g3m+h/r0LOwLagmv+//bZPMiXS1Wpb4R5j
pyWn+Jogm1XJZU/8oDUdOy/Chy+7Gv/IpTAWrPudSJEky2bwPRam4ZTNVkIcfA4WTTXrGiO4jvZB
emzPBztZ+EZ8iePcr/Zo6Gaj3PzpcChEiNZWCk1Wtj65aN/294AWVqkfcQYNSpWSkPgMeC+o5U8Y
WllyNKtHUeR9JiOEc91l7GmZ2sL+yL2ZUeT6tK16jjqZWi6GEMizcg5CWKNJzVjdI5dti4Iijevu
aJigX+eeLZFrOBARsCX28FQLON3Hf8YrQrBa05RRuHH2/j99wfFt0JDFbUrfFude04oUqn1fpsIx
gsF7pRhbyVPqC920lRL7H5q0/jK1tmAXsmx61fgOCCN3ttUDbfja/lG1AzXFFc1Ww1U7qtL1DEIG
z9l90THrlq+v1PVa5WzHqSs2mw/UhNrLJwMkSrfwB+RyxISPLHfPXVFZKGk1YGL65N5fpacTUli/
z4NWQK78H609jbjUJcQAjnYu2jOdu9NWYcLH5D0w5u1M16CDDSAbs7YIvC/Ex7KqC+wptXS/grip
ZVPze3D03k3SADcBoO7BUwMSV0oTKw8OTgNY/QP5V23gEsn31/CmZTlOhv4wNFJ/yJENzYpNNAe5
9q3ssLr6tHlLV0RgGhko4jhVzlBVFNGG3f+QQxys8bC7xuCcBLKQOxm3PHvruHc2xiX9hrREC7Nj
0HkXtg791vnZETYCFKafw9+1AXpM1htooo1D2RsFiWWgheU33AMUIrK/0tBjvG5hvGuKVRg7YHIn
vMUjEywreJoG5KD7kfGqQyVpjrH9xhxkXwxr95dhKpXgPxeWnKeBb1dFzYW9D26D4d5+fjqZfpSe
Zbfqx0D4bHIM2tY31VmJWcmVkhNGKBdEBzVEaGCn2QhPmUQNzj1Pd1WzelWhdn2clmkYVfyEeEsF
Lj6OBx51cacYDgZHuDyA9ablAspnm06/IoBbM9b4qMknZWpOCYk0EEQOhdr/r4AKWxI/+qujjiOX
mwXYRt+jMtOqGhQE//Gmb2ZxTc09pN4C0ZA3DzGcRPpaEm8Z+B3vH7O/19eOV1iFraWXN/ifFygP
kglkABWhMKhzqFKzYF4t6WxY1FAnkqwljzLfnMgm/UgqE4t10l1jrO4tdcR9HDT8Aj7tOGD1dFbw
GWbCT115/xZ5+6kiZ7relV5jRl41KuGVlwmWbf5pWVlX2Yq/if09Zove4GHLkioPRiGn39OujK6s
wtZYGONYPnm2K2eFNzmBSIYRRT2eymU1Po3zJ7n6InK1M6q5g6NLhee3ilCMx7hie10IU6/QXCIA
FLZDGN/cARESYIV59mFVYarwS8JcWIpknw6Ufh41qp7V67MSOv7IfZjh2Qo89CEU1yG6cYMqQd84
+JES6N/Oep76hU5VWKgVDVPTgck+ea0hCy8z6VTTiAxnZvGMQDH/SW5fMVajVC9X63SNv8GnRvC8
tooDHeXzyMzg+HiUBOKUm2tDNligWeyjWlQ4HuehuawAA9Nr/NXFsU2TB50F96eVpgp7r2ipTXs2
Mlu4EeVj7pJARz1oVfilQzhmk8p3SbNbFaXfsZniazuCpZKXnPgVhAGFkmFgBc/AVwgcfLPn4PI8
5uvXFDL8hnMeO5sG6Usp5940CyavKwujpfhOCfWqccnNmYso2Y3EJJMRXsUFG7IcGLzomTufDFRI
KqXZf9Wita17kGID9kaEgtyuQiiJuw/wqwFgZnc5AQH+UFJnI1jzNjzY93zuJwjpWFdDxFsnk0Sh
icmVlUE3jwuVw+7sn73qGaUBS4z1RASfC5l7Gc1FcBMXvE1i8uvudRaDlcak0KCe7krFqB5BQqKj
+9p1q0xV/BTB4rxBVqVDrcFzi8YcHAOGNOsujgAL6UvBXdpraMrP7C8LqZw56oDAcOM5HyxKP4uI
+QQIhPt5kGNH9Y55Q+rTgCtcIMTNRM9nrpphFVIwhOeH7O7Te/Q5DtdOByDDoE4C2apqELGuIF7l
2k11LG/kEO2DkQx0uY6QSFp45fMkHtz73DNbF0kIcsvYzVEy7gTqPdPw6IDnvnffjsdME7KkaZSj
d011C+PJd4XEyrDQICJf+mTYBmzMu3+GXSHYFc9WF/J5l0JlpXZqHLwXf/A0UK1c9tLf5I1jymq8
NaRwNFWfWSyjDqHcNeK/+hZYzcrCZNsk/+NyfUCSKonKEcw5ksXqrsgZSL4ydwgbIxWO4VKsTtRp
eDv5M4j9P8K2adncqNXieVGkpDXo36hd0+Afv8PybHOvaBL2vcfrxwpwOrvQdJBEp7Jh0LNSNhct
XUYKen9evrAjk+4wcYjkZFqcw6DZu07j5OCOp109rTXnGlPQBzkXXefeS34szsDQvXqUPUUy8ua6
Esox/IJgtkQEt6dnlmyBSOm+3f5CTaiJziTBqsBfLDOYx4sf113XbvJ6RhRyZI/ztschKEbiAwxi
Jv9xEUF+896WgFTISGco349B/dxGsNekLstDjcMDzTmpzUfno+312nWrcK+Hk+RFM9wsLcoKbdf/
q7yk5vM8xd9lo0jmomwRn4NVSF9nq6xU+AsI/oelY6cx0ilrWcr86uxaWg/AI3RfOAhyON/1VMEd
+zmo3gkvEtWjnYTys6/ysChFN7K/latZO+joosyULBmq5wRuYLgnmPUhFfGiIw5k1yo6nhUML8OA
2UEoXKgsIFxuUjUlSvlmAAZONMuN1bZn2j3wqU62BHV5YMhSOO346HDmnpavskmnkrA9gy7MgLI3
QnNA13rSLph/NdUCpIMCm74MX0vO/1AxDebzNiyB4VFzHJWto8CwydMum78978qKrvaIvlqB4Irc
8FjBLt5XXb259ktUFkXxmQi/ExAhOBYDcoRHKEo/ZOokSimoGQBBq4wis2SAguMHbDmjLyiK/5an
AwGzTdzKAgv9BV2plswPyMZGtMk1J1BV7umxI9TygXadgYcbS3um4S4B7adzB2ab2GE99pFb1n8v
IsubTrdtX4sISvo2OiEI1bPzJq9b9AuaZIFSTR05f8vgQZgOCPDk/ns8ocIyrj/AI/N5klVV6EwK
UNNrM63lQSSopPX+jFN8PjaaM7p6jDxJmI/bpG+nggmhOrOmRyqF3kt/6DkhZhbjmJyZxl64Emvc
e5GaYWvGwrMwKZcwmmynLVjJT8bZjDgDyzx8tSIU5ng6/cRr31k/zomeEQobRjQvgah5EOd98dtn
ILm/z94TaHFcmWvNZz2PxV0FA0i+DOh6GELy/oqE5SEznNJErSPcZqVlchQ83VJod9wiiBwKtPQO
lGOKuEY/Sdmuyq8kyBUq28qzFKhtkA4l0cO5c9YaPAJgLgvwR1qJbT5CodXRu+fhnOoGvmtbE3Q1
RF9m/6mWP5LqzJvdn8SOr+rDn/ZBuGufDPrcfKIas2UW4BgZFb/VJocjtpnXvf1ZoGMljYtFFl6T
vuFvt0GU3BO3OVobgXFpZ+ylWdkxuA0hDslrcEz+IiRBWGi3MoeUTUF89J1Wo2tpRAHuARKYeMoL
Mtn9D1+UySmKtwqcOTRRv2ONQGqSO82Aigmv2/wiXz+Y+/RtgHxGOllAllYd2JW+CYWuRYs+JsfP
66Jmn1a0GRLTYlx3ienhFdb3PjgSilK/OLCRdrZ/V+UwvQxrY0v1dL5xgDSuJVBUxHygLcVyMLKD
z0CJShZ808O7j3amkKdocLnSgJBCxhMuWvKZNg4ZZhivIFttCfD6Ce/sU38/OeZ+sHsz0J8Lzlno
duz4sZgW8V0QSN8/soVta165Zlft9VidHl7uYU0qVvOyL+5DLrNTZTAmC9ajsJPlandSX2g1tsDZ
EnCmFw3vS6RHYfRB2/FAeMOQSZe0U7YuQeZYpc6HCyWAQLfYhFOkKyXZkHrtp0ZsHVdKYZjzwSNe
jgjmpOUlfZ6LL7i4t4hWm9P/adns4HzVSyDEQOyuWhVJ+HIqEn622O1DmfEg5Fm5BgaL7Xo82vYd
fircvn8W3CYwFdaoYGkLGSvqp5rZ9LXur3SdhvsftDIhXNNs9gU3wEnLYDbB8vbtCkgEgfrgTdYL
Dghan6VD3XEyNV7jSELRGyIjPT7tk+cdtKbNnxwZ/SVpvLipr/ne79j4WToV3cMfDPDWjaI0yENs
f4nhEkTcmbn+YeywqEMzqO4EKizHEgkDCaHYZOr0YrdC6kfrVGZlA790GW6prsQtzlbYobcTvFHc
/DogUxUPeleJH7HsW7LANPYV9+JWE142Fz+BD/bC+o8TM2Fiwu7QP2RxVCv2vJj1FyxX2JZilzHc
QCFLIfeRJHXbNQr52UGKM99Q3xg1PqaM6bh0tZWcbNfCXU9DNV/g0l9x7Yy/Ak37mfiw2e1fNugz
nObDroxPefqZmeXm5WW5GIyaegH5fgU9/Cz3e7IG6CFsPupPqgGqvJiJ4pvHSNY0kAr1XuLxvP8n
br0pzmq4sybrwUbJ4bZYKx5QGDxEo4D+U7lLlLUrr97T6d5UxKzHIC9yRUOCVZtp0OtllQEB8YC1
8QaaGYhNCZ/HR+iu63hOOu7/0Zu+b1OtUj890C0um3KexvOzah19CbRFURnvD5LZzdd2SQHZXr2/
hasoWC5xnsXlBZiDW+7IHiOymN5rjUq3m394qlbJg9o04WzZiOLhCNA02AsyCprfH+6SNszWlLki
UTFPvUd7X998sDCrZ5njWqYIeLeIlo60kRZ8azmAWCvC1U4gwy6Ril/a+4JjEn0g7c8OeOlgencv
YBDSMYUC1BOJ5aQRFsSPhbv7hcN3m4XbQu3urjpauQFZj05LDA0sWbKJj+X4Cl722DXyv4xl0I/T
kmwFmdInFPOQ2FcvHetMxX+VK2zj6luNuqI6bpUImUGsDwnQe9jHnYTo45sLyQpm4dqviBiSxdHH
udHgAjTjKwUlZX280qXFmacliVz/Z//xHMJxgodRlgmdrUb26Z/9zt/5Ck8rYe+8eoCeHYcieJTu
dynZmMz4i40KVEnY2G7iQ/vd0Voo2RR0S9g0QTmwot1G9qXVScMCpMNcjKBKwCKAqhgJtOQ/lDaA
KdKnkzhXnSxwqkgt1nq8UJS5w/s4uHAFjd/Y9SrlYTCZqGqoEqdbHauReF1DTaAI6trxD9kP2M51
6RozMXjx7YZFF84RrXgNvRroMJO6qGAgQGy7iADQz766syV6eJug6ptb5QzIb6VmXteEtmth7GPL
jOqF01ewX/49jh5LpljwOL+xsDAlcbUJnTOlN5TiBo4+3PAMRLjDDHl9tFRqrV5+yEL0gNnqEdIZ
rTfX/sNFyp6IorIsAntNW+wF79HoW4uJSOUQgmE0O5ThOyTAW94Y4bUKoEyyyNHt4MMIwDkv18Yz
wr5+2pTczeIFMf93cPvaDpvEuBuh2lVzzqHKPbOjB6ax8ZN9aEvxumnOiClj1SUeaztEUje02B2g
gJPt3EB20w4ZjulUvZj/G8S3mXSk1MroO60gxAH7cxjUb7usMktnoMPftyzzOJrMOhoJZ/vA/i2T
xekB353mhkVRC3Ti6x9Z8g8AdRTYDTIUEyixx2ezQdfE5Rs1RgcorbE8V5P4y1KH8xBXRs/ipH+d
xZ8lRNavsBYJg3iYWtl3+R9c78CqjjG7qVuwAU7r9U/PgfHGI+FEX9hI4MdWduJlPK1POciThwFD
4JY5ukUFzfvoHzgH7/dFCbSieJJnVre4mcAmhkzrJBIdwF4f4lw5F2Wxt2mVqJsUFSn/WYv89QFf
QVFLnAcdmhv4mDTndjRypZJS0ikC14+iogeYnOpr+7zn5k5vVJzRkro5BVHSAhjmDw8beIkGthNn
CtdEkVmYgXv+jH0nrwEcXCcL7q+wHnRQO/VC5H7QdX7yJf/d9Zyxb0+tdtymKxjbZMEtKcjxioXT
dOI0ki35D/Tkcbs26d51VAWp0ERgbd1vBGZJ2GsWfd/PYlJnTfaJKgT+8ohtMQr3/GgSwtYBr1vC
D1+GT7LzkpeVTZGtF1uLvUx/Ne4iGVf2KfEf/Jlq08YiPEClR9At48ca7KpilD4257fueNz7ZmZ9
FmmS2OqrFo+uRc9IM+jmmhWdiQ7E7HiFwxz4JU4Dj2/PY+1lDFMrYAUTgZfy9iDYG/XNKB5rwKoM
+xrlVXSopHQxPhLEwAeEjVS6hQYaEOOrSemaSYPNSic4ObqRph/mthUmKcWndkO8ChoypLAN/Vjp
jFaCd1yCxNtWWXl4YYBKwys18D4/MfdeITNDYln66vFFAu66qaP7XD4dGYM8zJZbuW9taUN/V3o7
5ZL65sQIC7JWa3nMmZkt93cnEE7oPz+6uuqB/el8fopy9vPB7HZyJzvIDRw3mUC0kjKDpiJ5B/XF
zdpIymlRWgVj8DWs84RO7M2V/6pfQbs3DcQpciny1Ti1Q1X2Lvrz9mXIapRAryTHHlB4gMfuRcl5
v9QT4AbgXV2POJ3xT38eCkKnmBw6Lt//KhcrnXPOPkumC7f16A36Dut63hLljVad+lUPALQBwymE
xU3Bo9fMgegB37ZtHDfxC1d8hSlLJdQ6X2d+LAkcL4Ik8widqGMA7uEbRRI0IVBSGgxverQGjPNH
taksTJ4431Tv1WQ+x8IKfT6AgZDjSfjFuxenJSMWOC0bMyzHgZRojsnL+aJP/GPtiJXArt0JWQy6
WF2gKVMq8Wp7rs2KzOfRlQfMLlOuG2TmofBIrY2cZwOEedxsNDKKiAc1ZCZHEQAMA7Yyi14kfmyM
PNUlBlI1AFEZJZXDeoK8Y0aJR9o5FEZsLvXav9rLZ03aYTxVxsVRV+oUgPq+dYT2Q1ZqqnfBdNZ4
boXTHXigMghgxsnRBZLTu9oMLyYTQMyr/qfy/ZMxtF8EY9zfEsqgETYE3DcvcA/t2iF8cWRHtERQ
UvjUtiC4zEbSZeR2Mb/APNow85ZzfVlgHw00dC0Cmh8I1zyZvKR/nxIb4D9MKT8ZICg1qa8XJ5ab
7ITpVenGSuLYj61Igw3JagXDa7SuSY9uumGnf3C6DWnJG+zwF7KyxKNQl+qqIjuxoaBV+BzvTalT
lKcUFBw1zTEbuzCJMgtt709wtd+JOj1SvWoZBq8tK2WulplQIRnOTSZ+lYvgUJje6V3DZvJmLzZm
TlPdaX608sxhewCf2PKffuPbHdyGeJ9cmdvnON9VtdZhfXu1HJwXSflUToJkCx6wJW8iMxQxVToy
ry2Y3p34HQiBo+yWbaySGHMhriQYS+/3jaOA23cczwzKVMT8aKF4T2CCP+d62ZJYiueGvG6Pibrx
qlPtHXlhr5cXJpfYSgQdEq1tIgVOM3vS7xdssZ6e35fVaJJUzlDgZ/nWendH6ExMQHhjnWUu1gQ8
L60j+rxUQ8sjmdmJsjA8Q7HrbaAWxynzJvKdZZeHSiBuk+VaevNTVZWize/M54lancSpgzh9PoRN
c7OUkQp9mBvwmEGevZZSjZnlsphdnPEhy75J29XA0btS6ietgLW1y/LeIDJH2scrCZyFAuJjZzkz
vaO7bu5YhXAWRrlebMK9pn3tsbKFJtXDcBayXLXkutcozoTNke9WgZRrQTfC5FakIYrBNCEyJqt1
JETOGCd1PIsSd49vxBiMIdIwdyLPjHKVdzsTPqt38BZfTn+PkDAUddRaOV+uMVqpFNpTZCB3An+A
QCvuxt4xQZC1WNRED425ZfUFGmhNUCx0Akkn6FautvF0CecxBJ9QYi23xlUBVC6YrwiwhYvDna5M
ajpxy3As30y37giJfLU2HdyeNOoKa4WQtEH8qT0KZSwSUit9Q0zRDd4vSFmPGnr95yQe0oJo25Ph
R2YjN29ubk2TKg19Iund0Wk32+t1U3d3JNnno5Y2UPcgKUiN7KmXvftix5HRdk1REOBPP3XRkb7B
qf5LLuh4sZPEoF5qGLtleFJgx+yhxfIcvhyU5KDWb4JlqkqlLA72ELn0UwXAcbsl699F0C+1C/i2
2ZhFI7FFrknK9sAKiyWWS2NbYiHEvEOfI8rvI1cquh+sAo/tx440nsAJFcj3M3brzUsKs4jggeo9
FvTKTw48LVAcTTz6GFuDWEOc7mMRb+kaH49bSAqLeUi8U0dR7gNyw3LgVN5nLWv8Yv2Cf2dlIimA
fl/fPJhz1/bxm5ajkaWwjT6zZvU7/SuP67nFLyx6VHiPTAADNJjIzCRQfSvoGLplYs3xJTezJXK4
ZOqimC1WD60siHaQgn16rL4Fuh7aIqWkL9r3GFz8u5xAyzGjGW6Vkm/aq4PVRwrflHGnWasxPCk1
IqIfmiw6tmVI/udAmQHjnSn1uYsQ2SgqQ30xzMIif4AQ9N2dguP/0PkUJMC20yIokeHQHTVHxES8
SISqNze1m5O8q3/EaOea4yzNhq8G56QM9eSq8OGx6q3m26ZhUpsarYfx1zAIOZ+6H+3xaTHPCmID
XMnGdeyh9vZ//uw+JQfVIyy1d2vMVEliO6wQ8TZtiII8o1qHMaQsmdZ5P77U6QgB7eV1dN8ZaMDM
LvCOTC3PDymbVE73TOmtugWMypIU1I/zCCFARoq2skA35rxhM5Hv19A2Cwe6jzYZHgfLeI9WI7AH
4a2IdTYrb3stLco0Jf4MJH2+CWTcQpORVz8tCN9ZlioUj5VJgYGA4AaNho4rF7a5yh3kbDJchUXT
pvRKGL3B84mVRLQZufqE5Y7jWOuAh5i3uhkTn/IMrB5+Uu/J3ANcyLhlRdo44b3oLy6nArVtCYMD
aeWnsREvEHnxUZZWTKU7qktdG8VEE0DA83cHcvGnPSqtSEu/xq5SvKfhcBwgjhpr9zIgAGmHmclR
chrV+tpg+Q7SW5X9dYW/VZlWicSn6RqfC1P3BGZGaFQgTvGeIZApxGPGxZ6ftaNnym2EvPcBmEGu
9jQxGz31hxWmSNPpyPLr0cEyvju72sxj7YW5FBns0+VXA9ib3uDSNOazfWtl74sVgJkhq0BMgPA5
Mo7jwmAhZ5ACwOuWloVF6OItiY3IfJX1zbH0bbuqOf8wt/Mg0LIEamiH3mOENqjVnhJ/JPHpXXxD
eHhbEdh51eq3CZINyrAiLDNm9ENLCscFhKN4qKhIhsC4Zg1Km5JDM0AMoqobmgH8Eu2Z4Z4YPXtF
dq+r1pzlxFvL1eNERWA+m0s7fru7SOeAtYJ4CRom5eQdj5eSp0RcG3xXvKz4i5SdMXPiyxJQYN1U
JyjvrDMn2fJlAxYWjyjes77Xsv+hs3TrS4p2FqAZVArrREtf3DF83mIaPPah9BQfpO8xth0ldhLu
8yauuIXP49/jCjiBvndZEaxcQAVTj5rXaYT6WO1l9WecynC/GN06B9ZWruCjMFJbGU2CU8+blKEN
jwkgJbZkAJ1uwj/GJYdxGAaUFbIu5GdCAt3u49ydjZNS7upG8mHZaUsK23AOvZbE+HtchACsB20B
or4ZGrp7mEnHEbYRjn3/S5J+Qh98vzESq3OxtnUyc3WgjEawVGQlpZUYQMfFtIAUAabp+q6kHx9C
pyL4tIwik+3Z21ghjizX188rDu1WQDVdZ4+82mWk5p1+hAMyxawIA8yUuz7ChxTkw8nhGb/weaCN
++4rAYcJgm1VgsZ50wsvjfGqHqNH/Ij1T+pLyV5k9UpKYI9TYFvW8jjqBXq5h5XT3a4MC+XovWGN
KbAF1VMHjCIhJ3BDMFLf/QI/fKqqUMD8e0e4bIPuqg0mTqedSgAnfBdTHZYLJNZxFzNrf1VeDlIW
6TgkKVzXJ+Pd7dM9qB6g4993R+/hegXOx2lKREo8PusFFGBmQs+h2P/bIzeimehwxdYcrgq+tlyO
mNQJ1qNY/anrFEijHFn5m9x0CfSTdZI5F97C29b6wpjj8giPFj5R7hSuxHIB1a8fgFyu7hp2aOwq
g4gCA2atI505aCvb2HSxeh12CvS8Ld+c0z1Cl01d0mFlG1EtiNwuscNCUnVHOeajwBHIjdBs4sxK
8qDIwJJj+76QcsAlwcm32HyJxZKUhK9l+SnmOQDAE1nmW2OeO1TfOScPPCdwbbp2jJ11T1M3r9rO
kM+9HSyD9hcWBITOaaUo5A2kcwnWFTdz3hi5P0tD20o8dyz/T1kGtIuSftgAwYmgY6Ac3Haw9HOS
5Iuo5TESa3KTlsuzSxzIVjEqDSqA6tY0F0DVbZ3Nell9An+bo8Ibj/EqqNb5Ne+CKUhy31CNnEPX
U1mqQqdAb4ChwBOebIrOuHaf96zMBN6/FzUCw5ePbk3lTAHIB/Dcl3pkydR+uU6fEvCttbDIONJ6
7TAdAtzSbE4nOqVcyARUIjXfLZogjmrJqyDzIgWpiRKNvfMWrzHZtLdAxriENTG3JRpRbHREnatB
xF3IR7WcxBuZke5foI4fKADtMI5ymLNskPc3XjMKbOXB34EiE6719XB1bd3I58h2DoAZDi5gEl0E
ydnxBtdm39hcCXbJtYLWDGZILwyPqj9jdbibnUsO8JhmW/0yNZTxFtQOKLRUiqaS8gAErUju8vnF
76jOwsdmDWFakP6LUiTNNYQUrQ1d5rK9jhmP2VQQB+dyjtxXznAiTzweWn5COGuUWaXq+nsjYCmg
oNYhNzyLZkMdctexcLzNcIzyVl91lFC3GHlQGJ3zNVxzuMCTx8liH6imbDCbEu7mAhNkok/6vMsv
Ec2RDTw8xuSifCyCIsN7XWe2J2iJOLV/QnNiGbhudEPFr3dQOAy8LIejQmgRMuwWfOJnF11QJqmd
jAezdD5H4AC8QDcP3zvUD/1QJxSLLqqtLZwUeoo6j+vtvy5Z6bD3If9filsU/OfdFgU0+kYaxkyk
ufVss+KXB1dBu8OrDVD3HF6sRyedfsySHhEEuOqKtYXuzcDKyH5d6/u6yDytQ+CtRfIoMUdlGIyt
rKqxb/ZK9pzN3Zof5c3SzIYgS5qZwBU8AjPkD+jHjM992zcvC/QaUNtWoQRvgKtkKSbYbf4rNby6
NldIioGH/HCYjjcYyK2pWZn30jI7vI8LqFRNMwx6St4omzNU7jZCZFnikVN6rEkMhlcsXz4KRE39
5bCzKOxVVb3Vsn1yagglFLHruQjD3HPF0Bo3SvjyKQD0zOq0WKu+4hcDRTSQmtqxhgRZ52SPUyap
WitrZ257SAE+U/1vcH0C6Q8qVHmueAQXCzasqDCAisDbmPdqSCDw0hqzBnW0yjOWrWe+EtqhGIEk
6WYtm+Z1/5hY/UOUsbjAFDFTiyA5nVFlrMq72guAglob45v0g7lTTVLXvtJVBFEXYbpoqhgjOwi/
sFZH22VH6LuXhii4udPSArWLuc4kxNgHtZ2z+skpPbM07ZRq+wGKtkFvHfl8LcwvBsl3IjkrShDn
TdFkmBdzIxHTmZXj5V90pvoiB/V4Ngl4pqV3YzLxPIG3oUSvbOqkPtp6dqrwsdkAT19MTrGh0+o/
ioJMeUNi9AyRbJT9qH86eLEikki16iykZB9z5V0UD/zGq0Ec8C2t3tQJVinPps//Lm8B9JGyDikL
Oqy14o8o+LBtRXx7QCpcE5w7fLuRWCjqfkJb6+pjb/dHo2OnL38sEtNHHK6p6npHgb6ACWTml3ow
YNQwyYnIZgnw/WPGDeym+ijQHwQ5vqagLgFw8fn2zIhj//MXn5ScPNZ2LEje2hLfatAZHlo9RjuM
vb5qnJV7MCuPC+rzuuCxZ2QE98M27cnOArBpiVI105mjDQmpsZckIDR/azcRKIeYeRVPU+SldS6N
H7IbqvBv3Kowr1IM9hGHmaRStKewxp9z3mZiDJKftnrjBZ70nO77aYvqYysXuBAPsEORgV4V9esm
rzDrLzawK4RDMWKhpgnBuqn9CI+3SE20/xDiVYU3fEZ1FQZ4Ir1CMFSuy8zla+tuoDTfXUrXnuJa
1lNHTDfz0Ovc6eU6iT4AcCWcrkv4ZrvXbClMQh3y5HAWtKohTIH2H1x1ZjrS0kUbTS1OZwdWEUaV
u9tr1F+5QuMK8vO+jud9LW0JSyZzDWlSgkag/XA82ioYzvih/Lru+/wYMwYPLxBSA5zRna2bar27
4GNHunRAzedXMEkAnVFFT0+vheWfPdsrwwsuGOFEtFYdOExCTaIL7eX9u49DqUwdujPlu/VEZpHI
nfsSxj8BYAJGRWdGu4Or7rIr7GQUjS/2q6eWBEAI7vwenYr77OkV/PmbN2oBydi5iqtKZA9K/8Wc
kbF5/5h+dL6/kGEnKN4LfuCDLoqdo38JlB6ADznp6DdILGhbjZt1idSZqca9jI4beZHJuDyjCoOd
9i2hvMdgYVk3efA40MLj08YWYoXnKszItacMkhYFlSWP9MyQdnOlpWuqMbxbc/gNf67lv+fFEqcD
CqAeJ/giwwfpTG1BuvnrGAuh1x3B5m9m61UrnN3xmlcslNUX6s2MchCNPLiW9eqx0JKDbBJwwq/T
q0KPf3Si5ItFtxHAVW7riHPU6IPkCTSsrynA3y0rZJpx3700hAb0G5cuzMdd2BbZtXkdzk+WPHly
OvBt85RF2kkBfBAfvi/BCbGnV7GTTyHst7idWP8rHzne3FsplQnbkefOG2j9n6C1cb+aC/wNvrkX
bpgocdzsJHXTTKPqkbVuO8MW/purAV7CPZ0pnGbJN03zJ/aITWDUkyQqQZMscnc9HztOtBZan1XO
E0s5v6cXQEDhG2Kt/wmV6cL6DDYIR6NvLh/nhsluNfJKB4qATZtQOif7e3vXE9/VTgFr7zYdYnnQ
Y7s4yxcGctP9tkY9qhAoEK6Z+N3ufvajdPS5MuOK82IxfeANrxViS3ngNiGDeCx96w+OUi7Uh2ta
3w8La7FI8g1hDfGW9zFPii3oG8Ytv1mKX53tnVuQ/z6pZ5RvN8tyy9lyZt2QStDvFk8mPTHysUr6
GYL14WqThxXCmOHFGUTRDPVX577/osqTVzrbEOqLBzqTvSAk8pgTI24oUD7P9m95HFVYuQo/+mAD
tFce7ratWHvjLdipv2hNDsKumuRyzQQH5mwpRfcSuPJLzGrDqLhkQ7eYKlUx8OxK3X7O6O5aRo38
/01HTtk61Q2+BKh1rduf8JmzBp11mVwrmw0Kggyvthr6/D09Ye3sGeqVa+hO6on+Ebilt6JjCU/r
5wtGnhqiIzku8UEvfWX/P72ZZ0sDj+5tw+bIDyNUQwS0ZdBzgzJm9Hgiv3KamqP0aECQFg3DyMpl
XimgGK0+OGlqYFF7fAuaRWUYfacLBeJecb9LvHTKwP1TzzixDxIrPdwRPHJRq/AwW9Tg/WPt+Y/p
qA9rtvZq7UKRGF1qtQOPehUjYfiiQzFnP1jwFhRO7QJscrjuGUUZ0CPFSKmueFHAOw7biPfSoHO/
a3DIcW22SHH4Crjr+VnaGgCVZ5p6WooF162RgFg2+MpYkW9YNdkYfNUxRvv/2VTT+r+5ZlRJ2ALV
5QbBDeyghNJabT8YMl2Yip8Qaq2FXMDkEEwxa6k9GQw+IYQcZhj3rM+TwKGwrR3Lo+xSqktvGEmy
aldR3F0X/+YVwHXdjpR0l0wR62Qro2LxsOZZQx9GVuaQhL2IxhZ7QuQ5NWryhCgxlGlQK/bNIAvS
uUPbjovblNpwKQjtmjIuyWt8ZuBOn8EiUXUnkQwRSG5dDyxMXPuAnD3xKjG7jVSCY1hUehenMdgv
XSS1HkIR796Pqv3dp/4uEwyP//c++SmI+SvgjVJ5WXz8tJEF/bW6aUyx9XTF8FRBjLlYprc9m5Of
MtX7wpuXnipvecxH39LHxL5+uGibJPOqZM6a4tNY71GZ/tjAcOPXtaOyxbhACmZocitIw0Phmh0W
t28h72F6RD+5GEGwbd9Hcgkor5vrsQcBKLNxXptz9Y0Mids1qSLdA4JANQNQcflaolfFndZO40eN
bTIWPgHcn3r1/+J3utsleBhkvfd6iOcSQYiQPA1XFcY51y9NL7sh5II1Di9f7Aqg9wes2lg+A4ME
0yu64ED8vyxj2U2/0cpqrp5ai9Fc7LsRCjLHM261wnD+8Yx04fHhtBMiqqB/ol5bKVqLS46w9fue
tlEizGVkxaiJ7enkHL0V+nTyttV/lOruPj3F29aMh0wIGidzsGmOHKOzTmFwUdTL86ZpEXFG0AVe
Wu4LH99WnRn/51SITG323r0YjpEpAgrYgXWFOvszvpoeeU2ElG5h3Uu18Tm3tpMj7Z47QSiBCPsF
eg8nuzH4BZidwk1ki8TJLS/+k3937v9Dol+1xqMQK69e8yVil/0wbMGa+8rTfGBm7uvR6Por0SwV
ylHPSqO5uF7whItBFfQRfsYxnfXGUu7o91F2GWzzHQyaQGlZM1I3fxRgyGL0bF1yOHKDlOAtjmsk
IC6Rrj/CCzOpFNpFuBMkKpdU5njTRJqFbeC/hIxavjJAx0k1mOjWbqeUHwcCiBeSsu+ayqYGX/YQ
nRMhnS4DmUSD6FJrwEkJ0BTIvb9m+DkDJK1yDgG1FxyQfeme1B+RO3zRBA/ryVjGtFdqqiuFj0D7
HCepPv95kNARmobHh9ef2NiByQ5Kbkk65Vv61pacfiVsDbb7ZWkM7BQDv5V27+cGdokoPKQ03xEL
LS6MIrMVN91kb9B1SAo4hsJG2efJ9iw1FyLesOQR89mLyvn9azRfzoYVmEXO9xPq/Xbyg35woax6
+DgHcinQrSfVqSsQznZ3c9s4wqh5c1MDjChqmmMnmziDL46jnK6IPPbEyMOZy7VheUPeUB6yWPPU
UDtjxxN+XZZLMnnWrDnQBICasC4Jt/rAe9lyqXvNdTFOUMxWPpU+IspT1IsgkKawAkKVon9Rfwz/
Q16P/llUZHDsJDaRpGYwr5M5X2U2TLV71cSCuidw4KexiBd1xTdgZhxbziTQcJzBgtyWeJqQ57Cq
lZRo5lPhGX0ql+i6TzQOE0uF+3gS4/NuU/OoDxEyqnBJD7+ys6eZ5BukS1+qoe3gITwDwXeN+tfN
H4SyeD/vE5GKYDa3HtPjzxZNflpLvt2xs54cbFX8k3Ln4oMBeWDoRc3DtVnCH8yvdgRqoGFTSgUK
m1eWCyEgr2+KijG2LWrpAQ2/4SBoyHRpn68sIkA8Fa5t7CJ97Uc9W43Kh9XnjcT2rovUyBOBg/Gb
aaeWwKXjKW91sA9JN1FIM8EI3rW/SNMjyqSdEfCfzMhaZF/tRqG2d48K5a2SFlzX3SLG19o9ihj0
Bmi0cx0Ke140K8Fo12ClvVGYp49927yEsiMfKg8TS9uyZgbE65o5/MKlEMbgKorNKkWcvbCFT2Gd
UbWRlXHcfVvKcM1ETY9E3i4d5SB/cm0cHOIFDsQhLoM618naMY6rpsuLb6xfp5t6hLmV29FbOwpF
44wuqmb4eT7W9PtL2rNqBMP5sS2h+8YKIPmSpCZwU1eBcwcre8C5JgoJguv8BKeEFB6SCMq7Dvr7
E1WsOPnIazSrVAi9f1to6g2E30tZcmP0MxA9hvQbfwSWWi6cfrM1RtDBGLe5ibkPd+xAYcqmewZJ
506v82Xllh7sujTBNLSo72nH5GgmG25bLkXRnofDpYpDVRMSg37qSrq4u7Zx4SKmBuN+bO5GNDUU
ccJIxsNKAJPrr33wBNcy/b1IoyRMr4tajF5XKwRhGqYvtlP8Sa3GAIdreFlY6r63qy5onZfXBbjI
Fpik50YgYDLkG548lrsqjqjMw3YCNHs5b2bjAVZfxadvvKCX/NOJ817zj45KCE6MGm/KpTFuoh1G
eOI+UfL28bPmD/GwUUXbMLyJjTxtINVsI5/yQhZGX9zU2zTGqCIYgv3xLAw5AZMoS+koSa213mpr
xLPG92Jtg7jh5RMguPpZ/XvZVpuQl63r7WmAHSKoXx0P3wXJEChxaYMV7GhrZC13Vouhkictit1U
ngdccPUpJn+4jMHiwWjvsH11ydh0suIbHFR/E4+wzPlDJYri3/0Y4l0TY+9BorxthL9IRTBgalwf
9xAZ92t6IzsFU03jptogs+nIvSQ9x3dpgWZ63IDWeU7Aw7wT7dS/syiF4G/u+TGZbBTWHK3sipvo
8p0cNS6n/O+lpTcP1jIn1LlNpFPrvWzKocyve/N7XLYj3TGKoMN8vpVLdZo1Z4e+ZUt1yslu8tzu
hPLDIFGDmc2OMNm7APMWCNzaGF71gqUBBdTSKG/S213NbAo2dgImEcC3HOKglKDFYIZN5pNN3VTH
vNeMswRSgyfHpbVxdtu1g+zTreklJJVsZN7jvXwkwGgMnhhzs4Ii2q67ErWkQcO70YVjGmLpRlID
+uNm2oelq1sv5e8yNiFCanFHPTiggs4I0MK2pf98wxknoTMf3PDd/vAVy9PzR9gKqeRERZVF1+JF
R48sIeYLgy0QzmajP+fDLPUKl6xqoWEHNXw7jR7zefarL5yQi98kMdEi3u9Ot2k7wgWh/VPJexHG
lfcyCiGQY6P5UVbAoKaqUfdZee/+xP652lH2JZxJURg4XFZ9DbO4L/rA5pKprBq3fBIthMFq+VVx
lWq59h2Me+4Cjq/3tp6Ka7WWK/qIypF1qVda4IB4wXxSukvg2sm8KX3/UrVcLAiFGTIT+XF2fDd2
PLulNS2ZaOfCW94EzGpgw4Ftk7RgHlz1Mx+hRNBlHQZVnvOyESjbz/5LtI3B5WzLkO2/yrog23AR
Rl1tm5BEHrrmqmYfnp1OjwjP6b7QwAr85gglYwQDu/YOjZXyQynPgYDyVgNchmqVGHEUQtNodAzm
BB8UJ9SM47pwX9IKdzg56MEzatj1zP2JBbrvgTf3o/u+gnxkr/jQoNU9qVO2KX55dP5r+Jp8H7A6
5JgLacYZXWV0gllngnrXmKF+o0nfLuP+yj+zFy3cYnLSd2sXe8kiDdjrpVOmxzHsUajd/ZHUyAbc
GKs4RmUO8vTWZZ91153BY6PlNVC4cqb7zVOQPBVJdAkAgbU3b2+/CPlfguVbbTeJs7xaaZ/woU1w
m4C6CbVqjBsfMmAYOxUIVAPE8dbtnNyLySNFJJtwVzQGsgSnNzenWD/BhTf7lFT8AOPbA/agQdw2
n3oAg4KlQMtWFApNjwXXaT7f/f7WHqSoeQCo9Zj9vX933gaqpZ9UIAxLQgM5bo8aXXg2oLpymRb9
1usdozPOIUEpH08iWLXddy1DC6FqiaM2JhF/WJ0Nw+RHJ5GlRqzOBgURK546telz4kl4Mla0Rs3c
joRexTCeK3c/68cU6F9TrToelsFXsF0Ry2vIwduKrnpR4M9EgjdJC+IBG1brjDY1NIaJmYxIudOY
RvNGCqxlm5Z0B1Iwv4INP7Ts/3kKjOVE4oy1K/XKJG7as3asRRbk26lr/RTIpT0IkmEwIwKKPiMR
7aSCgJOAEFk3zEuTa1prbexumS7Yr/zA4H/z3K0AlUWSA5cLsOGsCCoYZyPH/Qd+73NZ23eoZ2i1
OZlryPZ05qAjdl4bUX0gG+5xxcD9CnwvqMrBQ1hNWF/HHJTHjzsxolSl/Ko/DaDQlfGZ8qgDmx+H
syurf0walBj7r7cRYYBuGppqZtO+JqeCihyvKQjrKO31XGt78V2t617Ouyo3TOO8P1sgRtpT6Pll
frAxf8ZRYgtfZlkcck0rS9BVWmO+ren3PT9LNvVEp3JAEvkCnJo19tfbEnCpbAHIe4PMNeBR2rYC
xIMtO8UohhqsljoJOwlIM85FHiRuGcaM9h1JDYmo2ceVkTNKRsb73igOl79wlvQiQBgZJSGTPn7i
VcKscy9ak0oNCu5KWO4+4byNVJqcPyciR+HUQpdiIuWnCNJG8c/GPJ/E/+FSvZevwmz412hP74gh
cSSSiJkBplHCm/MCIlcZJno2IG5nfncYokPrchzy2D/fBoGPYUp8vZqdGp2ivEv4zeAMM1nueu2p
t0Y9MC7HsCVmXz7tnPTdSEiLqF4b+VpaZlNgZXaoWSLbxIfNyXiQZaEzXyLE+gM8E/1tJn44RqNa
nm+++7zMxfmiAqJKYGKScgTRjxB1wQYPV06P6EPiYu7ipPQa9Wx6rLoQNN2j0uF76LJLAIG5fhuO
qRgdRcG9U3vPsnxw+8HREcRXJjG1Jl4UET4+D4ZYyj0la8a/mBjcUwXOBu2EuV95x/aBSgP5Fluk
PmFBIU0BNGtD2ozhi8MpoVHoG38tQlhEbz6uhOfPiuU/f0QHFpgriY5Ljtp08zqSAEidei+gruEx
6K/fIlVRWCEZQsObVJBmEJn6yQxv3ac6dzywuu7LtupSrRSbjpNgRNzu3wJim8nt701ljGztdQLD
/fAvxbXTQboGzoaBoFqAw+X9DLooXfd/7/kY2wZ6Ewhwy5yb6QmgXzoQR8hmSlpt6P/rRhKaCDYS
uTSXsPcjRQmAZEpXsL+EQcKQ8+b+zRm9A0WArCRSBMufgODf2pzLgYYVVws1BnqLXNWjGhqyEaJg
CJiBaynf1yMPlDf0v8rtchtOqrvaTDAhF38CHMOLbQrbErRq5MRGXMyE3Mw7CBgYmr3k8Kl0ax9m
JlfoMxWgkMKThpbJinGtc1sssXAMLNDcgVql9mNWjwTfKR1qVrxFVxcEDJXmEqTWp7h1Z7jTrkW1
YkyJnVg1kPNJ9TvWhelqQJagDScb56W8dmtVECcQTwTSYUM5H267A4u9ye0ZkYOpiLRLfWnfvyf1
fosGXVA6DnLftSnSzAkFIPVm/mm1de5pAg5VB8YosC5cl8WnjBhFXFEQKE9MMBBlJak61qQotDfJ
g/GRrnYhTj6VMVsiuUoziSo+h1ZLPpDvkj9DLWgjmjGkaO+4+peVbxlUkDvniyOmJLE3HgwQWfRS
2o1kZ5yH0kR6Y/7t0eDLYgfQ/VYr+CiOk/7DDfP0GH8lYPLx1ad+FNaEMkn/wkllaflGcXI6isla
yQtQVB39xYQ5uRwmHf3gw+Qzmyrg01/M83Bu9Aj4SsLOMidbL/N7wGuD04XSSOhL3JqOqcXBc7ho
bVCo/g5E9ocq6+Sm6+TjL+V3u7tBDCFweeqiWo6yCAAHZVL15x+CtXFJr0xesNLRMZ3imfYJuwav
CCLfS6f1NS9Yze/YPsehU8/Gkf8K4l24Vja2RhP4sRKvQMs8Eox7BOmz0+BZz4naDIEY5Bf9OPB2
AJZHWS8eznx5svUwx1N0x9SbePvOeghrIyANtcdqB1KVcaewmmTXAWd1NjE0QeFDg0sVtilqLS4o
lMEfUtsVb2UWO3HI95M6s1RFUhZoX9Eq4XD9/S7Xqyw2xgmE6ohNY39/qd6bBLDgZ3is0CTuQ5vD
o7vzPykUxRyBEXc0ti5i7tJLZxAFJyptCGwU5cj4UO5+HfW/yv9EJY2vNX3I77vnR+7pWA4ZDUGf
fnpgSZgbATY/XuM7gKGDSDGpgSIxmBgSvXtI7KicOB0+rFx0kScPgIbYJYKozK1DaSCu9UpWDpRI
1y9404NW2kuy1ga3NeWBnpPgoPhxRKbsosDYWIENVxFVdSgL7S39OyBnnDGszO7cu8CFkAi5G0gR
8lH/U0gt7Q9ELqkYSUdHBIHdzSPma98tuS2iI1XGeoGtuBAQG3lyaoUtuXTbYt7yWBZY8C6etaxe
D2VdkCP/2o2p45d80JMkHMLQ9GsaHt0jw0mrsWoaiiI+v9GnDjnoul4CpkXRrD9iACciGgEv3ATt
SNn7k5XvJHOz6s+qIKUvB+Ou4KzLd1Tpd2yqtMOYjsQ/ff3qQ2NH4gpvnTuMAKIyPsQjBHOd0BDp
3Ld9YACMtyrZ1OiSNNw5K65qj2pKfglF09iH8cN/hzScyXKxoqAh6OOcIYF8Uo8/5hVdbINtyDJk
c/dPAoVmMRVXYZauj2M3EYp1hCBcDChCMDrejT7L6tIl0Xb9vEr9j7buVkJqT3Qzi1SptjERxFNk
Y4nG0Nm9SLLSMiIMH+lgRYt5r21HTNaMfsE9M/u8E5mqgQtpaUnbcPUUj+TSh8D6niPxnSxJqkF6
OLUYg17DjON3Xx2pxxg0nviCmNHRgJumNyAeQlZpVhH5SUrV4Ho+ojsRxuHg9hjWR+TUrgEN6ZCb
CJtJdYWX3tgsY87rS0QftVars6MwFfOP3k35ROLt7d/IYE1XPUqiXVSQoUoK3vTvXNrUj0RliAAi
rigw2jq08iTr1FQwMKsQudP3Ar+h5pkbS7kp36wvwtqICLcaAjpWsFL8XrFwNrABLdvS2BMnGXKK
8peEWQYFvh82yYTnRZDXYgQeWvolMSWZ5qBVNZE4ZEhDiP8iIdinrz1VHlEgyYcjXebzoiGPBqbo
TBlln54hzdm1m6OAdYAmW/Nc8dduSyuUIdz31GJm6ygweRRVZzkSMfuzQlN2/iVSp1nxUgD4u8+G
4vhCdsqN+O02a0OuNk82XfcPdX1ppMrcrDAj0md4WhwwiYS2fTGUhkHmzWn/zvZ0nH9hyhetNOWy
V/q8jcwbwdDOgrA2dc1pbLJcgkAQeEBGzbrUzRPorPnY4Sv2aIjC/mdC/K9JFLte2eQWh2ZtssJ4
tl8BxEBHmTDLEnbfR6vmiI4ad7mtBzK5XVxTrCgJLmEZdbNJLjkmRbHdlV9JALXd6RhTemDjyPDn
Pi11ovPeVW0ccxYnuO5n81wHQrfqg8DxVRqE+3SCk4qW8WtNLtIdEbqNrwBNV1xBnvMMR1sNv0Q7
goFAwp5OQ0iRCyYcNEVqDUsTm9AVnPiHpGXitMNPLIM7q0O8t8xngfpW2RPhF7ZsTVjGDy9aNSdI
cV2R6kZ+jb/JsNEbK15P7JQsqrQeAN3bo4YZW8pK8JYEshmSBctYZek4pJY7XualF1/u5b2eN27o
NNMKt/mxWw65UJTaCyTZc+OcknBqQyEUF7zz/TkvselczYwLsbAdUaQlDc/85JqwqWm12yQERdCx
I7Ydr7yY62LSkjPofLCrx1Aq6fe5w/W4gq65gRrLKue+lqBZkpeKSLdB/i5enQl/U+Hg3dt+Rkp2
jXdBumHjt3RvJpGWa7xj3BPzVFpt+pK4Sh9laX/sAaFwJ3+Ru8R4TkJuUYAaCf8Tr9pcWBedwTpj
uXeYQHUWGX6q5M+ndsccOsei2xu8J6+DTdnPYAS+kMWMZVbVpo9N00LLtrkwjAsKj/v2qLi4l1V9
wrYMF1TpK0p/kFzCRojPqHrQbOSUBpnuKl6q/qa5xamAJXY0S1IOcMU4hPjQgyedye2/4LuI5fqk
EJdGbLTthySagcw7lGpfpAgl1jMZVwjpvcjlb+SIA979srM/Xwt+shaFOctbyJkRdCwXmpn/Ph6q
MqJ+xA/fS189Xgeu1WwnqsCSertKzescQkJ5kozAdE51YMxYF12ESThLKvo8wE3wlbTMNkgS8iMc
lUbA9+i4DnxTjtiRdTNy9RwaSyd0Vmg7FoXYuvO3aFc1DIqN+FRVgWdHlWIwoCojWKQbmsxP5uU8
nB1h32A5IuPalUwv0RRttgHn65c1KrM6Czg+lebXB/JjQycvob4HDdKRLk3vF3u+p8po5RsSwrE3
hC1TEWwHfHnDVRGfHWVv5dlHsC343XNSaP8LrVKYJB9CTGIRX4DuzMu7cE+cWoSXu3OA85b1J7Q0
YdJX5WSq0rZv1dXihLfaRVrlMrHsc6TlTuPOBPeWR+Jxe6AeavV56rApmHxvTGtEzSpYtTmDkLI0
wsj4Bv27x/HqWO7r5c4P+EzP2qBR60eohc37gJyKHXmVDH4kT6iA87IgtvQJ4/L013soL2LiopHo
DOzIlDBUazPqLAF4XoNy96NSG9omUjdKKaok8QvDH3Tb0xe6naQ7Fu/PYV1CFNGgQpilp67yg+gn
hqlpHdFJAKOQvHFCIAElLtV/5p3dYlJMshBJzFnR1PY4b8Th1OkHqJ8Iv0p1OlgXSF3Pb27MZFFZ
SgpPzEEsAW+FapR7fXKUS8WrS9i8LGh9bbziDlpKxCycUC0/5pnkYp0qusXSK7uuUxIcTBjQA4JC
3I2V8Y5CUVeYegibivVtQM9w59VIZuS+fdxoVB2Cvy/GkuQdF4RNgf1zvZOaMrsseBNqGG9LF/GK
7gtb5fEi/nqfUYVryIUH5Lt/8XqN3WhMAlGvGx9UInRbjR85I+YBWly1GGTX4eEDIbXDkp1BCHkN
aIAFPmzi9dNSnRIhf7GQdWOGifOzuJ+u/UJnusaANU2UBDNbWJ24MuqU2lY7ZSZ3Hr190hXqSQI7
Y6IUvA7lB/eswy4mUJuPYCQJiVR50SoJGMvfcOSo+IO+GNJTyZgMlIgi003ptExTR9U1VDfyv/fM
J+wjMs7aZe7qbN+mJglrxezbVbQy8wD0BlH13WQ/Np7O+kXtxgye2fX8/HH2ctXG/aeXMiTvO2OM
R+3vMWEhMNFOlyyDuv4STDGEIanvqASnIFGWBSO7yUjqsFjkSJSKwUG3hZSN2Jn3Jc8MkC84McgQ
Cq4Mh9ju7qZjh+jftYUsVmH6A37FVLbyazEXZCubqVeaPQ3p2rtzRFqocAGxOuzw07uhkgmZHVOs
lDrBxRC7We6W+jDu1cDvlF6Lb3Y3P8u7h1liZL/wMrSSwu30BLuWHE3ha+ny87Kks5De3NnLDGSw
lryBcovyoRfZZ4jHikMt4ag7dPYZBmId/AHKLfUe7XG5JiPSIWzeY6GZrQg2V0r1f0lHqtIXFQ82
M4O8HTjAFhNrB2ubAzR5lTHsScMRwXj+T/IcGQuvlaeSbZXF8Q7gOtUKA4WhN1g7hbVyC6YOyCn9
8C9GTq7nezdBCGgYKXw3T5SgJhQT/AfzdqYb7kdHUJfS+jkSltcgwQ7acjTqOOOqmLgvRS+fKIjA
5v067TzhCz1lvtyIXL4yJcSOB/5t3JesBwqFp9tPBUYiIsvsuCqOAU8b1Q5Vs7uhl5Zk27ZHXgxg
UTc1beV6hrLdS1SLR3A2RYcdm2APcVxgsDMYQv0Y7zzzqyQCULS9sCWUTjWzR1K6VUyuyh3qPC4S
NHyUkT90BDiYa7uC7lmglkJmgzesO75lro6UbGJL15K0LOD5XndrpmDf/SWeTSb9n/AEcMQ8RUrt
RchtlKP4tx/irmKrRMRAlH2toVxcEfiNbVlZ7Zd1EQmmB7pWpSmN4Db7ERmk2B1jGKGdBlMj7Lhn
Z6uUYhWVLZ97vokG5k4hC9Aw/waB88PtL1tDLm995a2GbSrKfFIULoShF3Jj13RCH6WtH6bArXHd
YB6xxruAscW5K9P3lOcBvOHwMoul2iFlp/HOgyeRMKMY6c/48tZSXzv2wglkwIN1GXsdc4xpGMPM
IdL9KnAPCDagVJxWzrPd7mtwP/d6tafbuieoOi99i3bdOhlQy8FG/5+JaqHgfc3om5AhzKiL9Sr3
7XF2tXsMCnTiNXWyjQQR6Rc1qjxch/1coWUj1MXE0LHjahV88Fy0A6enHlfGatnOMYw3ZVw2Iswr
7cyo22wPEEARbFYh3c4BX9JYMLcUgEz/i2vU6oPnKougQWSbZ0grc+rcjSTOCkCp67foVJCg/ftn
0N7w/oQMgrrtRWBJNN66s+wfoRkE4lOQ+irpyx9F7ISu5OzVPaOlXTuOhnSFVl3bwuFbnvF+etCx
mxSZTG/gIO0Y42yc1cVvLqGff50bJizvnIJebtX32P+ALsJ9gwsuujkMyv6lYevuKq3KquNtGoBt
vqM1zXDHC2KIhgcaMzf/Cx2fUzwCs8Zn+zjXoopWb4N7GPSLO5P9cKGGQj9Yn8bXwihkdJQnRk/+
hoWsr8BeWr4uY+G13m20GjF9lGZ3maBXg3h/lJAHaZ8ajTv8LSmCsdQ8Uo33yzeyKXAvG29pR64R
ps1cf95MTIdjROE1z4sMQRlXHbrCZ7R7WSpjsY1Zf6QVWobD7fHZJkYEYOVQS67dYVvqxNjXhv4s
TaHz6GkNGwG1hlgKhKMqEZhvkKFXpi3Tn05o2x7rfizlNMu0sYcTEyyRBsr/hugfTfBfZUdAxVaU
8Y2J5FjHAOzvLbv6BLUfEbGoH+Gn4H7LnW1+VUTkUv/s1kIXIK69fazchZFQyycbZou8qQiN4zfw
uy2qusCcjp81wfDp5KF2jf0Uhluzy5N/XWJvkhjAf8Oy5Pfwc8XWJkLYM2Bo52Mb8BflgP7fAuwU
4F+LiFymYUZS7i99JvZgBG6sOoWodoBjn1HmFUq7FplX7TeVXYxyR+zpIMHzgNEIVLHKt2rp7fBh
XZnkxQ3fn3hFEHn9OebnaxrfyJhc2LhoMoJaNY+hSpswOebtVAt6H7SRVqfgVV3cq4+f2RqesQoD
Z+X9LhNQNuUzRH8abfe0cDdfd3iCrtG953LIiU3Zd4x1zgSFbGB2BUXnewyVRNRbqqw65a3et5KA
JZI5CkHwjP9LoQE3s721qPiUounda2Pu+orFOseHuNgsLQdfX0gCuWqSGU07JmmUtaM/jAF7IthM
AkVrJkNxoElJ9ogE4w7M9U6ljXNbE7LOoQP+z+L0vyJdRHSD23XCJvqB5MILT4dsoyxYC1tgaYB6
PCWnH1s4q72E2TzN2KvbIvNgAzdLPiBPIboM1OTCr0Qx6FkrAL/6Pr6VPT2mkxQk1m2Uk+ANMVym
u494qwr5o3XOCZ9ms9CCYd7OA7zkZHmJJ9xULkpuFi4gyqc05JgrMU/xE8yylkOp9ZG9A7I2fABf
0Ixrg47YO3tIu3SWKp+wsjHljb30y2SINvy4Z23zPi1HWhbMz7cCg4dEfWslExTGjg64L5967Pih
INeq3PXfoDmJZAWpJYxRFvlGPabeQnA74MX9/YSDOD8LoQz3SSY2s1yRbUjNZL5P/NeDfkIr5MQY
BaWEuWetELRhujqkM1k7RJDHz6OK/PBpwiZkQvxQw5aGBf6F2gZTjbCkUSaFfC26UxHVi3yO4GmM
RYVrNs1Z6XqHcJxkjmxJaVsEmhipMW5XpsAZqzWsjNGKcFyEzWyoMUVPVztw2+RN/hkzdFP8Ia0u
macONrF2S7mOz2Vmd1h15D6IWKjxQseYZqyaS8e/cMCygfgxJoQiIYSc5Wec5qGo545KR610NjTY
oiHclxG9D07CRPdFymmn5vlHWcwKEtQs+VKr3JdUgH9mcohORAVmPhxKzVGsy+sD0uHvC/zUCV1w
lLHaaHkb+InJwPPg5cDB/KvqPvdBIrhnbpVdc5m89EkklKABfbyQEBzJNTFyiRpnjFkAcipdTUN8
f5KMUl2CD6VxmyrX97bqCV2BQkDcO1caaU+JTH5Vt2ENTrDEXrh0ni3hpd5nFp70RNWWZZlMIWit
EshkWBHfLMpwU0nd+pSH015mM2TKngdiF2P5PqYMLoJIRwBZCQphyrZCTEthWHNrlG32qZ7lepvj
NP8+fZAv/4BiE5qyb2YRL1piFjJQew/Av8jVOYAClPMTblOHOceKvFAZ9HZeo9LtosHb3d+ieQHU
FXNYxTzuDJ4haZcApu8AjVPNjjWyW88CJwn+/eVZocGVHsC3Vq7NQjFbcnh7IxCCK3wOOExlejkX
aZPLX3DgYwyvQtDQl3nIfN2JPKh8+r7wwH0nNdFXXFaccnn2SHkqL1CEv26BNUj38jrjC2HUCWyB
VR/lx8F+tiWeNdlDqa6eYy5vX78Veh5KCiKN6kdL7fgod/NVs4nxulOhOiIiO/ZGLbGPXdl53uae
Dl90N191HRilNAtpLTbvJNxCf7h1hl2z5q8JNEg86T/AShAWE9MBJu0UhJBkogv3dcJq+ni121OK
Q/10T7oSaz9A0xEgaXkwlGqWc6nqDbo9YyCyl2ErPWY84+6wbvMA+tygRmtzpbt/BcRBENhuPCwh
uMpPYmOvJju5CdAuOY907ENNpcUJ6zJbddAmBgIv7mRpBpzIdRDw8FGWJM+Sl6bWI+j2WqM5JoRh
eQhMZOVnfk3y8nj6Lchhvfk9KE7zko3HQrYelJ9PPsqWIyMBRNnYXh4ZGlRLn4FGPXrpuHlQlRC1
Em9wv4J/7TE7VFmmCtHkPMowJ0atW2Rua6638AMo1/buGbfoQbAtuK2Lys0OKIRO4g+Z2r/OeQTD
J+YZm8HZ0YmoxdDzfmxxQuvqyJp+3uuHmzR9gNJ2hELi71p9b74KWvTpEkuV2B7f1kaCfmgf8LZ6
QXV1ds56F61QNb0llwAuPxLYKOD8PIHHECmCqB/lV3pHsQWkseMiwixoREnTP5FBNX/ssr97k7ZN
li1C+SEl9RNlkGnJIYes1u1K68PoWDi8lTn5DD7qtbGjXZg1poZLqI1dIH56+YMyrgPRvs30EXiI
NMb52NWSshmRoYpPHPrteAxo48Wg+j2OCjHk8YnJ/ZGIXzSx6ubOnetyZ+7v/qz47EbyOeNeHZ7V
6q+fx5E5OO5OXk441GUfiaGzTeTnbXDpk2zR2yekmgox8HsBWqOoxYGZ7iOnaNTR74obFAP20fbD
fUwSuNPGN+cfg4hfImtSCbr3OGt+wojysnJKdFdlOARKnN3GlPvWnQYkewth0C9OYENQG0+AIqqB
X/P8tIbsOwXnD5k3zzSf4vqH0yVoZbMCO31uOV8CUaYG8IH+CJRHz6ED8dUfRaVubeEQ07WxHAlv
s0noBj3wbICsxZ6EjL9bHFSlZQIRzpaFdo07HEItjGsSIYYXYrDodRmFC5/dpfCdW9+2q/tpC4iU
fmn/u/MoCoPdmqIg6ypskcVdecp2UDNASmy81xWY8c4k9VI6uYBE7tbYQ4vjHFFkjOoc/YRpdTeD
wIJ54lljO//oelGRSsWMaZKxpsyzOxEja9A2UZN9UIKhfkj1KQTjq31BEGxt2XS1TsIOBZ0DsSR7
whAH6XAXvkJqpU2liBL7y/NEjlWoTLXucNcz399WR18yBkgcCOzXeJ8dTYNN8CGnk1kSAG5ijc/e
1J2ZGXS3yB6zdkNldPxf/vIjNO5hMUo3YZrs8usQYUi/of4OTZxtMysBV+e6OcEf2sNkUEg6AZLK
frwMac4qtGe4S8A7I01GdSVA8H/V/dhZsaJzPvK6SkBlrIGB4WMg8aW6Fl6m6niG/I/kapzFDG/r
HQKoVFjfpkSXrmaTi4egs7eL/Et2VhEbeDD3p5P9Vvo5022fih6p7V+/5KI6rn1DSLnfa/9eOPJd
fslaq6aXKzvJRTzDB+ioH5kmJT5BierP4ydYTt6E+TkZu9Ac4ZskIMDE4ThnXmvzQ2Cm0LmdZx0p
qoWLZ/IRwKE571RfdV09PTTaRScDhJVR+DOCGMU28/bRa1ovu468G1ThDjln614Za5hOqXjxEgqY
yFbUp5xUD3caNgc2wXLD/imk7FxBQQC5yxsa03X3KHMteDrbgbnCrqT7rNsUTwryRynVz+KwElcm
ndfsIrIviUHEDzNB5pU0y4T44k9LXxXwBQtERK1kBvKo51ymqrGquwYl7crnpMzjQ+wTKaW5QRPF
kT/BsOb5NNeX+xn6fAI2vuI9bczpIynMIIs+4x/xpWSxN0/cU40UjEkq5rc3PBZb2bOdS3skWZ9L
K2Rof92V5u5gplJsVk7EZlLmL07arjkD6tooAWKhlZO7JsFm5DaDUjh9V50GtkX20E63sj5aKJxJ
4MCMcNdbJK7GMrEsuLFiez39VrFTa8XPveu/3MCWmJVgZiU7SiRrRTAFlXN9VepRwURtotmouj94
nWazry6qcQFxleTrg/C7W9e0PaEjAfCOptCz7Ag2x1PTmSoq9C6LU42zaEE9v6oqtxw7T2fZ1ZTH
C4rTpJrFjfSOpCeTaXp7LaX9Nluokwngv9JhjmtfPgjOpP1TtibocVR3RaEwWVN02V3RWdN4uD0g
gJRsSMBSXfblwXFTEZ3YlP3mq6roJpG3Jov/birucYJSMd61EJWjmJ8LYZhelrg11c4Ie9Ri1dAZ
xDkrRHbVlhTKauhABHcEnmo0p9bVHDGpEtpVB23auMc6nAMB0dIwdkb/fg49d1T9AS7y0Ee4ESWW
JwkYeHvczhKPlN9VH5RRv8OQ9gQwOF8K1WFMRDVwl3NZ0F4hl/gGNeBaRT/JIcO1V7JsUs31hWMa
2TzAYdkR714/630i/gZrSkcAF6ZOI3irljgzJIpxSHLrHtfw1f0P2R3K/CLJ6O8+YWDruk/HJBGA
eTKKzyhkYgW6pgi9QHlyFOFsOjBCy88go46L/RV3Z+B706vZKMb/cSFwS3j97Tyywkfd1XBRm9YR
rgN/iWUU6tpK8F2Tshu7I1OQ5Vlppa7HKhUh9j90/gfwzMzSnW2H9QTNuJIJZBBQQFVGvxEqyL00
ojr8GqdFHslc22eXrxTUZEJDtjHxSHoxX65zmD+Wx2ADrUfHA5qFvXpGUYeIj27dGTaqbAXvPJyH
VwKvzri1nELkdr2Pp61x1AaZAN8pB697T56yiRGmYMKA6zS0fScCRyPpXfcvkYy5lll5bF7yG7WW
hks82uYi5kWfRSUmIsb8KWClIrOpTFV6+AePpqN6nLMf81shgrKDLlvmAMc/OL7wigynbd6nPnLg
BM5oEZZlvQDoXFg25AUZTg/uSe23iio9f1SJdJYA+mrRr+ag1KYHNrgyi+j/O8siQjwc5R9Hq7zE
cUgvddnBo+hHjzFuz19g87dwfyORwKv6yJZF9ExWzPeXbZjVZs7UdUBj+i4sDZ5tVlC6KwTaeiBv
FvWr/fwryT87ZS5rZniC02KYjGHGUdIctDVTsJi2f9o5buDkaIJuOMmlMlfzACYclCwWu/KVia35
5bWwuu4/qeQeKeCuidX2juqPfvV/Ei8uy5gAp3vxkhGZvX32aLtC0eB1Ae4bb89B5mSAWaWtUFyM
VZIbBF2Bo7DYDMtbtxtz00g+jwwftAG5h3cHZIalEinp9tFn7KjLxaXvbn0MYY5BuxGPe+j2wt8m
dxmdSDobtml4oH+cb5TrpCYtYLpDPJcOLPWOReg2lLomPyFUMZZ7VndHestMlbl/wh64Xl8tQZDN
xfoal5JDrmyW4jdeniTu5ESihbKVq3Dhu43Ouqju9VaamVVRSKZY7BVvsIh+5Cv5+lh3uV3vYsq4
wJYKAyQddDDvv0bcUdRfLSwXZ81FH7xz18aPolBw8IlR+Uv5QZYcYwCMm/bAae4IRCr225YPSTSl
MnyfiKbIMMLmlDncM1lOXM4NKeP0xFWbYSuzll4jIDW5DyERXDvN6URYRx9oIN2EeiUBk4vQ9B8I
+ZSyuBibgFdzb8hNwprK0a96Saz0F72WMFL2HtTa0WE1DeiSnojfvFz1Yae7BATgkbs5CcvS/GN1
Uopt7Tzl18xJIp7GMr1oz9XX7aExgb4Lzc4tb6UIZb8TNGfXHufO5tU+jUMrCXZCGc4fLOBuVbwI
H9aZtpT5fW0XBWphcetLGrHhMgsFlVM7YhNISSqttOd7oir4u/HOlrkJycpmU34SKGVUY4KMskRD
LfMvuBSAoxKfKcQsSGwagxYnEJ+SOgbB/PFBAqbO1W4Sjy55CbB0jWNSfvNpCT17D5Dv00D8Y7af
TxcOcrDN/8TVtMQs39EtOyas9jAfLGG+dhgiFS/pWlptuVP3rsv6FBMemORpOVkn9OO9f3PPiW6u
wHlccHf+twg37Ir9w1yA9/WssFBxOuBTnXBPioIJdYk/f9SbwbEVAiETzx/E8gpKdIP/yUZxldYP
GFSbh+zANZoSy+/ML4FScLJ2++IxUq01Zd3TX/FI0nX/VWpM1z4CCmCIpUUxz3m8kRZVp/Zamk+9
RmwLniFk5myj4v56NhuJXs8XPuUq7H10YlGzUOmPDa59eheL/cFfhEaTE/Wk1k1f5YLGRWul+HP9
iM3Ld7IpjdELztELl4tAtwo8ac7k9xCnejjy9bgnAeiMbCpsNSPZjYQg8FGc9ksKCHRaQhWWeS9+
QBppQ7UDWLPAQHJ/QbAAOI8GO8AXbegL2hh4Y5z5FRECPw9DuoEeQRG1EH6Nf6gwpNba6JBWmPXz
LOEh+9MgaqJwP8yYcCgNeNFWk+TecP5PDsk1Aj4XJscomePxwf4q9sjCzDvlFhhx2+tmI6ARvdez
TxLMjAuQO6hOPeE4V2MAtGAWNwAZSm97eDDZsXUh5B/R/hxxDwjng6twhb1Il6oI3GF79vXv/pXw
py3EYJLLu/rHE+/ChvpcEF0edpYAh4Qu+pheEe8htERmlp7RDIIfbuwNFYyg95TN1xjxdQ8YOtlZ
1/jnUhdT7QCoNxby37JqE635IdtMcFQ5IZbGXqSno9fLQWvo44QKWcGcvIHovgHJk5FezT+FpvOe
rCuoVtF5ilAWWP7dQIUna/VLOIc2B3QJT1npCe7w6LFxznU9skwG37ReQdFp/0YgKqotHBEGvKyo
L8e+wM7d51oySTqCXUrLJCFFlSdzyO7LaT29d9+sGvRqF6EuxwtixK513Go4wv0n+0ZZ6FIh1Jvw
GNqEDhcfY0Ly3nE5dr6g6paXrDRTr5EdN0zmgodpy7URfkl11FH09IyHtEnEYjaC4D8xnfDsvUOf
ED2/k8ZrR5erkHzNfA40r3o7C/I2er0uxUF2DaS1ilQMwrEmbElSUehLe2pCkofC95fB7gC1GeMw
Pm5GKaehM+xzY6UQlRPLSvPxZ5VJ0yyBAzLAI0dG8JwsPSJy6pHaXY/17ycVvijxS8X0G40LjBDl
1AtZokYGzjq7S/FFnx5IV0o+7RA7GxAvAXFQzsuLIFONY29CrdtHFbxetonP2Cj0azaLieg6S9eC
Fpxsj/LzSKj3WqstdtjsRGyVlfIIbxUHtD/+2eNB5UU4NioZPm/0mrosuGtS8Dfi7KQieqVQkBkf
5INfotvXIXSLZhbjfOjs/JIEL6amFUf579+eNOLxeN2SP0ou1rbm+/m6rXvcfdtiCC0Lgszk95TD
4oxPDNpcQc9rQLY+l8priqHpLsCp1pC9CjlwApPZ5K0flEP/elVoow0O2jpy2G3lrYelj1v7VvMA
yVkMWWDH/Z/ViL3RDcL7He5/Xv2W710Ac6QR2LSdrFNo7MVlclWE4j3SR4sqOjXEnLofFCRFZPnd
57T34w97QmDkOnPilkXV8U+ETjdxqN4W7sdnPgWnUjyuHfLDNmIu6adu+biM99EbM8KFp0cGEXD4
ItELyO4Nhi3RVBhXKcmGkfXvNKB7zatG0XfMmVDDVnVsV/dFTYNeqzLHF6gWdaq1InTQJyFuvGry
WApQwSKEu2RP7gYbW2Ar2+go9IzUE7aE8eunWdaTnea7otHe79W/UVyB/P7ksJ5dBTYlALkjO2AG
KcoXw3iyDSpYTmC+NlCPg6YnkH4PJ+eCDOsCe8JQbgCfHMk26TfM/DNlBILjzSUrV5P9p4gTHA3c
Z306+0XFRc475Fn4v+WMHaTdtUpRVTWU6YocykB5jBbeZILl+DRGsTjBY60no0/BWmJm7cXh1Rdt
7cci1ZJQyEcTqs8sVYMX2el24WFPPrXfy/BZ1V42cfQ8OTiu/oOpug3oPw/7agsKeEudJaSxsShG
jYzNUIafESFs/9iqlHOQzXPgbLegeU4qpJXRZUsfI8SFwboHksnvNIfLGGxbzGxCEPWq3wrI8mPG
n7t6ULFiRRvVXTHl/AO6r1F/OHALgazHVa9ahZ4t3zCEhASYL9vfO01UYHCm9xxPZcjFjw73elnJ
RkkcY/gq3c0q7lvRL46RDxYbu0LjiVdTLIdRVDj82i8AzC2ZEdhPTt5dP6URqgGHAMHWz3FcsO4Q
i5Wl5do/nQbhRAZX3eXdbwDUdvwGu6BpuZFxUevhl3c9cL65fhT7Lu/OVtji53VJ75lFSMupikeh
ygNj7dNuGWXZCRRw5RNRli21IE2u5d8IxAwKwExPNG5Fcj36Wr3c6akFWdtQXXYxmtSsxFLQC81o
mCvUeUwQTXFyCZjr94KyK5G7jnmi+bUmyxVqBnby8t6tjleJue/MkkRD7X29vfc79pYfHjQzcQW7
pCAcWGThATIxmbeS6D8ZSCiNuOXSgXxl1Hz3aq9bECcsZjUX+D8bVkzikzByfD2Fxb6ZJNEYCaG2
B6SrKc1bLSDb9b/8XOCipStmmQlgaEpLkmTgc5wdHArtyWTV7Bho0WBtXoWsfPq8xuJ4zicyvw0Q
ZrFp0JoP4yuvhCb3f3Sb5zMsYhyf0ZaCvKLpgHxJgzmTTPozBZNlmdx2ENv950xckkkpzTrtevKp
Z6Jcu5PaUXCIhqGQTCOpwz5AgSATTdOkZCR92jv11A/qMZ9RqgGEYrTSoYOJJIMMgOWMYbdPCWhk
1LMG4xCMwYDYEwgrMY5eEqYdrqXIr8h+FVcynPAT0KWcoPMeKVoSh7sYLkju2RWLvQxK7mFbS+rm
QtKqPd+fBZvRWHQmUq+2PmfQlj09tdrRhwYhix9cgv2szoKONc2cb3xUDgqjq9oQEjA1rX5qQ9Yf
pXYsdY+mV45QQfFhoaNPaamlcjfNZSryu7C3ebSV36wVEsgHTWevw3khwHHGXYRGbMvVzgZDWHnW
wgteXI5GKPln2wzSLFyhQoXy3ElCxDiQ3O3KeFkOQNsZGgFOTjLU/NxjuZ6UyoyzMZ+duC2akSzr
ZLKeGxKq1mIoTrjadIexIw9u0P0RVI6lE56Hq5GCgngU+Q4o8j0Jh8aSZyAVyXCybtowlFkdseDC
OCVZKYidG55WRMlmWzp1c/VyH0YvpZvEErcwedQs9Vz6Sz1CkGLA49VU2jJI5ROLG/+yLCUJvgv5
y8WTbvW7Aj8nkWwdGMbNLxP2vngxFtuHp0SIwRiUrqjyilwCAgoyi0HRS3/EE8VU1w/H2vxxzCOd
0dHJFQ+p5r4d8Rtjgzga7mUkvfZNzZqkVl5XoXJwyxytY7OQAJ/VbXFhQPE6hMLViCs8POTqMntO
+0nba1DcyDxsdeVes7n5PaXQXh8lzjnQ8nECCgdw/4bBsScXZ93AcwwWOsqH4uxbCnxFqmyX/y0p
7YsPNi9B5BmesKn8RsSunFWBuL4ixX4jr7jETGsu7WWGUK+uXbahk/190NN6ZDM+WXeakGm1W1iQ
//3TFEvl8d4d9oJMPiMd3cemeTI7EywNI1766HrAQf47kXgn8QAouCEbEJ3yO88gGZ+SqL4T8bCi
ULVflkX60y6+wUunTjvJOyjYSHNuOaet18QvXbVlut38O8pdC/rrfRpp2G8aEe1nUFgmlNqIgyMt
LSTEDoUYlQ1jxomBMbEQ27jDQhHFn5FpYSPtmf0t+lDgO3XSAqCGKLWqzIsNMePx0FsXYxxeSAdv
Xhe7GSrMhgy8JA3Mo//pZG6coc9koyfqwoLmeceozGDYONLqXSzJMm5q8JWFWgCxCkP3AIqetXYx
tdJxOWm09teBmyBcYkHYb5RoiMA8WyBcVjBCiveytbqWpy5PXur5niFDQrpi2qZNgs3YHAZwgY3s
CzMP7t7wyOupkTrBldfCieiILCqZJY+kuS0HuDKXskBDXc6ckq8uc+UcFZerwXoQfjGi+J3KCoQE
KDrdaxTyFTRJeOhnF5OKR+kreP0XJ0xiY/RXSevIGsK63Sv63TXRpCO2HwuzCykOwwUGTUExTVLq
4cUd3YIz0t37nstMvAYI3/PsLa/93UbMZqJowSZIDoQA7EG51UC9+ktoMwcKpv6Is3KDhIhYsQKf
S34O4af+OSmS74lQ6zsCcVhagGhMjIJBTwJ6LvgFcfMYQU6sejKsoKBHmSTT6/2IdScCowVi/ac1
zLrEguwn0rLyu/RLhY8pTh4lG285+30vy3+8APnSwrBVdqPvey+2MefWjy0dPj4b22hQUCY51umo
4Z7unCU7/16tTPbB5ohcbAuu6CNeq0QwIoeusHVqXIcjSg1YS3MlyFrFb68pZ9A3dN7xHY3SjdpX
0r2TGn+i1sBFlYOjP7mooe4bfAIOe0QOHcxfIUkP9yYhfrTziDEFPwE6Pnrjje3moNaAemJzbuOp
hkT+/kJPLCyaGVHpMFCylk1mMlVM/Yi2GgkuFonjyPZcfBVHV+FKyt+nz9JmUbu5xxT76eKoDTBS
wjXC0/0IXRZpbpgOayKPxwhUGcSwfjwFhHt/venpBPHgVuwdHh/E7Eg336UVyUnCMHexd/I+xmkJ
hsdlL9FVqcGk3vQXfGSL2/v/qzl7XoSpLET620Fmg8GFt9JW7GcXjzVOaU7HFHh56Mao5lQ5nedd
a9YcxSqBrSrAEyQqfDYP6kpK4pCnM1mpckBSVHQyKaBR6KulzCBvCaPMRSZZ5Rc81cvfA8WB72Zm
rXObwRGdtnUV01r+kFIvcdrjnSL9aoEQrMvz+ToLAlIyaXuziZXzCTzdrrHoW8e9TXqWJwl+0EQj
E8sxPhMzt335b75cgUTUx8plJXw1KhPajzmCC0x4OId49lOnZppyzeMTseLww+yE05O9p2c5nLt9
r2MpI9PjAsWkQJLrF7i+KVDTtafFgPgAZfv4pAGb143n2fdqD+D4JaVd0CsHXc+eqbOyIcG4IvWN
T1TT+seOK6X/EnzXMUN/WYG/xs2YuWA6TYMN787EJtrmtVKkYN+zFu5aTk95IXuqtnnjF2E6y9iu
g3chbfaWP3uqug5pjrtUSf1qzMr9PK03cQ2mDC55D4+c1X8oxZsuJ+3mOV8aX0oxyp+q2vB/dOmb
tNT0xBG/lqrmpE0jmnM6a1s0vyZmjMFCH3XnWu9bRE+FhNKxsi0K+h7IBWCuhApgMBgHsVLuLUHq
o6QROoUQ0Idv0EXR/YC7J0IwrHPCyFm3+V28h9LdK9E3+uTMHEkWuWBT6wmT1ZZaiEWj+SIESuGS
3RNXxKmFD8Djj2Sk2L9kAb9xMZZ/67//woxi1A5T7uqF+CW7675VswMJ0BQ1pQxFNuOKCNzyTz/i
xAWPrqkwzdgdQna7IQ74qm+kDwSau+h++4kLEL6pv+EQ+7dSjQBSY2/ckCNcPtgQvAAGeQwbWQ+9
f1tCWshlX0Aepo6ZRXjMxU1mlMDsreT2nY0htwy2KHs2Unl066IKMmrtKwuQIcy0wl7wMSZjSMc1
Xlwuq4E1VW/Qx7Bncjj2vdRJ8xVLTHORZ1C+aIhHexqFY+81DeuDVjZG4KYvrdKq6m4FRVCPUzKQ
h7SMOPG5seOS0dKAB/GVGA/P2cSnAuU93Xb9qc2e9geq/C2Ohyl/Qy7srWhRvgFW9KTibQzvyLTL
7XLyHd87H+4raJsZSrzSAGIvM5Jyrdgl5+8B4cXmDLbxGQtaGG93EXADAf+82u+rFtOjsyRSw3cp
KvV+GeNvkR+lgqqymaeHJLn+mI9BV6LPTCLOaafar8aNBu+RVrS/vpETvHKJeBqDc1qhiYVhwUN2
pdS8vCC4k9uurbT8S55Pe0JiWj1uBZuVe2ydofXOv7qtH97Oft0j6AktXa9yQpIspSXLZrGbLPLQ
R/LCTo34HfnsegETFgZqdyv5lo61sNaF/qgAe162cReYCqK/ut9/jsymWCS4vy9GVzbfvayqMh+3
MyunZCxs/xptNBmIVGzhxen/9zNssXMwu2aoF0PJv9FvnS+DhCebtFZSPQ0oMmGUwrAVHAAVV37y
E64b2jS2REk3LR+9h2TRQeLYcnU/Q8kmmsdYcc7ucIzyuZqqwxZLxbWQjGYEbCltxdcKfiEKS+Gi
C61ie+N6J/ziFo0nOJ9FyYJqHYOcxauQT2qGfGe4qamB6M8OVK4ZhB2QNofBje7Csi4AIr9KHX3a
LQC517XhcCMTp/cUMGueydbgYYebmgqJXhw34d5POJujlzH0Tcw/OpirFjEYO1h23ygfMTG+cP1g
a0T1BdcTimWpW1NyuSOpbz5TdByapPyB6lRJ1VRtKvQ8Cl7n3bXH3a2Ssu6AUsTWLWO10Ht83DI4
20/ifDQnEg8iq6ylDRBKDxa+m2ni8UK0AE0+ve3X5iVNi952aYx8a83WBmbVsPvXkk0Fb4F6h2XZ
94zzVZlHYEeWwAlz5Gmpq7cFO1dRY8Vm1igd0b42WUesv3bJYoqxJVYl9ZjZWemT73I7qpDqHMTR
FG07wK+F4gwujng/YoGpjOcifV2ztJvfxxRT7XZBH1e9J9zBXrNCFHC2InYviVScKd3vxVzUIAKr
FZhEtRFogJJ3rtaPIGm+DgyD5bkAYlTRh90h755+XiiZqjx2w3d0Z0iBM+Vh2l4K8wAfKf8G67iV
p5cYYY/0K9HN8jGRO9FvPJSxS2Sf47AZwe9WRbi3WLWuA90OzKtBbeK/hp4S6OYJK+Pmq9+T7pUE
8UhH5ddZ/NELPCzVoxbh5HHcvjzKLTkS7Q6eoychpYcN18mfOX3+utyL/7ZLX/+JVg/sXi2ez7dB
3spD5lJCa4ErAew/wLR6OIeHr1bY8haaIsxGR4J+ZD79Hbr9sRi1EVY9vmrg2eanGNidiTxYPr5J
E0uJ6oOb/OZFppQ0/KED+/IySgkfssu1RLs7NFitr9bprYDa8NbT9Y1u9fUpB8BlJJ2PXPYIDhUD
+Jc1/kxN/q50VZQ2siY7HvQMmS/dxnGjW/lKhLCswYGjEUD2DrdoTlkjIYpC9MgH2Z3PYBNbhztl
9jnN+pwa7Al1Ey3MhMN5vu+VOOY+KnBHYgEzAxV+U1v6/qzX6MDn5+GuiL0tFfH3gQ2ZF1dJKr0N
Pgn/mNE4svvI+mSP676ilyMTx0sYBOqhSBXmshMRGerPHThLbtnc/A9oqinaRzS5gxgnNxbc3nkG
z3DcV1qTWS7MEeV8akn2HBpBlyl+cNrZ2kvxjhGjKvvlz+T7dI3vt/LFXlAQ1HYrx60/dE9/hISM
LBKemT8IFFs+ZlyZ5jeCL1vFjm5fY76GxpDW4iObI9E3V3EZf4g7NBFdPBat7zdg275fTl/WU0Qc
p6rhuo8NrYpjFnQ5Zqln8JxMI44staJV2Eaapq+1FbbQx5f/Sl21d1Oxz7jd/3YH05lPkZkan1sp
PsyuPHzuF7N9UJf2HkYdkrrLoacKlectQEnG/RYf3YZAWakJgbu9X0KDDYGSXaPuZQApRiB3Wxsw
xYDxLoLjB8I1UAUEF0qXc68+PffMxXM5cgmUUco5wA6vTTXAQ9maL/orpNNUXHqkRZsD2xgZm3ek
laQjGQcG5OyCnQnwTKo/sn7BQLB/iVzYoL2HbqVgIBZAO3VhQz4sCI2gxebFCRl4pZv5dt83By8F
EvhIgd4ZPYdg7J1JkV8K8hZxrjrwt8K6469lwxbrYFMA+RjPzVdQmfKNJY70+K46QVoCuiacA8ce
lgeibo7wYjLbd/jMsQWq7Y5Tes+8/GlgH0YoR5kccQDwS8PN4UkuUUENEuyLY7iu63C1On4UEq8D
DRX0fot+M/DeWOsTKoWq2lM0lrYABViTMapKjgrlhsPeuei3LB7+dzQTv/DJ5iMSTdG/7pjlf/qF
ZExdlDaZ0SdNkHDXBBA7wisyoAUSO6Bqx0I8jYWtLkqe8mWVezWvMcbVtrmgeTNXKsW87HROj/6k
Ms4VMW4DXDKWJamZt9jAo/h3fFMfYVso3rG4b552eF12rGaYZNsaoLjXCRNt2X/L3mLKpi9xUsdi
AYsDYwHmoRwtxx/KCL4Ta7aHHSKvv4OAO8ebVC0+tzwIT1b8pRZjqO5h8OvDWXOitnFKE7GREuMe
ut/o+9iArYoR8iaxOrTXnjPW0yG5+m54XB1WFBI0hHin7H+kiCtcN5/4KTL4jVsMwXieNuQbTnJn
SjyJkClfyMjAHFGG8WO2/+b0xTV+LVoNbuV0fC/m6Tf0/H71HeEOCKkhxUfMqz3y2ztuIuC1p4xM
gtQaCcfR4HlhbXZxSNTytx0/DcQHJmdBf9ao5QLpNMjwLNX0imiB0h1jKxHHdGIROP9iNMLZ7Uwo
2CcL9UzCn1onHyzLL5GUDvrwA+wIcdtHWF4mWQzARoIOXPGdU7MQnt4t3210TT/YAiUcJ5A+IxI0
DTCeZQLo9LYo2520xZQUnNNM9jSTVYpeFbRSdukzQL6pCZ0M4GWIiADN3cuRFRcdcGJNftDRBuR+
FuKsdEUdUxErHEGttFT+kj4geUPW6Dhx94lWyJbomkOWfYPNIAd7oI0yuZtl+CekxFM6LCBZRxNl
VnQTBrnhKJOijAYgw7kUnQih0lMYWtEjj+H2A1TMs2f8FD3tWmWWRgY6Hfuq5P0MWj5h7lYkUb5L
QruMfqyC/4BSNmS/JNpgO5ejxozlLlQWCDiRjRuuKPZffLgKxTVlTJifUDkqMWdMULrbWiwsXC8a
D7izjd9VESxLyNQ8ANt7L2g9Jj1lI7UV0XS8z1dimz9O6036YW/iULqMPJQQ0QsLOpbSC3JClxe1
j9ias05cHFDwIADnDzMtvwgl7iOjo7ukJZzohcfs+DPSlhMqOqFoYzvAMMYUQyPVQy3JFdbwhU78
MyXhzd8dKpzFcWWrax0VMLNLVKE3DDHdtktirZfT8TfxWU+86QYnhYZ9TJIdxrqrxn+cWgJ0vNi+
t35Z6zmf+jeP7pSTQBHnnYxmpSTLpcgKELzuLVB7qeT8mTdeQjUxP0DzXpSb2fi60upzN8dAATro
SYeVTXZG9p/n5lsZH6ol7WUbmrLf7FZ8V/rHeWjAYsumG47LERWsUyf+UqZmvEQeOnY7xHBw3ZiJ
42eY5+CP8RSXAGvMWDymvYKuyi9KWZNKzm2y887hySvWg1ddscztBXxjVmIlay5Xp+KO3a7NkbfH
XCOC2p6VFv/b5X/OI59og11vR0CF9xwNw05y4izcKJr/WS+MICiND/PfZoGwXzog2ujZj6J1aodA
+FR8yTul/H1F8GSM5FJv24i/zXsZNTzP5j69oUSL/WrNNFVPEoHmCL+pdc3Mr1UuW17acer4pSj+
BN/2YY/vLDODYfHGoKB41iwS6x4nwd4xKbg4UCXxA1CdA1gajTZURlaMZxpffJRU49CCNIg/CXpJ
gTnmSN+gD6dFWvcc5mzPc+4HAb5dv1LjPOJ1hm8i3pJSoHj3IUJaEJn7Ca577BBhmsZWasTJKK8j
sbqg7XIVpZkUXNWfoHtDNDpPvLI3KkuQhEdtfagKbnqJuOthOWDGmAu5fgbQPbsH76CRn4q0fk0G
eMakXoBaatTo4R7DJnfXUvX+KJJWraMT1eN5lUxlxNmNZJeyIll0nSPBeVwIXpUz/rC/VC+oZSS6
dIV+YKyPzhS/Gf371fMYyYbHJU8jQLkXFTRKWR898+jhEEuHz2KdankHcZdPDXRGHf6c7HXZRrOt
VR1cXmGthnXFpr6EEarissYf+j/GHJqB1OQyG2DsJ0KN1moVeAeF/EtSVoR1NLMix7aIur7BkDkM
2SIilbN3b9il7DjA+TggsZhkLN5SEAxGvvXOHQCGU85yjmIib/5hB7yNPSzi1oCRWO0qRQQ/nAJA
N2Qy9v1uImYLtQg7A1aH4f8u/SNQYNv3R5KENBR/rm5jdn/5V5maau87ei3Z8al1pE6BcEeGXNiT
l/6m2JyGCJmmJz+U6WEOs1XOQ7Miq72+2P2eXYx58Un6jKssxoB8wNihecGEGUjU8wM3ehD1Ivka
G6Jmvek5Jm6BiotZTDkP7y5jyI6YwFALRHk1jwklVmUYA1hnyqBpCAF7Ga3Wr5/Ho+Wdgjoks7Vh
T5Ie2AG96+3zOBJIVMFKedseIgDjgbbrUoJyKGzdIEdNM7F6NaHegSYea5/kleFXs4P4IbSJ+w5+
lLivSh0w5GwQecvOVlBT6ZOMthU5ujzZ1uRFFBNCBLiMvgZdvWXKtKJfUwM418vody7scxoUOMbO
u/5Fjp6Ui+FlFsuCqBED53I47PNDjRTV1qUgfvUDKi01AtkRoKxATWgEX0Db+8UvzL/mhSxgSZlm
D//EKhr6ZR2Sx0U+icq3X2pep8hrrOz1GiUCuJ+a+Ub+xQF5C1VhaAcgXMO54/EshFaIGVK2wKWG
55SFwMB3MX1OfJCVm8Vyh8kNIVnwcsa71/FCb/o9cNoVCsul3VsA0/jB2ftsUldEeAnBFBhLyqcT
/HiKFdALzEh6Yb2Ntep+FGt67ScXoVhXNMeBTOt8XskznX6Znsqd+ZTB8CkMVE/cMoxwHA0QE8rX
WNt8ywEzNne8z+VbPVRZ6etuGvChrrpRECnS9WkSzbdAihuzTzcnXfGnBEv0SLN0WKMEG45PPBFS
oXUEZ1u8xcoNdK/yRe0P1/5zss3nPi26IVKEIX3pyXCGB1seEHg1MEdQt26k8Z2WC/AeTzSAE2q8
wIPTjUjBhzTVu5HtYp4daF/JyVGhGSydifzOcaf+xMeW/YySQ7rw1muod+SPQn3qhLOzea10ptJN
E0enc6W7XH5IeqvcGSFEQQLMj7x9RHwAYaATkAvnRa2wego9TqfSvkPX5vwaXAWvhDlCg0nYFXUA
NXZqtw5len562AuwSLD763AmaR0xNoZ5Jl1YfYAmKPq1ofObEwlvfjofsu08W2y6qLK9avsTB0Jm
5Gul0SsTBk1NsXtVIxGkAfqHAAs5fsBbXHjs4Heby3cD0u6OTBCZ+9mZ0nn7fq1brl7tmoATsODU
8UokhHP9HcQ50ay35a/ovYajthAx/NII7yb1vF0kub4WnkhaEAwWZdwvm4GzT5qtuOcQKmgrzRzQ
asDPjnwL8KRAihp3fho5Ogiy+xZY5hmw48VsPobTClUaat9hqadxdIbVN0w5LNvoIghyZmgMA+d7
NBXhTE6lImTgzOyQeXMXGYREw7+uTz3lRfWSHA/VRTex8eFR6UmZKFRM1qZItpoZb4zYaF8fdp+7
MfcXg5mCCwZ7RNI1dkn6/xMiUfsLCkbiMST/XJ2Z5LPEtoZF0QolhijwKKoqosqC8TgokmH1oWOq
mxWjKX62tX3H+xa7hmPdw3teoatw1ibk8mhGV4z0SdGi5apjlkJGKW1DHhUCjpLt4teUHWDhQk9/
RGZvkJa3twdse4x4AiErPAvNcB4N2ja+rnMxMiK0feesYtocBhH6ej5AVcPqi0HFVknj9QVZZHud
iFG5occ02jTFNR5MRk2nmnvLcWIheTjzTupJkY2+Si0uLmulw1y3m/jOiJlfoc331s48xDVRvxXs
9xRjQpEIkBOM5ZzhtBmbPEH68YJXdPPWowfZ/EHk4kC3r2vB9ylxXZ1xi6JXn1CjfKO8okuiikph
iBDfZpwC0b9MVXMXWRoL8v2948RqXNJOGLO9cHCtmKKeEahWuODMF3CngRsIBBZWKP1sLeDppisc
lK/dZaAo3MXBnHjG+hnu81b2MbFQGsaU4abiEg7V5XtERpehTQq2icptpf1CKnUZh1mGB7qBFemi
5F8zIBwH5l1Ves43OLof0CbeWzD95rlbb+j9TJ7bdNQZlJbYgcbsh1sAU1JgmsAqbSYeiVTWC1hZ
Xbvig9qMFES0bGd6NfqkJHFKtm5hesj/T0mKrGg3iotHdHzbCpmlUfiCLzEh3azfYOb8AYd+rEl1
2851d0R3n9QquWWSKaeo3Y2d5g+Qjsy7l/3dX0dKGxNqgollMA4oCh9u1M75HrwH2vvEdG1yO3St
czC+8ZWMWf6fEN8CK6qRsqH9GPbvvgbDDlSvODpQ0BnrekeP13qsO4pTb5jdJO/3RxiukpGFERQp
RMaocm2UQNmC2HKsOchHG6KwTXbrayWCsNi8myeBtWdj+T3fI4c025gDEgS7qFoxLJ5JDQ3Cck1Q
byqG3cl9lQOksTjNwK0WbPeZ4JB9CVI7CpTaPDoXtziEGP/AJ7nOEGlMz/BF379qcBOy2JW+xula
cmsYseg2Vc9vVpy6o48Y1swKVbOIkb9l1UMmSwVmC035KCGmiRw7/QaSVjTV7LG4dZ+Xe4ASbLWb
aQlJgMTglKzNHCbOuBHZc48mBv8yDxPYNSkoCw0gWdY9HJ0gHCi/YmhjQ8h7KZxqiRDW9oepeYbu
uZsyYJikLSaxPwJZdW+4Y66Wvzs1zUnqfiYfb0w9TZcxXSXX6MCiSlZG0GQQIdaZKrTdXGUE5uk1
yTFlCuVRidufVlZHiEkbqjLis9jbVFs6ZNiHxGdrIJpCw8iinKrq8nnrk3mCPNkqODnmtMa56uRA
EKTE7MOuxkydzwPwK2x+jtdnN20LCqbGx3BoyPDtMzt+/w0z8p+GsFS8A8AsCYyQPECL+5FqJoVs
zj3snv2zjarSDOD3a6mu8N6F52LnYgzUaGovxCW5xDJWZz9DLsdeppbsiIfnRrRbNDtssFyzwY3L
Eviygfho539mhzuAMk8FljNQ/OLLLJwvKLAZvLhVtNTpw2KU+R8LdvIu5sIVFt4R3xiR3Y1crZVi
6Q0u04Ta5i+jMqPrWIFFmSzlPuVtfvQUyDpFdVMsmhpKurKsQfWyCOJeIj1LSNIAFKs5K3DRkfqP
RBZCp7Ov4K7MnBDLpEeZJ+grcefvHCvd4WzINLjEPmoKaayzAfrDxKGe2cOqqRTBz7tnlpqnVoZp
4+BECzZBnKwLgaXH5qp9DWZw6gnFTmJ6bwxdhzKShBrDcxCtTT4HMsj0aeBAvRtXENDlOXsllFte
CkRjGelvvfLzucHceWpfF9nSbgRqHSFs2u2NRXIB8IW1uF7/mhg3eWvlOhGG79mGR11yTlYagi8Y
WKZ/siLCtLEgYoHDtKA+ReP7uFMGkbaWO7MOJZJjB0geLpKj/nnsvUpfU4+tPSEN9STjxK1lkhMW
Ao/xpP36a2R3R6tq+i0vPerJZrlAdT80z1hImcajska/DwNC6iVIP25bpz31xx0KwRTya0yI9X0W
YSl5Q44Y0GavmVAWDH8EB2nV57C0nVgXj/23uINL4LQTVyDULFQQynKIOp4h60ozmIivIxbXXRHh
JUB6LNLUnQERS73CP+QzGwC/ZeJgFjJjnW3quq9vv9Q6soEec9V9ccF21sYkr/Lkm7GoDj5M7j53
xw2TJ/7U9FM1zJiX7coGJjPXNuPbrKWws6e6iqCoLDJnoPnOdPiH34J/DleTYwqovIGFJpE8ORIr
/wba/xqjdGsqIfn/ylCuu54qNjfDLb+Cp4boJtWwb3wrHn935mDATid7IWqagyasErkTQMwUWbB5
ngGJ9WMtnRWzfViUU+be2XtKV1/V0DqJ2mL7FbyLpqpQVH26HrXsK9iszQjQuXQSbjqELmjdbDAq
NKValrmaqLqSIA0yTwOd/iOTqTp7h4bPS97Q9pb4hEprOc5Jlv9U4rlOm3Amc5TBjm6isynhdc0z
MqdgRgXY1Tjs1yIH2vCoeBrC9Jot99ndAmMwVOCefyEpcBkQ7EmCiPqVUArQgM53G+IY/Pp+vx2r
xS7yhS33U+rBH28GCyveO3A0Pa4V7WE8CwWdO0luTH9J+Ha+yxlIMsa+X7vm77EZZyPy9B9cTcgS
zXl+nvIDGhv2tmPQkQpDGyTfFa2sgHUMHogND9dJKGrPLGy+4WuMzb4Om2pYYuTcBlkXh61tvSeK
gktnEhTW63vzXzEgfjP2pNCAYbCg0AwT69GlOGQ6JInTakU8cITmw5dkdOqLc1N23Lhakc21XCuw
BQYsM7Z9j2Zc4cmWye332K73BywaT3GHJ9jM5bW1Xc4ZnzqhqbYVYJWLiw9PuRxsnpM1yfCEFSUF
0bojiX0w6n4tKDt9i0E/0S3U4hmAncRP18leS8+sE93zkbnX7fMqv2ICss2WeKNNPSYev7W0HMPz
YxTC8W5WZ2JHc5B1sKwpwLD0Vlmjxo6Jt2AX3qGUCukAQB4UXHLj3ea2XmsaSiHoz3B6RxsgneKE
hYgQ3rCGzhqhsluNQjUs9ONyZcK6S89eYLWyWjI+OwqhX7T8iA0RPpVb3r/ANfnJmltBzMpVACJe
bAVk260pK1KI3pgr9WMy8HJehN2op+1uB6mBtgxOQRtp22HjIZ7lnop3LJdmjG1NOJjF2E+KP4Rr
DikoGD4qQOEEMZBr1df3peD6pkQUqyM4imFCSov+CDqIpMeDylLuKOBL//Il448P4a60qoDMAaPH
PvvcP4hEr0EVYYnl4Mr/K15AcM0EdzKFAwoOSK7YW1kpI6r1fUN4seen9AyVkUMZo8cMp/QixGe3
EJprT3q4CcAAPufiE5JlJ5l4twjFpeib198XRZZCwWkyiKfC00Hzez9Jd3GCSuyRM10xF0HaH2nW
k7BCZtYhHS4DV2iafLxruUSmLxsl5jsBuFDxr4/sBtpbHJYGdOGqXpw3S6bw0VT7nLNoyw1CSL+o
/KtLgt8dDHizUiSYdoxQLXpSwdDwEnfRqzzp7WsJgeNXDq7zHlxM1zpAx0J4sIU+tWydolEGyVRu
HbPfjDE0Pl2xObuagVWjThK4s/vDNrLS+LVIsRB+vvlwhAl8Exmf/CQCB00goL9qy9sTfM8H99Zy
UwGo9mepCUosW5I24rs+h2iEzvotjlxf0055nrY/oi43aYvrnHsN01HuZ/7QcH35Ih/jzfQFN3Mi
U2CXD6JiqbYbkXnB0Vs3zl+Zre3Je+t8Gylo2t8EsB89ZnA1UXcyQZuEjKbcuXV1HS3xl28+de7z
/+V+FYeHI8DOP3cN+Rx0eYYytOdvDYYnvg9y6zidzMWFgeoQrnlJwWIsjPSIvN31TJwHV5JaH/QX
1PnZOh8+Qs6zaNIXwNnwxgAYOG0J6rKzw6Ui9JRUdxjJec4pwFhu6e2VuPKtaFusgtI4OIW/5CLS
HCOi4w610TnIZD00exRgY3XudxARaXUQf0er6WMjtQv9moTVwmGUllo9WuS8QQhrJGfTqqZXR8h4
VkxP5SWJ280QMofucHwNK5peZdhx9rWS6KMLzHG32/OK9rUUA04fIdp96gB6iLzcEKXb6xCCGVCu
Du79nrygFmUT/R+oIuQ46Vyo/Vd9MvYnat3jSxU1iGkQg/cmpvfdezCtcmSsdsWzwm6mkJFGw595
6yL3Jsjz7ui1qFgpL9y7ArQpK+YXTB1xGhbKuTO5YMcYmZbTDNQzU0k3PdVZSECrCe1NnIMzVdFP
liRtj88uqILaKgfJ2YgN//TuJnp0GPCERQ8ib1CTNOVcaYk9WwMtXKrXMF5QTCPJQ9uKc+j8Tq6v
aaumWTJ7Z92b12PQ7pflF9ivV2bsJsUbq2FBQOT/kn4XcqBBy+yiMFmYnKF2efXsiMutenbGVHiA
jOS9nyaqOTXEOUBshpnyiACP1IbsMr5ULa1CplZRy2ROGGLzF2Kr7TMApge/cdnU74ctre4gp6e1
Gtq5Ocp5zQlIvqYDGWNQbMrg1NuzVY/cXOvnfjG4Zf1deSbb3Dhb734JvTfSs4CibW6EC3MZOs6d
A+xZfUEqmmV2aN7kcPyxWPIcSFD9S19dZZIn21/3YWp2ZXtAiHh5O7rqIS7m+Q+CNQXlmOqCXVqI
SSbfNRh4uR9cDXELKeIAx5iDfDXzSsL5QY8QYmw2Z4PverAZXCwQo1zRn4uBjZFs5kHRHeKlSrhM
qLxv0RDES4Zn4DWq1zXKiv7hY3SKPs8+chfc/Ok6EGTrUIKxS/lKySUtfZkczsXNrYuPtlM0/K/b
eipnoya8UChmHxFKZgAodf33HOSNb+hXeIdEji64ubaavW0OsfhE6RgdqchzfhPw8RD4r5TxIQiV
0pvWmVatAHmFjL2nxHgMP5jTzKln5+HtuoNsfW546s7sboDuWH3vg5T9tVCUaLW4Ymj1CNBgG4LM
Tu/ZSe5f56TxO4OkoQptOg1A6+6IKmdnbvB7bhRbsIFb29wQQ0lzvhBdOAuL0jLwxJjJqqfwXde/
QFpAjnniZfJ1EOq1hglmHqtypQuFeGwFub6wo+uQCAmRcEtO1gmpJwJ4C9EWZoGBNftclYrPKEUt
HU/GTW3i2HNnHMRO+D1U5pYeGmP5+/Ef0X1D4Te+0lrZImx9eKLBqiDNzmrLSdzevUUvxNq/ryPh
4hqCNtwxF1rFv+W4et/R2+jrIeMZmMFlzgZC1Bsx6eSd+SbROe29K13MP+hK8maumQa48X/znnQ4
lExjGVyaAQ7bGugo8IC/srA7mAjMR4RyCLC52nbdFGg3uHDaIAGLGn6uM21F4YpRYM705BwgkMyn
LYcA9174LGpGUaNqeQl6Azs7JUIrN9a7SOskfZzLUU97V+3+sUhBKN2ZzoIOAciBel+9ywNaUPmX
MtNFjulH/txZ6NbYzMS2LgX9vPgWW2W1nyRm6+dFwy+s7B4uNrVn6OCTePn5ZVM4+yrDIPdNRvk8
oDLUIOxTbeCiz/OJYRs1LunfVqjsf9wxye9AvpY6GZBb4havdwe0omuqnFCClAw5sgthF4zJd1oJ
dEUJxmG5mnXFXJzqrJhaDLViXfwSohpoWyNlpxoxwXidpbnskO5e0DV5aenDI5g5YITHqdUkShG/
GPON39AhCKXZOQI8RZv0tSo4kfw6lVJw7PhHB3ZsKb1cGDszrrIwFBwtGV+9xlTGtVJkM7NRhKtO
RbNOUxIbg+D5SXBJk6MhIeEI1Zg1cIlW9CZTIkwPcjpfD3hH/H+whzvvoK6VCU7iWA/4cdEzRMM9
hOvvdgy7x8wj0MSZsjk12vYyS52NRaYjmG9/igtG5KwcPmL82Nvdy9UFj428IwxgMAo8UvHh1l41
6YoMNkKDMyXzTEEZIiWfAWrwm4hfSQT7BmnLxKr9ilZpsNJ5jYnxmDWiJSUatCJ7BZim8ZJVPBS0
j08DFCH/oB9GMwKKLzsZ8FWkBum3nN48j/WTlgzRtDVOClFKauOYBribaJ5+QSC4LuCCd+bjWpe1
+kxI2rPnutb6FQe1pF8XdlfMLNgzd1u3mnSwyb24GmpEqD0Unj1yHyNN2/55rXYeysGb3ReXTfxj
CDcIBcU3CIb4UsAcHIWXj9Ga6F5gkWnLKZ57SeUnP7MTJgxBlPcbFfy6Q3J2zib7umsyamRfZElB
ZsatqzLAJSPDRjRj5Ok6pimxaXHvdoRRR6Xnyqv4ZyYDpucXJCAnFc4FkENFqQZchbZJQKj1z2ep
0xx7gCaNUgpsGTeYAkKBwGzOwUs4fqpC+PA7mWUkFn2DgBHMrLpRDr6FKTs08KPd/97GR42hjbiH
vjfT4fZgHjx8BKQGFrnM2/KzeBvEm49x901wt7YhmN8MOGJS/YebN+hafhHYo5qC45T+dzK38mUU
Ja+H3/CT/Oq9pAajJRTY5pXCZhCW6p/FWyqojK4ktRm7ySji42K1m3Tiyg5K8dX2MhVlkVIqXZEw
BCy1ETcdDwLs5+WAH4bWBonV1+OCVPc1Fn/R02Vq7BPy29FgdB6pmjXQiS14KXof3ZemAmLO2w5D
6pCu2pWgubx0p7zfNXT37KDykH2HwKdI2Fb7aH/JDYmxGmxStQJzJ/o/snz2bZR/yve6xYGAlc5t
DPsicuY9BydREK4wA1UYY4COopeqgoS9X3qZQSjj49DhD7Sxm1lxEZ6eTXRB5Znc9qGAcL1yhO49
B1GrZ+Vi0EMyJOaQzeR/a9qH1EAdVg4pMJXwi1YULwBD7BKNO+5qq1b5KKGu8el2f0ed76ydrX46
Gzy8TiEj4dfq+rol7+cVCIheQNr6nbLuOvGvCEcLbPZehElkIZ/pI/kTqEvY8GS87/T1PWkIdnJQ
jo5u9DiI8Pi+5pyJnUHbGD89y5Ik+LqkTPFOexVcKbkB70PRgXVHSUiqT5C9G0YYyFTgw3AjA9Qk
IgxnNkdVY0uucipHrJ7xh4YeSYwSWsWbPhlMCCwU3OtC9quxSskN1bmGW1u5qdk1x7kzE6Rn9Dy9
9FSXtww6ob8y6dqrEPx3n2fii3+69FppRs3QzrC8439fbcf1c029N/Bk9n0ivzDzTFwHJrGY0kLT
oq/SXs8dqif1kj0oeJb33/5IIAtDjqBCqftHaXj9SU85tT6u4tEIDCuKqmRmyUaTeAY2nz18FDV4
35wUz9A7u4Izh3K13FcINNsufqEGvpSAApXmIIPCuAEyyzMMJ8M0A0/oR0iMOhP9FyNFwQWtQ292
i7K5fjfrm4VYrCf8szu/fX95c9GG8qPHjzPhzViwoPRJELzI/PVM0jE1wg9E4WcQlHmyuFIpLONi
ZTkpFv6vybuOHLlkiFYcwkvKUDJ+YciInyziXQM3YDgPo/kTYIUEocYVbn/fbhOjbVZ8sjT0pF3+
bhaPHfFNdDaGqorUoxo1prODADQptOAPHmMzKeS5A9NYY1tDFvPtCs73mdDCC5MW3snbbuv0yogs
wxcU2EX7pBIUG1bCKrGONTrowyOyKvW8FUkq2bzc5M7+vIHU40YJ8O+wvOpIiTSfGA28ESamRCHl
lA6okcBcUFN8yMpO/Oz/S7VQ+6CXj+siSuwdy8OfBOdrxCdLbPP8HrHf8+Nz+5yeIdDVcrHC0KlI
o4zSSGf6Xk31/QRDDaAOZ02ZSN6vyaQmbl6ituHY/F5FySA8nyKrocTy8KMuBPt8v0Xr/u7wxF4b
Y+kcBqW05Mpoz8GXgsdYRJdwi9+GBzioHGL/mKvUvg4GJfWVYpnn5gekrviuZD6YEy7EFcPwV6pk
YMNdMcpMb8xfbFnIlDuqn5c+WeSYd2yfWOBfPZiqtakw244cQNMgGzjqfB+V52Z146EM7MwM/g1w
6hJjQPfgVlGRE/EG4mp8/OG9t8IiYUZlWE2KjOTYkYA8Z1Xa9TcScmhGTTZD60ov4N2H6sQWNQrI
Rib99ZQXzA8dtLJ8t7El11mQmjs5ZEQ6eW4MYttPclFELSn4Zpk8p/GuyaWlzOsYoO7exvPuXAhW
Lb4FATrfsAM8J/nRMnwFGjC7A2H+ah5D1EhhvjkyCbw3OdoOYFZHOiqY4AludFUeccncaKzXaReJ
vN0+VwokWepvdpxa5I4326oW5GsMF73B6giRkmnLkmszo3ggxgiRgDt29kMNbzPy+DYQa2bGATgF
VvJABqzcJy1CyOAf5r+Asg1WSrABRJ5wqMGnVgRlJk8i+jDGuD5KOL9BkkS5Hh8wRLoH0YOgI6mM
eCZV+FmSJ88FbecoWnNP+3PHyJiBvwul5mXAyAqbj2aKqG3CGAnb4D2LuF3vDj29DAjGcA3tMbzQ
qib9H0rsFhE8hMpN3nbN7l9gW4rf9WH1DAjBudzfH1kUQBisaa8I1dY2sUBqEtePOG1CmEzftst1
HqC4wlXWF7PfDMmkhPSFU7WkMiN1Nzqc8WBrU0BTh3QCmXJvaZO17vBgdVnPGJp5F8C6FfAb9SmG
BzEQN7l41kMl7iepHK/B0qQM0C29/zWOja8XmJjdZSl19z0VfqXPoFVq08Hje515HBjRq6FKRDmI
FZAq16loGJee2/2TXljNNxTgAAENN83+O0rnVoqyEbs/gb/JnkC0JafyN/Yc9sGT+a4+uZr8j08D
VZ9DxyaOD6B7LOfjS7q4YtRL7UjjbyBuni6LjOWoyJUmw0uLibvhosKqtFczAekQ7+Kx5DFjOaqA
OiNg9jW0bUZwz93Lxi6QMNKxmxJ9o1hJ7asCFVWV5xPYlOJ0j0WSIQdKZLvoqzQjrjYzUFudFXkj
Vo7vj5Tajz3b3+m733vs3oMVSZmc5pJmZMpbSrwOQZBqiszaO2p99C+ZRRrmb/lMIko00UeifHGI
01/SwbEPah5AdfkHWqwdzTF9dTaDLAlQrHdQc2JhQIZgn/4swN5EKDhfslWcKgI8+ym5laiNomHx
bG62DGp/TMNnbxNpOvV6TfPqKDYUBa7K0+Ffrv/kRpZPLlBXDkBQUSUKi9HkvU+95uRKY6Su2jCw
SbruJqkSbo4k59ObE9qX+w7Zre5wTu8xQj0zsw4bUfI+Ij7DCl1TUC1tlLAIWVX8HXM1knmqU/XM
q5M3at0O137KWwr3q8Gf5pd1wyBcfYEInaA0bKv5jb04BsZ4ZMytTE5Rk4oNHe7YLdptMbDyd4Ic
xvlvq9xUZ7E9z7YGOE7TGsyGc/uHnxhGn6SjLxP0+tt/kEx2iAS0W9B2ThguDNH+jl16wo54P6GI
QixyGlChWoaW4OMsFet+72cJBIA/3rC5Tv9YR2ybBlaDau4lY2nWbqk6Zli2iwuYDrzbnRmRQdf3
XKRWaC7jwc23dP0jhlmx2rBpsjVCYy9BozZg+o3wedYu0MwflRd2Vrepn0Q5jIQfWrzjqyyMxvU/
d9gWjEUL65JrHaglbsgQuREMyb8GehflGUrpWB1RbK30+c4o3KQ/eGZEp83wS/y8YdohWYZo1XMu
pmP6p7BZpWp20VYtk1086g7mGoJHv2BCZs94RZRRW1RCrEGaB+uiUekoOMjAYtq2J+cfhAPqKBjT
+2QLmgOs2xQKDQCcmrzotMsxzR0M2vp8VrbF7rBxs0s/fHflGvjO3DT7sUF5z2GcQUL76LgIt4jR
n4xeI4oOGkZtKsLKTRR8QJM4/26GfArpm6VxKpwViQZDIDRvZHaUsCy+vjYrNpMSSySqdP5p1dwZ
2l3OnGQX7NaATJifVpmGWIyMPT9y5GjCBgqXYwjoxtqzAUtDjHt/2GJCbgZhuOgkFTSHMvDu5ilp
1CY01E4U7+u6QyMbRGOUoraEwKC08QupSSQxv6+QO/8IopaUrst4tSu7w005BRDeR88ZiqKya7iZ
Hgzsu6/SimbFokGBdSHzoxXg9C5PKP7cJiZ7/7taLz0yhhWrLPCJOORMn2lbrqmCXWjnftFgSGai
Bbc+x9x/iN6qvLgVSSqq62soPQTZoMDz2u4LBt9zudv4b4i76Kki+E8DNEVnXclTPyLeXCa8k/pf
NunJ8KpBF3iUGEzz2wEG7kwLGJcysqIlqvafL4CxeTGc33HLHj5eSIW9RwdsJtD5kKjf9WUhkmJm
Ikp9/MD0bLgLKIDK8mhP71bPMLx6CnbxWLKxKm9Wav13eQJssLI9PQnGGf4qYQr8R3em9pWkXvh9
hicxCAonHdYWy6laB1blVfiQGIF24g8crndtIuAKRRnMXEPBdjHwNFwLeqvxMYmZyAbnNljdkXa1
vUK34fZp+/S+VwYFQ3VYX8/aag20wrRDeScUkf6hGy5Xw1H6DZuxseis36ur3nCjqBNbpBVDtHkX
AKx3/kpxaThn5wycg42SLfxaHddEnBHTFcNF6Pf/0HV08l/hxHuki1Q6dG6+WBvwNdbGkuDsvjye
WPBWDUcYgqZQUEbTOLNzqCr30HBIDmz6HYiDS2LJp5PCUyuUiYP+jfAlp5D8J8EFxW1ZrlpdzZpI
b5ejGL2a03bNcg9+AjvbgudcgWF2xTt66UU7LbdoHReftHAkwFcYv3/usk2JgRtiG6kFCCL4ajki
M1vsdso2z8eGPGu0udtyz9QoSDPqf6DCS8Aq3v/j3WsfSnkaGQifN6xUJEJA4Aiw6BpZ3CUBGCEn
AC3wbajlcQlDOiaqzT+BF36NUKMpzQsUH+JTuwbB4flBja9ZvHzIRCcx3MzdneRuoCA+Qpe/T2iV
OsiV3Znqz0jIDLRyHBUqURqyrVA077caj3YAgEErEms9jDvBiYQ6pF/qy9//yEJ+44CRx7OctiZu
Lk1kFDg3TqjzbrYVearVCg9XTiaIUb7xL37xf8ERrhRggIQTJWGQAN5Z+rHW8dxVWjh85RtVH81F
vo004NJt0K3Zjj5E1OBgqWeOW6SM9Qpsrxhe0+c8phMaeaUKl6D4SnRcD4oNK2hZO7gWgzHq+vtT
BIb5aWH+18JJmwplBcDPcgb19gqQpvN3lpG5Qr6VoXwWYRFK8g2o5GapxaYcgs5s1ZcCcjTxqIPX
8v2TUix0HYbKkZX+nPe9BsbMVq4yCHTJgK74b/Z20lO79TN+nIFbd7/W0dFpTyRDeYgimwLMC2ao
7SS1IYOimXQbn9uoMBatsiK7bBE2VTIK0GasR4UQ6eahG8h7bifoDqWutnU3gEr8uBI5TIMcwbio
UjtoWqFM0IiGlsiAKGyikIWCl4xON3TzwKC6B0O64LDIwNEOvMjHhvMZy9I8njwPKidoqISBQ/0d
2AIp2GvHkVHUiNNEBmUxIbmiBllhiVWXP/KTi6UIo5Ai799qST5g17GP7CZDaO05K53hykV/KD21
YGWrklncgSLqCiWfBhCKFjrlDmBVhLRE94RdisGFMGWkuSH3po4K3Gg/CheKZ3I4DZkVOt6bK+40
KNEz0ZkgLaXqWXxo5gDFiIC7vioLBoKZE97/kc/DOW7TjXinEsQPP00cJiST6XXCASCmGph1ppw4
hL+jvFIeqHOdfkgWEjLZzPOyO25eVMfUgo+zARhAQVGzSdvPwYdeEURRrYUAzfZ+uFn2A71I6+Vc
TfzPbRSsqNyJA1G3Q1gAtVwOffWglXroWskOQ5uYODIqUXchdF6v2vgxwNSHs4yjcGzUW4IhofXc
4RHYtWwjhJSQTz6ovSan/zPsbjrAeOS/85VfUrIrJM9Z+8IdV4MAGFqLBjFMnZh/TNPWC8XO6fJ9
e1pV2lB2aWRXTSj1n9PqbhzaZBt0RZ2Q+7IPMQjnMvDDdXMFKoTX86IlQRNr6n4Ib2Csp5jQf2nz
AtP5ZnN6Ek+XPj4oTSVKcoM0Ag7x2nr0KVsh1qoLje6Or42xXpS4Q+RV8ELJFrP4v5bCX/uNL+2u
RWAbPs9ZB1Ct/etKNjbS3eaxPPZrVWCLwuhq/Pc+cQV7H2atkL3Kj6kXOasMM5gYpAhYMFHgnfWM
0WG9RdUCA98PAIpw3NnDhHvWVCnrZruAzIE3I7zMWBBnNAyCVyYIA/5YfRmfNg9h9a9+lhlVI1lO
MdnMXSYpDhm5kqeH8UQXcovQ4FwWZpGEYfv8WOFCyPiaQ4KO68pixlKvMQA/v8zUAj4nz6H7Y4T4
5qXDZ8tNGcNL/D5ia0y/OouhhldglrbX+qdA0d7j8nD/54hNxt4xT8qpCeY0lLkRYnGhDRcZQSaQ
Dr71Dma/K60/wko3c6YbfiUz1EBAVOv+CTV4/CJXnI2VcrumwlarAsuFDSe5q8B/YtMMFygVaxbj
RJ09Y9S5BZSnjCO4+1PFpHv99V0XTDOUGCanUbXfqr3QLAHrKKTaXjOPS7TvUebOGKcb744a5Y2e
OmEkPtDmZHlOyXNAtxdM9wSKLhO1hftel8RG/i/ORRz12dzqxj54e/p/OF4yOgLtMyj8MaF89G8Q
i91LieUL9k/wXlL5OFHrvFavqbqt5Q7mJz+QzlQrRYnO4aLP/h6ge2kWt7tlGOFxGhtstMeCyRo6
sIj2nPBSszqb6By43TcoLWU68F31lqrawEBWV4/nShWUfSApzaD/36+FTgUfV4XNo6UbRJWZbL/C
8Cx3tGDFcGwN7kbMyb0sq9RJ+Bs7GxpwjrykMQaDOJokys4/LiGkFw4CRDD9bnfY0hJJIOhM8wrD
gUSyxdE2gEBE5MBxxSUDVtg6GXfRl8bmJJkMh8rXVzx9I95FZFlpSj+WVFXrmpoF3BNiw2BMFI4Z
v0ocEgpeRKw615BS+c9ULG5xbWhtc6Ain3RxDJDD9V9FSDKFle5zxXbVD/O3HEPO0nAYOZ0Dk8Kq
/eL4cMRkMoJKA1UZ4v0yN1cEVtf8+XEb/dP/guDfNQfKtJbxaqdUHsJLyQUhL7xdZtHDJD2VTtuL
14av4eyp6KtyRTtU2wR5kF2L4Ka/iokLy5h4/hMVUYZ9/zYqeeAdQGxzVFxSYJwGRD4eBn5qMNLN
6WjZQJogxnwrHs7KPHKnHcnyU3LGV8ZB0NxVH0SKenm9yhCqocoO1Wfet1TPANt9sg/n1KBbdt1v
3H9pG8wArXmHFIkvYaz0Dw3uVKOyxBF1ZRfQ1snvVqsdSR4vb4I0sWJzvMxM+jc0+nkgJew1Ck8v
W6yqC+XPvJvhNVHUVHzY/fyzaL31yTRHfr5BuLV43inPawwzU6CZhBp14nC6vMOEZBd/CA45LSDn
F2vuJUVcasFiaDwcTy9tnRiDbNUy/lgQRCFS4Oz7I5yPrxddVXH/+AbXMlbMiVZt/P24DCbTbUNR
qc3AbVLx3HVr1gXnRnINtrLiglKhLZh6gJRYi7MFTjPUm+2C1q4O7kNASlH615RdAyZPIanB9NVu
xmD4m5374pcgIPW2iJtQ/p3FjrlajSsw10WUxmcF4ne93TSRC8/xlbdGNZ7U1VL3g3FniZjT5TKP
q/HKX4VF5mAol+lBWrPa1zMjVriavG3r/40ks1dDLIG3yuPsX4/89Yj1M6pGvGV9FD2gDWeZh34A
a30ffNYvklzLFvibbHYO+E40hGNtPa7wQfq2tqCofjUfSwt/qNLzATTji97uvWcwY/Z8JJ9twLIq
J9ZcE5eExB4ZN2In3GfkZYkXx2I1vJjGI6EYSzfkHlaNvln54G6PxXhHr5XsQT9yPUdKhkapGGAt
YjArFM+U8YpN6JjV+adEfI/tZNd68pOxBR5E1tDkGF+tebAlNKLjjkJFHwQknZpvlj0wXaw8G7mW
6ZIhNWrppTLVyTRh0KRnVJxHU5rir2U4pQZa/40Cs6/Yf7LoVLZMLvh//OgXOqyCd2FwoJXp3cRr
yHDMtHbDLldojJ5g8X0XHi07v8ExbLv20Mcl0pkUbKDMNd31gQ0uhxJbTff430eYjxUPOZSfm92w
bpJYYsyG43usbyh1UCLu/P5JLRAlp2BeYmnn9dk2kcdYPF2SYiBo2aGgF7Io07pbDhjGxibPe6+G
f1JIxKHDsLjEWzu0nPnb7UYnJDKrvc0IWoPAQGvlRZ55R+i6drxobZS2LZ8uAZ0zZ+4H1WD2Xdwd
NcDkcj6aM/5VhaVQ87tqnGvFwKZr469MVa8hHvvm3W1cHH6xDUJFmF88LdD2RB3OKbP2AZlAbj4E
Q3naQnXzVwukBnBMYj6vyxF8Vz8ue/S3BiWArkCPjmIDHpQUYme75uT18YqMDYeYIlggA48JRhmD
0W2mbMA3lejSEnw5VBHDZGFnN6xUO3aoAGSPZ5fqJn3CNjYhebTw7lA5dJPIL345SOakGAAslXm1
MvEUlTS6hiXiusAKL6JCpWosDy9wwTQJu/5M/fdoQOsXRE/t6jbR3dMZLKApuH8RE1g4fvV6KZDm
VqdcO5MVT6ttem+nyxwuU0FqQRD15YiIR25SlYnOfz/AONpTLSDO3CCbULEYapbsPnFfhhBXJ5bt
14kTlStpQBgVsrKku2qE9+NK3W/KGcJ/a8eJy0M4olWOe3Sxjq2AL0yLID4lOLoQtmr8LVRJ+YMS
r6k75DvoR0hCZ2NhTGrFbC2VB/OZH3ya1Q2T8VzfbLx1042nvFNvPBW52Z/feHfdgn3B2gaEEADj
4IUob37mXfc5SQWGztA6wQWyANfEm/KrLK5p+V8Q/vlZDQqmKkggzaloK3M+DfD7Ow26TlFy5SZG
BG+ePq1W4QO2A5ADRGYhC0jg5QiohRj9WKJfUsVlHasqomG2+SgFQbimX6SyXOOLdoXnFclI07nt
/xsXPOtbSt3sx7Xyx5HC/RWpkWhCGCNU3zbHk1UhtE6xvH1JUzUnngFqxZBmWH4pkrW4QDcMquDv
wNQASV6Qaq3Rv48k04OrLe3V56yA+3me1qOu+WKs3F/AzT20hNtvDr4mLTgMrt8vUewYA9lASHNK
QVcLawuiHQky5qIkn5xgzpASSxHW0Hjoq3goaNFchDbSKlrqJvaYAVGq9K7jw+UG1G2v7NLBctpU
33IAlUiDEcmk3qNwh/9t1cu64Ke/gD2BGF+hzInga78n9rEE/gaGMCc+2o372Z/9XsY+Bc4rq4Dk
jGScnuK/6JYwKBL3cHDCGGNGmeIAKb0Q98Y+KYaBY1DE8gdnSkQ/DI4k2vOdcnFRIVD3HByZgOzb
nKONEaKSkVTYPYUBQImGFly3ql70aumgQaAu7HnmWTGMTv/srDfNf+C+YBqteo5p/ETHLi5Mu0ej
pm9A4jedRti5edxFPdTpQQPehxkDFoBzaogRQI0/BMcOtwHkm2R2l8Irct+JppbJulnlTsSeJP2h
YQ5kD2FYdQm5+aeHSboUlk8cWlvQIIIDmrkAb+YMUWdhLHh/L3ezV8WJ/l7GXmnk6a/TR87mi7QD
gIofi0Eu86mg70JxpIY7zCi82wpFMn0NVIagBlsXFChcDHW56OeoVr9ZCsPrF8tby8uiG0C7SY8V
jJ9U6ssXHj1q1mrbtTrvWdZ0HeVOhpJuI1dS4y6Hi4ru60z6Xqo6x2SImes98Kg1E7JEaY1tYsrV
yhIMxVERX2fgPdkPB3CPVxP/Cn+r+kx8V0kOgyhV4lPOZ0cSm05ugUTIrF2w+ElMI3Ke/o7T+Bst
NiYxZVylnupziJwMBaJVdkPs3VgkuhlYWwKOi0+q5NhH7MuMURzAO8oVN836BznYBF8+pybZGrVJ
LrOJPhSkxekIoBjaxc2fgj3P8nSF3QyOGa2zWy5IOaKLB2a0ttXsGhLxSncjDZ0Po4xzTRxCUqnj
e2LtYwzAV8yNWv+i10SOfw3oZnPvfFu80BIuUcCMW56zcB5WNRy3tG+qjWIay0ibxfwmbHb0Mcas
S6qbNA4wiuFU3b6huv9mCC1QlGIbRWyyjfShwjRkt6DnBCT2zt+9O9XijOT5NgZVerf7SYYOF+S6
2QEwaKlysD20xQfFszvXOYJa2tbcU/tt/zlip0X452EnCspF4NU2MWuQIkdqoLuFOjtY2kwZ39+y
rHMsEnLLvnu3dOr2E2tKOY+xL0PF/kSw/VR5zIiemnv6z0zSGs4nm0Jyjoy+6zbS34A42wMbvtYp
rOqCmz0CdaBd8g7nmGqmmCeXdXWgq6cChWuNsXmQIog5PYXYiZxj6KIEf/wIiFF9T39rjodtsBEY
nJv1ECDbdAdDccaKZVvu7a41h+JZBaJSUWsM/UXwdw5qpRzbYYGw4AJMTpB5PEsqFNfyGHIvorZE
WEhT4SaXHsn11tnM32/Yr1i2srVeyVRb0Ns2HbWN5IUq5lMb5L2qFRjy25rkvbrlZQWLLmSh5ME/
NZBAYJQpgrqkjZkhTypySwvM8K7vHSjJR3OZSbxcqrZJjyBcuwpQ8ODC/me4hDswqbfn636J0Sh2
AwnaXhgyxPLxJIkqN+0wComZF/7SJc2iaYN5VpnzQi+btmK0KpKQb+3s4mVCV2Bgaj862aL0jVLs
ROusR+UKw50MSKJXwzcbuFr7nf/FAT4a7Qnb35Vrg7gXVjVQijd0IZ0B60sd0cZQfQnH2QFfYiyd
uL7/jXY4YBZvOl+4fUUpL4H3pZ2/CJjgzBkS1x2UOrBFsGjbVVxwl/hbha7M0UrndQ7v83m3s+L2
VteUMdT8M1Q7XLf8bhOXgZCfwv2hsP9zYoeIoF2r0W1OnrtZHYsTGtAnUn/zVavUKeq+PzkwerQN
XA8Tcre0nLHcZl00Pq+6Irx86EX6CW+sAxTABvj8Z3TZhHUn/9jd7PkxNZyij16OehzwUXJu9msn
M3Ks542GkWTb7a7DqScDwqH4QcLZcyhyG05XTxOXEv3apikAcTD5xzIh430O6nB+g5ZaajAlbfUu
R+PhJpQtwdw6WoqYAcPyfwGwYgzjc5tfa+zsI3EYwFeRdZ2UQKZByfbDkEaOBdIfW4BNYhlZMhFp
JR2uZxN83qIH4QRJivMFL0KfwxPJBzEveAuXX8DplU1QhxgWXltgVLfr2A18IUbsXkIZrkwxFGvv
nXi67cr/ViqNHpSL3Pd4vigaVe4eIR2UubDjjuKdC3Fl6cuVVPk52yZQXBNXjfTjtgsnGrwqj7nd
rZ+ltZ6TGHuLh1YWS6DH2GPzo18orh7dShKrrqPA0/ykMUaZJIY8ZZRVP3Qjj5nnCRySkcrb91xI
KfcNDDiSvmj9iPKnleUDNn8QXc1UCXqRfipU+Y87+sX5EjmEc4AGB8SdlA6aGP3iUSlCTw43NkE+
lk+KESSM6uhD17+tl+NrejoIimddbKiDUqsw1aSh75QE2USlUv/kYfvrgZ/abG0pEZMFbe+RUI0S
PJPWDLdhl5y6IlwtZ8cEDthVbx9kpkRqqmkeBF+dz76qta5NzQFmAKNQ0cf2g2FvNs2cAYXX95pt
xeuahd++MRH671Bm6e7Qh7uzq5Q7sx7YwLBCXfKpkQzsqVK7bQ3V4IHWxWwRsVaLiTa8QYlO8hpD
J+7OcZjqOHzjSgZwzkv8179WlmrkeG1JNYGtlmKbaGDqlNZcCWxesrXhmgC+t3vGmZPD6BGrwNn3
VItNEv2H4Myt9KeZXOg5MK+2zhVGkjeGe5SGd+hwOk98U/G11d3xzoCpO1Z28JRV07c6S5hbFVtK
x4+2Cg0K31i7TB9hL+ixAS70t1kEj5ggdZbuhM7TaitgSL2ibfZ/A1nw3/dEe8EzU7/8SPjB9z1X
WKe+Ql7TIIcJfcppemFlb4oAWB0xQgJH3cWyxSQQJo71R9bcaWLUXURre0yJSSoAewACLj7nyF+E
sG3BXzZEus52fbZ9xbcmSQF2l0AVGgY44SRERi60oeEa9HsOF2WZ2ienz9GQ53ODVyeaBqJ6ioGx
F2vlpRdjMyIY5Zwxu1s1UGBkdnnY4GilrAM3aLNJPAFy+IdnsEcM3MRcZqundHgYSLh2T+CAg61w
jAs+whoafKdqZpeMyi6Ok5tYBxEeSrxnn7vuNheSX0S59Z3WQpukMrNKNCvGKKryZYIvkSDE7rc+
iKUmHV94nsm0FNiyC1cHYrecLW0eqqI/B6IPieEXoEJxGSLT32MxGql+ISNoyJL7ZUaSDLRltkCp
DQa9DSRFXbYFvkuadMu5U+oNH8Tj1k5EafUvuLgMNVEjYl6xpX51xGKtQhhH448HHUiuEzTUu3FF
wXBZ8I+JUdoTpwAn3XA6/H+mT0TCNKte5qh3XQBnkFnnVd/JeDmPsC2aVeAAWFQWVllCCcz2QYP/
OHku9/eiHocKgLuGO4YdX+Q8/r9X9YYDCyP8rInx8fuMf6kXZdxK8KHnQNW3taNtXUdj+d8XK9x9
5M12TTSgmNRSv4XcRnEC2kRgckPrPWELiVS8Tu+RFE8FBSmpMYgesq6+msH20h2cl+5bJ8XpZD6G
YLIbUDcdhUgTVOBFfe7r70AqW7k7cBUC2agFjsBfe4jEVSTKdJ/9yesdPXj585YY84XRjoL0SZ0F
G2F7u6uoufWBKJ+/xYPM2u/Y+5u7vsXjISGWE1HPd8PEl+3HKVKsxynG0bH2o4GKTZo0BUG1ed0o
Q9A/zL1x2HElUYj++I7lL2qrI5a/AFp3KBTJVuA5KTezaFzwA75ey213hUPVURTaaRn96ySU4Dms
D+pU8Om/sH19IC/jYvargzZuZ3b9yCiyS/r6ZWKm6jVKpb8ZLu75vBLWk66qJyyAPo8Rks7WAfJT
nKRyKyasvcGNBAjT8u9iJGVkAn64TGN8cmWMlIAo19g3HnC8LMhYVqBytERfMuY4BmvIGgwfArHf
Nu96ME5rCqdBf8o7dafivfcm1I4B8iSG+tX6VNXD2Ec5ioNQHchlcyWg5R9H4qzm95Hi7DzdNSum
Z3A6p/cllYbtMeZ7R2HN+nYoLj0kQafr92rCvMolAJ2YntrFFUiu+1mUsRCIxsrNow2XF3LYFCQw
xz5DVgOuDyV//bgyFb6/xlitrcx3B6qVMFRuVIFz6fcsoIOMIfCkCM0kIesiK9JD5gTlF4E16b4i
74cfypjn7I2hhUS7j+U1XR62hhAehLTJXkXwO1vInShCbHL9MRoydr8spDtqoCivlBr6V96SoF/1
gt/Wgs1RjyAX5hpzpQx2YceBaFvQOobbtKSLG8FTHZf86o8H1t6FqUYwzcA3xbgUx5Ff6Gys/OUa
s+I/JAgbfBy/giW8tyYWtBdkHbhYXdKuQ0XnH8wLLTAXIIxsdEaAVlEhwEfeL4SSehMVAZTZi0Fc
+NhUus5L+jZtWkicorbNUgGIVS89H2OUqccgr9LF2+uJrs1lkp8SxhObSxK5G62IkbbN3ipKxfPU
h9Owqo5bPGQVVW8BY/5jf+uAO4hJACE+9rWTdZRR7H8HWDZNx6kFiikxnJSCc4nBlH3H/mTVSe+C
x60N4Kt8Ta4DatO/w4yNVWiZo07rFei5HE5av3Mtrog+bx1NEl+JIWgDdnBb22dEo/fDTellDmIV
wU+nFZLhoMTqopu0WBzdrL8X7nK2WFCmW6aud11EpU81p1oixjOgsCRxABAUqCGj0fXSpf1fYcbq
6BxD3aRD72Pu+Q5CQ0VVyufdBEtsJ0ZIo7RYdTkMZ8YRl4qGRmLjaKXszgUTyFo6wxN3D+Q9oXcJ
KyyJ0n/PlftOrbBGBmfCouGSIXH6XmJEcgXjP3+MF0krJzrQ3jL/EoF3tr+qKtpGe+8gQFqfUXQF
qpZraK5b18AOgjB/adpLNrnQsLhh0dN8IrvYHnRT3O3POA91ZsHKA2DlNEtXDs9KlBUQ9XRCKV3V
KN5d6zFA22gwfUHK84P0yhV1uc1of6yW1dU94TH1+D7qosKwmKWxPUQPT1TzmRRRdRMJC6snudkc
2gLjuAcbW10apaX1J/v/KWRMNAHmrVq+SnxAFkGHdgWWbFqcYDS7FUMco3BRtRHuVqj+mRwhAUA+
ugeyFR+zf5K1AqOs2vGBws38hXmU0VMWfwM9d3Mz/fWYNgZqCv0uzWi9ilI7r3T5CO+ccyLqy4Pw
b9uzla45YHwgAc4/afTeYp3HSm/FRo/vmugvOZ3FsbLwDQCNIhct2O2yQq4kXDyueBeBg/N9ThOz
6iK8gNp2sGzENPh84UNBHN2E7fpogEhNju2V0SKBO1L5vhStvuJz6y1x98AeNBzoPTbjfzjWBMwg
u9OuykXTvmDhkt8uR9RtKSr7hcXa5sUDPeFUjNfCn73950DXj5Lk13fO35J3y8uyNXiO9UR408sF
zFI3wqTPSmON+wKpYulgp0zJ2XLaYC8uFkX9ByVZAHU8GxRpNB/Xyeqsw2rIgGvmquVrgDBl3jtW
OEcrHG++J1oJf5bKS7kcuR84sBRBztj6MjM1QAAtTGF7UEMrJwVbJO4YkpCcFE1hQzGVwD9eEb9h
SzHaud7S65/j0aLQL6lHCUHBoSkwNo37MlGkODh/GEOVxmgfrtQ1gCrrdX8s36kccXx5fMCoL+q7
2KvXYGFPiai2LjDmxEgGgi/rM2fzerf2WnLEfqcx9BJkmJzJ5Sy9Yu2Te9RWvekThyIIzDqTXsZp
qcueK91f7tMp1Ne1bx6/CwCM5WGo8nNdJYd2xWZ10P/DV8AQhbQ6iZXM9HnvvQl4LSKuFL92Sg5L
usw7qC5bY5+PRyuA6QOZqhgY0ETHuN51Lzx8e6aM+DQbFDRe74qp1OnSWh6tItagNaE5As0GV9BW
PtcIXmtvwWkl02TSVSN/zG3uRR4rIFpnUlgoKtPZSbYyj5Z0w0nP++9eRE0uGjPTaOxBKJfAHLPk
fUaCb8gJ/rN2dpEscmXNy44W+EX9XQY5O+csO8qrntXrxo+WswNtvtxLcLCXK1RIsH/pvoVBi280
KMkGy2k5vo7apdVEprDkt/PjyNgF7EAjd7nNdZ5FRkGvrAsgRgiyW+rJY1PAw4EeP8IyZW25KGHq
YQxFEHqM6MY1W41zukxYP8AFXqyJKSEPtvvqW1iruQZPePCwsYjhQwDot+wHil9u5toP0+N02DdY
DMeXOPj245P9fEhjZv0LKkqWVlVKM1hlcxy6ykJ/zxPAl8z1RqSYw3aAjog/AOL8NVDw6oy4YHa0
qGkn4fFTjxH9JQ+xZmemaLzC9Jj6/+Gf9pP5/j3rcXVqob7ec0WgO96axDKoeo1GJQ47I6wRNSLF
KCHRk5f+n6w47H8UWeN9DaiWM2xcA1HKz1oHGuNGyhuSJl35A0p/MEn/2JK9kbEjMWj9N7WwbQiZ
SQi4ynvSYmFykLszS12Tr5SDS3s34/RrALE+r1VCkgqd+j4vXltsP/oqRYlVaAQy4EUJrrdnSL/l
Gk4Nq0SNk+ZkLOALuXb1l14XL82jFNVNZjc4uyr2QO5N6EcJ/B+C9vZ2Wvr1Acfr/+0JQKksboja
12JSRsCEV/g6ZXiW3qxbYGUybIop7UE5Xpw8Ugj/Z4Bk1MAQo2mlfI6Ajszgrx/qFNmZZhaAuRNL
Bt0lmkyhe/1Wk6OPlYpLvR4fSIItd+jPnABNdn/Muh8S/z/cL7OHSXN5MTxeUXfL0HVO4Mx3E3Vq
vFdI4elVmhKQ6U5cFYOxyaeyS7HVvYdcVix54dEm7I+pEzOQiPFs0rC8IlclGVSi3hAj4a/bCGbq
Aq7aucbov7OXXDKbFmk9hR8jxvH70LNiuTkx4dgqRnH1AFil+K/tT/ZMeba57rqn2URW/iNttTHr
qP7oXMb4uyH2qXTkXVHrBxx0e8Xk1o6mOxaaLz3DBgI131OCgL8UmdzmHaDxnwjTGDM7v51mVHpg
8/40gcUGrZ4DyeCWeME52kEtajBoIaghDsQPzEsrXGFozVZ3DAQ7GVb3J/XgBx8lzmB5LCU05c+4
TR8P/1asgi9hfWezoejucNtbkLlVYkmUghPkhOELxPU3kb+HjH2xgdE+g1l1iFYOLdWUQBwIyvJo
et9yB3I67kuUITFe+s19/gnHTnJPaQ194VfDXdz79PyMV1qEUNU9Sj8bX+eekYGndk2Ngbqvyx0H
UP7ruGPBnPWyvCgR07RT1dl0cq14A1MDgvRc3VLHiPT3PcGfIfyAnP7nfaab/eUjvZ0k249t6bTM
NIy0fLkgIuEmKbRhzg4KoXKNzh9WL4lkZM439mAgLKkLQG86aw+rDku3mX2DJUhE6h4zNA1KIuT4
L+QAesNtLElzMBADgIeCp+JmjR2ZwPZSSj+SxMLMbOpH1Lu64gXR2jLt2ow7Jf+2Siaa371VUNtO
MuPq3nurSWu55BnJCUGTjTesLd7eSQ5P21FADxNvqtv7HyF7ejubt+IU0Jwc2dcMtoDEnd4jwM2n
E1YMHQWGfSZwF9kGUax2KhBSu4vCLflj3wSEVXGlZeAeOtxvLp2EotLZnstHFFGn/CQ0RIDQjpPK
vSbRp05YImj1cWWIQ+giJlKQVCQgtc+Dl9qT7ra4kzIkeWUZkedPEuhgwnYx4jozH5pWKFErHq1e
wAZjYvlT8enoP2ThdDDR5wlhaCkK3fhbq7X/93gcZ9EDAyNA7lXEWZeo8VtbvIJ8oJXbK3uCtNqF
C6ANlmhkULJImQw2yChQVZe26AF2fbQar5LW9odXhtSWw16C6dKJd80G9Cj77hXWdblmuZldsmpo
j7ZMdwcGI1bA2XRG8Ne6MrYnegd78EGKDWspR+eN62VuofBwZzHPwweHDCO3c/3OfbBqtpTCy2Lj
SPjU5PupgEpy0FmNoou8uoGbfoFiMgi+ddnIdWWxXZwg8CAgttIzWnnOzOgRU9DaVxtIpFGYkt9q
PkoyzzdWMQcGmtfWWF/lOMAZf/Ec4++ainGQgXx++h1S5M+L46QSWfYEURchPX+6z+OsR/VYt+jo
Dp1XHhCZZrGmkMp22WYIy7VsHoutou20hbEGVK9AgWwOfMS9ZK0Kef7+OCCE1wmoYzThvx86HntR
7v/RqhbButdHpjPLXj6pXmLSOLsUijPoxK/sECaWkM9KvBZj2EJVIHJVAkR0hou8IxD/YKw6K58m
jacNGPv8L7NAZXlaAPn/VhkTdED5aJ2TYaCAE0t59nH2+vRWrpzDMwOp6S7fMGzd+dHx6KR0UMOY
eGzSGoPurRTroKma/2BKD562m9ImiRCLoS7DWWs2lg01MxJPKMssWFaEkjaTuQSu3wAqulmbqX2B
91sk/tMtEnmPT+Sttbhx66rFXXrEHjNg87dFH2pg/KDuz/uOev31/kBcW2gcXx4cROMkTY5Q2/Xr
zT+M84w1Egs8DUz8R+wAxnlmr/cSbFoWCkaylSQJZftGBbY1YIVWHhnwsSbACbjN0ltj8A3c0o/+
BN4RvgYyl3nIOaL54vw62V4zPEX5/77LkqNBFw7bX1TQf874R/9fdFr8rv1ijgaviCxAM5azvVKT
1kAQnsWpyM6wRIxAfUTFZ5VhNw6MxfzKDj/A4XS0UJfuy6QSZkZp9KC9c7fw156dosXi0C3UJ84r
cywbVJctmOHwacRDzipcu5cv81PapmE0oa3ou5VzePywIYcCGUcWNzu4aGMOJMjGCsVSBrehWdMr
KuZOJ/9h4GQRWu1mfDWBm18fUJnAW6humSB2jxPFUX7hunThBYa/QHgZKpBlIrJOgv7qmae2xW4Q
uK1kD1kMsPYhQj/AgUtv/WTILQ6/+4Cqg9h6xZ7VudI69COrK2yxWKnn2BYpHDbgumKwFHM6Kh9i
EERKnneXyJxWcd0jLGDRhg2EBbucwP4/I0MWsq/OA2mnEzvWv4peNLYFnHZxc1ZSzoDnnKJBqy1x
zkRjNd5KLoZOava7aVHJpKHjt28nifNpcG5He5qllytB6AtLvcMwex6KiNtk/VwzWFVxHWnox5H2
ZDFl9Tur462iTuAu+VthiQ9B0fsZM4LCnTYP476Q6oKb2mksOT/JVHdl7Tysgixtn/a1QCFS75I1
O1kLFlfhC+5YAK+vEouoqCDgsqxdI95Atz3ZsKjZStpYP2dDmKfOCwcLbECJfGLH9eLSD6DKZ8+7
YY5GRT75Hk5GdpCCf6zWtahOJ9qQDZ0WxYShZo93DHaSf+G7yaozZPFrf30nXdc6K/pPHkpo+zfA
vXvdnTHz8tEeJLi5OwxkHQPd0PztCpui598Zo6T/nkJ9MJMLkZjVYBFS1e0Tgk3mdd4k1zwGs77j
pgq92BSd6Adv0j2Xa3FX8vQy6ty7OiZ2Bf0dJA7I/5HVFwE5vpHsqAMYQjLXLIypB+LJ/rdyCODv
AljNcuLfXqSXvHZmdTW9d84VzLaI+JsiaQousgCKUEhvSW1wD2X3vQFdo4USqb54eaOC0l7fbDtQ
kjoo7YxIzdzZRCpRc+QYP//3P4ioS3053/+trFfbWXWZixnl950L/FxB/C5rlC4HzfhNx9FStl6+
pcE1skKh1mcreocIYBbbMAaXZWW1Pv2i4eYCJ9XY6/RYU2wuOkCUx01OhFXOaxJSGiCcapIOhh1f
rpi4ggffP+se4pflP7PyTq/kznjyD5A8df203rSOciAOTpJg6RhlvAKEcgKGJEdBdbiXPA3mIpZq
EO2clXUp9snuBg82zvVIIvMjwxBmkMd3G91xxf/TG/nnGCrNSCTQr8KUsY74CTT92AoeWu2AkDrv
UxGxbYxz3OAEJ2VD4Ku6OCsNqWuXvWytMOt10hpxxa05UTbYz5dWqtyHcwI/QJ/KHKvpP04zCAZk
WYaT8UQxs1pKRk+QkXReBLctknEGJcBzdEZpvQP6mLFxefN6rRrJxEIkDdwV5W9DjvQtpcYxPe/5
R+xvFXpbQNYUvX9BwA7H4g67sCKUGwgHWS4JJYtSlmmdALNDhHIWBQD9mI1c+tlTw6AQPdfAkZr0
IRfjAVylluP4Ze3LLPq39hzdU92yQwntgkbhGbRqoQdg5ZABYCs9tS3KwElDIOw0eWg5dQvtd8yr
12CQ+a+sV4otk0YEnEeXz9h6GsKFsskSoUBnidcTt8ZsFAT0/USCDGPhhDMOLDyv1BZtTJU5zydo
X3dCPCVF5V2DZrE2sXq+r3ZPDrpht3WUcSXzvu9gWptNix4svh9w0VrVbZidFX5ZIvFIyCjGIoaj
2TG24rlPZ0aKSAfOxGmpXTg1mhW2FyUJ2L6DsuNNDSlP0qpASTNPF4u7EIXfdo4BeDDJnRcnzlPF
5m/QBJ3J89AUAYcSooi+5XjSp7sTu4C61bSxSuxYa0bjch3AOTAeJ+5iOWHix3ozgf5ZRp6xCITe
/0V18/vMk3Em4WvA6gi8QnfvfS6KbBkQfdQlnif6th/GpcQHVl4a2GOUQdgtllHOFXCbScm9eDEK
I/UZmjlB7w4sCYHtVrwckRMsLMXMhylqts0GVTNXxtWNxNJQkB5SNL09VI7wbHFIGG9M1q8SDOG0
pcCK8KO2CrLROjBrSvTLkQFo+9z0wgTuzROeRdrCcVhmeUMULDZYF/gcSxgQe+ycn+8aKCNugtfw
2cvXOse1BIbhtfkC4yVynb+Ey3ZLUDz5ylRoPfJQRu4i3DIGH7of3QcIHuS4klr4tOlOTYffWPD+
K+acNaac0+maY+GHAhmqYiJGFy8h60xnVBjvbFBppECVHw0dmZ4lDCFPxmE+OgHtQQkDS7KmP5VS
2bi0wZSdI9l0/C45+EpDsEuPXjAL+7VbpmNqqM5Uv7hYZjpW6SnH3RyqIYsl3g7SGCwCWB6+YR38
9wlFt0hd6tZgP1Pwehnbg9c68XC9KZOTAG2la3aONfpSisJ2Y6cVj0476rOyFQG0sRequ3jpTy8j
QMAI7y0EC94w63GjIF99KDd47yrjyM2yB1EphFb6z6IMvaQRNG36CFmFRH6TXW4hscHN7X2cV9OW
KH7zXDchmylwnx2jek0KuOcQpfevBiJN8AoQ8Nx3yzAv4IH2BNHU925BOmZN/GmnrrNvGcoTtpJG
4PDj6e2s/IrckLTe6SJan5nMWOK/8sEBWgRxCvt93ImnaUS05zosenjPKj1/8LIOe6UPkFVuZXQf
4v7Ed4Jcditqi4/B9xYFmK/FyZ+PJIS1KpBAlFnNmmuhm57rtYoNiK8C6tDOr0jQU6T3f/6G6emy
TO5vOjQH71fghKdAY72sMipvxk9VKzyYt5PyYounBPxRaKcEmJrIbt3OZtcxOC+muDNHEzXnDZep
2uMCCU+r/n+xS302Dhr7pCu6aiEA7d8/l8YMuuwiafxX0Qna6aQXqQ0fF/7rODppU6Tn3KeppePm
K4sJlK0QOeGJPiR+QHKM1AhhSjb6zH2dBRZl+Kqt91bqoCnhMTuwg6Lzhs4wQ06LaO6hUvVZZvqP
k6P5xvB/uifcdBFXhXGihfvkVM7XuYh9vpRIWCNM7X1f3yznaCHtWpYQM3S1snDWo8NH34ikfSFI
PskDHTsbUf+dwo8RvsDeDD+A61cQOkTbjHeUHseqwQE1ylInB7aKbsRWFeYIO+Zk2JZGc8tzfVs7
q9Pgd8zsLil1XejJl6jUTixwXdTTe2G6U24Z+xQkW13pE8AualdWQEP3BGkD0GeOFkAVLS40IEgJ
w7j9sePcZcIh2VFgD4zQTYrxsOW1ySB/EBfIySh0bHY62xIMB6oRcHXA61I8BmaLuzVUD6XNQce5
jC1MbPizXTNI61pWn0T5i2/PT6aq0xr1PqW1+DIEjhYl8V3lgEfDHMlAkY4cmirWTmpFBRh4hP54
w23+2BBQd6qctus5PdEs404T3ju/UlmOAHkTX0Q/lX6Cf7zzWXlTcgYeMXVfqH2Wn9P1FhIAarAG
ixWdBrFU3ueFQc6LSiGocvjStkeuQHi/TPxYHuD6jOB2cQkyPIpbWUHKG3z7uBU3Ejb2iaNZ5fll
ehIcg3DAdZZrSmha34niF9sl6/ljTENLIDml6Uxrum3jQjypEauDSxcFSl+af6Z5qBXq1aOifsGl
4VUEdLE5NS/B60EURcIlAWP50ltgsxNIebUbpeOFZRrXqLALc2w8MCrt0IgCuw7OX0OtkmJvxbDI
Ht/ogsQDaQ2Y/2TWHzELuVy6LsR8FpyqLHLutyVXz7VUCFfXcA8PvUSAqMIh5JmuscDwO+ujSsbn
iK2jYfDGgRZS2j5xgyY9K8GqMTt5OJSZUNgg+2isHvn2nBuV2XpivKbF/JZ09KWldPYNru0621iI
yrfS263tiaY6OISX/Zio5biandmzD1DV5JuU1ono5NtDcgxQcXaeJGBHc+23c8xEz9fcuNjrj3ad
p0QQf2q1hmc4vovqaSGQ0i3tQVUF/zX8hDQzturvuvlBU9dEhY4sALMNbvgyxSRUoXQe5rnFGix0
L/ncKoUQhWg7eCARsK+AvQlUnxRHeGt+BZlsVgXo1AbPKo4JD4RDWL7KLZI0VY2KPFLFE2ltXYvX
mMu8zkb9dzeDMVMlHBpYEBC8Y8u4hBaCrqnskUx1QGeUgxxbdBjMEKpYUhXOYLYKW+G3VQ864tnJ
XNoNl2NykHUerNRXMjHhGRV6+syvYHBwSYVe2RPXlrah9/lgZIZ6U0tfqJ1m1lXDyNW87Rr7nFeo
wEWFVrPU5nc7CdNfGugAoDjNZJQBjEKChM6vTxftMC9qCg2wC1YkQrcrVKObrBGHq6BU6eQZrv62
fyTR8RoYecUie4IXvbYV4GMp9SjgJrmAkVpsPmm+BBxgdz9R2zldRnUSnCHJPRM6IYgIpbCnAxZV
7oECkTm4YT2/rAYobW5KTWUdlMLV9hbEu8oHCXqAUwXaxbYgD+RsYCBkw/9aczLZNlJeNSZ440lK
IJ9zLe49SXbmiG7Cp8JMZVHhJHxm60JlN0OYHB/ajQVza87I3afgrkYFOiBOi9G5HLStAIkpr+HI
L319VCh6O+Qec9zIA/eZE1+aIHkOM4RZnLdr3Z8WZ97wwRMcFqKBqVq2zZL2TwRr4kDuWPhN5ZvJ
1qNjXLghpbKbcsRQK0SUZaRwRgZxIK8fNS1QIdjU+GlTWpZHbLskti+K9Z3z7C3zgHlc5bI9R1I1
jbUR/VvjCaBklvrjwSW56KhGAE5VJfrxEhIaXDDHbomo03jjLgPYpoiDrXWNOP+5VLuxgZ4hwU/J
gATadycONgT95MYBmUhQm5jzL/ndMr9OHJlKqi+tcCzqMrmJIaUTcnv4J7OYcFKUnm5mBpEdQgUQ
CrGuNTWZDF29Vmku7YxyM4y9pDGrQYgYslaErnjeJsdpXlRyxhhKFCX3uokA88RwXAScA6qbGDY4
05QQalVY6UiwDpKu5CuJAQwjDKlCSjCQFjS9uMMENiwCJKkAb1mUpWJ+8B0gBrCpkJ2/+2Quhb0d
pP4REjogjRZND3rj2Hb+PqpsVQ57VLKvxKSOWCq8zWKm9HvlmrPafJ/7DOmcTX3jyUIws2kJiFrS
iLD6UVeyO/23F+ws+5hWBc5L1coucqwJ8h1GIxvO8W5c7HVlthvrpWBct0kaXASxlaXZ1UruR2Eh
wK/LbAPRj8Ve2uF62RWZEeQZa/FBNYgObO88BRJMjaNzsVDqdTwBi6d+OjxRbBEcR4znA5pjTgJw
gqZuBDauXxbvAuQXFLx4TnPQOvtfON2clxew0WMBkfapwwSWRetgN8eZPLJALUbqyX+xl3x5I2Tl
feK+Adq4/lYhjESFlYukYDVd/LsBLnh7fT4EY58r075ibDRzWTpmjgdMitcH6xjWgPtvtnZN0z+f
6vTfX/8bYFK6970on3FDdtf7OPT5nuI8J0z/MkikeduAzG9b54XFE3GLE0COAqxGX6ZRiYDgJAp0
lIb784OzDFEXbsFWiswac2U32ofTwektn+yCtEQ0SwcZj0rGqatDEu9EsosEt5zWWwcsfVO3DqtW
UyQPCrRKP5WNwrTiwrGsescNEyGOeTZ5UY0RO1Xz+odr52rZzSeH8qqJFg3IaOR5EWgeq/6BBW1G
wZaH2dZpw6fTLSXMR7dTnJpgxpbN/+SrDVia7+d4DsNQaeWsYfSOSD2eba90qxjyq7MLxhrTO86h
C4pA+bujn35AZtJv8eDEnrbgS6i4X9rXBVskun6eODHWB8Ub47d5F9OVhKlIayDwhNne8dlVSwc1
cn0GgL1Zi5pbJyBydz67uQZGgQy3JyL9JBmI2yKosmgt+i6jYqyHqxjKLYSQZakZsHWuVMca+75R
G2vxKfsMVKCkCSMBS21h+G36lRB7zvFK9FFp9DBMnwCrqoW1/Ka5YBOugi+67MnZvVFz/TBp7CRH
DLZYb4/oxzexuijxynoifLnDSJvErM8fApE91I/Jb1pfueZuvKcYmgW+AVBXkVn3/ls7DKroSTQt
JtPVd0xYHmA662EoSgmnyO/bcwW5WiAukXNDM3xrx0rpopx/Puy22l63ABDKcJbFQchFCTANCxj2
jBMJnRVv58iAPcsxBmZ9JGM2gsMbn1z+pcQvTB7KXcTrnQlkGm9sZt7wBSCO8Ipm6Ga9U/J9HIsk
r5Eb/jCLXPxNBMgB5r9ig+mV4vc3lGJ/BvKgfDb14quysnqCz2hAdIh4Aq8avKxBz5cVgxV8IA+d
jKRftn9mMSTGzUNZLZA44/1bXRGAerTOgMDquXABOCruy9qDJTFp0/7i34nusqm4yJkJ+DcS2cQ5
qMaLPgn6UYWvDTYcYE1PHGHktjsqI7SkgGPpjiDAB43Piq3e26/CLrgD5wDY1lZpbj6AJ7hmuJ3D
CTUylE0pUq9GioaAMTXjFjpt9y83zReHHfbq2wqCk/3vajfy+B4624PCvEngXvaAeDKmtQoj0grx
oIrtgYTqDzfzlMMdsQPQldqtq7AAIIm1na/7x4iNPP0AyJnnr+OZYO0FrsINaR1OBnviKuu3h1dP
rCkBDP04738RffqXuSLE2BOJMkNx2bXS8K0ATlw7O1sq6oZrOgTCKz0XTneqFAVpcvYc5yQ7PoTb
zUl1LjLKEgeLw5w907BQRBCXAUcsWeDzUSri7VnUjAyiCJcNXrks5mMQm1rAKTQeK0f8OtX7f61f
WyZg4hbPImNrf9e6yqEK7CMA28o3JmEeBgI7dMZB094uvzO/LFq8ooZTSFelrCt16v+Km9DNZQg+
266muWV4E7hLm2O+H6EAoLCgedn2KYplNq1Tqk/WSy+IxyHEnZy57KG+XqpWTuTgHvSNlEcrnxaR
nmIZWkVO6vry1dzuqJ/ZpV+mNHGoBIzS2BqjnzmFPUKoP5zPmuXcdbpY8V1jFzmd6iF978l/ngDs
ABS2wYRm6akBl0JIwRAc+BndzVHhoxz55IYajjcaBDiU1utMR5HIP6A+iLTmDNYLrxh75Svt8100
GgcOyC3haUNMHFYUJlifvQGMoiKjxfRe5JjcnwbWxHhh7Gp7YzHKcQEADu/aADQLTgktDuP2NSBT
8c0/GFDgp7xocXQCnLMCyje/NIrzPSQI7wLN8nLT2xvBnVCaNVnF0A9uk8jPwOd733FB+ynkXW1m
vHvLQFjKl7T1025VXgbfpQ5jmgmYXbrpDXUBZd3otZSairklw3Pk5aFs1aQNNoOkS0TnrNN4Qn4K
vVkCafFOAXv717LBHYMDOdV5EWeNoTkM9dakI3RhrpzPqdW9oS+wxRMxu0qnRqT9E1aJXNzaaiFn
Y8LXUqcVrPJ43ZDk50MMI8vNnzidjmRR/DWzHkT5kGdwH1yLyjhKbX4Klte1Fn0+GF+N5NF1wmnq
NtOhYEc1Y4AbaKS1YmXcSN1NR45Ic7OVWIBANFhbRNCdvWgcFXdPCPYhRclk97TRoo8Unyprmx8q
7r9unepzXLGGqxStWQ2cIB9o9lOhGfiT8rGyJYoR/OsmiS7BVeFJPmbCEyrGELIEeU3cc2XEEAvI
9aOI8BIVLPsj69t/Jk7kTUd0l6fXZAyEXEnvOL0o+X1SZD0vKQ+a4VW1AseGfYIL7ZBHBhFZvu+E
HbgCcODU/sLqzMMVi4CJjeWNtMW63pMk8HktOZ8FeXZVu3VF8ka3apPTkEiweil4ikSfm2ChgTci
hKPUT+bp6dJ7qwvMneD2LStBBx04GP3d7f48EgNLfWA1nXQCW9gTNBzcOmnn75likq4bT4JiAU+P
tGfm3j5WkBB4s1maGFzA9vDtVwAjw3XnRXjhSWhtNA+NVg4OQmnRSPD7+ekKasCIsRDFLhDQs94w
oP26MjDvLUvyXkwTRWUUIlSrf2Fz0OStbi+UPfFXkO9tV/NGqU+XSmBcBFiWs2LwvbgBpoXQH7+M
gwuOP/iNQNw0L+FhDw7kOoDjSL3rYVWVvJ2CU4+wvfbIv6HV4hb4AlZ6WfP1zGR1/rmBlVgHR84e
EAqZINded/Ly65XlXmAPT5iDTpFkAAXlbXgKa431vd5gaJaN3KCrFDzulxwiIbFRXBOG7vaDp96W
VYRq1QQg7NKXmiGqfpkR26Pf1EJdnFpYE0+6cENgTmLNO1bzcdl0fU5nkg1WVhZSfnBKANSsAsvB
v49dlY9AluT0s4I5V3CuFrL3OHDAnt6ah4lQXPqLb6IuoZJC0riEmynERvCJnSiTLpzYIHzc3B9D
OxNOE4sndvcZQUhF8ihwhfxT05tG8zT/8rTvO39D7hb2t9T43RojojolkMzqWvlwjFtC5cKk+n/5
CDKh0Ewt7t43NDTsbX6TEXLiM+urMzAiHO0VrWpPE9VQqfaRFCjamAbEfK8+qYpogn3+AHZ+8fQ9
DL9Bv42Qk8l+JkBRct6AfH29rSXlSkru5IpAajlfPCBo2yqIGsvtrdl3/gmCyLRfuYe6gHXZVj8k
EBQL4Z4grMK/bKWSXAow28n+H49ibUuSHOeHd9FObFpWKS4xEq8/hIVHPgFr0OxUwtsHCS0Lv6DG
fn/lrcrM/Pt5QBNIemxVHw/DeOEDQpHLzmkwdQClDVW3p9E1tIHxBFvidW5dp/8FijfHNV1G1lrS
kmfl9rtH+FVO55GgYmwOgFW//VS3qRRKrAa37NkArWYLQ2SPxoGgsYUpjzLWAd2FPJ3vLlM/znq6
t7gkAwOJjB3WoQ4AZLPuFNdAD1Oy6ohNY0GjkbJvpABSOqAfwZLrIvEPxzLT1QCJh99OqjuLZLl8
7aNEvcnHluyujXrXM9ZsNDAgcVtzWM+nyG/6O7/mRrko7bNHLfbeUoV5tEp4mVuPU7msL97Mu70j
FipIeMJ9PVSCN7z+gfstmazGrwPh8//beCiFA8k7kjbhPrO9IImRPOKxsy93zypQtVV3lrHKIF40
/mvFDd8Mx0OyPG1EunyLyFtjkW1qYXI8PCiJzcPqjNcsJPmt/aZfnRP1WqhQTHcco+Ii2oBOoGhG
PACzlzHj9r3djlKJk7SfJ9V2VlEKbrMfnzX77QihissyDs9iW9Y3kQZfrijpCIMRXPhaOo4Mum7c
e1Us68E7j9Y/JfSRBvrKYjnQEE0Dq8BWrG9Ve5/mtNHhqwA83LYG5abPbm0YQ2AYb7H4+1ruREEb
MUB6pE5W2xm+Tn1px0f1HbR7zaSJayudyoQg+gykLKag3oxCw7CfyBOPJC7Fi7CFcZTA6VeYq/s7
xTKVHnpwS9c2awPNH00/ooTBbMLOk/7iv/mFY5jzLlNWaeReU3yLi1u72i14dc6siJeENGlfeZGa
TNvbHltqXqhOrQ9culQOnceJBFS9x1Q3fGok7AWbuk8AohqiT4AQH7iwIYrLB00yeZx2CmVdQpXE
rYtZozJqJrh+xeK+nRxIuY8qoati6sfWlz+B1QG/JoBTuwjk13J4Cw6QVnZvJQtYZEDIUleY/5Ze
JxKw09TBA4VyXo6PuvM6Qb8mbLsK1fN6Og9VZq00GeF8dydY5QpQ32/ybiFjIMQusc4wtm0Y0GLJ
iC9pQVG+135wwGsCVyqlxEbZMuTLDuLnmkrQyL8Zt7Mq/IF30X8gFPNh2oLbH9mDX4bi2Ux3r2MK
hKZ0ZDDJbvwoxnoNoUq2B9Y7zfsOXN+DO5KaBBfeQjTktFNIq3UVHfiucXRQgppw2Rreicczbo2Q
ZKK0e8WLqmIr0bNL7/8Bi/Hl1laMUYvVliXyP//YRmjnBwVbPgGqlIqRSqh6+H8jNgXgsuNw3kVw
t6zEK0nMR6IFlu8QXiCh2bQSMyKJfxDovqKI5FB5DZRJvS3jkwV/q96W+q8wwT/JpOIloy4/hgr8
S+lT0v6I+/I9bKj1ky0HXPPxFq/c4NbkyMxLu3RZV5FXSVnkfO8l1mJnTPvktc61tfUvXrbjNz0C
hEH7Zhkj/y1zoGDLZgwr4MQm+if46hxZZqyAlvZj3oFANoH0fc8yJ0KFXRTUkTagAy2CWEZd/CyT
4ALekhq4UZonZKp6ZPRDnAfS05El2mepEdVTfzOgPU/g9tAzfVJLF31cbmiUCJnOrWrc//dBunUQ
YHaQSGx0B0u1k6COXdMhJcCo+vL2GWazZAnjvX/mo7lBdZAIzQwCYraxRjLB2RP/iuuNFBiA+hi6
neQTtIkFngQjuGqUzIcVYOYgqGanzSF1a4jlvSKre2wBMPHw+49pny9Vr2VJYTLOlK3tLkKgK/tS
kK5YZsDD/e3xUuZjxr1t3sYtwHtL9uoUA8aiMuyN/HDBrluAgoSZz55Lhr7oNUeVpEfahOhBSUOW
b1zrRY/Z/swz3naT67PvfNKTwocGC07Telzfkb1XKVCKO2oLLFIVEUvoWhd2/86MICLWkia4kPaq
C12QxtJ77AZce3W7w+C0MTIxNmk+dodzKqqkSFkSR3yr7voW+CF8MIDlJKm44xp3GDNYiZWAlzOc
/uPKPOWuEfuyZEcPmghe8CcZXRoWg6f3LHsNuVe1SBHrkc8tvMeJzlQM5wyArJTlFJFNj9PS2an6
deFLJ3zTfDjpPXWpyz3Bgv5bvd+w96GHg10e2CgdXa5kxFYgW8l/g6MxVGj8eEk34XmFLK6RBjTo
MMvfBhzRk6iZpMyBGhE86I4wP5C+n5F5mJwiMuE9SvM+rxrZ0yyFG4kvQYO70IkOM5Xplu5t5FSU
t67B4uLsvz7pR0dC8xTd/ZRRMU1IU2HqfnQzpBNQC/IycpErmSbSyiijwTPf8t+PROGk7jHdIk9S
t8cXDtjeiKNDbXDXNnXH/Nr4TyMz9qpqstEuxXvqjyAGogiiQDbupWUzT8F5GMAQb7KWZIUeX/Ew
5GJPOiP5a/pZ4D/YdzWc0tQZTqmsJI2pj165eZO+yf/SvhRGN72k8v8ZhZYGkDMfJB+rnMa/oNJ0
KVG+P5JeiXGzyCVmbsLyMgyn5JEcJ6CRhkEtaP0DwqnazVXWv2ir9X8ZPm4r3+E4ipN7MFCQaFgi
Oc30RkzIWCGVIUhzfOINI1YdDVZxObcJA/kISgBTXWo7f6GiYImw4I6lZjSagfcQoGgDSAoEh80e
khaYxveKjElHe4vS6kcXb1SjikKROyoGIz0h+4g38OwWaJNb6s2hJGgyGPQ6e0IN4HfqWUFfmVtP
KwnSZ4Wlnbbwg6KCM2UjHoVPSiDdJWnCHB59bphY0qtXv4RgVLsVegj/HTN4DySP7iR//UA4x2pC
ntD5hXa9PdjHpyNnZ4Kj8vDtcGQ+uyVVIzz9vQdIHF3M4fET+OmP1pkq/6/aPOL44ORHpB3WxULC
JN2LsalWvyHZsQQkZk/8mRkUObQm/nMy2aFvLk6rigbbed/+JUdzNeuMG6J3V+T5wSa774qtfE/E
tFaxUkyEFK2jN+FCJFtHa1AH7re/f1t8h+H4QBjzY4oVZe02Rxn7r3E3v8jrMzS1JXXq8sxXm9k0
uC7Uu2IG/K1JrOVF/qBpyKuRUWxQhT+CoFPpVITz+iXtDrQqi/utdW/yY3zoblgtcTwANgHJiHoZ
J2chwaVJHMCkd1vdxvBZkYObQD98WN68ZFXKgMf7H9Dssg20jCLoLUJy6iXyZ6zMudfwIGWbcbLy
Qj1M8n0ZJi2bZTl+P7/n65k6nJ8BBTbPvpemdhXLhEQnyfVGwhbAodqNuUL0p650cI1rraP5YcCa
0VhPt2fh1YttRYNK/NYfGDPF5DOyEl2HB970v08nrF3SHbtr+sT5f+C72Lbk/+brvjYQb+XX6t+N
e7dpTm2wMj9XlvKvVIcpul9nGcPiDz2W/a4BbsdXHfcdgJd4AGdvcorEFrASe7jRR0yv5Fs5hPTl
YZx6IN01N5CAWU6pbuZGhI1Qbx2QzlJ2dm5tkVTaH3a0JQspEkI27HCSVCtUr18keP/k7nWr+RA+
chEWVkh0pFfC7TKpCICxjM4qjL0TqJ7GwJPFc9IzUA06nrz2GCRk3PREf2xthoKQVW/Re4VA9AD6
Qf51w4mh3zsgiqfbESXyPTVj/cReUNDOfF37BOk5W4kxyjG+u8IhUXD1ShMbnKv9JNM8WiZ31pEI
xw+HCJuXXqAAPgZiByq9N9T3IMkiHAyfqG25pp6X1AODyxVcGtsF6S0AztydnDu+jyjUn6lgLSzY
JP78qLSjdrrYNm+hmxp4Zc09VcoT+6WdQlzCdE6j46EZPHfw+f8qyrOzDmDev34lrUqfsJg7nfN2
8Yc8gsLCp6HbpedM9f/vHDzFMLJqeRl2Wy+/olkPrQYsUkVXRbHdJv7RYJfxrz/RIs+TjnAYD7TC
ojaGzdKA1T09BmSty5I2D++dFxigZbrUMxLEIlfmH5FSfhizkGVhW2yEPuRktuKfpC9kPP/ih5Hv
Q0spZCoMbkkP1Jgbt3XT1IcK4pXUpfAv+ubsObLLPEjzXXN0oLOJXgt92d31mrN8kUltO4Y5hEsy
RhTNNWAwN+GgGXdKcphUDCzraQa57cXSQc+WlLFW3gO1h+hoV7XHs1ff6PUJgqyD2LzHiuWs/+xI
5EgTXZHirYrLUj4CSaaXArDyveMMrNkPyRc18OEDTXnDfAjFJDgWo8Pm7Te5LiucIQCsRjq+ZN9b
asErYTvVefDgu/avjf8n0WGawHxAaQXrttzE+Uur1dfmYmyDcXIcGakR3qQI3eOYEG6ToI0M2gBd
OEiYp9dfB9mUDOpDlrs3YyyrrRtoh6DAglrQKnmgUtkL99pnzWGgW3AWa++v4wUkmviEqtnShubG
EIe2nWlOlOvNTxnd8lLrkiSGvceWfUK4jWnt0mijsEF7oiOrITps8xqcNLn+xsGoInNywgo/7UAU
A82rDkKUhXcfOHUBPCxpSNZ3HnPQzqUFhannNfVCrn07l6A4xiAOPIQcJlzp0REAqYw+nXEjovnJ
B4Zip3jdRuWy8xeLgoLZ/mWCbf2tyKb5dGt1Oal6mBUcYwdZZnwWInhUtiu6uYe5pTrHFn/26eHh
Rk6el5pCIBhBV1M2yQNSLMrKESEwIc24x+r+TiIRMlesV/kdCdk/LeWfeUd5C6IX/457HgHWgv/d
hseRuRK7h3VcNNvJtknOlDQKvbnaRwro7d0vlSBtOeUPwwNlhR1hu6iqHmOnh1LrrHgs6E4myzXI
z6ZoPvlcGoNk/koxuFHAYcuvyXJN4LGPv6EKQjEP5z1gRlJlGIgvn1XqSJxMpdY6B9pUnZuqxgXd
YbAXyOkPFSQ42WjCq6HmZG78Rf+TP9gKpM/dsQyuc9I4cHi2ufqF2ragoCC+RdMiMM7/OBTvH6eh
mw+MTihsuMFXo+OVRd8T3meLF5Wnbr8JrbgIJodtiP/qleJJnW6g6otc58yWnO1Hh5OtBOA4zrJ7
QvugEy4IzHCmprAu43jiG6cSHC7AHVZ+0X0CopGn12DS9xT6o8sH281s+Nb8jaFwof/weUdJSg3m
TuNlgFgxnzlRvlK1pzJPvPL54bM1ZDSiwal2pF6UUVR19lPQ7PQPMm7OAVpw9nZMtSwAm77CV33s
wY+Yp22eCvwJy0rP9bVukrWcgDGpfT+qDCzoyuqFBnLDd/p1he1UICfOObUap3w/BizW5094Q2ef
17VwHZuyqfvZhcaXxaJTPRa/A9oHCjhccGCaFrmRGEHaLV3gPqlPyIuWp4+/UyL6d5S+njks/bxx
gyRq/xfyv29jPyvr8kLGkA6Ulj3YE40wGzIgNg1DzwJQkQDL8nqutlF31JkoWl1nWrwExZoIU6VR
cA2pK/Ldi1mw1mIjDgyMWBXNWQJkZWF3Pq2Lgx8e74yW8CHwRF+QEAnC+bWw63fhqFY7v48AsaMc
Feo5+y2/9Xmkvm5Ijvt6dpeu7dnI3ZO20AH9y3kUghA+ANswVVonj/wwaZGiw6R5L4IIfj/mixi4
l6+79UsMofscD1/LJaoIsbmGfNAaazVLzYrw3ZqfO710PTHcm9TRyYjFuUpf1KMui9NZGGMmzOlv
VUv0TQkroiYu3j5CaFox1tVIQZgxwyLZz1KHvaXRjpL9gRpQKCf11szbDTcmz0exfPNBnwnvWp8b
s0MmURyXwQxrqSg+xmssV72g7dpo7u7uc54lU9SI/oq2hwVLgXYqHnJfCbI5VQJdZr53arS7zgTV
FIT4GIozMWipOlbFRBSqw5SmPfEd95IHOFuF6lu8O2an5YOyUTaGy69EL3FAzQcXkQRjxtxkhv+X
KaY9rwRrBYq6CVczoozEB/8QOy88z7/flvhvcWA6x/u2FtFlTCC1eTWiYukA4bO/AhRRNX0ax6yI
DmX5XFJo1dmaQw9Z5A/SFYOgn5cCfov/eF5o40d07rGZY5JM61ePrx0w1WE6qrQTH3mFTvuU5vmd
LA1MNS2plMJ0S/KggAv6ID7MazMYOLcZrHC4cM26KUl3Q0G/bexMmP8ezpzUv4UyHXHs3C0FCr3s
u8u+ojI5le787PMojukcOvYw+YgSPTC+G9HwCp+FsAhgD0q6FhljxgD0vQSbzEFNwBltLoyuvf21
Rkk+Y8taoZmGexA5+i9ZnxrCuO99+1S4Qhhk0PvcQInbcXA1pODsZqweczM+G5ru73Q0r2oWLWUY
5sp5Eamyu0CK10VDTeGvVr5O0k0oDSVX+nRvKqn36AWlHN2yR+43Jdnrz3OXGPswLddiAehl4Wc0
0pqSOLswyfQMj1og+Be02B7RC6qXYtHALgFRp8+Z+fQTzysDmBC8l1nRgzVIY3XZTt0ohpSXJ9lZ
Mset6ylaAiNzsZ2wpyIn6bTVPzkzMZ6BvCityV2Wh2W87hqaSfl2gQ/x2vvDs0zmEil2AaQiPbzB
DcjVg/thEKEm8pWNYxI+Jr4Q/p36RCOAEl0V/BM31jHHDPtJqJCHeEWXvkW8gTpbMqHsMzcmWPMO
exDRF0/cv3ij5tiuSxcELtP9oJSLA1nVuG981YcRV0O2S1EUeo2R4JGEPqSr90SLkXVXsW3uEpBM
xJzloFUsF0FWv+5ffuMq7nN6NIAJiMdvyrNquZPvtzLctJsqu8D5fLdyZTCSAmP/cVZ18xPh+Yai
OPZgJlBKqStqHxRYaTcJZ+k8KGMkIM90pk4utTBdYVNU94k0+8YH8Z6OldIILCWAbXpogobDIxKf
DybtCmm4JzoFP3gv2vFDzst9YBsG+OhbVtJeloMPAAmYzAtwKlCDim6nNTkI52VYkAJtNsEF3jso
4eAdJcffww+CjxOrE3YoBWxwDl9uFz6rf+v5qWEJJXhQ6AAmVwNo9XDk+gVCjQz3eGZJuHqDiYIo
aQkwDlVbOYk2i4XncgA81/L1ycW+fSAq0z+pjHELXnPqPCcofJF+tQsk8vZ3rlv40xJFalNfhmlZ
3BEFdyGhoARMZ0xEFlbbIkzAkFvy8dgH4DWZLtluRPupAbhtRLoD1iyEpUyE3bB1PfkiDSrYE+Bp
yDPV3DklrUxcrXLiAav7rtUd/I7cLzlhNsnQ9PUIEl/ElYCbHKi+Syile91DkMqur1tyjhwmaTyC
5M6EUJ/mUb0CVSjMCmryUMuSG6MGBD/A91ZLdT3ohpmf1mPPC1E1305xy+1qybd5at24sTkzKtIn
lc5afaacV3+IrgEoXQpQLvMhNJP60orHPbvjBRjJ1i1lmol5KSKVsZ61c5kEW0nJE3jbZZQ1ZiId
meunW/HIyOxeRv+vnBVJPzQ4jNKT6LFdJ2++iCQFIQWqd3jCt9qwEwFIjgbMggUaBdxpxorWpkJK
ZP5m78vpnNJa7xt1zDhXSDCILV6BsRF7f73BcZesgQVtU0D1+NSyfz/ixBjTtGjXn09OrBEGK13W
hbLBsN0hpcwW3ZK0aDoCbmkn6E+WT3Jg4SgWC2ojfrbqDdonHOXuAwUO4a55ri4eB66Nyp0W8BuZ
XeeehQGfWrCAtMrEyL1VhLDlWbC8YOijbo/6d7nUSdco6jUV+Cka+tEEQ2YD3ere9V5p1hU8Hgy1
VAsfAUDcFTIGWYMdB0a7MvvcLm0haFGgOoKeLaev8/qek9L6sh+HyS6tRizjkHDY0kwGhfBa60fz
rNsGXMyFqPRcmIqKkEL3lZgynognBoel/8vVL0nOE4EJUVimNrD2AHDXg45eYUPR008/9Pya74TU
CuBdJrpFWAtv8+SPkgMUIReqZ+iIy3hFTWThf67g9U7aiVuYQmUf090NXOkRIUkAfPvUNINrjxAO
b2riItAe/2n5OqSSpLtVpUOeGXo1qmWtTkjYwlgGJgr4eWdXpAb0Pnz1U9fmzzaDxMCDeRwDtlCl
gmwoBsokHLlwBnxYfjqpltndnpFmimWYhNxv+wGeZ50JeLJEqQcy0qFIvn9Jxl7KtVMAJnqZIUVl
z1yZ4e3CeZ+RZBx56RXG3/BinyP/a5uGFZjTKib/vzeoERdybmXytdsqb23FgcyInIM4M82zXHHx
dApWSMy+dmQLUJbRYpqrZE4+Lg8Il9hF5n+49nOUpC9e1nexG3mxgGKI+Pw4Qi5+FDIDBqYe8JwE
eZwuFPNjF58cdj+ik4+P5KhATKx+MWd4yWRNP4lB2dhJQq6fFXXH2Y7T+fmYINzT0/+GmuSXXQPV
VtQcRQSSkCff3TXQggIbq5BYp8eu0aGVAYQTCOHkitkYPilovpgdoQPWCY2Sr3/BOzFz8Spb1sNW
OvpxjWbiFEBkqUXmi5GFyOIGiSqNy5Dc2Bjc4TiselYy9x2FDifm6OZ48GcvriZNx7xkMY0CT+nB
4x76AV2Y1IB8K/EsWezAcDoUDQBIceGTg4j9uz7LSnyN57WvdqeRhvOsAG7AX33gruhxFwgPaJNW
rx3cd7kKeQiM3nVu6j6ucE54Pw2otfj2jiJN9wgCzn+Mhm5fQRAc09fpEn09NxrAr5gi0o7Yqrmw
V0IgY9ozHwBBwtwsPl/sC2bqnU8c+NOEtoLuZLmzyTb9GaVouPNtS2yAm7WPRMbwU/+KXFH8TufB
reUdKyZmQ1OsM1VU596rTpZQ4GrVYVfFp/7i6Je4K3SCpI24gBbJAJ8qwLYWoyegRcNHMB4CjYTO
usTBn0n2U6qLNDplB09Uo58baC6V9NKFhmLVy4qb7fo/xYlskE7CbrabcTKifxep7WfSguFBn6Uk
+wVOwAo9zV+sd9mark4ODgWw/gP7iZu5hyROiDDTl+qfrTUSiUH6Q4AYvsip+8ouCV5qH9TOnr/O
AdcO2BNePiSmm5i0a1Ykofpq6k0T8XEJ6Q/IQvcj0MpqiPmqGTjF0rlkVrOh14VO837MAjn2j7X5
wz/GJGmKJD5jBsl6QXoTQ0MIic7fzz2U8cDtT0FzKufW58SPubD5Hy9bQeOy8JPhGgqQ12LGcctK
f2allFppHee8zqguTBbfWo8RNugNVYHrAU4JYnBa/eipnOFdj7XZAd1bRr11NYK1ufnhEDinmYK1
50xCR+EwMDO9STpTxZFGLR0FeTouThc+nI7x2QFZ0R1bmN/5xV6062a9n3WYq8J/fkFIgVePozjO
nh+TPUeUxtE4f35ujvfwnM3GfWLVnevwmu5VgGWADgpZUgnrOzk/kvCtGWLcV7kIBjecWt8Eceqf
UbiuojdMomhDDfD/4FhGtvCUIaNghOZ/rWR3Xl4r81o/glMLOiz+bYeg1DelzqvMrc3URZO8rU0r
7yC9/XqT45WcHQYqB51bggkzN03dasE3x/ekaKGmDUiNDYSUpktlMobSRX1sVkWgj4jFNnQbAZ3m
SfGAtmHXt1ad3qgoO83eR6T3AzcjWSvFvmCLNmqX3It7FeGLB8gcLyMXe65DEwDSYtCVHo6PyUIT
eEdaCXhsiBCarqiXgICg6TxeSLXFsdaL2KxDNike10QglidBNTLXcupAdiMl4xbaW8cm/NRzo2iZ
9MbGXg+qY2fk0S3dOgFCeNmYOV/NsMX1Z4NQuzVuTUsrmN4VJIwwWDMIHd5yEoSCYry9/LUigrBR
ybe6oz7+pP1TiW/Ox/xllNek8Tm09XN9vmr+jkDwrcL7GjEk9CR1rfz76NIwqtGT/D/zgvvEo8i6
V76OrNJnvxM9SWRc9dgLIi6IgpjW63sVtaqKEn7Z8b5aplShQKX9xVbSEp8wCPQEZ+3s+Kqf35Cx
rTj4HeXml2di7dqgGj7zSM/RPNZMikpml7gRaVPV+EnOHHHq59yojew8hc1rNW71A6+0FuyZI1Bg
WREDCTE0CK1HRyX4fWea5QkWZlyPO1afiuHR8GHaFP+pqoHroLyHJ8a7AFL4zOxSVZzoPh7cLGEk
2s8eL94p93U2M9esIV41wXMplGBCNvhPDJtNwgggFz9E8Kven/BXidYWp0LSa2aRgRuQOMsMm3ly
r5R7LRBtoqU2q0KOl/JDG5BGYHiI5bdxvThnno9CzPvEI0OlGT1eoDycmSeoVCOYnBIKLq9mWggg
hPyy5cuntDcO4pHI2DaE3JVZ7NzanliZywumDfkqsNTIVYX0nxRqxRG4EvleaZQoR/p6eYjgAtDV
z4L/jD1zTCnWFKWqkXyq9NqSU851XyP7QG8G6uzoYLNXTEysiDxdPW8MITHxPCwQ1GCC2W/JBwvr
+betVtq3t/LuG7yCLU+hZe/g4pdKUEHEs21rHvzU0KiZpld562Y0Xa1yLEydPslqbLO1bbnt0nPX
a/jnOAoflPvfbXxNr38n07Tpit1X+MGmJiR3LWBNRvJ3kra1hVahiVE8/sKjkXbrMvEZ00p0oWkA
FomaBdJI6z1UaYD2RPXEL0BCmbmW0K5KEalKV9cpXC93dFmB2a0kvfxBKob0hVp70HyPAIVMosA/
GIoWaeQWM6KqvO9QAAUpOgXiovG2Rd3MjbXNyWGNHGT7j+/sKvcg+xXFPD80yWByHY49ZN6HxT4A
I9M30px5Ybby+EJe+ga4GI6G8kHppVDsMOsLJs5pGoKWU/60zVWjdwTJIiTBODIoM1hs7CirGPbb
wW43QYD1Qs+01ruktos38PtQ1Ul0hQ9il/oOeX8UjdxZunPNFnz/qFzTtxIikPiLRU+8RguQtVQ2
OYJtCoe/AtSMIIAkv4xOcW9LyrDopf00E5SyKovsgTfMiuuQDi1UEDoDIG38EuWa4CXBa4z04Meq
kCIJNvV+xJ7sLFbo4xEDxKfKhqtzlp5W+MYr4CLsMhhhUI+rbboL0s0z8dO8ZdGyAzvteT5XayLv
WglxnwyP2Fx3BXtSEjgdGGc02rau9x6SJ+3YLk7Ja1lpjc/XG729qpd62Iqcs1m74o6/tfIjYZ9A
b3tBbPgeNpdAJKCKCc5RBlGQwCefs/eLukKNgO8vZfx2E79mBtUAfV4vJijI6BqMrGo0Va17/kt7
0Pk+XFV38hD5IQqeSO4LgxhrujKEbbGcjPRPsDOZ1JhlXK99HawG7xHewVVHHOYChhbJMWDb4xHs
KKkRVq57BbuGJ+KM2jjoRP2d5TYVTLi11Xgx4I3vDTY8Wqvz6NqCXE4EiTsaydUhtanmp7aREiX4
K5+CiG9DUH14J5qb2QSfCga8uIzGsNGmqoHLfLLEbGIkg2CRhQ6dbwNRIhRTYnzVLKvLFc9YsyJl
DjxlxUHt02nCe6aacUPi6Ve6Gqs5lZFEWJBINSx6ybNJw++fTQRzaHZAiP0bxRyewwJJQ5YX6kL7
jC9E6d0GP7C0dCgT8XHXlz25Ytuc/JR5/mwq+lHy9cmaRG/Te6F2fxb8WxJ/wQI6277HCU4dlp4S
6IdxzSydBXC/xu5VwuKDbC/ORM+Vo/Y8+Skz1X9TLfrK7YlYOxT60JaYaTCU5+7jtRCbZmcUWcIi
p5CyR8pssaXF+eoQ6nbz231lS6md1FCBVxTrJL+Xu2Xlg7z+Yd7UX3zOImQ8EiH8f/K9wZ8sODqx
qK7sd5LmhiglzVD+wMzHBdrKp7mZsFJk5uxsJJYf1cqi67FTAtWld8tVMjzxf0qNEDXYu8J730Qe
uj6txdv7vXJhIfAwcn8PCZXW1b3tEgaJzXQG0IFLwPD45gXR71uzlJ701J353EvBQgZoKFsJZiub
6+3Ntrhg9N11MDcHCkVy7TbMWCmuejBvX4X9p5+VU6nIvkE+2bwoSv5czwRrK46UUCqszmJ4aEi3
kLuKfJbReaIKLBi0ZFaHWBW6r8gQQgzOmQXmEffid0B9OjuIRiIWacctcYr+DjWhbDUzrRQQuBeu
CSro6ovp3s7Ez+fwuZvrumSpzx6KXDC+xUZXBOboUOMH0BHEQnJDbQ8aXeBKBEuPHfr2PbzsOZiU
39h8meeBPen3d2VfcD/eeNb4Y720lupHZ9qHkSgXCjFtSBGWf8gTK+8C8KFmrjO6TH34d2CsNL67
jxP+iQsaH682IVZI4hWdPAdfR+Nc90Lnp/rYQQEAcFIXz98cPfhcBleDYtm1fUbY9imFuj+WjWYk
VEb8shSCV2itXe9jdXPTWpOW9zL/j/1briIwaDHZAV4c0sfQRd8ar9a8kKgW/0Y27CF25ckcKKRn
nMbXtGt1jHpYX/IzhxSPOm+Dk359YBp8/E1F/mDItwPvzi0JVDJ+lRk4rPTXzzUdqR6T+A8gvGhS
dGJ3lmL4bZ1WoPuWBuUrDQiyCElI6/UXd9rNlTKdR71apLpYhy4Vj+wjTmRmZtm2xpkCLQq1k/rB
v6gtIoNhn9WNe30YqZsSJyUrmiXl3CRn9XUGIlykN3e/uKGKNFK0x6eMqXHCzQ3pRiouRbOnHG9k
1lvSs2LzTmpAUGwYF7qY93Jhc0KNa/zrfmzPSqPgMlAX5rlsDG52+3k6DOane/fegxC2U3yhQoA7
zQEIlUXX+paTgJuhkIgP53flMC42muimnBCYGCdp2Drr3eyBZNIIYVlVAgiWwTdoC0KgIhYX5ME5
e9nzAsisdKyZQRZe6mdmxzxKMYsmNTe+vE9ju4aZhF8+cTQFpoqPl4Q9lD/0ekO/WXBMgKzFITbj
79pCPd72lzJUmnFMnwryni2NziASgS8zPP5+rbswbM2fqvO9/a2tq5umnKrvp78w9SWvHOpqd856
cIhkMQcKt1/6irARRWDyuZCq+oVLSBdkEA6ejyzDH/Qyx5rMwL0qttYlYd3KOChvEpay8Af2yN91
F/8Gj9zPwh59rgtpU2TtsLiE5MrVL2fxtMU9UvOEdB4wtxXFSUC3yDxHfFvqbBYgxLbEfgzF7xWl
LnHrnvi4UYF2Nyic9UEK0HNI9lD8TL0IAQxnhID0PahtnOgQHYVFTVHb3z9U03UOoinkUJ6qtJPq
4+K7oAiLzl0yelqw/aopEmI1cLFgsxJZQ/O3AFVzpwfslePIeBiu6jHNc36a8yaKDgd98DACuxfU
SPSWDajv9shYX1ut9o+/NXzHAogW3J/IdldclZq2J1MplEk2Qztucdwhk6HLNmFgYz+SUnKZ2MD8
+SPLtcBhd8JJVxKJGyB97+F4XffCazQwrD9OFGdP9ihnK8kPJ29joS/skX5ICusc0l1mggvibHKX
UFkPPAB1dMo5/aLkTtOTi6lq7bmnTy1YdYHkVIjyxm04tYtEk03ti7QBMLPNdglqQiZl5+HjHEtD
V6bX8WM9ldWToYcS8+ZbB+zK1t5umkPjxrnmt+itYycG0GwtYzkYxBL3DHsCSsap66v143w/Ion/
YTjwQq8/zqQhdfgjpNv5TnGxUvptrbKR/OMpl/RIegUtH25Q9xB450HOFSmDnt4m136h91/kef5O
UlXWghfTXZQAg6ypC/H9Ru8Swz56TikXQkh3M9hIW2mYwRQLWepx0Q0nx7+xVnjPFlzUnbY1f5Uc
m8Cg+PAJXAW7tA46NA0DSGbwLIEhn5qn21epqJrqNDhcZ8NRXjHjbaJNVZOfpU9J1ySftrr7NsWK
AfPvWysPMFlsh5JhgR5qGImYLZ5VZEVP5CClY5ihDdrO3tvUtrnQwX0IaXIY0o9a5VGUB3jXlmAy
XxFG18PEJpAEaumDjvBynvPbfE1oKG2vnqMzQ30kKRq4WQaK0ucgkxrDqDSe6BYrCkjfQvIlnw/R
BVj+iu9k4ctqnM16vc3LfOxiScAdZsNORCfIZuckoKtTC8wYhPs0ZrvA7iJApn3i6CZNJAXIKSIp
9t5DgJSeC0KqGHEuuF6TXo9SbHh9SAyq/+rzlaGIvSgbKrV/9DONKTpWyD6rvero3X06Za7t6yaJ
/LQn0/biaP5Pe0CetPUqO+2QhyDFMWQ/4ohAzcNnPcVSmIE9C/QN0W1LlDMtbS5fgpZsTLtdx8lL
yAlV1uyJd2GgvgauhnoCuJOjMqUYNNdXhUmxN3+hr3hdjjYuV7pMt3KZFHG3IUHT8LDUCySnVosj
pBIuF72SyOwfBBuajA8XXuoTB5y5C+LowBVVQr8UJETQdbAR7AbOOmSPtSr5YCssiMAm3jhUrsZo
dd/TvIvUfo4QzK4Jvh52UNA00+Phw3f1Ww/0ZbfWA64i/+uvC2/zcg1/wt8eEcl1lTc5oC6Drovb
7FjACVzQes1np9DTYfw84xoxopUs4SDCff6JwK9dDfvkOqUPnSgJpWz1kdzIoW5PfE9DQUw7yCO7
t0J31cpvyKGpHSRNRdnkPWxx/aDPTBoIRmzY5hp5i6qsas05HoqYy6vSXjv0dll2oLdOoqodml9J
PeoOWBmq8+JZSfJksioLwQHxoifvllZplcuao4Maiya3hxfigVqRVOUBzDBmZZsgPn7Pr7x8W42G
QLyUjjc1w+pGsYMeyNsTERL/Ul1HPqYeGBLVCHHLAmsgIPavQZPXFSEhwl/2KWD4mToZv41OjVsX
2bBHn4tMrS9xUfQQBbuhCfPhkTuMatu0t+WTRijy+mnfyC0n0eO6eqnoPTn0cf51iW8VkhFUVcai
gScnDpb+0HPIL5fQrHgExFtYxsww2PbsVigwS9a6ytZ02Nm9psSAOpj/XX3vvUxDMCdqi2lC0IIN
NPvt47j42RZsnW/bt9TjQCksRsbsRtRHVhMm/B6riDO5Kvd2MrIJWkF6eHqRWCiewYKdVGPEjKx4
7hLaacTiFdq+IY09qjv8maOwhkQ/vRBwfr4BT1FZEUIQLf+gEVQZOJW1pEn5yIEJ5l0XTZYA64fY
HGqgWKGVPc4txzyVQMvG6CWHXghIiSfxZWshbun1anlRPiKvHERw2Nl9ufxhjnUTwbbZrpJZ2lNy
913PDl7gxwQlWHAJqdQNUA0D+j7B96jXcIJ4gR8QgS6je4TF02Y4ZWFRifFjJN/mQ9iW8z/X9KEH
pw7gjLcsUH0sP6RcmR3ze+0LQCGRGsXMrL/xf+zNJPUa1R+8MZrMEvxI2ZiVzmqxzjK0qIOTZC1o
xE1f+N6LPpTXwsryZnj2w6so4sR3T1wzei/O27WGPkQ35nDJ4I34sKt4rMLFP4HQg0GxWVa90wY1
dI6TG0V5CsP9kMKk04mSMCB7diC+flFSVos8XPr6/aw274yUi7mf6ZJZonsQ4o9k68gTt+zOAzKA
ezJpiI8sPFRQcgyyhhpv/KLUOcwtSrnaFKR4YTJlkwbbpy6b1rM3VIli79Y6d4hHtXOra+oFvKjt
qz9MX+0MBWkxm/1KmeXzR1Eq1NQTJdpSZZUUCtFjCsvIpxMrAgtESMv/H3U0LLpkC+4pS49eKAFB
dmV4iqXd2NIcxwrFIESE83Bpgnf5WvQpZi4rkrii9BQXwvbWJ7YYW7WPzSIsB0HIWmzLUO8EWJoq
CcdiSCOYJAHWk3cH+Cxe+YhGBRrg0BAcYL4WkjdBRuicjLFN3jUi2LZkODrVHIIP04c7JTwnio3w
/tsUPzJSOxjmxMY6VADoZ9dKXr1iTVycbn3CYpLWW9gCT5ob8KdTcaId2vYdJDcR2g0bePaTymUG
w31bs/aMVO57+CaNJPhYGgGappaoJMW4nOfuTAVu6Oj0sijugMqei0RAxP5IIl5wU+BGIN3Y32VB
W3Jq2CeNPLPMt+Yh9hmkgAazqyY24Omf2mZ6PLdovnytJ9TZq1mfefguqxnaNlg1k1lcVhGK5r1L
5tPo1WG/DsWvjffwMFGDvjlGAXAQG27tY0/9FH9qpm39fhZyfMqjzOakFGD8Bkii1nRxyfi4BZ+F
Znf5+DZdJi1+Y9MBMZJ9nsH2XNQsOWhljkclVRCGzB6CP+MBaUb6YbVSfIVGrn+S7tQpkFEMnDfE
CfY5TuEbeHdK+C3EXpawZubev0BchQokLsw2ZpGJG+vA8u1mpVprGZCIQR4WmEFu5OmTlxj0sH4h
W43xW5QBWvtxrFBQP8a9ERj7fQntVVIdx1U00mny1B6iQ9DoXvSBW4xkr4vbBkKMYw8iKKuccbwF
OdS1P1jLSZxmher+UX364G+ZYMu+njQWEUmGLpvP/aaKOhCP8oxPVq4LTpVBgeMQ/RpHJeCOCNnq
y1jpfFKJ/+Dpov1R1bhTkFUA1P8bQEfebOwykyIuB+Wm+n9gMXhWfpQDlNN8ey8WSJiS6+0q2tRu
43SDOitEDQzd/B7dppYNXE6rfkuFI1RHAZVa0zptW+PAygV58a5EbMKnRDe4NNKRosJjadP3jBS7
0p0QkXTFdJDTgDzrVzG44qnsjM0NJuOxwb3LlI39Gc9Di0SBKdb3CdqmzsRUsE0j7Y4hwDkbLuSy
hOn2jq/+MrQZ5H3YEr56EEDsQcnrzfg2BGZ7mBIHAMqf5nqI/RnxiUO9BoMwXMB/Eeb02SUDnCSj
0nBwAtY2RXiM2VVEUC+IHuL3Wj65YaBQWv5nvGX6V8L+NXLOUu/S0Q8QEIjbz/iInyBCuAQaeSdv
Tiq22Qj+tqw7RX7A0NAxqMiX4FTTgw7jK+y+7fu1Jc2K6c9ZK2/gsy1HAHSMoM/JjvKS1V9zgssf
K1NZZSj8W71gR7Kxdz4OAlcVDJBBgm71PcHQffYvrBLl5XvB0Rp27SqhiWOpHRL/WtDNl0cFbO9D
hjNTQxiLsEZKcsUv06NMCaNl4cQVrryuVeVsgIYK/QbJr8LPJHSN9XBzxKz7JBW1qILQGAxc3Ye9
x0blSwLYG4a5pZNapB5Z1iEOh/BAioydEdu8oExMFYPs39UkPsmvdIvBTEC9u1KGxNFt4jAJL+K5
vRxC2QpdjB0MXhRkKuPfIxdNwiX1lqz4Mon/cFCTInRFA6Yer/D4460/o7BZmEZd8Vc546ZldRv+
/Xb8wjzCY/r59y4iUq+QeuORGdCp375qAEmSKqc6OqP453jbiuO3PdyliXnQWnTTF0sWeozNnVrF
VFa0PH9YOsRm4935NZCozqmK5EqoW8hXgCt9TzwJt10aOfpn3tpDnjgG2vYCNyM8zTSC1tXOqXzs
yeUUEPwmKiiWQzSiNQGnd2xyHcgzKepYPK/pnbLyDKFUx0KDkUhn+D6MFY7gvemuzMMYH3YO6M8Z
bCa/b/lK7Xu3NAsUfnvPt7l9OIsxIomKfUARIn/2cBPJ7xUIWOsXVkXn7cZche0r0aRH+DKctGE+
qPhrgiiPVHcj7mqVnPmbHoEIwfBxNse/dsm50K2zech4RSBo25jfLrMHZFg9gVTEturZytdc5sz4
i45G7keTfOUb3GHlsqPxuRtwfsoSjvEGy9AQDhdjIzcSjGcmD7cGTq1Y9GHxabAtzTGlyemiClnC
RzsvFgeNx/gEq10gBw2Ylu8Sj7bPOTnhaSLRr5as45tm0j7MBZOqRuvlYrlsYy5RPBCKbzGvxP4z
zxEuTe6PqkTn15Y9+NGq0E2yBs0vk14d9pDfenimN3m5q3mw4IQroa10IaVzfSUK9MEWoBQJN/tM
StGjkmqYCtesUvxn+XoWw5yIm0rtWxZivRXXswpADhOg6YjQ4QwPS5ZPGzeE9VP34xGdV+SAfIID
eRcqQhxOxbv/D7+eaP/+qORuSPueEszrCbvj+YWWBYEHS/msL58LYeVI2vxEVDQroTNlOz2FEUuR
LSMOYkjgK3jxNVpOIZ8DnItjHaLqBit4rOYaY+ltBAH5m41nNq9UuCk/y8ZpW1XcDx1GAhMK/w7i
rGYzBo/02zIS+FZXxZ60e1rlonAm4tkkLLp8KtL9l+DXKnHHCMYIerFBPozuLBeauctpq5MDKUlB
nQBsTLJ1RxO6zdhcJ2+SjONfsrdV7AAuCdlH5EbeBDzsEFIOPbLBAR031pSgwlCUKPi7YHhPolZy
iaiY/zYAsTXb0U6SrDv0E92kIxHSrn0mZBrjXc3tSlMHuvCTg8AgPy4gbzHfRhsaZEo8wUZwwMeD
aFAgxFP2i5ob2zvv8ROz7PzMwFdcyve+bcm8zG/l44fhKTEA7M30CrWqbwzQSw+WwS0hEibi3gPl
VVhY0oFyer8jXB6kEKfIwvidAnM/2DUSq2aog80iCkjQQILRpbs69XR727jKRssGEMIqybwkwDUo
180YqixEr12bLlIOqGtrg/X8PxmmMYoHNapiodgShapGUWui/x/nnZMwDZxxq61vtJ00bDyTIlds
HBslJMnqMB70ThpwBSf1w4Pmsp8GdWteMWBDAtChum8hNPfNpHFpf0dhXo6Bi14CERprj1hkMpxs
wdvvvUbmLJt0pS+kRoNj2bCUdH55jwKlp9gwrBM70WrRHI0fAkyIxqVt9GIHGZq/Z4WiBcR5+TsO
jfRGqgqni5nUR3paAvqYZxIn+yHqCa1gD88QmFKIqiFLzB23qpLszkwg+Vgycw7rq6hGAkeFeAEk
2CVQBcDSzLwAN0l1PBsW0+ggkGcN12+kuquxgCbv0B0LteYz58NZXmGfyDbwUXWZGbmHHjhtb5uk
MdUqEa6g2cym7GvlTcYUfO9OsMGFaOyYzOIFVmJpwwoIa5uxVEEU5UoznI9HPHMWBP9oC/fsuJGt
vo9QelAHnjTd9jsi/rQAouCnKJZ4P1fpwap/qTGdEBctQ1075ZesyxR9s2Mg/okwpLZ+PG+wEy9D
N1XDh/81lx47rQVRbS3m5KPyxl2Yjof0dMsVd3/Wu48XcNzdOhEAY7gEYkLYiwAGtbFb22T51eWC
QsbA8dQ35ZcBZjvuHQ0Jwe1v4i3kj+9HUGmjFfqRqrmUEEaC8LcGi1isv4R6vpdfiSbu+6ejyeb7
qID2gghNbOlJnFQjKc5l/+mlBmZV4I2C7OAbNJwQM1CFHe7QzHrKFUHuapOTg3TXpelR7kuEeNti
Sog4/eWxa5VMXbMmVaOoJ+dtkcMr39X8yq60vAcB3LoEiavbxCLGJZVEoZX5oyV6tGE8TPKapHfZ
V6QnCAq3ghB88+OFgrwv7/tw35YKn3zZhBFPdyrjXrcdmcEuU0W6zYdl22+Fh34CZG3STfCd+7ZD
M89HcH0ErO3oQlYVxKM/10c/0agrzp1ge8y1wFg9QlTc6bVWs0WG/5q7QbWarZXCBGxxM1BCUleo
NujG0nY5xNlx5yXJdOj4bfbgMpCqOFLdBIVUp8RMyFvSoOvc5VQr5Dlaq3yQjLCFyf5tTXCISWkJ
sEdAG5PWfgQCJAR2LLjqZnPuWj88SQ/8fPkRunXOXbEhg7FIFXsSOf6rb587fR7BoE0+2V86EDNS
rjRFNgzlq5k8FaEIh2j0OcCsBYU+xe1OQwjGprlP7PVMxt5aMiB1/+JbT3T94WQ30NkAVsFf3Pdg
VEfUHuQJQH5I+mlJuFeiS/xhcfctXmBXtf8SwK9TNLg3DMj9fgb6gBYwLQpHP0TlIVGqQAcwqsku
4r4gGhG8daD1AjAJImlnchcUkqEZZVZTNPBkQ/9//XXcffMEYfbBX19uB3jc/VIsqtmVcDhK/MGP
59iK85PeItitAfAD3krUKAWjlqyEp81nD+UPGPR/AFUo/rPOHVZmYHBAcZSwGLwZBg8RZfUAU547
PqS4En2j4QlI/gsgxVqvHaxxF2ODmvpXJExJ0XpW9LF9JFEwDmZQVP0w8Jzrr9KOBQH5Y7SLVnrM
vGVeUts3zhqOpLvHTEHHVePk1xwmrabyHSIXbgJtjTuEF57oJjOXd49gZHGj/baS9jSwJfKK4yDN
jK4JqkkqVQg4ybPgXBjaukTi8yjiSzV734C3djlXm9N31aii9hbnsV2Er5c9FA7NTGrgyVR6df+X
q2mnly4dtasWpbX1ftnl0BIS2S9Nrnjy6qhniIGSHxirxfRHWCxwsHwE5L9aY7qDsVgUfFlW7ahD
VDwQP+g3S+STc5TuAhoPIvdFcO3ZoZSfs+QawlNQDylYLMq0xSnsAKhcJQG0Q1tWOn1obIvg4aWe
EC7NlNaAz01zRxEYRIJrCYYY9DeZGdNLk6DEUSctK3OA9rFJJn8HCipsxT0FrNsCLSVlCFGRoAuj
rAwjE+u91wd2Emtt8RdJ18r3N50ASJw8Au9xGCQg5Nr6l7v84ynA9wU22NrEPjz8HAGCDZtu+tek
L4xIgojqC+RatuEP5wIF17hGL8Y0el7CaYwzVRsa0fq7x+jlrj75yEYNQzp7MBkLlZhRzm6DGpm2
OCgC+xijlYSMcIBQgcaoe78UNlX9zJiAm0EpD2SikdnPdfQJmrtaMtNg+i/XdicSW99PfBOwGSCz
ZkvilQHLQx2Yq5ZUdDFYSaRySaf6MUhXA/myyNZ24EIeULvzejy9nwrGULOoGXRLCJEmJdtsOAR/
Y1kpN30skYhtmQpcyyeDnEf41tE4cztfcNtTJfK4lt6Fq/4zIwmTOnH8hheXfOPbNNIKkHI2Khmn
Izc+ZAxbO19TxMVtVqy8dn08IyB8vWajWqNDbMpMtx+J0Am4c6BkuroKXZwBrL/Pf2KhOZhPO2gN
28lWBrM5s8fpTYR1F2GGF2xSlfWlCDrG53ielYczB75lWtO0CKbIavZS3rPgfKxTU2ceUlGgCj4D
FYCcECNeK+rHXQrfmgM8ajS9ybVQTjyoBFy2RC8JP4HlJs9sVlzGeui8kDMHhDpMPK8QUo0Ow9CU
+xx2RsccvoXkDVOfC68YEVlmUcdPzslkOoVNCpZv/GhmDyxbgdEpF/+i2ZJjVAAI4yi1ByhV3GIk
MA4yzLzlfWddeR71RLONhjOxNQtVxRIP+aMsverLBpTvIWgfl9o7yza3RjazsdcYGF/XROYNViH1
iVMREYmKHN/+fybskXvgpSBH30MzvrREJDSRVwGqHqgvWD8ud+EbsJHLHAIHykvm5mSBbDvNdx+u
whQ2Y5NgMU3e79E88mA7+2xiPWy0xA9qWBGj3BDsFFX5JMvmeAPlJ1pA2GF5lQ0zeeSMksClmQbt
Eci2Vo4CDzlr8Ce90/urRhCoK0Al61S/IGUnhrAQC81sjLRNcAYd3J2iiKAOfzec+2DFrjw+4HWO
s49/bXVrf2B2KlavzXtwwcghuIM3+hX0AaFN28AlCEs4ut465u1crSkhxM0sa+/VlXfEOhqK4s5r
GpTpfXqv8jcwIdvPTM1uV5O+CbvGqjxklhbqGyGj3wnSnNl+rU2yC5g7O3RUADenp/p++83FxwSC
jWcCUAwJTeVrQmmpe0AjVawarKn+9sB2O/GPBjDpGrA+lAyc+VzO+e6CX702Vv8aNbTgnLkBJibw
lia3thotebk3tOd6R9BkwF91pRKhs8liHqyxOcBhULSlidp/59XWGOZq86pP7Ho149U5UUvMV9nM
DoZXgqqmEm3sBcs2BJ2VjNSB3Tq6yjusCRb3KO03+uq6MacXwHSkdM1o9lCYrozHmW+eQc4gtNZ/
XI15vCMIGKn89Dfa2obXeeuWfAOCcsGlalXoYJg5nDiGriY4WYBFJ7uAmPZf5P3IChjGkoBS5tPN
qMrwGhp9YJ0JGaKK9U56ee0HrZOzrkFdn1q1mJ0LvLjFaruojA0aRifeg8e+HyxRWXWN6F9MjUNp
k/3lfL0rOTt+e9kWbl5zojBQPe4CKOhHq/Yowszj8ne5PQMxhEzfL+1rZIJEyeNPtAQ23J1vAf0L
047IJ1NLmcKyMdh0lDdQ6iqLeecTzxU0IRofipmPOS7RXJrdTc8TF7xtHM3Lb7lwD8Ws5YBnofUU
9ygD219sgA4c2nrQyKhrwU1GDKEyY82/Te38mty3/XBmBPellmnUdEP+RCah8doIPaMg2w2sE+pq
lqrAzqPw04ThGnArCrOP+TZ2w6eRn1Cl+YyB1PwUf4i+aNF6d7u2PJPYeOzh+JblsbFqQDhLOQqB
I3MhcRtCtvNMvHylL6HBtQXYo4A/KITmKA8veljAnZFA6OyGPIqQxUC4/cYY/5S/KB2OZNXUg8xb
JtQ7DKbhdcOCwg88EZrOHsbgTquUj85LSsDRuryV+/Khd/PeODrTLZyvN3kEkx/0qrlMsd44DnF1
wA4RzRt0jvq8O2aA46+P6zh+G5+k87IQSO1bJdMEySSP1UznUdS9SD1SA+83pHDrhjXw1zxs+8wK
R8eXgt+wrwBzk+IVHRLj+xy0dvpxjXMrx3B2dYzdoiXs2owBFLVqqXatY0WiA6Ib5MnVGjiXkdI4
iD5S0uO99ZjOELcQfVUxoBrALuMedge4FArSXJk48YBHxc9G5plbjdK+yTVLFEsjqACE2L8FoCpn
cRQOLrQNxOfUuKyYpdTJD8pMiHDLhuNZ2F7pWGZuSMv7St7bM//IUHkBQf8O6flihNryzIdXQjVk
pXRF4Oki59M88qDH72owxaE1KFEY89vGqQZdgxm86s+KbyAvZx1f+aGkVdkRPE2xbx5nXYZiF8+L
JIJHMRibcvEJ5BBghp5jkne7Wv5FzFfJp4BN72Y0FR9OpG7QH28sLk7SE42Lv/FBxB2fMntPdLOx
7YW0urx+zv3Z5x1kbdwn4O40sTKhlsj0QPv5APtPR/cGyB30cuvialMv1PU+YYm8Zs24cGy/+gbC
SZYF06na4ZpQkYWhNXhu0YMdAeP6fPtOMjZS6epCplVZHUa2jHLCHzpvBsigSRk6Hud3RvFrB+3z
Sr5vAjl8/FEWjn1voiIe/0N2FQff4uUuILapWr28M0410G6d1VslyH4/rV6UlnJPqHh28h/uZkg8
AjXOMp2wrxQUMTryI5Dk6Jc2GnnCx5iHlkGsnTJw5gFLAcMbAJZ58wCPN0QF7bS2xDbNRFs1/+I1
MObzRoop6q9HupRxsGNcRm3KkWNKTgQZQiK/EceLy8cYdh9f3u13CmRtcEjAURvfObN3jiMRVM5K
uL4mhCGB1llpqv6x4rW7o5Lhzbulf8/XSHPu9SNG8R+8X9A1j3Qb29sX9szjBDYkDNfEpgH0/L+T
jVOaJJocmPGmE/cdf3EOUSB0Baf4LfZucRx34o01r960kQDbNyUh3INdCHi7IyXZli8i/1hxlTSj
dDf4ANgmUbBvduNuIOwGRaCDpqHmr/jinyGoDlu+fsbTQ+hamd/gUlTGgzolexZGitkH9DSzNprD
WhNi9DUOSi3mrUYHHYHvlRC8Q9YsrVj3WgoYpoqAiIzoPURcAtQTVKtu1spZMdsPMgGyoa7byMuV
RHS1fsZF5HTCdJ/wPmBGgvkvZ8ZRRWhjjYquNJMeJU0S+rA4iwNd0T5UWdrv8Og/uYqQ/jspfk6A
mLD6PLosK9+gbdPkR1mnt6yiCUT3HQhrORQbIVsYvzj14CWrYyD2EjjCM9DjQg5yAuuPwtzvqP2l
TsmpzshPwHqe2jft23IFM+98NaFH+ckhTRbunGpgYczOfvq9y3ynDJsS+PzsQDDsrihScfSTOjVA
qyMD0+Yo1bVRQXPrKQcFWJ8gp1izGunFDKAAqKUOP5A6i9QKFmGLEkTsBKkaxtiAYQC1AtXVN/yc
dSL7YkqI49jZoeHoNB8DyDQf8LKhWPSmIPxwny4sfWaqVfA8otBPWUoTGeP1WM27rPAu5MXz4bjF
K8tUmsY98HOF8zqBqhj+RPWbdNkspH5BUBFO5pnNXLv0MTul6dEODIvuCZn6bmsmqplwG0BAFjU/
WJ/jlOxF3+Tv4roHqRK+ljr+ZD2qGPqxHhTKOH1Cqt+WUEFn/R4hHCvF5OJQpaSSpfs7NmMRpPYZ
KbvH2BAWdPIP821eOYKTKPTc6h9Z9B9zknUgM4OqYM63wrbhEpWhPxeFsypzFuJGtHw5Kk8w1BF1
3bYc9AtoNm/XCHCu3SipN0DqF+18E+R6wfGjewnV5fOH5SKHYhOHQOgBkJQ1CkqHFVMONWaEzvoZ
1FOnWYT5HBAy1s25wLlLahwQF7dlVbbGxTxqPdUmNJgByA73pQ0iT8cBAquh4Pd/lE2SJ+fuMl6W
Clq+PgmmYdN0wwz7uHV6Oe2PAcBk3TKhYq2zD/GD9Bo+2G/XNR+XVfNVzKTsKKU8SQ0oxnlbfFdE
oi+izZvw/pkvXI8WnBYrHi4Lpgozj2K4NtDNIl7iGq44nqWSqSJjQnV0TPyYW3tvIbE2XA3PF+S4
NGvdXda63eDzOVGFJ0HX/xPv17D/OJ6b/RY3sSvI1EF6d/7C/jxJHbJZc5m5BnKisrGwtWZFBQlt
bmuFPiMzfuYgWS7AEsmMJj5S1vlhcldjvnqsHD9pnCmHytwqN5NZSpdg/C+DyvKOVmSBmkNGn7NB
635i/8S1L+IaTzY/Yxh8vmfwLk5KDqnM2lwJE5eRRtkZ8rnY7CJTi5SKLCW1eUco4ioBMOuhXQ4Q
AYtwSeasA66JVribDQxlsenFLK4ims2KLhThDvBV/6gcW+2OM5acBNMS9HtRoG2jDFJrrHdhQ4y2
FhyjDRNUVSPJ1ORRXQ+BsLh1/h0yBXCrtaC/+Fmd1Wbctr2fhvI7PEklny3HZpDa/QMXGJPNy934
Y2cXjuAEVyIAblS+e7k5W7xrinBH6JXbxaL0ZVJ86Nhy7owSV083ypkif5+OMGxz9KPk/mS5N9iq
iYu0aGVl0zInkTgaiw36CVJIyfLEFVpq8d5V3O3hiXr5frB3rYy7vD11yttSORVru6nW2y0/Oo7D
2SjdtFqOcE29NU+mcD2yYFMN7WKz9KGTf3bN/HD3XUOnV7cum633eyLlXFpwZYDZOVWmD+HXQP7n
CjiaPPWKjviKviYucUtkMUZa7FfOe8Tmeh4BjQeTgr1kXaqd3zKcnnExoSzvcR4IVH7wFe14QCzJ
WuLMxwHHtX5ugWL1UbI+bh0ouzM7uiBN34NPvNoYvL7w3h86Tjfc9obTjeMtlwRDHmBBA4cZIeu0
4TCC2Q/Ct8gY6P0ZmfYU64v+T0nHh3mvuU/pt7ESp9WmWRweEElRtciyHHMu7vAIIzUvY9xYW4c3
JOM+4Ph+tWjVy4FyIniA8O3c6LSCU3GNfZ9sNfn8kVhtdYGRJ6vwitzgco6QRCVTKAkng77cKgbS
UvnaWY2mTgjjQ7VtlGoK9vg0PoQExaKjoI74HTGAPCJmgvex8zFFZ/QF3OtV5h/H72eiOBbWfkFZ
bGK4+aHA7KWcI3SinkmyzpVTf6m70T+AS/50YMARAPkeXsRD+n8HSdYR49k7SunrBh5ArSFFwIlt
jnGR2ksLPNrpgmLa6qw/JxA3wP0KwYxjuOVD6aNnhWHzNi6emBCR4HWrB0NSramwytLu/npvZvma
RL9n8FYihkfMWMJvMHvfjVwydJcUQzD8ko7CJrOB4NzjzhOKy5Hx9YxVCCW1bkMz7SW+7sM0TWPe
vtT5K/iuqsQikpGiAGLV5J2uRcdL/UqoNRTY9GpPEUmhaWbBtOFt5B+wn5xeAvxGp4ecINNzK0t/
iUinoYzT7hv9vkNVFVT+47vmIUVTkHNpdfB5i6gpcwph8r19N4su3SHntf79Uy3vnhqp/5jl8udW
wHWNoScWeHcicrNJY0N4PHlm7UfDy6kvt6IZn8EqDMqFnQMygaU9lR1+gO0/0XJbi3XmOp1DifDJ
6kQHRc+FJu525mWlLZ6x+PmXQAEG4BvNtne1/5ZjzDvhvyOKdHoNzgcAZl5GvJaMw8iLTuyiOmjD
/C9gRfuBOM3+xOPKjubAXDLOp4FYnaBNoBElhbuDm2AxeWh8ohlljK8QsIK5g/OF4sHxEvgwFDNS
zq1wXZfhSZyVXA96b023Ac943pe1SOI4ZVuRywm3NAveTN1S2mFiNfjmUYFgibTRhyz6S4vJYgfV
6x9EXhK7RVAl6SVO42b6armjoG9Db9Xyhd4etTTKnSK5r0MEKBmlJempMoDKA5vSYKhQEiu7TJfu
wNRI85ZDQ1wbzdylxKoNtBBeD6DOBdqsltkvA7iUBdQJCtvEkunJ+WcaCUQxyRU3XExWSdXubCtD
U0g06q/0z4OV+tFUNSxxnetPb+PK0UAgOZuw45+A3aOaFUW5XcgLmWBUtVrcXLZ/mTzfP6xsJD29
09x/QNv7cFSC6uWbV75/epNhZST2B7gp0Ua318/r0Q8tkiQW09iceRnoteoFKcqwN6gynNLweLML
Cb0Wd7XGhL3dVTaUAaGbJ/Bcjcpq57SrRR5KhPgEO+CC5mMVoHkmxbXPsGZIlzMVl/VDoM/3G1D8
gZxGCaaS8b8bG8seQhA89xF/3iFUR0AmIOI6Xd6dm0WR3q+WCO3eGBGY9t/2u/J+2xH0M7gVTuK1
8L2JL47mDepD/1oZ3KpyCj5/SXve/RZ/xm06T9oDtaRahmf4l6BpL4pDuwGpXVBwOqvMTWDRVcNV
ESdkQ5B81dimDB7g9N6vyn21O/sJ/Lvasv3vpmIVRsmCuAYafp911mrmDh1p/w0SRQ1o8+Lbny6d
yWykQcqRBoZEzWMrOslh8M6Dw+lYdb94c+E8QO1RP24jEc+7rsPrU7ZbHA8xTzwIDag0LZWyJ3Tz
a4PFqHxJwRsZzeI/Bj47x4sIjP4M2PnctmNmgYu3pxg7C7SXr3EFVyMmIHLTDKY06lA++Hlh+YZk
gqQwbGbjD6ZraKeCdO9HEmvh8G8ylW6Bglwv06W8NmAuodPnKlWp/PDsiqzoopDWp3zSwwVitJcZ
pSlNQ5h3RVhyrrIdAASNcjadKdPlBP7VwKMSO+uzYQDkB5dctDfWDku3H5U1KTokwcERKa528Y96
lGZ9eDhp9VWCq8gkMGFAcYy5VttoQ83AmNP8FLt/xad1Pp2SOZxnX4NZZWX1fwxHfUH0a1eKb2Oj
9nwJEss215sbfuXYfvmEnF9ZWALk81xBvg4v50DwHbDc95Awt/RdOBbCn2Tu6fvrf/LNgriGiV/q
DehsCT4BU378BxSd3l8nlA0s81mFMvslrVPw7RK01o43VjACly1ztYWyg4o4fSdBk98Z8XCHfivJ
24V4nygMf9gAIwuV/iXZBXG9xj2muJ5eosT6Uk0+JH1NNDupXpSza+CgBD2nrhIHbh4Eb1Cxvy4K
DDOetnooqfVzVJShom6AzvyNo6cXstGtOP5H0DLjpuuU7vEnG/bGHUGn4EDmfwE2pvEO6UAY1Qq8
gEYlqtYyIgh7UAA2+XNL68bl+at/dHEiy/dLNqmtDi68U+MDsbyQ24VKvgci6r8QhDPjsiAh3w30
MshEGZI4D697OcKbdP5oGfwm0F2sKHuvs1SedI5s+N1mlgQibKQrVTIpO+iTYgWwaW8VHYGXiAWE
q71J0vWW2jXHb1qXzoItpsdIJHhapErqu+6jTsLTMX6Yagu8Ci7xJUCLhYbjgc+Q60Fqm7Rl9xtb
Xa+ptfMQXp38Julbr7dfAFI3tXK2HZVXdQALgHF55tpGZ77gKf9eVcHme3M2BVgQeeHqxnTcpd4b
AUe7ROPup8rgoIOELp+LZlB297EbEJKQ9L+YReQW+ZOTS3caKB+HyrNJkfyEatjnPNrOXQa/Mov6
ocCW9my1rQ4RMq8wuCnuPi1nireYd8I/SRBE0NpPzTflr2rvpFALhSZFkkcw4Q4V1ykNDUiTJg81
STl4XvO9aNJg1wP8rg8C4Dp3ID42GOny3g928NdDJb0WiJjAiDC3LluaZnuCERgtQcY2YLszAxxj
6XtOZUq5n3vRA+wEm5XrDrZvd5aJ8LSBSY3SkpQuXoTciLhJF10PJ1IGaTu4pj8CnemFBWiW68sZ
5c+8ChFTnXJwirQ4+kkX95N6wHfA7Y1Wh89zQXJZvB7rk/93yCfBsWRcMMKUkTTig4SzTkmsfy6B
wuDHR1HHNbcR+c6Hh0X7GiTMWrcGku2X9Kux4kqbtjOm58kAM9reixss50dumvoKDIw4XUZRXUz1
Bdt4W8rvCVkoeWNvTYxM6WRJOAQiLrgoOfX+fow6T8qNGUiDFYiT4OeLHqionqiNRJJ2wIlprgTi
YD3kZFWEInpnsmYUBdUKYN7VlV3lHoxHEQlJnJQhDbJiDmEEWrvjDhR7QUi/8cS4y6KSaXNUwOaM
lGB4lUGRJsgVv0K/4wynOP1Rrp1Oe9tjcoRAdPDJumjztnIHknbg0USug/crvT7N6MCFtjrWdDo8
kOVdJoj7DafCdtB2/+PEPZbSZdvQVwxJY0EwZF+8UuBRGuSHARnFB/rGeqCNbkPvo8sDuAHeTnq/
WPN2iB5yg59PG7qgWFjfKXA1A8yY3Ob7PMfndbJyFLqtGAVL2bwhC1X8GLNwEIAopYzBhRK8Lbwd
urgWjIB14U9W2vqofsuMtPgEUnW5x6vkB3Fm0/eUn0qKIXZ7Fl3MwHE/HlX1jRHeIUtQ5gqDM58M
ixh2V9jmJjkXJsNOMCNsK0iXD/CMVMKUwuUSlGWOzxHBnnjvCVrbVRZqe4lhBBRVLKtYxuridZDl
o278h9jzXBzB7Lydijm0Y1dqjifashNRl+I9oG7hYTbtUWTXyMjYkJudWjFMC4MONKgW6Q+ODe4L
u9AMBHydEx5GEkg2OABrukvIQOqYgKUB45RZE3j+1yrrCXxQ57avFx1qDNc33DliZkY/jsbg8vb3
/xfA6s8Dczz2bXThoVQ7UMrWtMNN5ZJC8C36hOBkS1iVjOkrMvfWuR/F2vH3z7LldvISqoFextil
Y0sYsFW4jOmGqY4IJAgZGaW3WboFYNi5g6YobiZCVXIuuph/J24gOjy0romk10TFjTCyRJ4qK7zr
0HKS8HaJI2JEPmAnmuyieqO79KadyoviC2JOF60UZpeiPnI8zROhXHs6I8OPRh/41NLb0WqjUYvH
hKZK84phkgS3swHBzAIn5eZknARNVe2p2BBez6sULXzKRaw5n/s5O3d35Q7eKe6dIoE2FvsmVbDj
+/3IkmvafBDBDvWmHjubAONHBm+PoH5UtI4ZdB92gxw8NqEqOvxr24FN0LHFDP/jP7nF4QKbwKSf
rosD45Q6Gy4NLAkFDPEkMNfcGzaLv7GUAt4QO1DlGcnxVRKt6RoT8oMqjw0e9zWWzbyWF8nsUOBv
6QulA2kqdHPjuAdGQbQ87gxeGPdHjaF8EmgdyVbrtM1afr0UFXCE9nSUcWu9cFgQfGvK2ZwKr/i0
rbESaF/f99J2EQwiS9BMKHFqxi4EveLlb+fhvSKnfMW090nexcdr5HquKL0H0wJk0kfUPhxcwJ6F
+Iksnd458gG1G6sW/ZUccF6SJM9camJaarxDZmXtyuhlOc5qdAR3WfUfsowk8LqFu2UQCmUWjLZu
QeCVFcuWc4wN7YWnWlLVoUaOGPHYMLY76/DB6leOVGwCz2lriE7qieJUyBtpPeuX75a5z6J0aJwQ
F3y3BoS5q3J1PstoUcOEDhbuYFK5fNizLF5TqOL5hGB1hOyigN3fWjnvpXPtoajr+jCqeVWr7QuZ
JTNc01taMj7sO9kyrjOZCeXeoCeSBVVbd2LOsRetYH1I+Ff9+W0Du8Ue07JGjw09g0VnBx+VS30/
sdzqS9eZminJnc4WrHuNxa7tuSXYIZ/P4Q0VbfCKrj4wqjG04aRoH06dIYoge/taGEHmEpo9moSp
re2pgZhOxQYaTH3+Go4ouPT+E2dl5B7Q4nwT2i5qpVB/fhj0rzTjLfe/qTdOPxzfANtdDxMz+pf9
NKlcZfUl9XCJ38DhtdljiszkJoj1PaIIUWHrKwdeAYHuVd1VOjqf9JboRttNK4FuXILR9bOsVMj1
xivHzg0BQdpV64Qvb/evGoS+3BtWLfhH/Iien9FGw5avgZKi+9+Y86fPtVXr+AYvyc7LPvT/f9Dn
uEqIbr/g0nBPOvJSbjC9PhlaVGCsJUIMzQCR6Mt1dNo11vN1SWtmbQrCtT4uLe6O5aMMGyMPz4nk
LMVVkFy8sFTOE2uVttas3IW98SDMkFXk5KoRrQsoH7pHRDXa4Avo7Cci0qqH+jjKx9Dj74vxNjGT
vWKdt+48xLKu69uyOMFHvX6RAjvd1Jkj3HyzQ7onYEnDo8kp9iKieJz6XsfvVGlFyW9hz3cPwAIL
enWS58JbYbTlBLmO+4FH+ffyrtHKbht/EXc7cwQTu1/1hNLFICLDwILng4yeIwnGy+nnbeOZuiJf
ykz0sLxAywa0cQ4RiigET9Cy1ffQtrBO/8aWv8XUX5MRa+gtrZS4jA1fNwRUiVGpYxHxyYTTELKi
S/atq9xT9R0naU8TBcoQYvpzp51o4hhrsilU0vJTVEAg5VMB1W9Gddjc7R6zNf+m1vpeH0AvdVaA
5JuCwWoWZLJ2nMmpF7FhJS98qHPhbrOVWi0FnrZSGWANNwF0YCSJ3lVt9VkqKH1nPiUJZasFZNlK
NEXuSiBI0EMhJk2RKQq4NLMj6QckazAU/5EgyzGPzYEyl0Als3T4KZj8Dc++lVny+CCeLTtzKA/4
hMLWScPzO3/jycwEA3KCyzWh0ONAiCtl8E/BwnsR3tg5cshxX8sd7xfT7WDHNUTt8AsH6TcfOfTr
in8mXF3JXm9QiCx1o6JaF69Ey5Wx1Mh+AZNPZ0GVdOBnWQeggVtuNSiGf1pQYLtN4pEbzLStzRqb
MR4/mgug02xgAdRZQPIQxRlttUxEXrAIZwBiwNOCYaIhL9U7waOMpwAsExvBSb/bFB5cztcIzkxC
EL/HQkdMzAxXfloIg0hDNyn68NYyXA5bM0lbb2IRYeCufuGEiULC5PLZ5iq8FimUrLDVb4sALoFt
alYXrW4AblSZxNYatwBhmkactieiT6XFWWZBJNj3ZATbrOWUc/qZ27voLwH6u7rGLtXiG+zqxz5A
B446LfBs0dlSv6mbNX9R2JadMQi0fo7q62jnDAFOGbXg6N242rq6lT3qNeIiMUIvWzkviZ3i/VNC
MvRQUR30PtAvjj0o+DnMv7GSlZChScDf+a7suVh8zD/F8LVuAYUFOfhwYMcRfAO4ZV0asxZTehoz
8bGfAQpEIbz+8yRQ3FleDleLVg2ut2KRNWOxP+qvsQdEH1DqF2Q+FBwTxE05ERCWZA1Fdk7uB3Zq
qYgdW3alRrD4+cUHLuOLBJQtVK/7AlknwozXj4zc8XVQAxD3YYL6SCuHCFJGtnTa+p3z1ORiY3Vo
a2xDP7zDhDj2MxEGXVdBSZzDtJPTo2Ilqkk+VZ6E2/p3gfLKqraxkSXF3oMf1rtazWkxzacgvpo9
79UD5xs7OiwHIzFXy71NrtqBr/2hCONAyl4oUjRhTWwJ12hgAYWxogOLNJoUhqk3Bu9SbMNJEtNj
rjWve7atcdnJV/jdGFOeKiHQgaD+DUx4sGcZMEejD7BKadzQyME1ac6wdP1tT91fX6Pj00MP5Xc9
hD1n5uiBL45Ce8idjDzzB1a7dTSmU/i32uZ7EtonY3uqaJ8+RRFsGySxF4yPytGZdqSGeRuhQ0y+
SChpDKq/eKzlfAssIStDfLTX5Kr8BjgR+5jjsFVaMdmdo9udYI37AaQzEoEUaFH0LPGVE28mdJIm
hi6oprVbsnEfbeiiiHgQDXwerfTpB8FH7Is9uQNUIzLAR2Q/KhXGCmfmEEKVtIp603SuxBKOOjOD
iNBdAdbIyFDE7GW4Ae5nowXSP+gDnfFz1XThTf28RuSa5d0mShab6JR8Hy4xzr1r8G5GhKrHKuEO
w6ucByw93Rhu+sGxK0jTt22LOqxJk+WfEqHt9rlP92tCOiqmYC/TAhowdlOupfqzioiLwE30wKzb
iZLsq6h1BL6Ia8dqZYlKG24HExshre+UgEC5mLF2wrphiNmHf/uE6gTI8mQOuqAd8mKdtjCYlFlL
tt8KO58jdk7SCh7aCHHOF67LqFzwk8fcvGOR2EPhLvxNiFyVM1HoVvFvNMnikHKWqfEEhl2CqM1V
fqWnh433O2ec9HKOd8p6SIef34pgCeKodaBa2Iw4bjpXHgBZuOS3TCl97oAjJkbtg4QpQjwi3mZT
2NO7cY0COLVfOhCf7enWn6k+TjseiNIz4+Bx+RERNooXHmxEax3vcjwkkP7lZpaetrgfgka9Xcri
f+mqfrDa8Xy2QM1aqieIg+vJSHSU81khUN+h4IOfoJD3kSJ42q4ifJxrvYuC36oJCi4RcRlNsk/Z
7HGw42qhaJ1Jswu54eL0eCAd33j6KD9KJ1zn1Gpxq+DNROWIvff1/lHBcrYfYHgq21WFjn98bPXn
vnWhD2Mz/I7VkhA1WEsWcg48WNzrVz5doACaPzFxGIBC0f+mHF2l69kN8c5QpGmpwxkOF5/OAuwS
dAeUHYN2zCHsLIqIOstV/vP6C9H6tAaUC6UtqGT1Ocr9eCObEk4TJtQ+8/pxch7ZYDmCgBtBWqQ6
XpKC7F+K0gbxMxwXH6Xl0wy7u/K9rhkcKDauLrzzuv9ruq9XpIqXKY3lXwa0WS8x4W9oUddBtif7
xA3B037oNePvhNYUKLNnqb/9gFKblrKXMWidNmeIgw0zswMBghtnwzUjKebfq/SRS0gSo2UFtVLY
/0PFDKFi8RzFNFrne45L1VMqHucSfUBtiDZbWSoWv+1z10TYPHdqDnn2NoD2+SCx95y9w94uySKe
p2wXqjoa8NGrcJDyYIOPnEuhIXmVIfmxotfkzp1vyyn6WmFIj6m/Xg3pfGpKS8goOR6HD7AS4cKQ
8Q0C7P1AyQmgWbq4Nz/YG++iho2S3c/N+QlOiBYo1QsP54nBP8GrhIs1V4DLoak6cDtXlSg38bOd
rDeBxu7rK5RCCNM/ZaFzDlcDr9Uibk+3nnCqtj1g0coFHX7TSDC6n8ThzTgJixMlEb2bEY/5wF9h
VMz+nejhB61K16V9a/cXP959gBMHBHsfWqBa+dOePzBLV1jKEfexTu8psKAZG7IHLqy6LF5yIkaU
4WQw5QYlLmrT3WJ1n/jRCiDsbMhZ72nUUoGYnuBESBuTFrWd+mB9SS50qGRmWhC9TEBqKXvzI8Pw
wXkf6rZazLso/0EBD+Vmp86HNGqwdm98o3aWXrGRJ5UHEfNH9keWLRO5SeuS0u7rwe4EEm70gShH
rJpEPjSif57uRohVw/ewih2fTfnr15qU5XY0/jlPFDrjfzbuucA3QVYrieI3VfC1dzqCPeuOLuid
qajY1yS9AUkn2cGZnvP4lJCz8tCIyNXfHwUzu21MW0OsOsk7+3qRmblNa3Ky+u8xbndgaUvIS9En
H0ejyJD+TE8gKp5PGEKw1N7uN+PR5WjKwhErkxSJTtccIv2kjTt4TKL+M3pi8jbGH0vpoyHnoOdk
RYjpqzTVP8+FRaaJbRu/UC8cqJAd72LsewRZ3+Gr1/iH3chss+8HnEnzm0LbXFXTEGZXuzigKBRl
E65CnsRt4HRV2Bp/9P+SzLC673XuXd7o9v5gIuAFDF5vCtn0obeETvqCserRFmsEjvvf5Xjh0j55
Py7JF6OFroRpH7BNmd3cGUvUaHvSmRtvDVCDXDU1yDeuiPnXxMNf0+7+11BPx4m/CT7w3OOpSRHS
nzZYsBY/rKYPBny3mdIg/GaTkql6t3iY/GmHITCb5FDSpTErVlrFLFd1IT2JdIlR3rraCtENFNRh
crb8MkA9PmBYbUJ0ykAOK2zztWaCjw2YbJs6Ik+xgWgc+JZz20mumRvGXarvbtb6Bfspe40Gw4L7
giuTGDJC32TFv+7UuhyABe50+K4eOerykWVgNMhdbNqUtqVT1maCPhPtdXQl+F13mdJe7qkZuTUe
tIVyTwvU7lWshdE+H7nNFyGMxgCrv060RinoI4zsJjLnwsYkQGtUuqdk5tByFWXfZC8pnGcq+zuQ
8RljF9rjH9SdJEjOcvDGJ1v08SUUargLGGwYqLDsVqOjHEKAPR07CJb0rMzwkFbTMa5vcYoGLT8Y
nWBWDV/dfMViwWt34j+84TH7fAk2t+xSAoT1GJ8jnFHhg/do5b24yEPuEliJMiT9ysVDUss+OE1o
lxcA+4y/jgsMXqOOWT0m4ASNTJk+1FjDvRlQqbXl5VoP7cpCmGBBUF1VPl/beK+zrepbKTmsmLEY
FiY/9RKnXgkKY8VvkyvbWnG0pWThOUMmza8iDhuBnyorIYCAY1JEzJqN1gKe+u8xZK1Rh0phF345
K4221Yj/kloGNkVCw3WHxScniVwizM9++YtsvwV9p3FdiuyVwqKphSt1Zh/qFrtVz5U+C4loP7Vl
SejMNALUzZNHQ07lMCqCck6R2mQmX+DMRF6ov6crtDagsBucDyA5XhgHMSRLmg4S1KFlfgK/jYyj
kqYm/iCVOtZYj4CksvuK9UT5LwLOykHCiPZdLjkByzV073+3FhzLwYL+6rxNp35YuYzXm1BONwAh
XOaP0aLTJ5NYWNG6WP+1ezdF/siXUNCwxhA1xNc+3T+o6zq71x5aHwLbRHvJIQsKKaohZM9CKjRM
4CtTILTEx6NFOaSAi4rbc0DNibgFz9OiBXdco2c1IA8VYQEquBVGOnrei8G/4EdCYSbHD9mJJpZC
MSZmy2cS6mcKygyomNg4bSSXLPsdR05hs+4SeQoyr6d1duuOF/+W/HfKXQe/5lQWL7AHsQej5ctC
b/mjBlagKCgI/myt6vDIHYppT9VanMi7taaXG8Nse1BzgbihHVzIaLflqEDXE0tOucHoe8gVmKTH
OQVvbQB5JPs12iNoc2E8TUWJgAifEVwnxb6KpVNGv1NmvQJf8rexpj9mQCeXi551nPE5I7nmS+hN
rWms8BAO2O1G5mWNNhqY3Vf1X2q0DcHwekzZxBFejHUBN9/2gqtEeREXDQGNX4WkkSdkvd9XgtOu
/Z/43U7IzTUKBbamD4aX37ZffoXP1eLD5GBFSmTYeNJx92DO5w/F9G8gty7e8VCcL0vGQrA7+3qI
+9iIOXw+UzUtoOVyDoEFzR5pEVTkJ8p+kcAG2luA9dOpQuhCRlzu5tjQvaPet8ooQc0Nafjm0Tq8
jD2cmjV/xFYC0vm2/aXFcXlbZO1JVxEwvm0+kU0lPUe6H1Wv50x+p2/JiV/rgkianWlrro4mpIzT
hhwEJhSPeHsNhTKSwkyUUjPwXMIqGBtub0s2jlg4VLbMzFTMjbf6tyjK1g78xmjBgX4QVa+4+40q
pkW+HrSDGtJsY+DqT9EUfXaHyOsdwtHaodSKxh8SNtrTcB5jfuPcYWVD7Vd8bCrrM38hC79OwAvO
ugjpxonT/BrjOokLVUoSXQd2V+0iain0pdXPB2U7SM4LIPAc6exP+njzwhDuCHFqKQdln7hoKGA1
JKJgjNkEfThOhX2ir/ulb08P58aOwWuzHsh7oAPzj59SALKYzbK9Bypm06ACuNXHuQq2NR68vd9/
D+6d8iVFrW9jsWyJeO54EUBGExGieVcsAltOZ8WFp1/31jdIVADBBeQQ832jUsR135tgOZpgCqXw
T8de1EUv30wwxw/FibFrzBMRrYHWFQ4CPGzJWq51SLMMaSv4qoxOw5GmPz9P4T6Iy5I7ef1rYt9I
CkQVZQTE2FMalPsnV4+EDybx75JqADNrKXxzCwlI/qvWTnSiAUfqIX/ubhqbCCJ5lsC5hRfCsdi8
y4QHQO0cWtwZJ066z7/Zr8zTm5kUowkb81MBVPoJCuor1byUpL8r5FeZCEjtTH8k/3GS36dMvppc
sGlGJP/ylHdWIhXIcBoUITtm4DnBZzRJnGTCGmT4vp9IalAsVV/zl2xlLkK1I4YR4Z8Nhddp6Jyz
dYqnisz7io0k96FLreieFbhS9arria9Zh1aBS2qJH5KwfXzM9JYMmn7kcz6N0vIYh9L4IJ1VVMDJ
PkFPANCvcV9HxHfjLQhkBwkEUS4Lt9tzv2AznkCPsRIdMZ1+YuTGy30WixWglBDh/A1YKoLalMuz
GbBBap+mir4OFRwkDlTCQfCmOsFSj6E104nBfY8Ny3EvwWU9pE2hR0DdmCI3pEWSOVfCdxZQKHKB
PbhwPkIPnxzY4mJjVJD4q+qJKxXuw+eD21/5nP06+cjKHZ6pQjxcW3MBzyDxWBmHG34g54vjaPPr
uExgwGvx0Eor5oMxx3m5TNHdJJRQd+H3AWobkZLsyVUnj9YEafHqnmdOPzj0UWbLRKYtzDaIufn2
xGgQR/0OcvvQbj5oHnHdlUSQnO6UFfKVZQGUX5hVs4iR4Zreju0iSaXDEbAiHJauPqjF2Vm8EcsV
V7t4TrfBRk5pBfAPktfhsrKvoEdmAzuKpAPsC6hKtQtWdanPOC4ZFmzUA8Is8V3wpL87GDsdzExX
PDOipt4l+kdTPjG2KUvaKaJ3rdls5gEnZotTAQPOLWKtrBTwipIUl+1fgkCpJijUKuecZNloemJC
+tHsOkvni2wi6OB1zeA2pLnEmHPPZyPiVffoOzeRC/kK2Le4g/AReYyfp7jmx59oWW7wpzRwdgsT
KueUxPahSFeHVE+6mQZX3TGj2G0loyrJhlj1HnYFAb0l4OEPo87vcluHsCaGY50lztcKw4vX1aq2
4srRdGA6QKvzA8eH6NKD6ffF+E2PBtTTdcusuy/DiEc0LLiaWEV4BGyl3vI0kN5mamueIfXET5b9
xQhJOCXGTWTFUAgXwg9SbV6G6HG9oDWEg5vgYs9Mefu1gzsVMXKFGnp4EhzToWAH/1M7xWtg9AhB
2s7Q7paNP7Q6Wka9jm0eIbMT8AcpZ7pM9ejBLIwNgDfmiTh1jWB6tH91C0mCbT+7u48GVYwXO0g5
kLvmrhowry2I8K2qe3CLn7qN8Ty0I9VxjEWs+p1djkdN/Noft1pqHOpj92z+yVBmc8zNiikDAizP
+PFjLHbRHgAm09M1JOYmRnoAnAaPOBdnQje7DQPTh37i3ZA63zl7F8gHMEvnAfiupq2VAMPbMcyM
QbAZe/PeA4kD3f6JeXJLmLHOlWo1khERBZhQZ5+9f9O4wlcFd7fpJJNxCgwVntmnVa0x4BIwAoiU
DG+qsTI0nhCcyTzjHnREiApCnqKSBZiiFMzWvi31eHr8OJuFXvTbUOgNJ6YD4w1GpZ1uDkXTecrd
I2MNxumIwPdb6GQvwJcPhT4VJ21GZvLI2hyDzk2dy6s50ZeswH8PIStK0/35eiCN5MstQR73FRpt
ffzddk5uiINIx+R722H5VNylVKnd2xT5tPBSftFrhakUF/9ECjSM2bLBwd+zM72p+uL19fl/Mea8
5pL+cgQP2YKCME/f0vVY/LlQILWuVXemncEISVo/9Qakz7sLCxBtMDNqmaL1RNLRpCFpdX31fvyY
Qu7DO8XeTo9IkJi4ndlH50g6cWnPlBbPXrc13AYRRYXD5jLUjdFzHeQY0TR4DmLh/kM2E0rSefIp
7dN8qocKhCuXlzVZlBhQS7TPsuihdQdijETn1Tdz7e+ofw7kc/AZmZKzueeTC8lwJJvjl28tJnL2
SgpH2swULcE+PFIO0z3Wj5bD3iUsii+Czf6v69/NC3IpUW2CAm4rdCN16aMpE/qBhNnR3zKdTMEt
0TZjjln/adsa/x78IgzD1uPACFiOhfpqt1q0Kt/PxCaaxQAkmMWDlSvBTIB48V8OX+x3WKN/5ljm
Bs7x3xNaMWapFh7CuTNNZaG2BoqvEBwvIpyV32tbNgB3IDhsa8c/m2gALyS/3nfHo8d828IPs+ly
i1gGzp9PLmr84qg31VTrla6Cr1Utqm+0JbWbB7El73qyzXEfP1bTEzyPmieqvmZqgjz77JuB9/yx
HMMTtafTGWtQj3ibSiHz3+/KMkgjuFPAKLzm2IiRFpwp34O93trN+p960n+t7VhEmNHu+9UUgrLj
/RXrttLs8Gcchrey7KmD0tg41qhUNbzOVEivsvs1+R5/8sTSg1bHMEURAgLisSjZzYZuMRvbVy8E
0LYwuba0BANa8GInY9ZKpyJHeFk3YsunEg98avgLssGhynIDcFeb7LMdLaE7fP9nNJsOjYaLPgtN
3xSeb9qfIWeg5KduyxdKte9WRWuk6Mx8zmg3SEV+4DwLlZNQLVE/dXU5jkFwm972PHxTnXT1goZk
poMwiSd1mMP9aDJfozfhAK47p/5yoChlpkJrhHkJ8C1MZQl9nXd+klA71+Fi6fnRM5vOIVTKz6Jj
uMDq4kPtbrrSkFi+UKzjO8RMIAlIssuZcNUl2S6uE6nNoUEYN1PCWtK6ti7nbAqffpWYwxibQ87t
CvEH87woC2ggVrA/2sAA+ereBnCC1OScelWJMH1jeXNFfaF912J14euFjLFL/qOgtHJjyYuuVPme
alwscsstX0/trZv0EEho3knyrgP22iBeL2ZOVV6YnEgvawAGkkLlFQUxmhdekRf2q5BlXYaB5HIG
krF1dH5Opxsm3FCfazrLCGCffSe7rqBMvVdWYgeQt0EBjD4FjWUYnTfjgXxf74I3Qmfx1BJajkeu
o09Vq4LqT2xTZWBt5LdFUINYtvRa+Om4KHH2m6nXntYHZ2D53RpMOyNVwZKXb3/nNL35tZYzrl+K
0BRtfUbtzKoq7wpgKO2lDwMADyzLf9GW7NTuN+XQXGX6AbF2XNIOJh7ew1ve0Mwcc7K/LOMOBIGR
LhqnVad0GoohYkEHl2OMcGE15FJaei4UnAnVwFY1SgP5YEIymr4NwvPxJ0KvzuNRn2OP6t6713Uj
xABsOg8UiUQ9MMFfZv4HQyEN/7z5sB1PHCzz6AvN2q5uK6c2BwQYjXB0dFXrMFaO2rYTNqs10DFw
tQ84eTCw/Y3DH0Eh4pAdSTvyNF4iK7FO3tOrkHUJoDhN1ZE5tczgF/UVPn4wLukLmZRDJGqQPVtX
0dcpMrfYzk0p0atQs5JYFg5aVjXQbjPSb/DZjpp72SIQ20dWX2zYwHelwD4D0vDmZ07TE3e7ydsp
SUrZCW+e68R0XxcyxQD2nS/DGbsqDYpUB2bJVMR1r+EowR5zqIgC6VIbq94pKtJs0mHGRKM2sH5I
bITklyOiACXT1sF0Xyl+owiUfOJof/SSl8sVzewPW/DY3YC5aunT5/eF/8+lrmK/5fRCwtWyDPCi
lFQC8EDZRRNdss0iBk4cNAt44oUzmH5sIihKTAKrzHWceQT4ezA6NjUGpZum7XeU6QySgolaY2If
KOvJAzx682/g9sbtmchBw/l15vOxVPjznHfLhDOr5yFqMinZuEmd7m58HPFTEt7WQHYOgCYQLxDV
+MG4Ct8KqNj0QXq06EiCVNtKt0hHsCwa0m4p6+tvDzui/yA1c4mw9f5jzUjSmMeTBcaDCYc36qa0
vZ4rjtVaTxPbKKbUMLjOxbBCNHrUZ1ZfS8v4t0/9iw0kbYqJiRLzf3wjkdo061FPLKhdflTKsDP9
5K41y/PJE/TLo2NwDtlmR6IPQ3qPvfEPKznPmCkRQxQiRJyK9NkDMLLbSHrmNgkm2iELL9ccQTSd
q6EabpBbjGP1rmVq85HOqleJWadUStDGfwLaBe+O0zWRPar0c1s5ce7Wn81I08LUdKEQgLdBSM3d
0BiytWKOT+2kgFQQHhflOuZ2/E1LIe95YV8GCOkquGdVOj9CVBH4u+DULfSc565KLWQrln/wus7H
Vwh0kRdX6bgvglxQdRwjIlnvnAxvwq2EJQKq9DrZcN8B9KUOa8mOCAYlJzhTM/wNujTvZEaDZZFI
7DzVXHDLSlwA+u6gEBpuck+g3Yp5OO7TY0ZjxcT7lG3etm8UwBcqAmSGfb+E9Df5w4FPEsZS1HL7
AotbvX98NLm0kjoA5fmdbjVGqJN+rIHhdXoBQ1dQJq4Cb6v4uJ1ITroAqdS6ib/PdRH0KJsPi9Xv
AigkcIA17NEk/o+4eKafVIu6xZRnrLQb6jhlmqyjKNnMNX1CD2NstwK5H6oDKiVwZGAIawSK+5eL
b4Md6wEF5RGNjYvZ5jz8F+y5MSRhGXmXiKAuqs19AWoDckVgOf8lOAUlXuyBiOTKYZMGmSGk4G+A
Qkt9yYhQPRCrFnO+/Kbo+Gisw+dgI+FCI2PUtq01w7kwvThe/KNxDyBwEMArJvJZv9EmEU3K80ZA
rPgnfvfZytrAn4bwi7LDohkXkJVZ3udzFzaNhF64mqceEGjQ7OoLJkypoT+w30KEJhgiXTQtb2gP
XEdx8noqozSwara+KNRX83ymtwslTIfARi0sxNCxEldSd+OoDB+KZjdZhGjuA+K3CgjZfafXZMHF
dtoQA0NI7/WTnLHXDSarku1NyFcxBOQF0my1UvCUf6ghkhhEudB9/EZ3CeMV1F55fx+CeQKidBt5
OG2vzVFPjIN4kiHFqrgB5IOoI73bwTNT1QwJDyvFQD3Jh8s2RvcTwAbxkHlv+n3Q9Wam0/BmHyQF
EdTGVHZRFAfApmCGsYFG7FN+ckrcreve49zbXWqVZwG1WIHiyLx0bfOhhHqMo/BovLmWkUXr3/FG
MplU9RZ4qdFpJdp4UynyATBkd4iTiDNXfqyv+Ug0RzSPa3Dl6O30t4N6vWb2cJOlN4xrL9uZKCx+
2Jhnddy5LarpstxiIJiF9pkilrjeNgqn+pjIoQYYjBYoJnV3kCwYUPi/yB0yLNFPWK4cH6ego3zA
KaKkZE5s3ix3yp3dE/67OD4ELWx9Mb23po6nME0FDKn0NVa6EFs97simuw7nbEKrwFBFsce6fzZa
kh0RSyQbPlYWtN9cjttk7UetRdmnssFkF14LWQcJnZJuPRU9vFAYLqFo3wmEdzeu+uLJ2/rZeg6Q
THThQyh5f8GYDT3azjVVG3uBIl6IJYRQ2OP/igK4Kg6zcmkzGBqfJ+GMXwPu1b8vCQn1VnxR62tl
VTIOcQuvz45JOODrLabtWs1fFSPQ+9g7cOpplQYfTwmNZ8KmNFrVGhSUwoW6zshpU27+R0LamIEe
01Zbcr4n7/ArnKxYG22UxpEpoEkr88n//WEEcqVQ+4PXee/mqnGqxvkrcXkNyOgysXpsHpvI0Jlq
gNGWhy03Gb4EN4FqM79+asXuO2LTxFQ//2QSVvv/6j+4dx24b9qBEEJPMe9J66maaQIw1kDfDf+N
UucLqF5GS0GjVhtcUBhHoB7/FAn8iAAZuSjqL7DVtykH1DoF4M2L1p8tjmY0oSwDhHZoO3lhMlX0
0ezNb0qFr2M9wYkESuTIsn4e34T56YHme4T0UlRQQWyaRu5H1QOCukv+r3BL/SVSuP9VFt6d9L6r
uCQQ0Ecgj8rSWmT89QKXCQHscEd1gxKDFBWezdn8COf6ekQDrm1yeyk/fYfRsAYyt+a5FuKfmmCy
CRQGBylh4ZeBGme6ipORXIhGFqjwHhYVBUg0AvZ8I/oA/C/56KuMhTV2bDz9AOWYyqMWMBdfoNS8
FCDXaA3w4LD4f5xS8cLSI9fnbDityWdxqbzFIy1xA3q2mzuLkFqzrRhZ4ywohcPMzKkxzfba7oHD
ju00sd8rlSzwwetA1BHKO0HyHVyfM5npRy/4EH+dCQU14GwgWpwz54cvjrU6L99G6Qx3IRCrmZqO
AKbJ4VIA1nw4919w0O4TeQXo9bEI/lKFMy0KfnicuIPhmQukkOK/ojYL+KOwm08Mlpl2wL+QiXhf
V1DmpquS9InYjBdJdOE5iHVgnYVe5PH285fQ8gP2vC/RMm73LlSkHyCTsWdst2QD3cDwJQyJ7nl7
9MG9khbglXrp9aJubvVpNtxgfhNzHmDwiYGeW3hteSYtW1ehsMK4/o+GH94lL7xS7ZH22uZttDGQ
Z29l3ta6ESUE1Tz8Sj/Zrf6VJLDEKhpiLlxGDr2xl65vduCM1khfRSi3d2XQJXZd5okQUK6cPJNM
kKiqIdIbrX4oufOcmcTI3nBu+5UY9Sz2Ddn243QQVb1n2eHBS6BuqhNmuQK9sDP0USGngEiQxxJK
7EE2W7fOZ1t7cLSmoqC9HxguGhyLbSWlTEmRSnlWRU2XoXxi2ehzHZzRnMPYkrq8LzLPUq3cvZW6
Z16FpmQHrz7s/+1Gs/k0iI0+s1cmLdYCTS/Jx3B9ZvatLzILldTW9u8pKSNFJd0btUFnuteQs5lK
UQjaL+zG9GJWgPlYVHtR9/Gj+FSQt/LlyrDIhvDkTrenaPnRJWg1su22AqMnrBoc9ltM+qH2UqEZ
wwdoNIjq6coPh51C3q38zfJTJ/DcyIHOmbDadm/sSCb+HFuy3gOCBbZB5+D6xmMMVvv3vBrNjAQ5
73tGoZo3Rtdo4O6uN0zearuAgBnnF/QOhLxFYBl4YSI5+AUZXgQTBbibYofNwA/YH9uO7298tG8t
J4LPclOtopa7YkNC8lTUWtUpDjYrnexIcX91YhfxRkusDvRmyY0KZLgct7d4/j8kzvx6uphyxGHU
Yb9JMOG8ZMeTbOT7Mx7PNKkZ5GVgddAD2Ta3nt1uwq7jePg2gN/4O7xfaFu5BUHg/2iyO7ZBnpt5
CkPJcNWjHjtKK61y9FOEQMS7UEz+6NY6C/2hqxidyTxmJnw3PzNEiL2nTzg2EXLWUgZmhwLEG7sR
tjGJD+V8d/sgitT3rphObE5oXc/NXfUGtoj2Su3KREZ2qaBB8K6toxLpuW+fq4ckx7pyH9MLANI0
y0NaXZFp951hwCtk6weQkxqYOZCc7JZ/3mkqglNe40P4jJB/S2aTH5DLDyg9EtwuHzQeaD0iR5Or
O41//UJXiBGJReZ09heT9IOpGoHHdQk8jK2HHzZn5H42TP0UAJQhJeFjN0f6ci3lbfuIDMMQDRM4
fZ0gZUQmTqbOIcdsN8lV36SNxRkkId+bx50KeLA4cCJrpPHe0gQVWTQKs/zLtEjT72rt+P1TA+fQ
hbHbh+VJzPANcp3FpPRNf/7PAVgOxZX2Neopifk5KoTtpGeDoprd7G/8+XOqejAXkg9klYWE/WnI
Yma+EUyyXjJEqxitTGLwIi9lajgWKYJ/sNeBJEoFX5QkznlHbnLnzK0RKPZapJ5yU7r+43REDjMA
mf9miw/Mq2Y0S8nBVMUL24EjVcSHOl74fYivNSBKM651Xgl0rikET0fc72Reev/NS0liLwg26gsr
MRELhwpgSb2KuRfJeKj8Uf99soCBA8HflUNhPJwVP0DI5bi4QFaEQsik8p+ZYwr5Sd++BsLda7pz
VZAY4JeXvhHjq4Efa1RTUbWdiKq2FD7YXwv/alphClznT/JLfJyLtDPhIlUkH6ueAZMGFd2Mdt+Z
a54TR//ZeuyTbhheUR24jyIuMyjXhI/ipMLoYwixb1dmAXJjiapNg3byT6gJfABb6TCVvBovBwU7
EpcG3X6+54P+dIAZctjkiKscUCeoj4+G+tmIIdDvNrqLWwJr3P3ZT4guQBB0ju6+mtV6F84XazHl
RiwSHjmgosA31MZ0kKK40etr3MoXiH0qzb7cgTMuoboC8psxdW3Gc0LfzV6OzlCX0UMwUOxuRC8F
ln47U2JCUIypSRs8KqonVHnmp7Fa+GBE/bdJmAHIbEOTfJyReG7MkbghaPkrcClLse+dFUFZTg/3
JOBxZVQY73n45n24HPrB/6P150cjVTTtlq86zvLJFjupkNkYKwnSORRWA7IfIck+rnLU2+VbJGS4
0h6oBwvb6TmbIahbkOJjOZMZ4obVVhEPgVyKvGRoytBslpQxJ2KpWnOrjZHOCSTjgORzPqeCplOq
PoD4/SvA+skO4/zvLMrAlgJq2ompMQ98IjMYHHUODhd7b4/x9Kw7f0MBw+dbGYD8SLQs5xAnTx/t
zzL+16Fgt2IpUCjkrMdDznlWojVyCouX61jwGCCwcJtSOQjlBGs4urNmf2+24BS+sMxzPtbZUraf
FQOrjTAvd+bz16DWiqyPkawbyEt2Mlx1ltHzexNFH/JeRm3toZlHDCDcfOWOd9/jTsH+7IcgBCDg
4GjrVdSyvUyvs6tLzSNyBxk5AQs4HQ1j2kAaD1O5AxPejS6Lfsfuar+rApU4s0dFdsOOvZJR86H7
wc73v5LgGukwF+rMV5d90N8eJvrc5Xg9mWt/DCa6xTKkjhNWRhy0p0YFzWBTdxTT+QJtZj2xMorK
qdB/Q8VER73I2wNG+c737mEraEWPptgkNKu1pKmrTeZ43KonvxMaE0FN4TgZzU8cREQUGwXFF5pQ
ysgWHJy2e2o3IdsKSzQyvtx96zI5io6sKucJJCEFAs6c+jmXpHFum7kuo7lsHKNbPH8HGTEUPMGu
SyAsxuqrhMmy3pjWNFqh9W97AFgnh2ilx3Ejdh+s1x/xM5ITlvj3bRD8iU9ZwQwz8wcR5b+hA1Kn
TpJRy6D5W2jtNTZQz+3KRCttK2UW1Z9CsI4VLlNSQmZULjgCooxeCxWhVSYbME/e5LDrqmT0+ilu
/nYWkhyP8i4eDz6GZkAZ7j0n1zklW1TcdT4SAp4GBMMPoti8DqJ7TwUPKqXcvZ/3KH0h7qouBtLH
fGLlKmCv39qJh8HNA0Xi1W+L3mRTl8sht09HP4kg3W+6ZtsR5wFATUw6KKg2MBdCQ1WcHH0lFQCA
+VGDNxJAN6WdGyPtZHpuSXP3wL2pO/AlvMCSKvGwQ+1c1DYPr5MlWbXWKAa0WPV7KiwAciHSYJ+a
7kPvv2omrNgpAxg9qsYRGfRkBy0/ARxcD5v+n0oqDciBkC+b+5mBUSWYYzUIXdhc5LTRAsL6WwUX
9XNqiD9K7Y6iSk9vza11FmfwxgFfBKjHCOL57DwS/zp/ba90LO/wnUxKhOy5yqBo+KrgiAFtq4Ke
+G3KSF2s0lkgsIVbxCWLSQK8pq7Lyk6psgEBjV/BntGvFQM29gjyRkg+cTyffCGrDVyjxy+2c/qs
Vv07A0NgnMXNi01mfBbClovsvIZwvZWLOmkymfrxItEj68CmbeQluVGlZ8nqrx2AvxP+cAyv3EDC
9QJM1P1dkG5ZxKsuQxsYwT3L69wzAUp5rJYXEEeD0aAQEbGD4LOIphB9/vLHqErLwrpp5wPp/7t8
rlWuDmIa2m1moUmlggcoTJFhi+8ID3QLQofUygWO2d/n4k7XH0bkv8r5VxoFrItr7RiyLMlEi4R1
uevFJ9jRoT3Js7LBiuLFq3cSk7mrFh/ODcS/5vJRHOXx08ArLdCHlhBnoLmHE6Igu6SLXTh8WXaX
p4mzlwjJ+XxtVbNZrMaR/tBhDrUfRjJ6fne/1SivhxTTexjjcDui6fOyIydW2BEpewQEdM3HoV7y
deXpDVD2EZ22q4imJP3wbJbH5bDSJDy546N7pE4MyTwbQWeLP3CNpn+1zGdAKZxt8w1IZV6zWX0T
viOr+GSO/NEUeLIjwLtANRxpZ26EN4BK6+89kqp5xy8XNgzmbcm87iyAe/nxtu9IZbXIvj63gQIA
wWQfzPqCCl9RlhuKVMCwZyR0s5WOVsr9+pNP5cqDWOzieiBwWMVRgRmytU6qD8b1oUDA9DMlwLDd
cuoNAdPvfnBrBWISeep8P2yvQNqu6+5/fnYv9gETI+HI5q+XvHTqr4S77a4p2DFIIGs7cbrW2Ies
8bUn/O4FmG4kY7/t9ICx0LWDY73YDmc98LxSBywSBCU3iq/Q2bq06sGKvEJoK2eU/t9bPj5bQ5lw
cGV39KwMTjcte0px5PH/JgN637gibVh9KmICJgtR9gTI611rH3tGSiPj2lA/oQaXN5tsri7LuzkW
zORs5RkeEEJ54x8QIcEAvvR1TkIBsXViz9m9UN+AvVQ7qRLCf5+wpKsMjA9Cz84TJhQm6rOZyd0B
6/2yvivOZ9R3znoa9zCwOqZiVro10iWjoLUxyIljHAyr5QZSDXbAe+jRJWNllFJRAK+dCrVmQVoj
2Ibe2wmmECAFm3/mSzf4/iFayGvb0IvcHCHI074nDjPB8+ux+ncb96Td0jsEhX4zEA6FNMIqRuJ0
31wvUbSeJLnPRYxvbiT6MQ81TX/bE8yaWeInGzsVDlblvrnilk6q9g2aAqTivDqMchEwghNkJqdc
orMJqkhRFFykTH8SJ2TC6WI9ElBuVhBdRcR9ZZNciaRQMZ0oi6+M9wVYi7JohNr5thOowfVET6Se
829HdO7Qjkk1j8NiE7nygSUESSE0rM7Ku/NaS9N30PiLS6xJnCzvn4+bV1fVzrCtA2WKFe1HgBn6
luXT1vdQoKKCfbfZrFw9jO8JZNHZA+RwvrC3aRjvdrGmKQOC48ihaos7kbfsjYUkp8q55K5edWO2
zIRPRx6o8cpye0tpl5buee5cZ7LiDnBj8igSVHTTSaAQ0ue49Z7ePEKweUwoQv2kJ1btK1myLoIU
ilb/Mj0K0xV/pWdF4J7vLlyvVTJHDv5irSuNAH9Ptz/w8opJj1kqAALz8Zpir8rxjsHJshmO04DE
rlUExH3Nm60ujkN9ErSWSaPaeRdhoV64JtvVRJCxTmQs/pXrwcEasAxQXYyuEbNFw8m6JW9mmK3X
Qfj86MK4bDGTrWgKihNEqDFfgG4ymQ9YVOOPjmwXV7ogp2/nyOWClMwwdg7+2XwKk/+PtwHO5Asn
OdFacTXakJzFQe35MhdkhlRb6AcsiY0qpD4wWrU0tqRpaSqDyB8mNz1S5SQ/fYiH/CgS2uD6c1S8
DD67Wh+R2T/S6ExDgl4ertD0hLdwVCF3viUL9e1jUAlDv12O2fE3lwD4XeRbFszkuK7vQt9sMvZM
3vbhh3H/3soR6zhu+37bOWJfc5jHkidqF9VOcBVOLZV4440vnyXsHYGcg8uTaUf9XhupJDjC4nbQ
y3o+GW6lKhJ996wLWc/+otVqUU93esU/okLrdfcC9YKcqhb7MQT+vu2MNLuPo/h7nwfIBnPeRxHP
my0Lht3qFDS0CXON4bQUi1IgFoHm5dGvmjmzjeqJ0mTRr+FKkdF2D5r6odca2B8QSB6Q6iWNLA4U
qZ+LOAEJ5Xatzxtdgs7J1zUV543nt1Q2JhewXFq7cyWzdN9H16HQeFGJU6Sazs2wjL0lDYwc4Fem
iS7VDk9ldGNo4WRMPSz40oLWz56m2tUVae+ldimwuLeYK6rnpg/BM4vRYz1I87HnrA06kRBgB9Kh
O8xIHmTVIG6aH28KHurt3DLmHrX7TgcUbb1SXKKOCVJS+jbzwb9ct8kr/shhucuX2+NcpKe4wKqY
aDiTikc4XaLdbgV7zkzKqECkgIcm7m/lTZyRvbeRIRnwTeYMinzfJ7kr9pOTXTNV1vN06ubvfcvk
tdt4nWrw50IGvcpEiRcg6oAPMpG3D1e+iKccgmryayC6KLamcj2VzrL74zjYNCeVFi8ldfs43+kG
No/LeRfRBGdtFZIvEOHa6eWC/JGY1wA7zJiWdPGPNQOgHS7ZHLVBf4PZ2rZVfCv6X47yQwaNXVDO
xRdjI5+9NsEawc1ULJcdid+JFDOinyY5YZDDa7P6tus+waw6DNuBTLp5otsaQ3dhjBQL0bODlNVc
ztSzqT66U8RgXNHR4Sf9PT2JVJdtbKgHntde3Hc8YsRhZbiHPxqpJjqy0pLNcNbz/FWXffC5ZWfT
QPJ0JbINFILjcQMyi2s3uO3MqJwruhx2syrl5JhPIys5GWOzf/TD5jHjidGhnpUaokQ37LA3Oh/4
53z23cYO3JeMQ4v49dN3OgCLUZDRHCBx6T6cjgG37x5qwlrRC3t8194X1ixuXGiRMP/uLS41boDG
b2JdaNVF1KFu2yH4w9LSNX4i/mtX5SmEeXjV0vwuS8YYWN7cpSd1Q4aFtZDQkRAr3CliCocmJ2bS
uHruwDvkNc/sSOehghUb6SttpP1UDZoPjUG7NNOiVB69zrGqT7rxa5pTE8VVXNCl8z8Ty/MCCwxV
C7+zPONuuIN0eDtQMk8mT/8lKSac/eDrhsx9O2uXss1dhgf2q/DsuBZ3rYiwO/hiCTC8wUtD3XNT
C3PcUHBcnk9Dm6Cm5l1v5DwWNz0JKNt9U8JfG086Rtg/ENcZXWgmvUSWKJ9F+uGb9hy8SxAz8hz6
qG3Ayg+/WWkMc9FYFE89F2coy3oiol5in4LaypWczPa7ZwdSX7h07HHDusoozENQY02R1+sbr7d1
SirS2fGCE7e9bWwcRPK4Yn741oqYYsmPie3n6y09ssAew9UZxXuh8uUukk8Ck5vma0KJsEV4a/oQ
Igb8CJAE8o5vwjo4+wqrf3Mlba3z7gu+gbV0JjApGoBzjvbEU6iD1luz9udV5kx0lSAF1MdllVH7
MhucjNFhrONh46Tjyno1wbSSkotIyBS5I4mFecn02FTg5DRiS72i0PLczocP+1wzrsRRS11pa9O4
ZiT0sAMYYiLzYSE7EpC5kFDZMk/GLJYd7qpPU6gCet+c8V9pvZkVKTVFhjSrklUDbNjIDjGNO+dY
+ILlTJszbSwmIDNaudZgSg9I9urwbxfQMpUyffGkY1AoGBLRdPDXhuIQs26pvmDPR2Lg2pDn86nc
2SvAFIwLRTqU1z0jQUja/RfbufHCFGge1nJ2TRrOG0H/9nUoF+6ps99XWTuUTcAkvbgzWdIXA9Ke
93Y1on1ha8k6EUFdgvgeWhiOXwk58WNbqczEbv+GVmbVgLyhiT5sEdPVtDPrDn7oZvhDUUxX4cft
y46fPeMdtDu4EN1BgeV7OTyNpQVa8z1TmaFEWlF9Yk/fTFUmxtfh6Q5XUfR+BtkHLPwHETEr+J6p
+IZypgBw4RLwFi3qMqggC+wETPdTvvxswML/W/G6+hfrxjUKxZTPBzKxPO6uU2lCN89uVXKRn1Tv
cLNyJAjY6GKWZ8RyvBKnIIB2qqhKC0axj64rsDahx4TMJN2869YdYUumbGvj+j3yDkT1hso/AA05
DvArYGxaxuDZ+oZGufn0opq3YPLtUTHCgTHqpFKPWMctCq2F1layL8WksQJvviGmgMp6lTxPv48O
uKyf8S/2gJ99uJPxDgL4YFuRc0FUW6lwv5UBhtZk9mVLXW8PJW+qU7rhzEw2oGo79NpV9K5xkjY/
c69H6aOEleFEAF6AugkSuoU2ZIsbRpJzCsi9d0dRgRApQihKuNCgy4oeQWDtmj8PJrIXwREg/cvf
ilW0LjojNjtritx5Td46wpAiqVJHX2QL8qX2rEqnW91bw0nGafwJEyByx2w4puf5E7i4u+vTEH90
tsftZ125hlFzlwX7Kc0vyKooT7qXzRqpBqE0DYoJ6rriPbiU37aJF6EsnsxJaNwgF+pRkE1/Yha0
CPNOWY5/c+Pk8DcGqjUqjL1M1zMVWrwWnkr48lWZrjA0eD4Zh/1Iv/K9ouCTb1svwSTP08kWenfv
HSpHp4xTxXcLwTc5IO6V+RcxeQnjFRtBuVdhVKBHEe+QPfyT5/Gl6AWILj+8du3fBS6fT8851+cD
fdN9k+HmlYvmY50JzAQ0poeIre2ZrCgGSat4rIxUhV0K9EpEydwwsWy1kS6X4d9YAw5yZGbe+6hd
AoA0+S4ZEg4/QX4WrH/qjGFxFKhwgR+PmhwTrYUSKnQ9v2qHgANg53Lg3jGA/sepbb5ercQXh2t9
tPcG6UgKpnhK5wYj8PcK4T0oQckP4ET0HybcXgUjNYeUAhdDYr8z3og4oC4F5hLGa3Qg4cT3OF7i
o8PlBl09r0Wf4rYTzBi9I2LY+u501mpa3yFIQZcu4CgV1Tq1JuFJa+pqJEhpfbtJf0LIhJrAyfaV
B3CpEFDZ6zpGL7EI/7TnTuF4KEUiO4Dzs/JIQ3hgg3Tm7b3T6Pph36cato2FWD+gYjRd/xo2nrc+
izcl7BhPTgB2H1TSjyYvdwPyVGvPfHv32+Hjc6+mB6ZBQDCfgCtwSYb7pl7eyGBUd+IurDKUGpte
3Gg1cuaEkZHmlXs36zNK3TOiIrQsUPEaO8AZE8Dk5CpTnaYNt36/0T2YeeSm99i2Bk2GYXwC4MG6
3B/8yFAZnTTs3bn1okT1eemgF4mBJKaeyCTEsqzfyzsmJkEB0rLJebt+alUTkJ5yp8tgcHrvYDjf
97ri1OxJlj7JPNLy8rszkaAxSthK3bTW27OyU7Gnm2ylWvfF+BQ4pU0HHqquYYlWB43IWFJwT0ak
aUsj1IIg5qQNnN3Xl/cQFUyjDkGgZCzG/yJ01ZbnIqEAi1D0jPjXq5w/ohU/65hMtlV9BfCzn5ma
ECy4iiKPSAUfHBtot5c4U0j98cfQZCwOwSorBuEXnx/X4hZ1zmMFODUgDjTyD3vKBCaQhfmognxy
sWVTmRKEI7YrT7L5WPcw6qkFGMG2tLGDfQiinn2IkXqoHVgG6sFXRN20tkazJGZTiuFya9a/MWk8
PoC6hX9AffGfQdAZrTFRCWt7uXjesAqpIisNR8/hLIavA4DE4212YvM0WThkR4R2UA46B2RWaRH/
QfcWP1KpFAfFTNHR6LxFwpYekLdWpA6I2wyhp+F5ngtHm3KAY1P5ntYqltXAlFcoiOpXpdkHL6D8
GAA10SQHjFLkDGdUPIbQVc+jO/uL3TuRziPUr0JiLCH3mHOBxMGvSutgIyQ2fiZODHw51fp50IAx
wDullIED8nmQQ18pBLPe1BMgZp7kXvvBlhpzhwatZoemQ7Jow+v4Ke1IYRv7A0sc4eqNxhBpamdo
uGKgzCfQOiz8DqbcRWM3zpBuKUArHf5w3n8mehqRkiworg54dE81+GTQRQgGd3gPBpF2LXgo8rXV
2g1Y8ybfTv8ZWi7e+YnmBDetJLJWthvOWQLvCr3eNAA9xWX2vuij6kjJvszJAI4MUwa6+W+0vJIj
hY9iAo421W8O2dWQkQvhcefh0gchbqb6XDV/S0JkFf61ODR8tdMv82p2OZgOZQ++RJem7mRs/VVy
hy3OE7cNXt29/xp9UtSTCmNkMJ1qfi51pUAt/IhvbTU6LSj5RgzLe9ziBbxIDT7KkBD9hZbDH3GU
BhUToz2s3+s5LaM67cVzqZ5IPmhFH6QyD5/8rXZTkNZZaYp4NsgLLglQUq29fO1PWCn8/mgZhbCG
TK45o3XH2cVVDlREo2hXTYG8pUXNWS8S+lLRP+4D//2ATtxbYFDGdpxMV2U4sQ09+pm1LmPtWtCY
ijOZ/SnZ0KrVqM8WR0tTS47wNeJcpARRM0c5b7UqkRR2fIID9GxlPkUnMe7PKvmCM9GvVJ2hhQz+
GLpafviCCGxV+hl6L9Jc5nRP/Cns/pKu+aj+4x5W61O/2qT28yQ8epMT/WZu8jy1LpIlJczszy9S
cwXkzsBo31sPle7fy+YPNP/cZ4Pb1XcqRk6mwcOLN61hVljDrgBetKaFfgnhEQaFfoVSzmkVw/c8
/wEyg+Cu3b4n/QHRBbxc5bs4XONHdREwYGehRTD09OZxB5QOCRzVxdINagE1MHsoUQXxnhThRFz4
R1YaIKWwZODaIgpFdQ2TXzbi8xJ0Wp7u/82TL6ljl6YQv/YKsoKRB5B/J1gPWo/55/Ebh2j2Ix3Z
U68KNHVJCku9P8TVGRwJ/xtE1JPZ4t4c2rEjcQY8+PQrDextot197VwvlztcBYL7dIxFFAocHZJK
hf55N/sew28mr8KjcHQkdYcWqePbVlnQRTPlF0CxG+ok3xDw83zWaVFC/0irMKKpuLmheM8NwKGg
QQkAwxFDfH/AwOaCVtQlT9xLs9eHiaq+4VKp+iwxRweAwH5MHmlMnP/WAW3/YbKotQIsXOeS7DFs
braeIDK4ncfC+wSuzkBHAM6PztTjL1/hrcao79zT3UrC1kEa31S9MAk/qJf05bVejfADJFYdc4B2
DzJ+iF+Z60BoApYd3ICUkgCAEkis55IFFpZFhQ7FyyYB3IarvWQA/E/YlBDk87BxwxyVnNUlcr4d
++BfTqapzjRu4pTBeanAW8rbm0uRXRlTgfTsr440vg3TiKXdVZqEPcrFiwZyOZmfjmByc18Lzg/t
iUxpmqTlzmcbDTFtubMgWHU+DvduytVoQ1fAnQLux50ZXicA9WloaqSKZyvO/N/UIcd2MwUtwmO/
0gR9H5aDV56MIHw5l/G/9CKSf6ysOuhtlVI61HZl4qTZW4Oubx6wM+NQt1F2PwiD0EM30p3FFXYg
OAHwCfIOicyltL4V5z81wgWdJLiTGOCil5kWzjZzW8wGcXyy1W4OMpW90CoH//My2GxzdURFSEwL
HNOqwafFTFIYr843LIJPnBuamRNhHLVYvAYuvpvKO/0aQG5HBCCHcB78ehVRQlx1SSJrAVXstf5G
RUG6T8RJr2VUxKMd2Fz8KDh0/jg8yRBwj/qH9FUjkqc4PaS5ahfxTYQPkrjSJjVr5J1MnkUG1x1x
dmHWiLKBG7RR05H1MPAgHBVeSsCJ6wPEzND+7Z7murPytkmtjtU/t1tuEf7hxt6XidStnFydKm9U
0qHD8zbn/xZS2bSINblHtN80tJhvyk9BtOhCaKL9LKNtRC89miQPR5n0edsZXf66LQXmh6bNF5dL
hepYf/Inwx1aXfhVwD4tjVSIMDiz9zq/AD7JctxlK7fh8MOFtoYrkGogE6eZj3FvgHKFHelLQ6ce
MYuDdBD1NGtkOUPl50/Ex0lLeVAg/8jFFf4FFWPgPSO+c/dTkUuXDjCYFJmPkiR14nL6MedhyvZ+
KBqH8te/g69e4EUSxNGCeZ6LaE2ua9EyJCX9GLxvOhZZuEA1Z+57W/1RSHG8BHQ+upPLfJpa4eDa
lu39rnOSnxMhScmIJpA+Aqg9rd9ak8zBtHESbGYiVP0Paun8kBvDnRWr9gI2seWv7ZnTCix+QIcC
n5GQGrfsaI4A2a03mOeMOWeKcFbNUko+ywEXbMUyxpwmm1UN5g1PYwAzsgyg8rhUDegHxj1w77X+
dSr2LzU5XbYoKoIRQdu9ywM+pcSpdXP139xNR/IABeo+Ah3QQpjE66syi/RfSfgBF+CJjv6L+sXr
effGerFbLflPJh1TzkbmctUTGd1Eghew2OZdzOGDVq0hHM5+BvZ+idbkeKFLwzhFjVHw7xSi5U6i
hau1QpevfToRovy5XxwDpu+2DqXpqn2QcASBAlt1xtZ7uxBIGRkg3IUnvh786s7VSloBodCaC+/r
HRk36UrbtW/fQsx/VQFOP4LsIUI+Oe8oDznmfmW7K54cVJYGtHsWceJj9kXW82xmprdDQROghbpu
2X310ih+YgUQ4pXP4zrCgwhHxKQjsm4aj6MPTS4vvtQg08gslImHU+b0djXWxhhmtcA4UZ19f2y/
L/Nk79pMAllqKILOOtppv6O7hAJVyKB68dLYwQZ79wut52n2u9Pn4Zhf+dedC7vr6KU4uZD4hnZ0
VLlPJA/IDm6n6UHJ7UmY7bE2/564tLo/2gDYeLV6kMd4MPBuVGcUSC4ZdRioLfRpDk4En9Vpj5Tw
m164twUIC/oKE+BKFoA+VPJtQISh8h86KF0XZCxPNDdnlBHWiAWpxyjfqi6XX2EwylTXyYRmH8P7
1m0n6qjdqXvJj9FtiwrTr5BwxIb8GyAEtNNuJorBJ2BNIHaxRMAc9MmrarPQBzDNnFYCl7NdVPNP
ptfHJLwSBcVAWJ/hODMw1uqELCfM4hCTobU5LUrJ+gTM2IbfAlxvjXVGTSgkX+28VBrbjLzu4eKv
eEMzBZBgSZEh4zrSdnQBWRzT+uvlEvvpfTfxujzVqtfqx7ar7SBiiPyG2I7X++sW0faV+nPsvUBP
OoxLsqpEbjZSs034M22bbgmP+fDgOxkclhJSXu4rO2tKzTu2crYILJCcMhLa3MyWDZ+7vJgDw0Vy
7TLNs3/95JVU9XXQ6Uy+iWeLTHGHBxRLyUOAvopOsCg7sGcFWP6Qc/U3Jn2Q5OWojDnaV90CXuuu
eECiP8hOxdfVDUjB4ddBKUaDmim6XRDyh3uAqWAOJJHtKWQu8Z0R3QIkJ1kpfXGXNCzyrpy2ovv6
3LzGX0e2JuWQQyJ++aIyt3keaSVgyR+rAiTvtuCnS86vlen/7ldf3pJi215S+2+ZnvvXk87ZIfqV
SBf0QCLqVOSjY5pPIJLj4dbSlEJDkwLtHkkLPPpUEYkkHvXfXWsQSDbxaCh8biQYa/kW30ZOdfdr
bnWDGv8JMBLDV88ULuXUh7EFtMOTvlbK9uAfPE73Rw/ay5OdZ9PUp6dUtFX7+hz5ErjsyqUUhrui
ADe7Rdejyzq7SzsRS3bmCtdOnostq8EQheXJ8dYn+Ml4x61sh79/M9i8PHZwC6AxByZedZcrK+Uw
GysgaoQvjHiBhgTZqqD36qCn3aptbBxGsmQJFcST6SbdT5ADRkoyWnfmGEfPrOHJaxqp7WfVZj2K
OpwrgXBotJnZaEbjPtYXRCFDnZAc67h0ZfLVX7TA3C+H1N0YITXLpjK+i0EbegELqX2OHKWZWTay
i/OlEC6WgjC0MTsbnzmaKd8Ci0pG6s339B0Y8f0rXAV4LvE0R2l3QWpIUMn/9KETgNoVbW45YrNG
aoOtBZwofcORAISplmK+Ls60nSGXBeQid9WdneBYWCotfeOVct+uW9NgY9fkps+G8VCt0645Yrv/
xE9COjRycpubGmuIY+v8oSfP03DrZrLv2098wrCBVrFj7OM7T47zkTXk8AzPNqyeDZvQ0jmPiqUp
kCw33VYaO256rzxXeWg2pGnSFvJ1KiFVfqCCVRJHNJZM7m12xHMaTYPOSQY6p/Fn9oaWfRrp/YMM
b68cINEApBpIPy/8aKDi3smMu/atBii+bPN7766gnfMoqzbYmxeRiAQ+sA995vgUsWI077TRVDs0
eOWYtaGlMrP88c9DqsyJFxtP6726CAQ/fSYn/2a+hp+TgG1tPk/cTjDRv8hXm0k037IuNMA1Uvk2
fMmWnHCIoxQoMIZaISmRKP0Um5TktPT/Q7Fb/evKUf0TS+1g2JwuutVN251MaE8OjXcYcQLY8BB7
JOJgvtKy5QI8b699vmC/BPan1pO0LF+v6YlAI2hYoKTV4vx/L3lq0MkKhuGBz/etAo01CdfRd4p6
C6DSA1cqbowN3od9csbsvi2W/7rSqoCunjhCDnXO9HJ8OP6T2rQHbe/ClC9zR7iuKSqvdVyCB7AI
Y0EGtIdXJ4qlxqPwb3nY6nKgjtDuFYAdgFI3YEIDxmMJ8kwNQgKHiMYxQxpFE9BBWyS5XHroDXsl
Bfpc166it0+EvH7wiOJD1MqTkTnznWWO7e5GtBhZ1oJ7amL7b+xIHS9GSByD+vAkgsriuUM60Hfm
jIdmnecXSq8TU0cfmW2DDnRSqafWXJI5z665rR26a5eNLYDRye1XQuaISOqYW1FeQaNPD8EZxYDd
MEpateK45deRLx5kG1YOx7su28kEhS3b8RaeXQ7kUQ5jWVjdOOA3Z+kk8xli5C4rYnOjlqvZ336y
XUp0ryRD9bv6wItou5fraoiR+MXUeySCXuJDQcdcw5P0L0/Oc12zqq9XWurwD2cvMNFW5JLqydHc
oWeRPTZnT0CD/LSZmz3RuW7pYnMRVnIUfP9gWpl+ye2/WaNjeVT0251363RjgFwDnQ+9n2pO4X3V
4Xtzw27mYH+GjTCh7sG+aDCe4j/FyrVz7axum1F2SmFTtsYZUcV4QBMaYXIIU0TpEr5R33AT+1Sb
bDxUlmyxFTatKe0QPbMaaL8KcjcCFWTozMSR5e0f1UhvaSpsW03bpSpKbr8hQ+AgKL2kuIUQeh0Q
oD+fRFdxrhU2ZZlEWYkwYZJY0wzQgZ4uq6HxsXHAgtRZoNbm2oZSEKsvrrLQiEdaC9FoL8pY0WkI
/pdZEF0PYZAVvQ5mzk8ldXyQ+ILNSCp9KV/BNNxlY8uIhJglRXavdJN+GjPRFz56zb26KwvXHAxP
CYbHJUz+eGox2g7rGQ8SUaAxgIX3xroS0Wkq1euKNjjvh5TiETEhnbzUwRoWr6wFvcMOuyXYgwQQ
B53Pp5uI2zeSrtXSAlxX14EC51TzxdznXqA24Dt3cMfRW6QJXoFbvT6kqDJ6Rta2jjbvBFr/+z1t
ZQoZnZ3qUO3H0Ub+xG8aA8lEqu6jxFimDrmihdMG2fVOvP1VkeRme5NZvCGgx60+3YN1HXGDdD0S
h9k20//LWIF4F/TAWW6NWFcXYND7hT27QNqU0a59plorpZfkTMduNPVa7XOVDGwgm0HKFBH+dy6T
PDbGu8/ZGAiLh1dsTLgMDoqwOsNefrLGtTLPyaoD5pwfWXOOVY7jE0O/SKR+SmwMzd3mzlyVpyOw
bqfFd4XJ0scf9Lv3L14VAoR67ww/PtcCVgppC+6KTQok3V3Kc438faF9FZhdZDAO8w0pDRlG8l4Y
cLpuotymiBLpjO2CdU2fjW13bdglIw9QVMlbWBH/ocUPN7s/Ca5Nt3V038aeUICRkS2kloICl2f7
rMcUYGqFmUCNe0JRHxlEqSW0EzeUIQDz56mhw/FQf4LuJMj5DS+wARcVEp5Xy8ibu0rgbIQfajRn
3OQTYhs2PJbulZFIG18lAmhjAHb9oI8X7RUvwFmqfKOuSTvlM+uCLWyrjtCjIpOs5WQv+sDpiw8I
a7ROkiGoY9hxNTdWPekTxsfenaE1Q2FxAHjg7DTlX3owzMV20qzn5RLvUtakSO5ypqGnJOC5XAkZ
jv8mJJYrl3s4L515iml9D9rwQHDksvnO2FPO0q8sks2iqFlLeT4HMjwrSqxKjp+esj7gG4s6jpNX
au8A1xo9xFVLdD9ec3oHGxvpv+2ixV2CtqVQdIkuvJpmAnWkhRipO/KhRoxl1MhIR3GnhUMO1+Cp
JaeNHj1h6fcjvq4Szs4+j5E+GnOHlwvIxMCW5k/D7zLbUz83irmT7+p9xR5jamnjh0R3IOaaclMd
YsMsQ1KsJ1YhClbGO5AaB/Td42JKU+Q4VDdkQpFk+YH2ukXuhrGyAf/ecWGuLtN00/bmkWHictVM
crpknRb/yO2PEeqbD0leXAEDF8i8ZmWufvtkffHnsMb/TA5uJxTH0Wou6ILR5iW2pU/b6HAOiTt8
OXH1glwj/tCewHK9gOjlDK9fo4L875PNn4JsY2jkrKmGAwenlIi9nskEjhd8NF3BhLWQQiRbrHVr
iFHOUk0ZnRNQj4iWJykcONiFKFqRhwEcMPx4LDsssDjQxOJ1ZKWPeLusz95oyam2XGYY5i0fy9S0
hK/7HEnOsL5ma5MimsWcXq4grvx+X4aoheW+y7gD2iKW/GqUQm2hvx/bCjk92sek0qUAjkbxhrar
d+b5P/PAtbfdlI80pSsL3Qma2BDvKOfM/5nG6u+eVrVIllEmr9kPD2jxyZGPvA8Vwm2u+H6iMMhr
70oRVYG08SPjmk5uySzKpbaN+s4AUK5H+QyxDYDCZ/u79nPoO9aq8an5IqcZzV+gJox4r9QAm/uJ
P9FjZLC4DNhMK5D5HWjwluchtKQ61a8mUj23WYXMWg6RdHd7n10sDK1oWCs/5eROWTEtRxgGp0BI
wZumdszEARPOe1fhURqSz/N4VW1eGaKQS7kOgDhwhXydrKvYJS8ZXyxH095wMgW5+v3CUGpDTF2q
ov7EdpTMrZHEJ9pRV0f5+vnNQT4t9p4LgY0fNMS9ZUDPktPjADAqUcTv/b8H/A7osDgygmw03wWV
AerHH1AlevVSZhaF60Nui2BSLpI7Fkas2m7uixxLsD9nfMETuOSVm5YUuouL6OHsDAN2uN4B0xoQ
qW4Ie7swtA6vg8aqu0qnN3RmaKkOvHhapw7ro65dzUdBIf9Q7bNzW9+cSGRQ1HD/Mrwh7l7CKvrr
LaB3+ep//jz1y2TM3fCoL1EUHCG/m6NgP5PBHOy7oJLKhxfsFT+n1Umd2E4XPpOMfhLQ7Owts/7I
p3G+QskN/POdG+h4CEi6I+8O/+3omSZO9m7nIkKC0mrweAGYmcZM6OQ12TeKizlAj8db4OUBSXnk
ZbUmsN/Y1RCVE25i7V7KaIvqQHjP+IB0wHl0DLfeX9dIFcBe0iODN9OOhDEKodcFqrZCdDy6gH+u
xjceAyX5QJGx1WGNNr59ZwICy29zln/3oaJ15gY8JHEJtse6n3e1TLAIDWNtvnsiPqsasal145/p
M8iYZj+mHG8R9hAT+ZQKeTX6jzD4yK3NS+OxBWhZBEAhVHZ0ieAbquIf4duGrd6xdaONkNsofij5
a2TBvQjUsO56zZaelrfgAyNt3oyt/dwfcSGWv7U+CoFOAPusyRCpd7USg1LclrAAnOoagcOFjAuN
6YlUCjvdW5XwoHOFFtKu3A6HeCD7IhFhv/5SaM7c7wnnJ00ItInvbcjmqder9buD6RyirQbxlH3D
lDtXUG4neCkaffGF91qQFEkwjR4FnVYm6hemi7/mBK+wF4PqLkzjDuGa0h8xq2w27kjBfDMkebXc
MPPUEMjndvPn5rttadXfEk+fw5lTPF01plgWJOogfuaWeU1aDQO5IrMfczM9i7BcNApxQC0FuRHc
e6xHjwoWFgH/fAF+QpwKPE+GwmVr3IOEMrVVb0etoMR7MefluVjqKmMlpODSKvifsAtS+RaAHOBs
TOQHWUAWZMoqV0R3Zyj0nPwtDBswgLdRQUtseYqWJ27d5UBJWNeQGi1v+pWXo9yBJ/HXsscEA4Kp
HfKnAgMfFj+coWiV7d8soY+f5MN7qHPoZxDbhlp7j62auZvF4KdREG6SH0XvaDi/46BO1cbx6NKe
Q21m/mLAHN/S4Y+vLbHP7mTayReSArBrQco2Dxm2QEnZyXT5NmSRDcMFSZceqoNZOaiAXHJBfFIK
oabcermfy/p4O65F01WJ0x3mznr5ZIwJ5YtDm5lXHGS4gfYM1XJhKCuSyetNTmOojdzBqOrDpAz1
HZokcOcHGQxxd2JRGgNl0kKArLMkbV8acp1jyTbdXwi7N3rqisSnftWhQ6vx5v0Z/5R6sKT0AfJr
0f1/tUoCVXalaSzK40Smuax4jKtWPIqofHh48j50Hy+2fNbVsh/9R11I7bYG6gFOor0xKUnocYEI
r5CLLpCA/RTgZF4YnPBGF2lzoh/cvHRDyrYBzZpNmB1efgAezP9sRg/YvDMNRR/6elbIxi20hPTy
J3y3O0RJqdFGccRygjWxxkQh1pPGk0dD9OGBHFER9x9EYCZLlHVihDorZ09YkM1UT4YZa71NAdqa
S3tb9/eqFD3Prk75LEbadR1ijtL2QVV+H7qpc3bfFe9LdFoMK/SZFCtUx4dB6Ds64yA+MiDOlzN0
SHm2G3RWPcnW+zDxBWrmHt5QN3hYRkcBDp02erFvi/Y+GoIrgcLOA9ZIMg3sJe1Gfh2668CiW7oU
xUqK/DwChD2tQFXDve/CWoF/EHqkCMkv2qYYm6LBL5IaOjyRD+OH5q4ZpS+cr0wI1PeIO0cbLYG+
bNGDpAAuXXoMwJF30URkpbqStcqXLsRR2NpoSXwXV1kmqFIUGO/+wXCt5iKaMa4P4xlUwn3+cSNb
nzrbJ3LlUWiTnQrvmmOK/h2tiALtjokuL5wq0ue8OthRiiFWcg0fYB6hRm7yF+0I5g3Rg3a6lgWh
A4Xt2wWCey2BAFi9W5ImL6LetFglq/4HjVLHCp5JHTb4VI6y9GYqNQCPjqAPccQz9eGqAEtz3nFL
Q1LGC5HV7FNqVQWmistrH4uQdQIqVBwK9TjSf+i8/xMCRcl8snBnEQbw9EXTrnwLo1irU8dvuKnG
wOuLTt4TyYdPd8uUE5bE87RZtiHIUpKuC6qmr6qxxbM5XoVG2V+n3C7f0p5qZaZeoYeyBsj9Whm0
yHOszhf6SUg/ViXzkNIGW9emb1fP0BydqAV0Mzn2AZZ/You4MYJJroMOe1pV0o5xKDmbH/xR/+Xy
6CrUHZLDCBelHnNgvGoA85IOldKfS0nTDKkQMu5qJAqHuLjy5OGTlqWG0QZUb4FbzCQQHOFyGb2m
aA5MQkUY31Xz/CSfYU/c77sj6omk9exgxREFpH/phR+oUwVsAZUL3+o/D7dYQTRanvh5HxWyD/Wo
Q/D8NYGcjVs9vWTvREo0Y5+n/hP3cdeLfgRmocHGT1dElEEMztAP10adr5xYRhuglzfJw8VTUE+u
LWmrwlMf/vuO6JV9vliaYZEokastYRYMTGi9gtL4zCJE4iQL1rqlEsJ+swVVNMdMJfMTfFT5jkVN
gMt2cNOejWoMN7DCRxw8ZD5lIYan4Wf++sxQAkQsFdcaGbQC8wn8fL4B3t+xZfaMGtII04ihhOUL
v8Bp+9rTCCZ1IHUW+AVmuqoVFJisXqI9cWpwUvjoukDDbz9feDhX8UknLG5yTO/QLNcT5wUVuLCH
clKYNOdWOcexSfP/pRT9uKtHJeZMEuFN4i0rH823SeJU56S0R/taETBkffH8MV/nywP83NqVRPMW
HI98s7kJJV5n0lyapa/FaFdms7NQZp8UX85ZkAO7tjaoRxze66pkK98IJPCyBkxnuNmlAQydxvQv
TW0hBUAmWMMM72qG8oNqYFWsdHqPv7NkkYmLOTOMgt5I/+zx1LoRvNDiTyjUMOGMZoGeCn4YZhyn
yXFZHUo7aCxkr9elH651T3Rl6JxmS7E06l2Hy0zXRTf52jsmCNHSjgcWyA2thF+/mVgB+RVMsWOa
P2U51OlNLoS4VwwsaeelbkCK5mYyvG3h6qJYZcANvQ9Z7Czc9dfgJH0xPsxRMw2k6ShyT9f9KKxL
mPXYZDTS43GPjSbt3D5DiU2UtFIZJlwTKJwxngGL90GZ613caZeBRUjQGHwB8hsJlDsMZFxhGRxf
5LjoRK6IH1JqOIEJtS1Kd58zmJ0mpJQiZy9qEcctSWd4QFum5YGux2NR3DeDgYcAY0UNuwDH1CMA
nwwvLF7902d1bnNPAcbf6Z9hVXv8NyuO9hrn8+JVmgIWMYHPdu1g1dQAHevWBxz3dAxU4T97aPPg
HDMW2XBaV1qvOGJbPwF6EApXjy2LMoFgGQ95cs1l87FY0L+cCuoq0/8yqnZ55+5b0jK5vigAg+X3
fmPWhL3Z16PNOQpl+3Vj071+lTTenQtAEXzMChx9AuRpywDoe8heO+fxv3Oqg1kxFZ2/GF/4Gev8
m5ktWnwq0HTnbqkXU69ejIkHIV58NBto4qQjo/WtsLCOz4/oDye/7malRRrmFFmWbiM1G/E0cpZS
a7N9fj5usEk0+s+pICpkaUlyxR148APF3Vmz570NXOKXd7di0IFQI5dVCaehxs5cj7qcfCAQ77zH
UXJvMk2+g2ypV18qfr0q9yG/ofee3ZaMb+Zxn0oODtpLd1klqJ690OO7lJ8sXWnsi24cc226UpNd
52M+lMwYJPXEf5BKIGnmgg/lNBwvQ3ZpCIGUhwG7yUQAjKupQjCO17nqrw8LlRc5oh/j3aDKEQMx
4FnOMj9tNni0FuLKOMUNnviiopD3aZVFdeKDqIm3PJ6kA62/FFjqAT2hX4khoqhfr486LhTOO2c8
68ZZfUwpJUE7eYiufLODGRgKWe8IuJc85+cCx55fGRigkd9ksx1QwfVPSOHU/rz1sPRqJOk45xMX
B7ivLBse7h+vVJG2zuSfY3U+E2WidoPcPJEK7JsvOQ1Hmy8G76kCaQHCmeBthI5yChl34x38d1Tb
Zn5jna7nbfSFcbi340uQuLBOFySNZa9eoK/1OdRR/dI8CT0zCdWf28bbi95FUnfHI6sD5J+30767
wDQ6j6H6xO/0wyXiZq0vU8Mhz1hgw7QXBJH0bAUWcetbcoW4OBIK2OCGkA/myjYsYY6apdrTj/Af
NUVRJtGFAqr1AKXF0kquB0vPUoxPAl4VwQhHfDfIC7vaIsEWO130YkxrA6rsefmHtsNbf5lscl8C
Ih1gCOulttuBCYlD3/rNwUMJN/9KROdCtWVktQbtHtHxDb4Tukruk28LlJZvCjm4Jg8uvQfpO6Ow
J+khU3vjPniYoanLqJZlH4rt3x3Tl2VKHDGQh4+Z0J1XOKhdFduGopkR4HizYCYmv37l0kiHrwBz
PZaoSNPDcmXv/0Ku+0geJOflI/KukVmXvHJJ4PDG3HJqQ8s5LK7beVwR1t1rR8/xsUwef+Vs7Jpn
NyKIHbrKRnZwYi0oEyLTv7TQU0MW/b3W7c+voVSBcgIjfpTdRU3Ksj25ZLbtzxuTD3rnIHwrTtRA
AHL9JPTp5b8hTmjhksfRjtTPvQvDOgobmqDO6Mi3B879h8EZic4ENun7ac5kDA6RyzoM/lkLzrnT
Mu8gd9cWVDoJS2/qHD55n+/OteS2y9IZKf1uEeFKG/Q2cpRECspplyvlRZzGIBUkXyOaVSF5VOJB
SDXucTa6fsKhKB9hsTxuluraRQTF2/phxkQlNHCt3kt//+UpUQTCiTIfD/VjoFcmo018Hn7MSxdU
mrZwP9wknA3PpvUcHaP/cJovTcT5KIRmt3AKBMxz2IIgpGhM/+0Rt5czlf6QpW0YgEns0FKXFP/K
xt9o28VKulT7BLr4144dM7b9e98DlprtgEL1rfevNbga4tbsDakphWTPerrAcZjoELXPIipixfCC
gOrUaCKnp8OUg5dnxAvXyWgMEqIpTT0uTjTTXPCKcPyVNbjIGRmQH5cFSU18GVApP9H7vrmfAuCi
/Qp3xp4AwbmAKnT+y5AGWxsvAWWj35y72+cVkYIyJeUPpt2PT+6T8/vHy5OetWmaQCbFoW+IKgOn
jxnVn1YgjVQPXsWV9VqD6YeCo3Gi3aKNWLaWuzLvwjrOaEWag6GAbfu+GqFb7HRi5CQw89uDjQsF
SkOQ6c3rWmJi6DjJtOZBUI2N6bSiHhm4x4s9PDZHFEnnBVey2JttXH2HdA8YFkHEDVLVzQh8Grlj
HbATm35/IFeBBzRhfKy/OAjtWDYs8WMu6HVW518JUoeUBt7yRSo5M36bSk7DTIGlmqLpgtWuPT77
EbEvy8KtrTMHefyGUQqTMskwztmeJGqp0ZNzhpPZvGRS1xXgIRe4KxOwXJgXkir2DdlbuhMikCsa
3TIvbxJh1Kd/piziuZjgHsPH70/bOXL0dUxyTLsI6Uebch/H3O/iTgYJkE2sUEahqfCQQCMS/xGG
qaSQMQTxOaB5RvaMi2Rh8IxjVM5AU621wZdSqeBarRiLTDcdS9EuLzZBKLla5omAySKk2IgHzNYM
nv1rjFrBBuDuCHLVSMKZCbg5nXnLmaW8XEcx2/8p8oW4nO0woZ0q0a9fKCJ4LcfVvjBX1xhzsrGv
G5v5ZAeo95goy6pWCXWHbj+VSKPhO5ZUkp31IKe4nxiUH0ezm64+Ct3Jv0mLbTu5e8+Yl2drabD0
vhxhkiZVXt7Cvm2+apFS2AZ95LJrm/kYnWsIfjAYetBHg9Fzm00g2/fZqDAtfem/Mk+c6RRSJu8Z
KA5plPQwaDokJVGr2oAY0pU8EmxCureljog2CD+dXtqAVewAWhppvNv74SNj+tqhe4C44Wl9cyq0
qgyxClZ9HfjF9X7sPNaN+YUC3jJnni4wY3OYS3EYXo1BhKofcfPvHhv7J6oEiik4xr2wxesb3KSR
joGUgOJyOU4z07QfeMwTkE/zSoN1/lN/vRrd0ECo0JqZ6QgDEYdqRvveAy/+unJYKi0wAasW7G1v
owkVRAKU5MpOj9RSwEEF7zqFeOsVVHxr6oxSKllQL5kGpkgKCbms7PzoQGAR4xy1xEvjMxJRGvRZ
VjNPfgXgNDqZbZfToQoeELrc45NtQjOpdKSk36932y6mrn4IJVmwRhjZTxnRguWPFnDa6zu4c8K8
1rkdOknZnNTnWYiksRPdUQ0MfXHg6qKUIh+CJISQ/YTqwiZ+1rw0EHlY+QX3c+KHnJ4hc3iipLaH
/dp3/bxSgElA+ouaNitb7CS3HzfkndHVFSs83FWAPIBVMWuEAb771cxcBR0fHpufCS0SeFiLsWcM
Cw9ulXvEua0RYZehxu6H2JVETJbDCr/asx8d801P5rIM6V84Qt3/RvrsJw6mw4sEjYzIfG03y89d
CzI0RCslM6WAccUz2x1pzwFLktTlkAfdSEVajI2I54LMWGHG1BZtI26qFi7FHRE++eeGDmFDFTWH
QXNCRSF9BNeebepxaazr0lIVXNwtL/FZcuZHpaKWQheK+aSqN9X7bhI8kVsR/Y/ml+8puaner+ng
wmJ+l2AsCbA7P54wDVeMUjAkdxnr37ECsbo3ZZzfXH+GqB5o0KErdxY09R9LY4G03bwdfTCvvbhw
gEHJWBk0G0+uEeD/U49BK9lZFQpA3ykFGo1SwgdfJzjlrQ+gUS8DkdpU9Rjixyjr19LHQWkN7IIg
AYvJyNlmlzdCLcZPxMdjMxbtk5JX7W+4rumrGgOw4zS/d8ZzHZAot/wcKt+6EbVChcNpg4nUpdnj
hzJtZPz2JKtjYFSL4LRE8vuUBlfTWs3Any3Zu5HOJsxpbNMUENOxAV2RgDfRfLUC/KWBAj8bzkiK
a3qwFTX7sG3YowNHGODomplTCEq1S7cATut/4vWkbMmsAOoK6rFLxcy+JFYcdiuyV5MM/uRD+pKB
ymYei/bpSa4u5ugmEqgf0wfnGef97GYRc+mIqW82JxuapbAQFe8VNwNLYDPvVzS4DiUWX2HMGM8n
XMDfqora7DVBvSPGEvqfeT+mJCdSCxsYCZynrfoKW9leZUQZYVGup/EdLM/UCeo/bb1O/vNggz4t
nnxLHSsPYk4XoLnxOmzXOQCFYZZkdfadScaXEe+uIWroMRInJ8BjyDcHAYPu7ZQeQN7B8jEF+Oz1
XnQNuLDTpFw1vqLC4YNU6bJP2J+n2SiNRzFyzxAF0/SJD5NKtHS34j971n8iE1jdH6p3MbCCmVib
rmq+IB+tGTmK3COCGNNkRDtwbcRWhro3k2IDBeAtog+Y+dGJPp7Y1cb5+wbTpEYykL9DeCyYXP+x
LMgQUDLlDbItK/XQkMypS6qI87f7XXiGRsWDQdAi0KatfNIJW+7RsuxhK/P6C/7CeZQQpMitNcgH
MVOKQwDVOI+NvOMnEqg+OaRGTusVcuiTwod5WB+diDVWWk4Rdp5ObhIzmSSTnVGtOtGLT/hilCi6
fOcl6PxlImcOeSWfAMxHv3R74Z1DP64nD72veSug0X6LKbn6NcamS5JAjVZHfhW5gxn47qJapMn6
JT5mw18xk8Rj+RDqeWAn6iUPuC4+1sqtvGPqFeu8Xg9byBjlgxydJYIYnAYoaBkBhri6M7/VBWvS
/UZqMKUmq+c9gYL7F2TMT5+0+ES1nHIg9b0DX810pNXFed7NIM9sO387Z+mYC2z4N11CFEsWS6eV
Nl+OLLg/p/rKqDJgk9sgfwg2SP4Utz6aE17C6zwFTv6GSD1Imbew2maWBmi3v5xSf8DngbvzibnQ
ta/qXTeP4PuzhCfw6xdixwk8qWflHFh9Z4rDGSQaCNKGvL60/laQuZPoaRG0hISvV8tMyqPFEpeD
8UzWARWEItySFx/ny1WAEMs6uTa5Yd0xYx3ZKqs2RgQeiNpDkT5vn9oEEdBb4jl+GE4AVBXjx2L2
hD3rwEMo+7mRjiFQKfrGf/vpHvLyZupUoBCAnYz8OUh7PJnnk2qnVjs0I3oabSCtQVUfK5mHJmdV
qSBRAh2jYzbziTvE/vOHevIl9JNHIkWM0cCqIOzpCZJjgk51utsdbrgcuUJYyYMzSuYb/5q4OWbk
tpVENpfyURqNK2Betj5q3t3IL+1Bl95pUk5jzr+zRu5M2C2wYIY8ENKHLomnts+4c0Y7ipJC8XWG
W2batlA5x8ykL+94SSFvUYzsdKG0MTXxglrp9gFmoxWOrT6+FKEARW1XYdnnM6SIiG1Q3EaIEP9Y
M7RuZtPc6EgL7qVLJRN9jUo4iNx5BPpNSmppFOOHZLcEnxxZ29JrbOL/LyD1N5RSSMJCd24dEO5K
U7ve5KNc/kPa+Ee5nR/qQXT/uD/kWt48KFhIRfhPRP8kSsdymVjA8zw8J63IUjEdRAEvB/Buj4rf
I3OMOadC2eYu+B7NkakG61RrvEAGtSh0QEITahmQov24IQDExaZCJdTnLaFHq4QtuYUVWkBtKsOC
y55IuCG/Ma6+WY+U+ccIUwKe2FpBkq2fMHE00mHmH+4tqRmq8Yoqqnbobl5iQehqwB3ZRhWkatPI
iwEmIS2rLmwnSUIVVuCvdnp8DQnv8zL2bnXZ7A1aAmyOLHtAPJv3aiI4Ef9tietLsuxhkhY2CS+v
tvJa5Y/ceKigbu7m4Ow3Gg3RkXtbjW0OTjv3J66Hh85h4fXWJojD7dKi2Xy6Pw9Jbtva6PdsOA8O
wI+K42FHNG5MXg0cNPp0xvc9Uu4EC0JYmL63VdP1e5mUT/hPWfv3K3UyOJkhGw044dX4KAsG4f+J
iJXXrOujLRIsk2T/cSg9L2rdPbBTTT42z07QZUU+p3jxeDkvEvf/9qvLHrZNYgT3krXxvYWwfhAv
2YE25gxYz+dhLnsfiuQEz1YJKG+1QSWvPAuPWXcBLjvDV5Sgk6B8ZqKt+cEBOF0WIe5fyy/lYT3P
4jLgR24xx285V3xP1i/RAuiJRErxMPa4H947IL87WjhJ5p/0/ZOR6UGd83T0QvqNk3yiOje98998
BKRJRD49zHPTpG9St1DtELZm4CcfGm4SOHMe8mN0jbB+pzxXxfJeW1Bxrwt9IegYHy8sqOIyWIi7
8HHPDy5Vjy7c4HPJCWRmNpOudFaypEaRvPOlVjkIw5ShtbianWjge5vYR81xtrmTIe2j7v8K5xLl
FdFZphg7YK4nd1ks94baNM1HWEKecH1HrIX3dwVzoeS26ghccSGWbCUT8myiQporg3UOcO7wYmSq
8an8u7DAGRUHv+swkPGWe1ift2yiq/Etdzbxm9qd6JghLdtPUr/VivEv0fa448IU9WbYmKBeVHax
2DkUSndfk8GWE5qwtAvWFjGQ5QWJh8qe0rZwTthVZJ9Tu8ceahIDKgc2X+IhTZr6zWFEKaVNjpYb
9kTBUOIeeSkPe4ahY502rPzGWe1RB779olnE3vnNBcH/GJzUNQc6Z4o+d1pBZpHB2KAEpa7eQbTf
BCsyrVdczxLBBVbCdVO+cvELxSkm7e8dCxcK60/79uFypvWsK+PsnT5yaxdCOFDWctCJ2KhgZN1d
JuaEXXKOI5Sucrw9RLhzrHLXmjSFdsGtEZMH1eOZNdJVboYARPHLlbAd6dYNemrkVR3lXB8eFoPh
9JXPrfJzCia744T86cwaaXOf+x1xhYDzp/E4HcEQ22jISGEX6ivvT3M+NntGBs0D4KF7Sq0Rfl7j
lJ8Uc5WdXfII7KVFpL6uN8tatT+wXic/D+wsMmvz9YoiBToeztSSwrPxoH0+XMsBbfKxRZMAE9z2
nqGIGwDWS+77rlTOFFTM91sRKbibVtq6k6EkUSuIrBQqKl9Tn7BNPF9e4qrQPGHQ7sD0KKFcI76d
UKeD/LOIxI8uiI0CGabTGuzFYrA97ahfiv2KVysPf3fE8c+ztrz4gBW7AjIrzM32Hy6WN1P4jvRd
NNVMbpotVunhN3Bwr2inor7CmC5DsNvlrZW2/l7m5wz7Q7aBdBj2H7Ph938UW5mgjI7DBYAoz66n
kHDGTIbZ4LJaxzAxEP/ejHfJKIvhp4GqtJSKN7zKjvjGVtYKAGcGie/uPcNgAU7N38CGVGyHWi1x
QYQ4sa2JYxCD4lU9zkCs/WXSO+3kY6Z5x2h/WaLquqhxoyDD88ONkoTrTLCZZ0PDCTKELrrWcdL+
1UnxFKy6zfOOTepcILQ7cuyPWPgWCQRNN2jwCW3O7qM3551UjgoT/UA+MjHdvQP1uqQMhQidK0jE
2LcoIAFz4Ipxl/k/q4ZzfvHmdCX/gwgiosHzZCmPfiyoy8FXOUpN822m4yyBBWpvfIy/imrxz3GF
2WUuTtX5uj5c/7frmGk/edXIHsltALOxHIRlP0p/CqUAWC4r3sDCafSgPlyG4Et3puvlIA4EYDIg
hABf3aOzMq3tgeWlP+j2DwvOq3vDGtARf1sYfxW8Vw1X0xOBoSRBV7g9RHbyzf5rQDzzLQzR1kDu
fhDpriIXRMYwunNKsxT+crMXv2xihoNP7ji+yVEMdp4utLyjqiPQqjMPspTv6uknuLwpv0p+vyqU
2XrBJIYetP0fsL3WkiCyF+XQh0a0p0hSGVGBTdpd9hdsuyruJ9hMD0KD7I4JkKUcTs+V5WhhVGMh
MAfZV4tfuaSfUHe0rwqULud7tLIyAU3pdShDZRxRhXMfwDzU47a9FAYmtPy0FBiF2meC2mkGgC4k
nWrrNVFCb4au1Ldbd4LAqxjXWumypXn6EB8uU6uJoOxXQb62eVTMdTNERKU5wD7LhSGTSNN93a8b
sJ9YNotrB1lZ4Wd6+C+36KzetzniAC7CCm58OImI/O6q8FAbJ66ttbKd0T+AVxQzKH7MTFm7hr77
POCFTG+Wn6DpIBkAbwObj2PaU0Tq3R9Tp6r15YU9dr5npY3BwDxNIz3iu4L017zOEWkwHjw5YbAX
MtA2A+t8QuwyiUCflUk6nlvjqvQwcqwH6T73T6B2mIvieKXccnkXHEmPP02XEzYN8d1lMZbpv1nV
XKHMOE2lV0fpurdm6Tyn/NUfG17RZgUmAmP29xNH+Kj+2SCec+P+zlydk7aqWrS+Xbb1ElL1q4ZB
WAvBkczgRRqXdZTPRjQmlUHnIHiIY+8DUN1qBGFBjTAbIpPKOOwbFK5xs/JgsHzNBhK11QgrOAzh
/3Hl7nc5aDxq5EAke+Hxvr2nH3wtZvZRHHRSco/87D660zaWAbbEVBl2DPaSAe/v5ldkMH92ABNV
ktNJmpy3aZxR0zFZ4xToStPu3hjRBMbud7dGY2gyXCxuQA132Estdzf6kWi3iNZgHe01iWo9k0XT
DbEnSDZ1cTQBq9mZfKQ6fDqIbi+Ftx3JTiixSkkm4qtMlDqWOQosw6/D+SEJKjFAG+9wdnsoPi/B
UfQknr97XXGjJkCUfiA63mH34RqCOd+3NU7No+hYfHyCmva4QVH4SDlXVp1cPMzOZNmGA0Yt4oC0
DmCuLR0tbnfiiFR0toMbsmZRJ4wc8OA8YdqwqJM46ATgWQHcNoRNR1m2RcDDEoKsfzzteSU6liBg
DFmUpLbGj47HPWj09QzdBf2g2sepJsTVFA1mxkvAVCAg7CKv8g/VaEwQnDhcAsP6mbiA/OZOr9qC
RgqaHLQl5zNBTOZkRX1P7LY18eay5XiO01q4vtKy092C+FszxHrlcEDO2dkSOMdhMoQJ3fntHITE
f6qd8FDZ6rdHsosZsbdXAxiDDDyJF+tcebAb8UzoTSuL3OpGrHhhtmWTzs1DTzmMHj5ZYmgj4C7F
+unFZDEuQOJkfX5sP2/B/6fTtUbfjRh6bZDxEsQBskbnHQpJSYkSCmbIwp6k00sBB+B99hH7Sku5
OhSTc7u+w/5Aup0JNeh+gOUT6m3qH/poxJdMaleIQk1FLnbxYULKtHDGr8oVgU4z3oR++V3BmGZW
Pzl4I6GfC6AdCMtT9xhxmvZgehaNKlSOb/rMBhbDrLFVDYEC852ZGauRFFATbV1YcaNAIHB7wH+O
6xkVa6gEFjH1YL+EFxCpueFDgYAjtPNLCsHNsttev1KCwFVpQjfDYUsIZtmBPOSFJlWDb0S2g9wK
NT31eUu+jPMCa/+p7UwLcbveNP+/tDyVL/d8nk4eWznbwoH8yOSLhLXt+WGb1Ftn4sCSHM0/o7MJ
ZAwsn/1KFxYJqiLEdfQKVzqROv96QILMDmJ8HrvpNijMTWXEdfUr9o6XnE4sLGTiuM236Ek6ZuVU
H2e4czX4wPloSWAq2USGJm3GAIgc2c5+L2qPPxo1RxleRuvlKor4kCQA6YsxRoeexyjH1AbR5iFF
Y5KcGyHZ7m6Vr9dljjsDvRX+8fh5AHUjxszxcztB4lAlRaflUsU5J1bUwVPVk3R5UpJKPs3sEVQa
itIyiC6iJDeDr0GdUdsgVao5XM+H6OJFe/9FjuxG/80yYU930ck/SG/lUWAGEefGUFlSgHUvJJF9
d1DfuRKcE4GWfNYhE1RHIktjF8AX/yhcXQsMf1hyMbnzZnUaJnaJn0xt6w7KzLg3kfwNyarAaIN8
+yE/2kAhDXlcjoUlup8FNZr9/VEfA3BuIWPyRaCQMuw4+fVcfz3isAkO0T23UtxFVNdHHRKb8EPz
K0zbC1bHvoSwdqB/S7FP0pUc9rdtQfZalAjUEju4Yb5WwmtINvCypZiwzZSX17ICWIfoJ0SlD9HY
dQHkDH0mcUr9EEeo+BD6q0FBf6VY7/4bAqv3mznehG/HfPgPIVEpRs2fc6CWFuL4s+MV3MP8qM/g
QJHhKbsD6FGqyomQKg6COyckUQU8jn5/T9IBSyLCUTRWKBjokMlUWmb4kWosc/CHpaVkEAAgrLmi
KObeTaXXUeo0dLtcXBcW/RtVLz/ScWkk3HPqSPwqcxvzcPXbq1pVleekG6Pwi9b1oJD+8q/Lu7kg
e4n8yyUcnenx6mwdXwkg0SYRzVV3f7lskiq7MjxWaMLnGbM/PHqx914B4tYLQUnEl6+TsPO5BvFW
8LbazIPvxBwC8q1KRzvVCswOHoNq+E886yGis6o3vCSZewX8FdCoyyKPxZlq80haK5tSWEnzlgPV
HtZHNdN5YFGDzSJpLwkTt42UY0w2CI7nVUV0iCiBgpcFv8THA1j7GFI2TfGMMNg+KDln7vJKVSlh
+rxO7TxZFHFRv/FNVdC7M9HYv+wMol4LgjKBnCglzC8fRI6kXsc/nzdkfTOySSgkibxX1cJkj+kH
FjPSAhmnF6VcBp9JtBb3xHclXh7I6e+xMDjgvGJ1h/JIlZaQyXdPAk3PWxCJKcBJOXsq03DMdIUh
IEcsu2Qd9mkcTcipqtq4GMpUeur2BEjfTMwlktSmFQylZmbnsdoIpAc/aKC+hWBJkAAFfvyIaVq9
PuuBenzwrlAoKTwMVMw0Vi3y5x0FFHNT+C2W96bV6pCMQWW/Lgkv7vySVr3cx22Aw4/M7Nv5b89m
JHOy/FMjhEjaGdsS6X0tl8/qPEVlx4FxAt8+reQeSi0OjKtY045qvGZLHMA4veOFDReiYK9D86P3
EfCAN2dHIJirUUCpgMYGjPWo0lDEkApfhL5maqhFkXPJaoeO2J4ER/EtnIXxSkzr+R0I8+M/Rre+
W5bgCALykpBZ4Ag6b34syu1OVy8tWp7um7o3lfDhHsCpFVI5xiZljzJqYqPJkyJrqebcyRzinDOa
eQPUb5Pwm2zdWKfZVXx0K5HmqmUpGTL5o9Y8go10CyECkAuYfScJEhDWQmtb0VR/CesGuKoAmqbQ
ltvS3fHRaZk0NRgo7TMSGX7prjg/HlZ/uMJrru1R/g3HdOMBq72kV3pOBX7KtGUxgCx6A0wPFG/E
yTe0TQRqC9G+HhZJwaes3gV/QDfbbboTxC3u0HLM8hnGrjpzMSNhKzPplzhM6K2oo4CqCHLUv7pv
NE1mRo1ZGWO15W7zc1jw0AwmxlVphdIs0yisBd3ms3zT83s3fLRneWZSLf5kK5eAB23bVV5sM2Db
CeiHpVwyEAHW7U5iG5x306GxaznggTT4T0UfBfyzTXgycW7BlxuTZtyTPNlcVlaFOKsHS6QXdBLN
z8C8fAW0SpCTcgG5WEufKruBatTXRHXmOKKHvpqDbXOTaHo+88ISUrVAIU5SK7gx3aEtou5QYEA/
FMinWFdTk+6J7OApMDJ49MYwid/b2KgZ2AyuMIdMyERjpYDERmAq+8PLbXU0ocyymOo2/bY9Vj/D
meUC77w2LYOuG+cUet6rIsKwkxT3lIkLrqMXyBiftiXf5C4SUMJ3FUlNsaVcRw30nOuWeEtgHF7W
IBXti8Is2Qau9nNnRwaK1BKP2D5vKR29KPLaNrgaBWVW/9OVCS1Qb61meFaCq20avNRKN8YXdJ2X
sHaZSZZLrC1Il+h8X+AaMp1KfhTvnccg7SWhtyCVL4ABQSdCsfwbQN0p7ZX1+0Kcy6P+ls4K5SYa
2TD6iFRB42tS0EnzS7SfyctGw+P+QQUOBB//r4uw56Q4m62jmKeVRdNHmqgy+cVabvl5swG4mMce
uN2TB1RK5ZK8YoAO3eHlkFrvGdxSpD1KhpO2W7+TXDo18reAxYRm3Jsg/7UvtSgLl9m8EwLlt833
/Vt11fWQLwV4cJQ+FPFXcOKRYLQQci0soQ3vdTcXdbXNYrwRKTL8COBCgV89Zucezwp6mFzppLpC
eds0vToOlPbKrsGMdVyyTtpDn2YzcgRxpViremtBce6p3FL7QhmqFTp6wmLJLpIYmXYQKKwqCxfL
5hLnjIgy7ag1aODNVWrFjUokmHc5i8jtpOZjuymfyyTgVKHPHkQM1LMInx16k1+3Hh7hOZsEL1vl
ANRV9VhS21GhHr3lBSej8wg7o4OZK90XdfYCt/d7geWPQK/UxZ2h0sKqdUWhqrqbQp9IcppdCzU3
M6Pwz7DCHORKi7saU7uszo4+BDnYyTmqJFQzfeQyM8SL3NXQl7qoqJLhm87CvvupWDlcei6W2xz3
yvMZLb2ovgSW0SEqJx/Kw26NoDaNm4Fg2HqfFzAu6dnTSz7BVbB6GRFNiuj7JphViJ4Sh9iN6Bvs
bFmSj35oeevuaRjCNvlgdKiYwC9fFonYM7LrhEzz83T5kOOsiuUZcQieyG3eooXRSV1TLrlFe+DD
CKGsiivEQ13eppiZ3LSuULzIypFg7o9UxzXLkO0PqS+T5chEwXjCr4EJNU8xzooffZledzdq/osz
e7kZqCBGsrkF0tztNax3WuWBbZRJrsyXHOr5eVWZOA0N899Q3V0wuqRhUwEH192JyYEWX2WSC/vU
v9tYK8nJGkeTbkZNhVOx3vsaKlHO+fDSCXGQlacd4SC3xAhR1e9dUsQqAnO0KD97k1DR0mjkvZ13
dA4J5GD+QvdWH7rM3t8jlgWmQbVS7HR9+C1B3+KAeemuPiyEL2BXLfVvLHG+rWc7cKxR8LCfEJ2B
j6ouNUp2JaxYGWaXNWXCOiGGzS4KTl+uyozNg7e9OpCTZ4OJE2D529BG2Dji50fYfIYKlM2+fE/z
ztwV79sF4yuINVexUkJ8mSj24kISsyvSOnk7Hp1HAVDy4nv7Jqs2jc//4Is94l096ruATne302VG
t1Dbn0pOI/jfpmXjNPweDfzwFsXElPCMiVU7fyfgfDfrhyr1i/taen/M2vEZ4alEJxyknmm/+8o1
jTTj9hlhL1gEKAaYYNbLdlDtr7QkMGjctiGKUWARhTvo00ZGoUyLp4XshCZUD3DdR5ar+Yn0trne
mfTIUYixP0OdPwS2lO0WDrE5MM8VOCZW1VLvFsgHmNo+4lNOnqGBOTEq64Mr/OIdnqjDGOEoobvm
o2GQMcXDuq6OgS6we9fUMbUKDhBtUfXzIuoTTw+W9+xES/FxcXHCUw7GCvQhE6c5pATIo79sAAke
B2JghnHRxhGkR01yxf6uTzhLY62YMmN+Uy4iF0yFvHj30PWxmXC/9Hhps8WUr3XrSc3VpljIpE8p
7uEX3Bcojy26wVzRXtkWW1J2jEe8W+0IVtO5O5z8tPVHWXdaoCYKrVIFzZDX7er7fcHAuXdLlHGn
dydVBOLWLzidB6O2LVcNjB3dwKFxF7u8GmCTuKFcOe96DsV+RaxWeTabutq1NUbcibNNUeC+9MVs
pOEytkNLR9Ec47mYP5wmFli0A7iwPcsKiHDolnACkCImMfG1trcITyzKMLPC7zNqWd5vs+M+XqIt
K8cibSnt3L4VIPJE6qGw+rCEpx5ZsyLpY0ayqsQMG/5fFIzR1fTQXl1OWXZNu+THZ6+wjZbm246i
TeygIfliByPAhXoP7NZ4DP6p5EnDPhQAoHMOQ2R4TFxyJCzc+TsUiCIwundzgAh+6UBMMYjWMhH6
LGGGwz2jEuLdwbBleRYePCIbL9y2qYos0CZzoszeqpW/kwdCvIxBeAWF10CDHZFZ+cDqaic0xMJ9
Kf3OiwSBlk0dSCiUoZWMSV4r5STSPNhj4ybeZAK7nYHgYQ8DZKIaRCcj+gToYvhK1rs22xttsBdW
UvSeu6o1lrZvIcQmJI0B5EvrmQVlJj756pL1Rb3DKZ3gG/OhpkN1avaLF2gtMnzxgUvrCJr7RC2t
J8nzHl4OdbpUNXqiqjFMGjXsy98dxdkEp25ExN9SBBneEXveaKbMb9odPWyD6pwvw3xP55NV1Wo6
4WUHg9THgF0m3efGz22CToJ3t+51XHH3nH8V7+L2U4NZ1qCOh7Tz6V3lHNbWnmcsyBa2ksg2Aizs
uXel35BG2x46Md614HZcJWGTXFAHJOO4ytAo8OQQo6ztYIUJW68hB937P44QDZwe751pF8X3Ovnq
jWDQoKxvxBDtzWx0deGC2kaawClPXnUi2TmSpMpfJ7gsfbvmKZtttyuvqJi1B8mGJtRCO8pBo4GF
Oc6pSxMBFO/qcdWuoVj5pCwG2alXVctn1nUg8cD2y/GgtUMMx4zn6dKLD8CNoMIOAt3d6Ckv0ztj
jXMMfzxqgQarQUJ4fwzYCgnnlCx3GCpdsxTLKHFsGNY1D+xFdTengghHa6eyo4osangZGQz5mNSQ
kkPfNc635X7QTK9aByyazBsdXAfiV6qlirZQ87DWgG97KT2JFLqAwpcwcmWU5rKFnOrAMbdJbMja
uQLxJpvchg9ZKgeP+0t82U3RbS7bLV5uKuS15CKarz/M6lAN/RH0cDi70qk9dYQKpVZgyZwh94AG
wyYhUEKcaVQlbitbJODTFQMYzkMegDVG4k58keacWXfUjChFdQp1XK5DXU6hLY+8SIpyECdEttYG
P/GTNYVuhekqQDNc0qh/yi5P36lJJMiCsjx67pHKunCzdu3Egk123lRJGs8tLv55xwPJZt+t97DI
3aGQqpy1+dxUyNe+l5SlwoYvh4shDgNA5sNdQK+ujOA8vUcsFAPFZppjjdxLdxoHFnDvA7sRZadP
hIRLVXmtqm4XkZiTp3mK6TWr2M/nsvNTVAcfhVmC5NWRyPNRqp7AKKSTXA2/C2d1wm4I2/C5ponn
KJq14mMPC3KXdLFotpAdQ0dlNwp1GfhexjLcONYxbB3GDWW8D73tLDCLKNlKfWAELdpNfWoRv6dh
/LeOdvyycbNsO/oWfvuaxXRZSl2G76vNJcETWbaUsw+uucoCpVSWxv+EDbrfazHO7AAmnBJLf7vK
ikZx0OHGPkvXPYjX4jcZEqE1u9jgQvRLANnicmXlKgYF2jz1AJrNmSmvgF1w2Yj7sYCek7VWJsA8
ulnRfsLtqPbj6Pjfra5u2XJxJNdr0PKDNNLOWBMK6yGKMpaq9HNv8OC6P+O9l0M9T6SGFXZ3/Kng
Wa4RhPBzkid6unmn7a4wrpbkxwnsftc4cOjoYpYvIO2E+ky3eP5hbcwUjyNZYV64d3w/dzYhRbqr
mg8oEad8cx7VpS8MCPijXf1F0NEijNdoXjynElbUh2wC838xHgse6a+9bAO0NpfZFLrrCQskeoB/
viS1sclr6oRJlwU3rAMhpeCezaqUSTDEu/Xxm4wVZlH64A+KNcZB3T/qOOAxq6WbFCl7F/AZpWrq
El6Ii7E0nddvOKT/rNGM7ISUWgoBCWmOLFMiZTxbpzWzMRbjcK3S5HyystWEZJYpqWZafIlZ0Vd0
fiBb29g/ciYHax6U2xQr6Mw6oZ65NkvxBOE1Ll2oIf5urnTTupAlcNeImxfQo86S4XI+RKKu1nUM
7UuVDs+Mvi/lBkOFmuNrynurBIW4wrpRk7p2Xoep6RPaSm6Au4685O5k/kJ7mfu/Uhg183jZmvB0
gfIYxlaJlbPbKy/peQ93JFA8wLKw/l4VOKxP6iD41QWHKE1oM0pGEZlm9Ax8yxIckRHQwDhbV3G2
QoRKRhE+Bq+ICNvTuxoCkrl8vUw955svQR2Kjy0InVwOjpFVL3utB2pqFVFOLTdanuSvRiTvNvoL
KcZf5EOOf/L0J5J7FaeZn0Y/V1mY4UjOs3JfK0lqyMXT/ev2JmcIRbd9SJGfa3bc0rdsuup7UgV2
jMBGlvKYxSMlWMV/Tiv3g5BYmUb8oDGE49mM0DRlg3GovrFk+Ldv12spFnA/gefsVdibgRrKJCxI
NYyDNKIu7q2xoBPuigRuQ37M2g0NCFJ8sQJ38OrLVxOlgyaE/5wE1t8ma24psSRf1+6je0u8/mv5
zK/wgJxx0kAnl3XStyc//BUb9oSl/cTaFIn4eHwpXZWPpr1I63ewe8wr05uYi3hmMUORMyL0AAOz
Ftd560YdmbZ40QJuunr9wgL60cdWK/MxqAJeQEOXszxh8foOHebyWuzwpZM9dTbgPeabPY0ngxyz
ieriLsYT5KdAazv6+7dC9ZqwjilFtvSB6nWp6xGyQGbnVL/lH6bl95OO1ovhK4nLMO0M5Ez0klRT
wp69pluvHCgrS+Vi6CwdzDYOpr14TNFdSIIkDXfNFEXM86Qam9toltWDt5DlphgA5DCr7eeSwUGl
mqh2907C5eKMM9YPr0z9EItZcKZvtlThyL52xwdcvoV88mcsXgjJZYW6W6HjkZup3pRsuBzhGm8s
vzD5IBlr+tasmq1ql3OXMJfJO9xqYxREKKmo7/W7CIi/9vcDy7yXfdVqM4SB2K53ffVu8MMk69TI
ykPB7ak6u3iRQXQjg9/Ef1ula4IMB0E7+u9OqMDD5E6Eqcyd6Yyw3BbRivufVUI9DKEaQFrPyjKa
E1S2igJO/VX0nHAx1Hq1MqC4egWKUWfuH9IsozLv/dBw2WUe+ot72xKfqHMuaNY5MECEd+BWbjNk
AJNOVwPVtoi/7toNkWsl7ILp+2YBsqP/CkvilHx+Yskd+gxy7Eq0b4UTOpqyRbJrt9GlVzfX5ibY
2u4H753YDQradYP0nlyIfNhSSbrNPhvB3veIJkUd9ZOnhSlqgBRV8cMUDqhjvcYETZvBatrXqN55
wKFioWjvCQZK/waymku02tRGHXuK0yf6XB8Lm+4mOpl28SGfv4qjyEY71fRl6KiVsaU//KIzWW8x
YSJR4FC1YHe6LZ2FQgz40bOlb3gQ7pnoSR/yI7jZicwB2q5PB1BG1DOToBZW1BtYJl7/XyX5Ctn8
Ateq96ipRE0WjK8X0ybCfNn+eFP8Tk4MHj8INcbNnGM1JV7yEmkqYo3zLSEPtH0tyYK0Ah/WAOBM
kCKTzMQoDU1Qa8rbuTSTzXjjSczM5n5s7Viva5Zu+W9fGoMHSx2iOANUU1Cjs2hCvprbksuWdWW/
YDn9bQ8mQkIQN01SOLeY8f47/I5tERbTblZl5jQrjN6kr1RgPz+hfYl6Y36IEM3f06uqLcnWXbQ/
bm6ZedTBopGxbtmyE1qqj5MdO15RxYkkUKpm+79DHaT6GEJAIPU4iNaxMsAJdycWpnPjaJcQ3j/N
pMIQvZ/OM9Dgeidfzp6zCCw+mtySwLK2QXzmbG3PnZQL5/lKtPYA1oTImUTOE8TdOAvbyinjzQ4B
B/26i7stOWd9qvjslNjak65a6s8nTtEnus1ovQCytfbLPd5xeUVTrvbMmjD6AAFkAUdniMghMh18
iihRkJRSdErNKH2Jmt0XJ0ApgQHHPJG0N0PG5gEBJpR/HFZuPrff0hCy26zjn0c8ViIpA+moHLts
Ur0a+LIuMSwWygEC94MGjT3LNUcX8NGelyoPOXXaxTqsvhXqhNnWLkYVk5PtHO4IhjWTq16xFZfe
mkkgCpuXDEwiKFgdKlf9UsxVZQBGaUMCV6IBoRaWozYwGkmukWrd0/wJAcCB9sstfjlJDBPGxx20
BJGMAYEZVwmW2Xk2BWoihYS3yAtyWE5oS3wlLuVKz2+17ElHH4++NEwmVBf5ivzPO6vW2kOf9s3R
BhOEzwzhQOxzUBS/8IIudx+RL5Uf+n/dFMRv06R/2DIYdkk9TgisK5hBmdjkQlCNE2c6S8fC/OQE
0zEXXJeaBUZu+v/18qt9teqd02vlrLvS5WMVHPXXC6NYkNn2Aiz4kEg2y5ZxSimVbE/iRteKH9aR
9bwoOvpHYmxX31okjQHrzNeIc99nNh1l8UY4cJsvaJ4En/bZQnJnGzo2JoiEp5q83Z4Vf+5vtoZT
189Y1oaIwLa/T6Q6y9CxnjWi8QoCloZT0CcJArsskRw83cippq6ZVUnuSItLfEZkPNxH6NqHGYOx
8+lmW/iV7V7GTW3VfoBje/q3OVmrrGZaikl0k++V3pIVUo/yqeyyNYxCmSmb04+4QtNyLeBltFhd
Lsdmdu/8Z/3btjMXOTAEevDAmrOwgiAFoMiD3T9fJATJ67KteYtWE718KULJMpdjxp7auA6HTqBv
0VzSJR5V/GsjSd934ReZBf/dPrQ5Vukcq0jlbf7NbPm9Su8sLkP4dcGbSXPmiRjJUSqEgeqSz3XQ
cfyiaCUNk2+49oPA0Y/Qb1cUi8yNdsx5s71d3CHZ4iGRHRu9hswPxWz6PK4s6Dw5UZNqOAMvXi0O
gWT//Eng4TtxtXiHyUxsQG6hpD6pIWY5+2kQvfrym2+rrY2JNE/U7bJI/N6JxmRbq17muTndMxpv
iXuTNqwsmmtdl4KJmkwjEqCTbgW/ZeHisVevdYTiSDZ6NtVpkijhp9hQ8rkZOfpI3pc33tuyANaj
XmzbQGQTzqI4U++yvBjeAVd173AWGtWdizEvRzkrbrInQGz30NCQdTlRQ7/KDskCgH4CG+UESwAl
btvJP+UZwxda79wIMIsGFVct8avkiSwiT5RfrSbXmIuyqKCFSu9WRRDNySHnPoqWwP6VqaC8Ktcl
JIExCyXmC3O2reFSonqnGYNxktKmNQcA93P8At+Wn7nOcNFqi9LbWygkpfFzRS7jv91lE7ry5OCJ
TnL+dPxd/rW/sqevLEVk/mor+Itkh1scvohlzGynWFXh6fbo4rKGuNq919ENZcZXX6TLymDjjKbS
D8TFPrygE+JbXblihmofzrec0EAoGbSwVmYgpdZ/kOI3AgsB6YvTrgXctT0ygvTgvRKEURMQujWi
j08e7L/ojGWO4KAhO9118H8RpA7h9L+fXcYd6DteeryQjUAPsGZWsepYC9JlLGpDKxBKZ3b/EURx
TI0aR17jAIyQYVcvVPt5xJEqb4xShYET+SjfeH1+/UKzGbs72AHySZ1SIkpgnOcZDBAYAxWHVvLt
hO+98+z/CZPAr+NGyqhrpVo34Rg4OgYoJHhda1PjY8idtZkBY2gjKPOKgDH3y5wRkLgedzjtwW+i
Ws9ges1ZZeRVoVQ73NXJnH3g+zrA3iaaoSf6tt1yGvZ4+EUdY6Ols9mkEq2cEawUXq13o7jy0tOV
pOsWgkteDQlobACi4NX/iGxkv9cqYpCwlRwrgVRffdp8/Qz2DgqhUbTukOM/1PdLVUY08vWT8D7b
pbkBDh0KuDeO5K+Q9HKBky3LFcPUGeoyxUcHSFDb0BABqGAv3Z96YXltts3Ea41hOb0JPRvJ7pBc
6k/ne+KrCjHyrEu+yYzGoHLom8jLrdwyTIGzpwY/DDKqBVwQ68V7+k4u/e64aWIvb4TSP4U7u226
xZlk6C1pvzX1vt11DhR4VEsA6D5cViQvYdhCWeHhNuz1Jic9bo7CbdmVos43uDee3gYhi8pSE9Oq
zfNbIdsj8N7qjzaYGOeGAZziN4+KiCGecTaybOPv29OSzUZOtOutfnqdzdj5QFir8oc1GfpsVaA5
AxryshHMpYXpAl2cwZws0QDR9e0f59aW7D0CWMP+PPRW/Zi5In4G3oqB+oARra68ZYB9tmPLjdk7
t5sSPGixvvqf/2Lm3+cQBZmuDWifc5R/ME84aYHD4TdEIXrEw/ewbbs2zxe+6KcKoxGj/VnoXYn/
PlIVd5n9+Cpwr5xMrabI6Os6GPmBAWkMAy3ZlDT6WnuWmtafc6PrQbbeAD5IGvsCAII330deXL3h
Drwect6zNKoLPK1ZxDCesRtA4U4GfGvGlsSeXMPZbwpGCWLzXN8AQNwK2lndjwjR7e2X8X1wvazr
yw3oEY8VCqag51C6rKbWa5I5t1rjElL6bLF+MgmNywuMRqCk7PBaEpq5FOUktEh92u0M5Kglxcx6
RqSATsUGQ3yLByt1O+WI0hMIqsrYFoGyFGLqjvbviy5Ep/Oj+ysYN9HrVC2y6iwlJL/YNn6kPpsO
UgBy3z4pXUqpjqRzGJpN39apIlLihUIhGY+AouMX8sYGbBuwqRuQuuWaxRBWllSnNI4xtxIsEF97
lYvgF4OFEC9m3JwjWd2yjtYagxqOPxSsTw3WS8QOhO4s/zxP267ex3nMntOgii1bPwrt3/RGupGN
oZs6SIUYnBq8C5Ng/f8ahICNIyoM7amctmp+QdlB923y+450XWXYWgDEcLb9j75Ru1ylGGr7hLuL
o+dmuCIhmxulWmyt3urxEiLY6RHdnrI+cJt4wPjUBDEyZZnvRllWn2nVViVA8r3P/HmDRD+ZmPLG
P/uwRfopFRyIUhDTq7DC/Y1d3fCyMUSCfDwjTNVwtMO4uR/WJhCv/bogn8OGd6ERYydzRelxgswJ
mxQkgz5ghVjyZhe3vzmOL/F5fBHEFPnBtN7fN4QoraBdbJ38v/bw0+m95xTe1dOmtakMUHzM4+M7
zvmIMXHq9BhfOEmtGFAibXbNjrghWgWNCHTIG+IoV/iuHWrNHvFsaJgH9bZA63oWTvcMwT2bAm7q
+yIRK/durNsdgZJNwdNy0laEcnUMTZ9MdBIguLUkCiUm3gXcDCh38qF4F/u7W5hLjqGNgyZbBAse
3LRqT0VA3Fo8u3ZtP8slZeEQHMBSEpinYg4OtLgwv8YugLapQzE4d2T4nOp2B2NOyYyYaANS9W/B
WKdQLn5Y9zx525KYWJCoS3FjOkEb76ytSmLXeS/Z66xpg7ZqIjm0UL7QWBqXqfV32Dt9FNQoqjxq
Ge+jTToZQR2+a4BhJUKCuAH/IWsOvVuSfXxfrSeadExFIrWFPRhCcdTGfIauAPUzNLAPifRn0NWg
FgAsA9HW4rhmBbsiR9NAex1ILQiY1ozIFtF64q8sBWXtoI7etmQ7GZ9x1/za0TEaa5USXvyXwXD2
wDwLqY6e4tGCOX/FURunAYptD2ic4K0kSDbp+2vVwQuJ/JQAFP/XValI61JJNZ7CeG0su/eqOW/Y
+9IaE0QgPfkyoaXkDPPfSZvTMLUQSMwL8rvNDMBEsrtk3DR7CUthubEEV68xVQ+LNAmXmQRUzAi+
5imJA6UcrIajWcG4brQv9MIDG+LFIEEOpOMd+EI6crnzbV8P7rU/+eWRfdStb/VNfVjsFhQAEY6p
i3HFzfk2KcqhjicOko0ZIHrEyaIVetrR2gCNzPow6uJqEI+N6afr5Iwjh1lrJV9JhXQrhJzfZaMF
vc5xfxBVPz+AsQhHTALUF4yjJdIjA5cvQXPC6GNDHeIJRoFdNI71pc0FLn4O2xr5gvYYInMBURWe
Ozemi1hwv3AVcvYDnLzoXsOh5euVqNBCTzujskzG3SDudyeN3UC7n1FLMEB1E0fQ3fBBOzji54r8
bPWYBCKSDLWL6SBv3zjTwFFdt4GSEJX6r9jiHTTlSaGU3HqCU20vd1pI/j2W+MZqeLUamoskHN/S
FoSVwbrhWs2pwIyzu6jRgttbxQQJkF2IjcaETZRhovjfCDeCjHPxPVzPhX3rDnCtFqoelcFjQng1
Ye37Eut7hyjP+Zr0zjyKAl+VvQ2tHgiuc723U8nFX47NR8NJQfzvjPx6+4yz7IZk9xSKXW3PIGH1
bed8xzpgUSMwXue/PcU3yShIF1XZNRib5mfY9u1iFlbO1rKlUdoQtVhAEva0Qa7l8WjdkRUB472l
/H7EzT+ylruv6oUlRmqyorKibz8K+7fuDCJ73FL6OALNdHhl3nlAAaojzY+Qgiofsui/KRzbdslW
RBGPsaPZI8+U2kKrmxsKum9sNsgGkbJH4KKNUSMJzPC0iPyYxgeptEmT10zFE4rfeco4G8W9yivB
1m4b32njlC+VrZnfbfhH22TQwTr4oiTj0RqdpW6oD6ID1DhQBNL8bYLU0wEIiUwkTooNOE/F3+eL
brxplkPCgWieOSry0q4qWe1DC/YOpxkoFpe9cBhVrkJ4Du/BbN6AK+lcWKKC8nic+Z5/qUCSNC/p
Hi5Wpu9KAOSiWt+ZwQpdy1TC9znF91U+6Ut7TSLPaAleP8cmnqyBpBEy21Kqvbsi0fjRcA9pNBQ/
Tnd6nIqwDfzbw/8WpolCroALlMrLUX/GtrUbl/uU0OJV434xkvkjPIEKVU/8wigtuEIl1OTB5m+9
i/sdv4dIVyEuv2Qp+PcwBXVsTWXtfpRwQBqYn60QiuxZFY/JRTWhbdy6te4oau9fpGjHCs7A5dOg
Q0UnU4YCPXkwuP1nST1pMyHAIJ3LI1/Vs6Q7WqBjjpWTOGmH6yibIpmclws0ipMhvPao67A2cvG2
+tYaX15G2ahC3rGvGRQjgXvZyJA55X03IboWMaCeS45CE4YxtA5OOCncSF8eADR8oN1ik77UZKLf
IlqlaOS49qcLoMOLVOdh0wQBM3NDg8h2VpMPpb0XHXa1Kw4t0SneA24xTdtGpua0mIeblmU72Xk7
rpNNKMeTtyGZJj0MV5+ZFSlK8F2pgtjDLhXCc8HqvIISkz6XDQscfGQjVcrorZ6dam1sHyvnP1Px
8kt02n2sTHMxyiImcuYakUBExQUwRGZrJRAb+7EfAp0fDPfxZXhQnCNKpdXQD9q9EwjVsKmoBYu7
z0LwiGgNwo+qTk33JZ3bgR/vV9XbwTy8NIcXHm/Ob19+o48qNq+vIEb8zbC6jB1IMNpNG/+8BaRE
2j9zCkG8+qY6sao9+2yF8ATgTvTmuJL53OqnO3YIjuPIxQdSklCpwPygJDRXWKfkbMR7U06Lw8oz
URbIa7ukayMWlvOuU646VXwWn3iXwpKn7Oyuw347FPDfqdV0FDM5VH8Qbn01JJ/kruvlRQCq6131
5vxjtonJw9qnNu+d7soLQDKIysnBkhUXDTeIojUAM9cYO26QxFdZRcLkfbUrb8LTPU6Y0EOhE9vU
8hv7rJKu4s6cX95jfJBX9eaUfKtY8Bso+dLrBTOB6A6oLqb5n8a+fJYf/QmPEKP/1c3qvzdOkbY2
QLGoxpesjVreC18Kg6tTUlsmY+Kn8SN/c/SmltrKWd5O7h3bxh/t2rZAhxLLhHjFm1hVVagBc43m
5lCKbFWL99pvXq2rlRk/9ubbXVy3OmAJE6n2UeouycHzErZ9ICv7MCXtCTaZHbcdd6DZ+Tr2+Rx8
x2fTiy87LJe0MS38qxipauFJnG00iX+WuTjGj+zNk3DbbBixkD3HXVTT854lyChT4+P4l8FwdjPb
RY/F+qWNkw5jjn+vTOJQUHfL1GNbmryqU1gZMO0r3lnRzRqG7YysPvhR1tX9aouEdMastqY8e517
iW2vwDaR5l8Bc9TvOiilxvPPNbnCCK6MF4t8ERRVLHDnoOhMTJPkG5TGP3G04M/2bS7BOuDsuYNV
PiZ1BsSF7HPZyYwWSGP2hhjZT6vjzj8BhTttS/a8yK55JiBBcVjglRdhWEuVpZ0udXcIS97iqnT5
e1JFIJBCPtOpPrW6AgaXlpYpINWCl47ryU1yyy4W8w6B3xZQOGHd4qN/RuNVqc3xbwFin7zvWNB8
qebCfbS7PHOavrzG7KvEML2PAwlSQy/pkOlhcFfk+fGKJVjOf2fc4FipQhBKHGRAYb1oEMZxM3Bm
f+I+LuHEM/s/jkX1m652mEce0Cw4ZfgS8ng76Rvdm/Z5yWV+vH+LZSYpsua4sHtOP0X8arkEXNZ+
L+vKNHRkLIff1PMlof73zzkugHMzsC9mcHVgp/S6twgJKN/M6LalVbbqRV3ZxC/prb14BmZpAgfT
Dev2B1puweM5O4gZXIHbwjA6gcvevD+52nRVX5h3dfqSQqWJu3SJfPvbhZhCiUTWiHwrvTW80lvp
htQ447YRq6iUrposDUI2cfCSq3C0Ni3hYeLAU+/xrzTTc7EiCgXSB8Sn5KxPB/yxDez/w5inlMeh
nxxfwBlrsjCP+K8SmmT+QLDYQGDuJn1t1OYiZDb6PI4pSM6fXoq5klDNQFxRE5Sc3Z82K3n+haba
n28ktnBre6mmnC3u9SSm6QfXgSWTG6E6zzVrQZuzcI+ILo+jODLn2w+LNw8zWy5mjoxsT3UMMS3x
VG7Ieg81dvd4sRRDwhBJnbdhwyIEEUw84ISt14PUIpbeflaVnh4Xt3cvj8Ljp7gilXfn8Lov8EJy
TzyZCKiOVTR+WWF7JRK5g251YUa8gYJzASmqT2hcLmWuKz3aeZoX3wlDmvRFfnddgcH6L9hhdrZ5
oY9Fh9IudDF9xdmtBpwi5y91YA2txO/htyy+uCow2rYCxk6atQ2Oos7dY/a0Va0BuLqZs2OfDIgE
Uz5TRQIE5KSr5hxDWGok5U0ZdxUQZTPt7Fj+82La6KgGAQM7m5uFb3Dej70yJmzThdzDMUzF1rey
IxoqjN0I3qGuat6EKZbAinLFqP6GcyeCyzcFt5Dqx0SsH3flyTQuwOaQUiZ87QLonVFCvN0F60f5
56VTclDVkRBzy9ty/2fXp4ETbkk3CtPaN1sz/ZZo73L1/c1MAZP08TOyqUN9YxzOdpRvUx9yHcRV
T/xmP7hUl/z0LzIW6NH08ANd/NNwrw/RYHn3ke7jCQds8KJ1RKF4Ep7rFBMPKQMqzMVkLxCj0fvU
V99aiFU9sZbe8JJVq5e/DMbd446ZbsRw3BjC7hl1Vg8O91U4FM63vcUjFo/akWvk+/mxU7NAZ2ap
ENzfmVZ24FVwADWp8GN46HHQY9h6B8d+jHXMu31xSIAuzVkg62hmqhRvFU0A2FH6vqkwvXbA+5QF
tayDAPmDqWngX9EbOLaF4NTkqqEh5Ll13NBUHhT3+Z/2+aGPaUa3FlRBtZL9LzhC/G88iIa2d8AG
Znn92WWCUNRG/qNi/DIvdg/PNFUlk8QWl3EDP2X/BrDR5SAaOAT42u0wszuetkkIZRabjWZokdoJ
0x2DIUUFMkEIElqTd4ZGSxmF/I6+LEKbFxfpxgr5eTYwhXTmYocSlZxLrxGjxYdr06yqDMyySLFD
tO/j8dec1xyd/dDRLhnKSZE9iHjGURkIftmIN6kjPsPjJOuady9stobmgEZlPemx7Us/O/cOLAQN
Bw77oODskC9KOQuuolg5KIaNaiOCTNTUBsp1QKa7R6SVe2GaslVN79LY3rwgD2di9/8gEod3+poM
TG7dqlxz1oTNODrz28XEYps6sjSM22i9jNODuu5dAL/z+Zd3Ny3RFjutmx3i1hHgJNgLbnmCcEZn
58XvpQOtgLKCTkUG/Tnr2edeFCwZMa3fkA75lDaqerf1nOAb+i2FGmngr8GItFW8XDPiFtWXSeG3
6Sm1AVdVzjZY1/UOVm1SVqv8JGsYtVuLEmvHmGty8m/Br3YBq813Wt71j35/eJJCg7z8NuW55Coc
RqRjcqE6oCMBt4/QV+pNu3AwJG2qRK6DJNqYDgDpWMbBxwNbgKtuG3NNaNO/4z5ynQxLFla/AL46
CD2OekBkszaq+UzYclIzwiKv+FJv3rc/v3nsCrX5DQLY8x8QL3LRRv2EQtC/CS6IO/HnOrUCgEm9
olHfZ67U+q6n3k2ndEGOHRr6zScfctfnXgGkNsgPXhDkg3DqxeSYjehSyAMjR+OUgtiMf1tvbzxA
rayTPObd45yZRXLwL2T0CWuFCNc0yiOyPOXvZAohjER+wFLOTuEXBlv5HLlKQAoUHpnTeF3FV+2d
LQs5Cryf7d/H1W/Bu8oN5TMqookCCWZpN7bQu2bY23g7owgGx1pBRuxs/jrJRqO1MZaRenhx6LRk
YIByhHryBWC5hkhxcgdYopRMFZZe9IAMk5wN/HcU/GhIqde4zLQIa746K+plzNUSpF6gwCz80Al7
bv5kGsmY/4DiCLPj0bVgkW5lS6ED2pXRHEfM6jgCQZDqqPMih1E/8/XIUGyVsQQwDoq39VJezngg
W3liGS0E3YGYrQrS7gi4lyxQfapHgCxr3BjeBn+tl78Y6RsiO85kETKR5a0cc7D0DJWoZtdCfMxz
tJY7GspTMf8vSuA9kA445g4xoONWSNPvdDdyuWP7gCA3Et3M6PXacmmvv0CSndTEdvO5VHbeIyBJ
VJT2bQOqjLpnM4pd551cZkeArUgwRQ5QsbALXENanMmKdtEk1fTASMMg114Yod7Q9OljJZE0xJbi
9az+c0yBV7Wn/Khc6oSqzYYlMfspFLwdW4JZBsTN2ZfMeNg3MyaWlnwP1igZ6gp7qtSoHYACFUJM
VL5GLgMpRYeVLOkyyYif1p1AFgvy7S6nLaqoed6lKx7oWi0qmQQ3MTtjtBNzpdvVUsfMchqv2N9G
pmm3KM78Y/yIzglpGBb6uQDeadxOX/Q0lH5vFkZymW/iq/tbM94ES0QYXicbA5YxBMF567TJ+Gv4
WSBhqKxcvCCEuFZTtfMpcEVQYjIcryrm6Zab5RiUu7Yt4Dnff3jOcCaxL1SzgmG4/Y2T5xuyB10S
lvslR+qS7m57KrZAxnHkSP6WU9LgMy0cFbjRJstCuiy3OuT3HMWnnpKKUpUVrBiMLHIWxYfIuweB
LgKsaDEvRQV/kZsnNXIGxIcdzQLhgIyjeDACE0oqywU5XZpSsp+BdvnGwMsENdiIyl+F3Y4MSV1E
CCGPm3jrJX9hPGy3XJlcPVVJHMSVneWIHKhSM94Vfrb2f1d2ljPN3suw7DywEPZD6Ii+cQWF+PuA
btrgK3bj+NE195Jj9/Rul0eILWQ/HnblTcnHAr62o4FbaIlQUJpGF+xJhxL28ypJsWQqoXOEI2zD
PWgf9MCInpG1oZiu0Rh8g+aT82P7nYwtUKXB8+uFq3Yo9j7VTToNXXzFs/uQZK6wmgFD8czLmDe5
ROQv9xOpd4VucYY0n3iKvAizhqTYn9CH+ydAeMyL76aF08rM9GTnx7UBw+/qb1/cRxkE78aJu7LP
SZJxYBFVjNA5AkLuEyFBmvfWnh3r46wXH7hl59ZKGn1UEoqcPONTuwEdZJbZIhtXcGiWofoayylR
VRl516fdHnFHe65k5fFJcqhx86p1v5298bpUKuHvbM0qsFOaErXCdqA4MqjxlsI7bdVanHPEgRSZ
JENHv/BwqHQ0KqczMxpNsSlDEeW70e7e+kPFr+loi4LiGhOaDoDUUoikpdrjaz9K9BvrzzPxkNHR
Us6iOomsJYOIkDYG7D+JUCFYNdnVYmr7Z0tHFokxZyhCbrMRlSWIuO0tPgeqb9YBV41SbIVA5zRf
UvZxo7bJVoyHJLUmfoP/nmaVgHMC54dHO6nB/Fx8vKjyUUTT6dF/6klN8WK8MFZKd4CEJRRSPp+p
RG6LZrANxeAmvYMZ2//qXuJzdHvO6v6nZyaOZ2tvGR4FN65jJ8iUyeY0hNroFr7VlhqLpqr88xJJ
e66M8SdwzWC4Rw/Jfyk2g4XLNWabWMpXomwG3WCUVaKQCKqs3Pd6D7bmVq/rixIYZJv3U9TL5uDM
dyixKkEyP3zht2Q5d70j+0QRPT2PEWP9Ug8ZLh4Tg1Fo1IfOAKWG8pIjb6TTNG2jnYVaQIQDwK+d
4xHCqc42966Y6SxcIuEk3JXOPLfEyIvPF0NOpxxpVXwXhv7v+7EyjsczMrHK53f6LkbKvGyMBsDf
HS8q0jn1dy8GltFacwApgYQUIA+RlAoF+DRXKpF/Pv0uHNVzKegC9s+OzD0UJkQkGkCagcbX/oGM
WWHhbmidoQojD5B+jEYphlMQaKJDlW7xLos4TRWz+nwqY3J859dTK3JvaWw9LQzLIFg70kwGZcY1
6BA+9dGGwe0D58lXjcvwDtohy1WFIMC8bx6vs43S6JGrqAFtCNu+iYHbYt98TQtJLrXNTzqPdJuH
K7cULoThRKsZs797NT3k62TmXC8UDnhvILqj38paVqgLbotbGfFBFtUXhRvQET0EmnbngJpYlZIH
mvzn+2VZJnLfPV6D54kUDx/CR00EyTDNDATrIYFVVgg4Ssw+fkgBzidDrN5bCvCA2m8g5y3gpfNq
XPGrxeckOs8SYfgC8/cswT+/1bnx/mS3G2cHS929+33mo0vYAPNFw/xyCLuA9nnKUzWSq2H9Ob0A
aP3LkCMFWsrJr2WIBZCTLfKhrltfWAuuiPcPC0XqBCykCX3udade20SIZWaCV6Ang1a1M9SVRFEX
FeMNzoI9o0othzHeaonVELkwZh2g7gwUa6+x79B0kU126yv7VyByMnE3pVhOXOvtHidyoGU5q60c
U3h+Ble2ioNOaJuUov0qrLAiBHEuPBsoIhmVAjEjRyFhfKo4EAh3mRPySkXHAWS+8qhARRfWlqK/
DNuBVt2C3ISTWoeDlDJ18BaMs8nhFcNk1VOrf5aTESJMnIhKuZA2fgzbKtiAfZAzVHAbdqtJu3Ul
TvCnneDiEX+4eX/kplUs/tAT7DyZ/ufjkjYlhIqg2BEoDzPIhU+H7fG3aTUYe6hKGXymfJmo606b
emg+DlT7/RnOWRygwb8RTKYaMhSgS7pnGTtwF3GLZTJrB2CD5v1MveR7rrBTsubB83ad10pY6y1d
DtRPKOl1+FBfHNXKISsjZcjX+GSr4r2t8ssZCLLTNg48EFBs5bHrZ+qlXQwJrum4FWo7og38ucKB
HqMMBlmWMuAQ8qe5dgwOr70otZD8JZZTfgHk/r7veaxaUO7rkyXWr/PckHBpYjpXe0dsnORQdMrJ
1F/rn8hVC4sBGyOS9DWQHyarBics+G0bO16WJcxP00GftACsScI2wolOE7hh1xgODrFvLQ+WXB+F
6TfKZYGMEYkXUIJLFAcyR6o5H/0MiQnUDziXzvOM0r9oKGeQltZVPN8EIPG3kShdiingbPK5xcyc
8SVtNAdlTBK+lGCeNaJLzN6ypQQ/alTvVl4mn56VoflW9nI6Bmi0w0bzXXX0JLxhaFynjAmAmhlv
9+/UQ8c8WqA3UYL0rchkCJx87khNGHmwM3RyXa/ykeZhfq0FAXVKB7rLu4MuGvRoxjWDnRRcP3kn
98f+1hNqFR4bGpei6vLebHwVdePHyPakJvd5xJKRYkyw9lvTVWP5Hg0kTiWc97wMftli2d00TaDG
jXiSQhD6lvUaLJqgMiovFyrskhI+xqb5/JWc0afkhP4VZQUPfnf9ukkhSDz2/9ET8bfxJuy2Bhrn
LpI7YgvjfVAeXNvexnd63s0NBtdsDcmgZn+34mhy0pBSjuV/7MXfMDG3bgFPKZgy0VR0pCMw61pW
U3a2ZJzBu6JZWFnbWlYZ9WkXXG5wHtOF0QYjRljJ/ZEz6G2HEBMba0R4LQSmXs274z8IG7ao/3x3
Kw4vH9s7JNsfDkfDsZUc6pE1KqPh4KgHZIVGNAYWPZYtEqSMZU+V/QJNBZCTrWt8eGECVM+Uuxot
Oln2HIubvY2J9Z4bo2HvDyH+4k8ReHvllxWtfHsGyAOSYyC8q/aAYHDmQLvrf5NBybcFJnQCnetG
3loEiUkErUc/BWYmVDsGMuJZIxXrl4DNLmkFe7naYsnPq+Mw89INrpmP6dmMG9K72lycQAcGYHQK
4ZJGiYPqpPUBW4uq1NtS8NxFnjHgmMBB7upRFJMFSwW+oK8X+ctPzPLFFHozax6mMrGmvh4P2CdY
zhateJ0IC8DxE5EkfNccX/fL9fReyQHMQiOtQ0QzyfkubVEKIghb9n4uSqx+Cdpdsr5TtRKWCvqw
I/T1o5baT60H6BUPQ6FFOuR7x6x5fg/6OUCseOav3sF+IobOIwu366Xg59N+zYiE/YubDZFUtZn7
4vl4oHR+r3VEQdIVJkcCagexxaycSWdtKK3ezBtgwsouO8f7RmNuXDRtQqoiK1lUJw9MnDhvlCLF
9d7ijiyZ4aCGQAGnTXtQt7uShqdgGP+XuXwqjOz5qHljU1s8Iqo4krSqZ2GSOtPxK3CkyECMjjpe
BFokGAzMJvey3FxB90dF7/43umypWDLOGHxs3pLokMLhuclW3BrE8pAOkpjcEGXWbfKaANnYovko
uS578LB8keMCQvuX5Bb/heqKRrXl+NLnrvHhYPoq+36S79lwWbS8fKaqU5LT1MKqa9Wqt9y3s7R6
jBEe2m9xRNbC/A7LebTsRccdoyw32hjJKlDfuVHWxQVjT84VFi/WZeHe4D7nqQNUV8YcbzlEkK8V
jj2BCRj//Q3p/joQLHjqgCx0ex+d4A5tv9crJVM2a+Oi1ayL7lSkFUyu4DkOFgt0qTKerDMiKna3
QqRlBaRACPHDMiQIPD8OZvDMoP2G5sKu1md+iOkF7glTY4gwUam66svzhV8I5T4ZQciTZeJttSpZ
ufZS2hxtiKXHYUzEm+R+cYlmBWcTbxZvisongt0ZBAHJ7VoJ10yVWexAX3Pgz+SYSTx98cqYM9HV
5pVWUfCaN2EC9HX70Di5bNgwnbAojRFl48ZTtFEk98y1cP6KWpC+SRbWoIdJTTkNIYHs+cj3NQV4
GjUzwv5L7zCNqaI1L7tdjJ9IPdAAFCaYNuuJ+UTOE0uYr3wUIY/nAASDqxX5JXAtu6ATZkvhv3YM
bT1dmqaEt2/MNITEXCORe58MybUm+Ln1/00wJgfDO5zCUIMvemfZ+Wx3SiNIbE9TuzbjUG9w9tjE
agC01jcUZ1Rr5HPTsPAXQzhA++DeWQfVCIYaI69fnQposq7Dzfmjo6YlOuetU6VUbRn7J2ZcuVGL
hey68wu/9jMi/DYlPZ0ImTkRgybyi9wIW3FkaTEHLzARp227ZzWvaQo5YJ7PZsim4p1SAwfoImhF
Tk6+64H7lbAkN3tLF/3+wnhNpX3H8XG9glt9kPPn+pHJ45TMRsub+UBhq+jy04sYAlthIENscJOp
YTVyjvnJr5hJDjjP/kyb5y7ScZwflRVaTTMRfGiMVa9MgK6eHhPNAyB04OdSNF1Xq2diuPfNK0OS
yzrWqWZ8HlYAL+e+kCLREanDWl6UNGcmfeEDTk/q6z0Oybsp8GGfZghJ8MFXhA1Xikd7jSUNOeCt
htjgdEhhi/O1nPP4ZushIY0uaeemvt/sxUIzONT7UNfXFp6qfGMoM3i606bsHWBMT7RBUxO9sEm8
Iwt5XPQZJFquE6VsusfTSeiBMJXHO4j3yPymO5KZCGGWxzFKBXnsqzynKmJUuPvnD8k3KclyM9bL
7lc/nZ1CAU2zaAW03YhYFdMd6HKNJIFv8EZbMzznhbWrdG3Btw0i5gA3+CUg+gYeTW2nPlNuryHo
i9mcRiNpsEf0iCdy/pIABWUWm2Gd34ONSRpWhMrbZ4qu330RVYaz/i6Z7E4nfWiztMHo7Lqiz2e6
QB+axRGB3WieqcTIXS+mL27O1TRBz+eLbSOy1JsjAmcUgU4QfBhsuVEwBOU0/0bUvDp9S/t0rLSq
9+fWycsS5qiTgUQBuDaqPfqlbibnZEOfmgswECf4mCxBDEqYQL79f98JGnI5Ynm2IVnVyTQ7Dcce
VxQ7RXYxAulnus9wOc8FWxlLBstw7FWIONPLbxde2DdzJHaPTgVCJOc66AEbU2+4t0WVI0y6Cx6h
5IWqk/XtzBiHfjwHhINELTsBEIqJpQQGGb3CU7dipGVZ0iAQrqdJSDWcbcy1tFZwknmqDEHFoJl3
/69gmeA8WuK22Jz2BQZ5Etof1n4XQtXcyn/2A3iaDoRHYZlqKEKQ26Jk4rFx5ylZgTbMVywIv5CI
BHzWWYqBHWSB4z3Qj+Zuk3enEpqgzWzD0McCcWVWI5pJpW/cW0eMU1BmiRguAUoo0Z5Dz70uLCZP
IL5F8nuMbrgKsYaBqsPemb7jECD07lvMPBswudi/znlhc/mUEYJDUK7P1J4Qitnk6r/y9oGHEkxd
+njST96CeYLCJx8ToZIwYNo/SsVxjlNgvr46mX5A2dXEr6Ac656Xp9cY+ni6mpfUqVCALVO20ur9
frHm1zcwDeJsbKaQqXwznYqQ0baIgNqKlHgRC3CY+JFdgMRhoSWTldhnFKlNV4raZ1tV7oqF3FgF
J/cFvDZw5nGDEbwe/0Oeik6PEGpDRoxr8G8b8epOmuuiicRTHXy86UvTNyDy8GUpri2g8wbvXncR
ry6i1BxvqEj52l8j8KvwPSMQUenJ2Y9bWvUtkXz88lw2Aas/qrmMyJ6+Ve50+2HpywjnjD6wO2pp
BbqpcvSGJ3VA6lvzkLuCinhCwy4tc0EQbI2vZIMWuDkNg2/VDNZE4Y+AscgPNNGE0QuhcEuG5yAG
Xl7gMJFNTQoqJPYz4HtSkslif31kchsV93vsI7TfAcAijoKEiMgrobBvbMBPSJKxF6sarYJokwWG
0D9ZKTVmnhHQpxcsSdQofH/juragXWYz4SVwhso6ORWZiWYbE+TmGFCFptTGLE4JUweBysPbBaJA
3ZZY+kjvI6IuVCcxr3TOlfRcCz6RsFYkloNzLodhMy15lwRrNYbudG6cDM9nzxjVD7m50RCRmuXM
I78R4vitYBW/SHRi9ZIJTcDa0O1gks0ve8BlwObJbZ5Th4qOzHLypE76/eMwdaLq3z38SdFvvBBW
gXfqTZNDOaEjWJQN65MLZkIK6tRvkgL7hBhXoGHHnksVlY3kprspgiGZqTfPpLPuu4YjPlgUxzi7
4qCbolZtKZ80jIZYQaSC4paEcArRSnyIKMCxdfx+m0SXlW2KV662c+oCvEfziHtMqdpbH6b9UayG
wdKLMIQ6K7mi1vvxahg4GwUOfw7YrAtYnXCc+vV0i0olFApgsh10rSjZ3WfKtF6mwybzBifFR0SF
AoqREBOgKr69iQkF4Tt829O2VY5oegikoMdXq9zQ06hQSN47WLouA6I6wru3TtPU02mMQY73akad
l0Vz7Vi59x3BNp1oQGQzqrF9UUxkUcg6Nfw39XP0S6TcwmWzNtCHyuxPUpiBe1BghncKaqt87eVC
WjRi19FS01u8bUX7JEwjMGCRtDCqezZMaRy/glqT5iUatFSXxtLgv7OkxwHOwZ2YYQOul2FFqBUD
kjD1LmZlMAGAaML4vc9yecMi1GkaF5EUKWyqQL1xmwSXQsKF+ws83LvS8SUEc6ux4Tqapr1sQV1t
YcDp+ZX91HqJRqf3xSq7yNE7LuguFFi6DSxOHZKhQ5UsIegoj4KDyhJxFvwTTWDUaSpBiAmbj8po
WkkF0AK1miLI6z2s/g3q2JZ9q/ehIncQSxnFfvIDC+8EP9eFOgdOSqYQHwLVHyXJihPzgt2IuU1T
B8MTl34EQSNIXP/TNIHX0XLGShSaPR83HtwsW3RIA2uuNu3K3GKXkPb4eDhijXGGNolbQtiBgig9
ZV/nTkrfPjrk+35k/7RiLEBKm9hgTJgSTDWl7IUoAtVfGDS06lM16S6VqCurrumj/K1kNxQxHVLA
bMG3BiFKp8RyIx4QelmefE0CL8zghaBs5CidAzgaEy3tRcG1w0NitED6u1v75CySL6Gkp4FVBA9N
on/EKtB27vLDB6JMNiLpeYFD7CCr4uG46RxwA+BC4qAsHBRaKyWeL/V5OugdSt/7fKdME4XjlvZM
SmxrKdxawdG8oGf1majPcD742xIg1nLK4VuDhaqDw7s01slVq86LKeYF7ZePlIKGp3mu6wLRQ3P6
pWEfJzg07ms9izeHiCziNCGpDDLjySnEccEkvdieDitgb1Re896RrAOIYSePVdXk/L68DJsfKmsw
bEqmGhz/4/rleoRjW5FdmIZuM9/QWLrUQI7/4Q6JTcil/mGANUaeNAEP4saDklh+hMVADly6IUJ1
hLYXFfx1iD8ZTsX4S8Q31rXVOFs2vcxZp4rQguxso63gUgv0QM3HBaqXaS2cho7wnfbc6dXws6XY
Mb7vPPPl1JK4sy29CBttc6bz6lIvSKG/FZnSa8JK3LZu+ex0BTliMJUcI7RgFnhYJrssCGSg+Bxp
5m0rLdRDmkdZJxpZYvNXV4ivobe4v1MClrtR0Z0zQDaXqSLGFiY1k9AYCnVF6h8uOrI1HL76e7Vh
dl1ykWd2Z7cQIIdF2y2SV62tuPHzOY6MwO559RemySPrVyaiyG/wtqlH6cDCDAGgSBRWChZf9Me6
PeH/Km0CwcDVxeZqpq3/qqkJX3QmOyoZa+L9fjVzK//53307ujWzKZVWOH8NCMND/5wbalH4CB11
bzmqxU+1hxYUpnimj7znLiWn32uony/nDoP0wJVd2LnzccU9aEhWlAm8rYMsku6cMDCZ1Qz38w7V
KCQxMmp2asWZF4evjrHeUwtRhqI8BjFn/l3VFaa0tZ99xyL0tKMlZJGxvbFIe7VDX77hiAqTQO/Z
G3/ils2Ltg6lx8IYRFYcu5v6V03U97D1mOJB4TU40oPhfmpBV29HCP8lwjWXfXmvpbILbaW9zj72
7WxHNG8hUaInM7Rsv33hCN5wEnrrKwaRv3WVleM2Z6Q/3V/aXzA9MazqxbOs9934XVGrq3Oa1yfM
2pBIEQ4vEskhoBEY4nvI3Kd4+UsEvq166oDjPjCnVdMoSRpACblDQD9usCWcQoJmf0lts/mjtU91
68Kc6lE0BldpDhIvhyWtQtsLudDw8NNPwEAhQjV4OKBaFNF9V3pwbkCiyCwM/kzLshKT36zEs7WX
y3OprdsfXMY4A3U9ce30KM4BylprYUtEF4B3XrEeRqUbkequBK6TFu5ZYb8xwYtJJfOdBDgrLN+S
WJdSSFzmNUrhmu39z9LiVKvjmceZAlkCG/K3yt/0DMOfh3syv8JK1HlQStHp4PJQsxLisDLs7ije
UILpxkFERj9ojp87m0KtcifzuyXkaTRB8CzFQ9FC4IkXVRKbo3SX9P3h0Qo1YmCe7mIUc/wh/xD8
jwsGTcO4dKqY2g1py+TLO2vuVGNJMj1p49gMecizBq8U4vbqNC+tleaegacxVs3WjNRDb8ViOm3d
j0JUblyp90TB+VyFijhu4ujuQI8fw4tr+FeqeVqXOZ22yyhU+atnKFA9NhtwEMxKGG9J3G/Mb+9u
FOYD+gL4CFX7Ivm3/xboNqk5+U1WfdqVeA2B3kX8ZbnOCJ718nSxsmaRAA2WeCFqoC+c/vQUrUph
5C1YJN3jjxxYyHbQpoecK/v4f4umxyS0xRMMnp6eduKFp24ojA+kzbW2KEs9OyZci9vY30FHRioh
ZNml1g+kpWWUHy58pZAbInCh9+q6HBqIUwqZ+MfTinA0xfI1c9r0M3Uv/oMqukQUiU3SDa48Q200
0JWdfHmQlOdq6U1PEIawebVrjkcyAyr79p7qXomlmYcxbln6peqL7S4aH0Rs1yVip6tOHnL3pvc7
OG7ar8vLDaPR+43CX9PVp3KxmIXFzohtdMJR7TDe/DkT4i53IinKll3Eu7Y/T9m2K20Cktowt/Ox
FLSxGm9nP/5kvtdrXrP9IPUWl7jr8l3fTVT8r1yIjNLWPfvPY6nAN9E6nXReIAfS00fq6Zr1f3UY
rCtog3gPJzbe4w4TPo4CpAssF1QVH9n0OJfEKHT3a/42ZiDG1a8Po5K5dyBL4I6P85YLsYFsfEaS
vt79hPvOMgBn9u61aKSbfr3uh8elYDAYXMBtsbC8VAPcrYC2H57j1PDnVNP9YS19qSE4s6ztH1Iy
8D2h2C06GDHcvp7hPTgba5+kggiEEyhWoQ2Q6Ih7uE4r4Uvo0jVKdWv+T4MpqtxR17dwvo/G4JYs
K2ndQA8Uf5gDfopJ2caj5S6rLVe5uObOtXnyTGXOBSe03HFq+V9dq7mSkfprrDdDeY8gPMEX3RX4
OHX6Rzi64947d4MhpZQ3jfwQwr2GQsTy9WltWN4v2sXMiOolIfkCTihYvIvtdnxSf0xwZRuROXPU
83HuKfS+bA+N7DJdlZgiGCuEqLJ1RFwknSDcuSmZclDPbTAOdgnNsTYbPsE/QYOKIUHSMKkHg7xf
NUepEZolUX4hYNpcoVzwoVj+ZJsc9MGwtAfdS1AiKN4MC+5uZaCSJloW7ynI7Hsjy1H4ERROommI
aX7U0HbYkQXBuC27WrgRYXNppe5ux15e9RuAdtcSCsHscH4XavriSdFeNtIdquXY7EVA6Q+RtE33
fm3g3HMo1LIVDtbmprqc8Xmcmp0OC+Mqaf6HUXXfzMZr+d0K2f30z4mmCYXpibIAq65H2wcY0nqG
4DowBsSZECLH1CXwJQaxm/rr7jbpczA0foG8LBb7ooAI6/fLSFoWfjmO34axMTlJYlyJRnvn4ME9
O1A/Ib6n/2yu6MA9eku8IRAxJOf55gk/SL35WpwPtQllPplai4oU9n04x0wU38A8J7+tYSgyH1kA
3/4eSvBrO6mXGsYxOGwYydA8y+mT1I+dwjh9GQ/32i+WkYoHAnz6EI8YZ+oOlS/hJuNSPZ5wJK1I
/H+kVk8eLwtUD/3vrfJvePLaD9oO9zDj2zD+jq85eBaSF6wmmQGLVvl50colFs4FPotOCsvPpGhX
NSoCEbTznVillSkRWb8ZvGL585HXklNAZ558LVRR9hTtvjc69IHxxi0/sf3fXynaUWZbYvHLxKAW
o9GZ8IcdekQ/d66pr3XxloBL3242A46YLxqlVPeuPyyMojMeEjZRCSGyqmeKTfiUWHrhAnW9294p
XAUP6nmv7vXz8QiJm/a9+70fs42Tkzzs5GTYYqg5UBSBuutfB/Edy0BsfU1Yj7lsmzsFJfDxc8pZ
mwFyJl7pCvK/40VJ+/bZw3WnoDqIZ7YKHOHtRK5TbOSiMYzc9/KQgJM7dHY/Eim0zTGY+P48vAFo
+UE4ks0DFvvv08M/4aIgRbD/w4Cl6jbr3oclMsc8akkG7oHaYeRJRphV27+Xtw10zF+/CcvJQ2rR
teuX8n8fxiFVZ9SZieOJnXcCA4URUV+bGe0cG3bBw7uuuE899qnqpzD825GZ2PPnll5ebFDDPUgz
A9ipZEjXG3Z7wEY5QmJ/fiRPoqrtBXr1eAgJmnYFq6/OLmvUJYhdg3io1hpo6yyI7TddjtsVapsi
F8F5Rteipo2qbSro0Xk6QiVYVShRw94t/74D2QlXw6Jf5Adh6llCZBUk2TY6Mi+6afuS+X9An8Md
zklPJLwtWge2JwXCOAMvnu1IJ6FmY2iMMGF3Ap2iBXM6zWPtNH+fuOZ4ETmXPmeWaY9+ufb099Sa
3Z80Wm2rmfIGiT3eRZg27xxx+XbUzubhoOTChtwNA0EfiN7Jkhx248I/p+UFFQy6OnyHXCJw8CJ1
5tKb7OK87Y+pwy+ZGAbqRS6UXeSXd/0bn8QyGyYAHE3Z0yTwxvCsIJqgu0Z0MQCH2ANhAItxwJpN
UNRDo9sWADoSCklKFNSK8HRiMxorhMhX/yRY1ldIiVijmBq5pRGlqndrFN+u4dVe6rp21gafngS3
fxNIGKCSLIb7vo4r0ms7jI1SS5CSA9lyaNa7HJTNusGpWKXode33ixwktQ8QKT18r1AeO14x55TD
U6KQQRCgQKycQADtPJQ6yg/osgpDQGJ7ZmiqUp56M372T9uXLJKvvwXL6qanpB/05XuiIrD97MaF
RNuFMhuJiH6WDelnr9FdULWU3mnBymzS7UsB60pd6NfvLunjP8UdCgFGknjaNt0V5n7XKf5yZczF
jl5SeNNXd+CnT70+bvNM5bQOUMm3u4rXlrP/DwIsIBplSB/BvOc+AQGojmjyVIdamlhiOpKBiTj+
ICf9aJ1plA2LFac2pGFo+Fyo5v7QcS3zECWyaG2SPy7XRzicq9+QqwQp14NVVOnLM8A4E26p1JQZ
7/y3lV7sJNg1NyS4iZQu3x+3wHnjulkQ0kE7ybXvRFAJrx8j2XRQtieM4vw9mhgRNsa+HBN71s7U
CQot69YxRIW/wjWap5q4BmOu+rtDylcQfSatS3CRD13yTe2kuv/U7HRE4WOga1f2cDQi8zocj64k
oWK7bCgtl9TDn2L2kJKpCoT9vHvRkM0bJ8vpPAoJ703q4/mgM1V9nTnJpyd9q8l7oSbbnWgabfgC
r2VD++Om+U7pmqHcK0GkCv4m4CnD5q+sWKncPnb/i6XoCoJHKf0WN48FM7mpHfB6uL94YefWlxQg
CQiCIlM07g1OQklAXioTpgM7D9ZU4f3GEdhWPDxC5a2tmclgJx477XtDbsWdzrweQAJQTv9Dk0XF
cj4EdTyXsbJLQuTQ/lSuRnrnm4pmgL/Q2pZoZ1g3vUmdnxzh0IShHBnwQJpOEXaFdhX/zfunYh3Z
daAa0fQMUPzm0nnDhEicgdfqMNwCWXlkujolpCeUqWw9LBdlN5Woarnz6n7XLM64/XeBYmwMQizI
JiWI7loH5DXOjsH0rJpkZSVW91vC/80AE1Xc07kx48BCqFdMXwxuuiOrObLEId0hmsdtl4ktZ1kM
ttNBkGyH5FBTPE/z/64E1rZahT4ItWuzDkNYShGlKc5w02W1SSM70K+9lNaLuxAo8+r7iH3LnGDT
ovwLH8uL5lC8BXoAeDPY+oJ+XAKaybVn7vn2uW5tqSIWWrx4UlRj7LACfm8npTjLEw6nc1NStOod
zB4XEyl/2jgIQKm3HnKrM0pOM5lanY3OyVW0PoiqhNYgADnQJ9OHJe481s1BZ29cIjr4KxQSsBxk
O/2inrBZ2X3yCN3wO9r7QS1pJbsn+OTXAk8fCpc56pfBDYtVDqYRu05oZeJInNrYBYUwg84WZ6GP
7afl06rCuidPeEad8t9JZ22EKuY2lvNbppSPaZffej4Fb0zOi3wyDFvsht1F1XFzdEJ465Zjexzm
y/oHqdyB9xjWZLy5RikXXew/2iw5FnfWPNsazSNbo/K112Vsey2lVoPoFp3vav+xQtDDnXlm9BFt
gI4lz7OA4Tz2CNUsidkuFoJEJc8ZIBgvYC8mt3PPC3/Z9jNp5xxUhZV3AEz5t9oOHFVth1J8vYct
Ife2Z7RMUZaO1bmTHlxeSRn2QUUpec6ggFwt2WJ+u0btRf0fZBztHzrpsP2O0826VFCjZj86OTeQ
chAMRYCmoSxohc66+FdAAlHd+YwlRizm4bjxoRintt4C4ea6Ek4vNQd3k07KNY3zrIN5DrGWYgKB
d6ff/6HkUKTE7Al2mfHy1zzXb/dhlUUzBedpYTU5uwKgfWW7Zace5FSLlhmMhRsLYAN+4FW3sXG0
CdFrakTz5dFJdsDERiPc0GW1diC3CkvtHaTtRhcgGfgsvU+tJa3JjPzb6cdeXyijTzCGwclq4D34
uwFQNbpLGhnXPoT+T0WYhReMms7yEl73VUYRaPQQzEztX7v6dwpRze+Jl69qEOD8UyggFn3EaPBe
1SeQS+oP6PZEuNEa+dJPFuVmzr8zKak5VDiUvoJQ7xq4N2WNvHNznr3NqRIiQ4qk1xMEpYqivRGG
gahp3PYXdJPPyubKKGGcmphBoBnQ27PiLtLBDgbI3VkdGkLKWywqFUdv0idhsrZGF3DA5o5O+4VS
2t7IEoAIMgqV+7jGAO2W9RpRS1T+q1XHZNUNLyC66CYTzZNWJqZZplQYLNyoTCQt/eGUlodrvP/0
ok9ZJ+3z9TdNg6LrCEsINw/3rIg372gnxz0n13LccI/gvJonM6UzkxNr3eYck/0gx9FtSRZ4AS7o
2zTVYmirCrbHbIBhVA5kzth20IXl7z9TMr8kWtpg3y+XOKwk1Pn2f51CcAvuWDbEqzuTjKyFE+Zq
22st4JIdNG4mWJZR+mBzrKVLdg1ouLZji9LExz3J0RR38LBPJ5KKTXY89iMuumtOgtHuW3syMgtl
bebJXbBkH/T+zDisATTygMQmfPsJEjAbtS/H3RZN06LfWn4fd8pV2YZQjClPCBZmsVPUK3XS8sEV
M275cmQ9XzZ6ibVJgAlwZR4EGn5n6sF1Ezq2rBEKrOXb+Oa1kB/tvyNB0vlFZR7Qm6xBP8swNJGI
o/1hMJZ0HZuDs5QlUME4sbwJ8RrgfS5G+44yCDgEN7s1jUBDm6BbmfLHV/YCchFWZJiYhyGxCsld
UXPbSXCgvwTJP5UofPOWdbDNqBo24jo194D4cHRV3/W9COT60FPLUtdiHAWr/HBTlvuthan+TaAJ
wxGMbs/Wc15RbGzPxXZx+qHoEsNoJ0yKSkwbvSf8DyQEmBYurXriQU616RpfR6yTbEQYaAfdOtRJ
JkmwDeRPLlznNRSlme0Fhs6J35mnjGawVnekWWPV1PemM088SXKtnIcCrQ5mc7vACYuV633Lx1rh
0Vcvj8h/YvUPG4PoIE8ksyc43Rnbzoow8G94GMJhSCTK9YOKtQEYNEJNkGE0vjWypvrVypqwImdt
ZVrJql6aJXgznuWoDCYTMGDMCm5zP5rh3yU0/Xvvow3OPfgO1+7bKlIxvqW2h0cUvL41PStpcTOq
u8gFQDwQvxDIfK1MEvS6R8aAnsh2fxfUn6ELAcuMM5wpFffb990oeO8caqn4SCdNzCn9Xd+lfc50
MciUCJpcWP46//tknTbgyzeQAbMRDUaCQJ//84Nos+84YJ5OVACQ64eBXHbFS/qyUXn8VPIYHOml
dSeCrd8P1KB00MK4+CaOXJpaYpsF8mkl7+DrG7hjFRgNvhmRc3QMH2foH7CjqJo6UQiEEzdxjxEt
7YIq7y3DeEs7EfyWD91UOcnKBy93nyS7RBvup/s16YbN8+RO71JAqFJcqQEbc4P+NmbekQc4Y7fy
PX8xM9bqaMczLF/5qa8SIYQuIiC7BzdV78brDZUQGP8MV3GGMMJXrlt2XVn5Lwxn0XAEoIiYob28
ms6N0uYjun4leWFOqLgL3y9GH7h+wFgvXu/4rPhmbc5Q3/MhRVzcsYxQpuVNGZ8hO1QSuFl/0TXA
KMsnXfRN7ZI2mV0Hll2FzymTdJmgB4bDGJg7yJPEQ3+Y8TktGjP8cncbIr6YpvTSyRQbDu/TLXKH
1u/EGDUQUApcaaL32DO0FlDr1ts5jGkVIDZDQaKopvX/lnQCn01nSPVWJGDOTf0EIoMzJyX08Ry1
a5f5HxoelY5UjGTKDuBLD0s+p04H2r8UZWFlZ5cXcLU8gwmrUCkG+bKlAi6SQAQavPgBfLz9cP09
vnF9R3HTMwV/tkuuJ2Xj52D+73G8yzsk4AgVZH155VeunMWZS+rABYnzHIyPZ8PM12wu+u3/t3F4
mJ1fakivMQx6g8yIlmWTAg80RnkquPS/qOyYSRtXLmDRtjnQa/ZCpbUvH5kVzbxOUWMw/8WVYDwm
y1jy8d3Zownx+Y3J/PePYlyuBxNAuqXA9AkVFCMKx2c7cA2QJthxV2B8DNGwQpNFyWp6WVlqo3OT
A2qr1yWwY5fy0w2PDMd9VrpoMky8Ptmmw/IpMCDx4tB52fNLsEB17MNfa3OpLz3MRYvx0XdL1URv
ruumKQJFXV/soG92G6tpkddy0pUcxieTUwHFjjd1keVxafOpS6ZlrV664hZz1b6ft9rm4sWHKm+R
NAF4fLuv8GCrS+TsHUe9X7r4SIVITHjtNMj3lWX8CN4hMKlXd59CCfYPP5gWx0NHmJ5DpqnWaPz+
l65DReV9UPQ5u5/ITR2GJXAy7tjabymAMtWMW9aYmNs2dn1Uxgdsgsrg+uf1nngDxW26W1BIgiKX
GBPsHAr1ODSMmZKHfJnifxJoD5pbtY2AD6oMtHFOKpHJIouml1mGmtejcyfqw2GUQXEMZ2GcoZ1S
zq7OkSl9X9kJtIcMgnIjafbucjwB73Z2BolntQidpcEyjPef52wxKkOEyNI2JPx6GX5+j+KakHWZ
CjDnBOGD1bQqVX/fkBZBl5WsHPfkZ32l+3vBzOprltMGFCzff7w9r1pl4zrHA6MAsGvBZtRu6vOR
y6WDDBely7VAWZoLr3D2A65OFhFBXokIGC474cmJajrthqZQ1H/yLPtmZhKCbMUSu3GfInJxAiC4
JuvRyskxFF6spJWnZhHgZtE+yqDae5N58UcN65QUhanJjd7/L/0FZG53/s+BN9kllso+m5lqMf6m
WhVLpddqKyurCErgDVQvkMLDY+olur++eANnvpz5Ej4civk2Rj6TCVhkU+QZLU20dLkG0fW68V1A
RaY/2Zk46/xbQ77EBzu9fWQlxzSHKPJb1uZNAhjM9DuN1LH8jX+9VJyTCscP6+p6d2o9aI6KZP5X
nbqiM3Qxv/YX7S5Hl0zagq8W6/0oSUmuzE4JX0vJ0rnKlVv8esyMA6XAaCMeTo5I1ciN7Ghc1A5o
m4X/Ro9BfAfW9zNYK1jGOaCKLgz/X9FBbuysvUGCz3ywvH+wjc7KVt7sr0u1cPWKrmrM97z+lQQr
ZJlVMA2mFL0JNPkdNba6gKfjI4Sp6BPps/uuo2yMVWxBrRqwFbcstXI21tngoAgU1RJyzOCAokHC
327J9g4KsHedW7juvNzXJ4ZN8y7/L7tY5NpJx/hLfONNfiC/1APVb7G0z06iv3YdJpMO5W+qmmRT
RHbJN7h/Focbsqo38YfuiPayoAANVdF5BxhTxiHf37eOHXGjX5YF2ibXr0iA8Wl0UH8WpEHwStHn
2MuFDJtsRQxeoYTbfnAS7o7+NGsWrFuS19qa5UoXnvC+cnz7McHA6gJ/Q5LTLKTv9vvqQCe16VPB
Ri9m4NwyMF6I4+rvfUGTFd6MbvdayYFxYSiMuhjcyDpt4oNBG4qxYdjnd1qwbDPc3YnEUkN29rfu
ZQHRy1bnPZ6yq5w4RFRfnYESjz1wwm3Z2cVgbPyj12Y6NsFaLY74FVB7Pb8qgmIeW4SwGU+ebdD/
xKzBbO/WInmc89ScvP7USsckHGvARn1/rcd369nX2YB3hz170gh63lO3XzQ0AOyDsCzUL/LLTSIG
eJhXQL2nqKhla9IJNCy/Wma12CK6EdGvztZG0HgT9twnT1V8v/H7rxrHAGowx6apRycbY+sg+wP0
eoRlbxYTNoPlArrb9FuiRb6JtGTbTa4Guvk2uL0CM5AxS2FsC6X1b89kyW+yyNEbeu1ELi1q2kJT
eHezCl9t0Ozlx9Ini6Lc6+cH/NqOBDQnlTIGJIwINnGuo4m6ipXf1D/8bM1bvQWN305Kwzt8M3bB
3Lvkt4x6PQAW0MBHgOXQxcRx2RscMvqgrpuTts9bEo/jEH+ehquJ7nQu4r4B2fI7tn7yTJFmLIFA
248s0kHo4wS4p9/GC11on8idP6oGLfFosTqiK4lCcePR81bPQ9gKiWSNKtUiumKm4JvtrGKaRp74
7g4XIaln0GJwXVz2WJL6Q2Pu7Th4sFYbYBo1lxAhVKEOGiPuEX6mf2UBnRKb8OWeia8HtEyzfYp+
gkkaGDSCuNUJNSSiu5GQg9J9Z891zPVVi5l5PEnR/8VNBfG9XmbO2qnck1dV7xdGxc0kYShg+eEJ
AnrYMfUbeMxOfgZMXlseBwNQPKyRyYEfkiVTns3hXedHO5T0Nb2JnGYYJJDX/M0AwSDtyKFHYrBc
nq4um0Lh3Xrnxy+8mD2EAho57PKxsWzzm7A5T9fPHxJILJHJn9ZcdkSds0fQ2Wl8CXgMN8xg1Pkb
VUXctyIAPaQ4gYTLTxgsUJUX30Vc1NfIu5UecpPNulCssgQPw207FauSDuR24n2/f/bjnVygEh6v
wwwt989DmtbW10TCNKWMOOz17ilEiyj/6fKTskDG4VdHyj7DkX2crs/njg/yQ93JTZ/ZcBjsdguR
ItHxMRlxKoRGAhq92pQf9gCvi9x5miVcLD69+Kvog2EyqNGzGLVqRp9ry4KoUBviDEcTyyV8WyJJ
Iliqs2jY0101jPrL+qXyX61jUauC97AM8LhehlR3q2I0htBqoSfmbaTDyRNncSvmCcMvqIIwn7bu
OlFueUxyGPvrTgYfoUDhICeeRbSg9nX2UK1VMIFZZe0H/lLj9MdlNno6PmlAcU46kYR9Dz3C09YI
uZtTrQQkxntMGNd7cil3a7dZ0z2oNacYLgbgkFSXtX2p2S1GJFWL4iJzRu/TCBQV3q7rWOUq9q93
gEIdD4/5fw8IFUZmy75IhpK4k70LTHIKj1Tf0lOkC/ELr+iIcJLyAgjyS0CQbz8cmaRZLROMqKVq
wxgZQmkowQxerKTUIE8tXui9a1WlSpo9oRNIpdxCPtOyLZdA6JLNaR2J5m/CJIXMggRTJpXSPXFn
I4bPl/AZwsvj7JsqW+epXhD4ghMFTaRzk0y7UbtGTx4whLaF4ajRNU2o+wg7pyFBUOY/j5+47Pix
NKDWi3Pku4CjGRrd/x/MIYVE51nDEto4GTwHflo4U6cGM7Yes7e2+vRbkox6Xxx8cSsiaOwHNv/d
oSYIf8jyVHOERKApEyxcxm8K6hPDevB6FVBLLro2b9oS7/vS/euvX5Do2SzT3hDoKuGbY7Gfz1pY
weOTaECiHeQqJ34B+K/J/aEMcXUKVlzIut/MlPPuflVgQdlwVoJ5WHX2xv0TEI7O+Gzd9XH/jLzH
iadabhy832rijZ2ypujLM0dHNsKpdV2xaA/VckwYy+ACJIM6wZTwd1vq2RErDGPShGInQzOFcRve
1SEFAlON9K5YbmOqngObKnyW+JjfX7xjXbjAsmUQonJLXOIYNjbg9fE1EaZ94ANmmf5LR7pPuY4R
oMomJ//3rkISfpgE7xz5m02tjgojUXdbP++JEgazMF9xXwL3ooYBrmWy3DS51sqPqZproBnbx+xR
2/Pm4Bar/9aWiID2DOl2dqNcyg0NQTAFZE11RpxU4E+YBwEyyWiiiEilIcxc/9c4MmStIK9qxjG0
ps5ajG/A+nOQpOA4K2b0oVNsoj7O50cPzaS0Jc6ndVjWQvSABmKkFLK4fhwGhFrLakHAJC2LZL+F
xoGzT+EXM6vmo5Xk9uMXtG6djjcdr/RIvbqym2Uh6bzxH5CketmnkEYE7bHF+gw/SMZos0AIpufU
p1Fg8a8gs0VO5qYOU7TcQeHdUSMzLG6fPpK5LxH+6MFpwdpty4jcelJPCHXUbnRVx1qehUXS/mtW
Kj/2N4pGlHri7vJUkOfN7EXK3cceSQub7NsaLq+lpemVVJ715bibnHbdbULOaTaGml1tnUPamUDk
MsUh4rWRKAG2mxGb8iAtrhTCrbAc50bk3YL8Ui0Zsj6kK5KC1PCPSPm6xocGM4w/+v+3UuNpWxbJ
Jj04LfzBcyxiRQZezszBCPkV6RYC73sg41wlYDEJOpPi0xEhnSSnbr1a7rBz8MbXu+M/DhK86jQT
uCYa24BPnIbAYYoyY/SbqeHORlgPl1TsU573YrDm2eVwihnRQ89cART3d5ptFy+Cszwdee3oo8by
J0v47dWP1mgyoX+LzbUzdNbY2EbEkQXgibcDA3ruY803aszF2MdlYBIXVBE4oyAYhtrjf6VfCF2o
5BZstUHgkVt3+KD6SSKWRaf9YNaZQKfUcLTn27irHnUl7lbladDH2UBJng2jJREvSHl1QpAA1mg0
CwFoRj5ZImf9/urPNvQoCi4LbtC7yUKDxTpIWSpdtNjksMh5m82VWVnN4xC5vY2ktckKQQDRlkbw
lPUVgZHQBgeHfieVLdN9za29+E/0wqHTTU8UDbM3jvYvpNZ7+Ca/E9d2WuNFdZpf+cWaIOB17d+K
NmFX1qDxclgjst7OynK/Qgwfk+5FlnjOjVmPqT4Ny/mnGHsyDcTRSwHkyfCrKltvdnBvzzw17t50
Fj0j4+R9CM8J/YaQT109SoMPcgGjQzoOmleT4PXCnpQt8kiwact0xNfCgaM4l/hkvH471fVuxYbh
Fw9zhOz/RJ0ySz3xhPVZuizoovAFg8NUV4Zz7s59AMHGt7dafn90SQ+t35YkFkdDxRJpAoC6hv6U
EqQvI2HocH2s/goXP6QAzxPm5Ubh19CHSu3w+vqgGOHn67kv+zlEl9MkKocR5pUkxicbgoWhSxQM
JiAlK5PAgAO0271Qe6EkMp7tyUS5ekhuT2O5JYhqUz9/dyvVi+mBywz+FmVR/iq7Hr82/xkGPpUT
ekMkaPZyfDBC/faMGXF0dvL5uMN8BdKibX4w/6ciigVwqpQZGWstWTt90w2XYY4XXC/lgbAOWgTn
edU+ebMnbTxkRyyxrxsKXKYH/Zcd2VhUP8wFi8sDc1CD7eS1HNDocAlCwe1dIPPZMvtsHFltLuLy
+DVKLF+3ZkeDswggKgHKrJAuDSI6sQ13iiFHiu3RaGiE93OM151Mi0xRe0xHJhRZtxV3TyYy5dYe
VAyjVoUI+jBglDHqvnYJGl2k31HHHXVRARTXc/kYls6eE1My/s67kiYBYvde7Z08UcN9whMA6Smw
5t5UjlwTGJx4t4Zg/kPLzhXUDFmFvSI+rDEXA/MozjMdy8yQQkTc/5GgdHJNZMQi5P7+cCzGFtaI
WgVMd6JzKhX79IzUo9vM4Fw6ELyC4Z2O3jF/km5RHvZXnIhw+LGEqfPFTWLuEKJeeyU0/hRY0gJ8
5L/e8WKtODJJoJU+q4P/WTbFvrzVEzRx78lQ2SyN5bQZ2UtrHSjW5REn4GPFM0iNxy5kYyp3Fe7L
nl+l/esKPrw3pMEgeDmU3Ag0c0etK4arCrZUEkpRq0KxwZiFvesKQdCS0Xur2ZpYoOO0tQsKY5Jg
dD+spog34dcds8jpYEFbIrN+WnZ8PRd9Sn7Inn9aKtIKgHOErH2+ArMzzfpXQxA6jeQYWC2ButKB
RGEzcpG984O/snI9Y3p4WL8FzEYn8IaEU+pafvkSVFFfieYcS5PW9wgS1mqMT4yDttm6ChwU9wlV
oNXCRWaenUKegPEx4QhszJC41CcCGbuuVFnSgUnpdE04fhJuzuztmCAsujc6MkbVNMIdSroqBVYC
mgNf6NtYSZjwShxDjfnuUtCUc7nXENSlvmCkxMVMGJyVIMuKBgwUc0g4WKAmMbPOd0zTuGm56yLI
tbX+9DnqfIyfJQZtTPsoX+w/X9ZWlblfQ/guxd7/U5H5FQ1u86Hq/D4PLBxJ8RR2i1LWgFryKqfY
SqnYGIMc/4nV1iSB1uqJUXVbdf/OPw60I6jlm97PGGYXdH2fLOUpiOaV11Ibndh8/nXGQpqxHFTq
qsZaqwHSfHfKplUxtXZcegqmbpvLatSxUwmPff+GKS9xaZyKeqAPiPrcBVT4ieSu9UYfv1Rl+9Tm
ZvHO7y2JIqBYzg4WbJ3vg7FEJyzju9Q+AsYBVN6hfIiG5qLCTh1tBbVB2WC/U/wU1ibIWuV4RjuM
Uf9NWUx3GdqYjDNeyxVYqPAicCHgX45VENJah1/N8UUmNTXO7PxRDwxoRtezuSweGBqyWeEo7b0K
gZL2RmVPnx/wg20yD5AWE7U5hpB8L7jQwDQKJnMRuEs1Kx0mnQ+shE8qPVU0LWJM6yZy9AY9f9m0
UoIZsZmRSvCN6vFQWMb1URD8fKYet1vYTe2OD0DjRLtxzjZgf5bdd+UvK5R1cOb+/PxLlDsmTjK1
ct0nQ0lRvpWFoNX6QN84HW2mNZVHedXUnsvgRA92DERk5gQWbjKSs7CZJLFN+K4IxOVeJDDx+O4d
lbbxTI7pYKwGnN0GB/bVP/Aw2L8IAWM3vGY83tKOw61lIt6G5VHpA4zM1vsKHkPyeNO1IpCWKP2Z
RliEsdm0pbnv9nLeIMNiEauT7K7I6VGhDSMPMqmE9ctuMEYcU3n+E3zmWl27E48axVzEo6UwAiZu
X67ku783NrilBOw+Yt4sefNkSJRbh2vxRMrbBj3qq415IikyYYkpgUbjD3SnEBDb0dTZ0/q8a3Ro
eapQ4pcVUByCOQjN6s7JNwno6OYiI6HzrHjNfQ6OQ9BKdtSxamn3kve0/meESqUsVoIlA/gelyrD
ZZj8dUtrzdkBVx46ZwNudIBNlSBRr9C3YwivKysr/foPeSeFp4eWSBtJwaYlYbxxxz59Ax5bWRKh
07YptielFs89c0xxEvZgTK7Apg0OsmXGvdw2SbcomlBiC8aCvBWj/OO4lQGvovSgRzqdg+CMek9U
DHjgvfh90SeQyDUjHb61/yUfMyH/9duCAnQqfa/9JU0EENdP/+PZRuN2uGjOJ39RzRTXXIg/r3bR
U9qePK+n9lH3dqNP0UAG0mdeanMdGybpeSj/WWEx9F67WVWUnuYl7qpWuKN17YQ5tDHlX7QhW5Km
Rk/mBG4RcrxypbrfR6/brSs5M6Wa+V7n7HkzTsQsh9btKtvU/9MeAMR7lTYPxT7UyCjAZ5ZQWgE9
i9KtUdyQO17vzbU3ClfRdO2FiQ5HOQeWuQ2KpZQG7ytDdBXJzToplvK4ZgFrG+jmWihWIcwZgcNY
zJCYNBIdu9CFNc6jdQkiLk3PVt0mYdA8MpxBaeuCkhmHp0wKjLwWTZ0zFacTlb7+O2aFWt32KEPX
NGnEi2h/TxDa+leg+G/8Fy6zhv8ZXa9KHVCtP+/QwB+lGzMVi3C1ywjDqA3Av1j9++QcOomGRMqi
qvK+271j5qawL9KypuNbxGYozX9kZOKR4a/ychRalzJZyMaG6tBxRB3i/icHBfGEKrRzIsYcw2da
YTOr9fQWsD3ou8pvaPmvuPlPBDSas0TVQpmLfijdrNb5sjB777Tb5I6c2HJ8xEEacRswuvK1xjkq
ps0juVnFzkTHkgkahWI9jXjsNkjnS9z9tuhxT+LYI348yeOdg5pj4laOOnrlsvbbseO0oeOklm5g
aD/nsX8z8F5TyrqdSsEFGBOWn5vVNcuIaeh0nE1QcpMJ4SDtBHZplwOLbR3Cz8v2ocYnU/OcF38I
pvBDoRnX9KAZuzIQMIxvovxDpuh245pcZyKm+PujCl/CPKHGNce+saUDsMntxrRIQ28Gq5wCUdbN
qdXm9+3IzVaXDkf91SVgIDyBOhDZ4Li3WtUZD1NdJljeXt9RTXBFjP2lWaB0pMlxFOcC4+qbFqTU
bzs5RBBHjp6iqf09DiNOIisygTM34DSO+sDxWBNVSn1toiQhGK9T4nmpgYmPIWqn2gAIqKR03say
DpRuUy/zqyWtt0xF7mbHk54SzRD7bBQXq/u7h1RGWJkVC8EUdemNTH5wiCm+DctihMnZXXD5Bdsv
sJCOb6+XeBU2d3dh5xKdCFn6lNu17M8zkq0OMyZR+pbMwHnhMG/qpxuKVfuf4M2WEsldGd8ksF74
dljJXNmWK6AhjcOPJRE8wOTrby1I5w8f10bKP1uc+FVHrsL5Y4WFeQW0z0DzHADN53FaNHZ+O24m
CYajxSy3r6v8G5bDrQvHfAdfaRAD2Xm+84K+vFGceP4BcHjZ3HWPXT/ek2yyYT08xRpkRu+mhpgJ
l5T5fhXp5s2ie/k5enXEQeDIvej2SRgF0I2L/o7xOqEzoMK0bMXd0k8CXQObtyd0Ab3pKSBpLJjD
/MUEKDQ0zszYX527ZpLdXvJWlWPuPex8tZmEHLigjiI3Iavs8eOZAuvJB8OR/ZaWLhsObzkfcDfc
NmsSIBmjgBV9Lpf1R0rGLyhu0+wuKnTyIfGaNaxprzrvzqK49iSAUg859QAlIxHbWdvCDj9MK4mf
n7ZNf/byr9OF6HVDYDbQ7HpMOxiVc71rRAUVdIrHfUixcPPjm/IpPncqNo7geqpOfVX8hHgenNP/
0COsa/9oMyq4jX1+BE6ItCTzQ2zwnSGKUIsAdeaTLTzc6g5pAqMzTNguotLX1VVRallYxeiUo+yj
ZI3lzOe4N5YWyzErzShwNsQJ6S1z8/A/2iLkAXBmV/7niorMyjiy9+RKuzjuuSnDs3ZSLohzJ0AG
d7+hwIzOjQM6nY/xgWGeYPF2ynCx7H/e1kIR5CF9ig3CmCaGFUTDETa2Le5rcOWwelZgzOT33rtn
lHk6ndRde4EDgQD3g4X42DnjVseJBBofuqQODLo9RjleMpFjPtepXSd964BRA09WPuEXIpeomGCL
AvOQAIwyYaPBqkvnqg3EYnlsMT/wfiTfl8gD2RJmSSnZ9FhMBr0qupxBSsSeC+Wn7rEkGj/V9OuF
OojTY4u2Hz8+bFxxAAksDNOGyuCyMXzdQrIHXBQHIn6nMQUKd8HxiKLuW/w5utpDeqybcl+Q+fp9
Af+NqcKg8hyY9uvWntKL+M+tYzsp4U96vbVgW5G6WEAr6J6d7pdcAfTvdvE/VPuwRqOWrVWp0Z97
v1aDFFOvGX5UfrjE2W5xauBTNb571rpi3BRhhwXG8SeoIMgiyZ/IkM86rFgkJaqmlUWkVo/RKZ0l
HVQkRScObdNnYtLRMHX0wJGQXruYg1Ieygw8L/M4uoRUJ4OTlyzlquiUKJ+Vz1jlOFfdzvFpsgm+
9IaZSU26+pqXIZeovaJh2X3C9DW8czpQBiTVUfVSHUeAP1Ebem7+1PufjJTdOH/dJAcw62bzk4Sd
iN3aDdtJoymzBDNRX3DKspGw/E3Y5n6D/kqj5/PydUvrXcUK+9RsZg6gPkbQh+i8jxSFJYSf9svS
1df8YbnXDfaRsMWgsFsugPi20PuOfOF3eF4Q/O+EdbyQx6jU9yWvYA2juWvjNXEgsFCdjHay/mre
WcVNM+6hF8HKSFJQX7tBwd6vlqNPtije3sG1iYpbGjyw1ravXQ2bzQPdVuJI+BZLFtGoGUBAUMS1
8KxHylLiNnwDB5awINFJ6/LfplMQZEcriJeyzded9yDT+RkSDOeJezeeo3Vqr1d2ch1RNU31cg2q
GuUN+/x6pZ/FMtbXbxeIxifq10DNyS9ZUOXPlPw38U9do7wHOuzhryi9TZWqXGK+IYOVnS+jjjdO
L7EoOZONhUf10jv/hl9wCygvOQDWd1Fz+bX6T1MO8fSTrC/fuuO3tQVrvFdetAalOT7dhSZSQGmw
PxjM+mDLJDOvQ69MufXmzegnVRIyGdm77b6qSCtQWajpgn9Y8OFzX08zZrRUcY+lQNwkIuesKoWC
R8lS0PaeL4DhDtz/LrgZOYzgj+I/Nku1zY7aX1wq5jMUGB/TF84cvYCMy51qF59Y2qk5snKM2l5L
yqndYXLXdF0v3gTNuM3DzCTKfImJQ8g2QhakwTxxxjWXWfTcg905fpH+KWkYFRNW+8Ak6Rk5CGQb
GXAEiVaOPO88E6Etrd2TvqDA/7rt0x+hVTrXxJkFZYf/A1ez5s+Xq6jhEbcIPxHcoEh1qU9m/WTo
vVsQ+KQ4a7Q5IWmsx9fAWh5hpCOjWhXWyDBTx0kLYepkMMr6pNuWz41EoOd2rt7be5yeNCwvhpxF
UXvloLtxQHDOZTLcicdtIC9d7CIxM1c9hOgNkFTYDLjpUqtp+BGJ45w7jwecN1MpdFWuNM5yyPDM
M61ss55aTeipzwncdjpc/rcuJ21VeeEHjwVvOaIS82/iXYpLt1Qf0wRorLoSRo5Fht3iUZoTatkT
UKIIKRRP2WCEQPiyurwcgLV9s3SIgl9dqjxd/ZnCS2crI5iN9j9bUHjm2hLEj08q8m5LFcbuqTCd
PmKsODlLg7TIORgEMwjJTT/PFbejzFDrI52uoCLc/RCa0QRUynuKckmK66KqVBbE850OfZ8MB9HD
GSujznU426OwUvL+kvuHV7IH/Kx7mC9ttRRashJ/9jNbqhstQygXAW2rBlBPt2InTYlZRVVIB6/r
i+CC39M4gNRkFMb171hzUCmEjQUOeVkjWe8yi76WVfw/UFr6ufCHCxpY6zJFiTjKZZ0D8aLZH87Z
4C06383FWQ4ml8d5Km1hVmrtU5i3yDO2y5b2/aux2U8Ebnylg90afbU2Mm22mnJleje92jDKidRo
AqUY/phDwU7QvQOCQb1sx1uXbB/KhqsgqJEB2tykQUJnOOX0m70C2jQQbp5CFYIX72iREEGSSNhY
u2lGK7hg4I9QMT8k9ADFCZpaWGsn1m24P+qTFnWp3E2xYWyZEaG3WegK2kAb5qgl7UK2Cp0ntHXv
BcPSwhWB0LpJqhgIVOQX94+gqbO84R6NPUCUktWN/xZOs/ULc4j7NcuGS/vz6he/pi76mPikP2Uh
dMt45SxuhxeD9S+5yTiQdu5ZAuY6TEKn5gryL3GWI8q73+8PeVbHp2/5I9rXlCSYqZp5im6tP5kI
YigiTjOt6ZNH/8L0QG+ta3Nc5Rl7sPsyyS/HOWjrcalCk1BCLY5IGHzd6uZ16YG5LCeL2onU+Ay0
GryA0t0V3uUkEMfNXMhqrK5X7/giZQH48xXAL5b3FzT1f8oGjqAazVoqJv7cueQu7KrICjSm9cWp
Yya+meKs7Gkjsr9i08AiUx6N6CtR9Xb37aUGUCk9IO/PXGIswxZeoE/gNYIPNQdUt6gLzsW8lvmZ
LaSHcP8HiH1SgNamC36IWSxn/nBBLkkBR6UlZ2KJUUSDRtEwE7JQQbtn7JEkyLAVQAdLLeEug+5R
deIgVO+uEYFmf2IDrzg2FUEyomXLLPJnlvjHmB1TlrzCckZ5/vmPVKL4Qsgrl2Aw+VVNPdh3oBHj
zFilzOakLTloE58ruBXLLmYIop/Oq6FnKuMSHHdYQR4dphiFIocupEisxrnvwNdTwQhOpLB8uXq5
NUCqoZYzbHYjG1rT+kOvAAAlrD25INFUL6yC+BbSoVxhakOd5b6Zf3kamp38WVwoqNT9yqUamFZ+
2cbikcbbVrc9wjPqg1Zs2mJezi4kbTfVEt+BfCvOhBfvKbLR+xDSvVewLD6KBYW1K4g3LxFGyOTz
Dhv24hA4hPafRpd4ZU0Jj2WbqL/OgR7RCx5xZF7Nz+dt87fqWKwzWQp6XTiXJmALSy1GsDRr8kT6
FQxN2QuCcL4G/sJIsKUYeX4ocEzvPcRiTOU3UImrdHuuhhZ5D1nJZIM/JYQe5EYMS/mPBg8MiCbz
3zCQlmSTwO4yW8XcyNrRjLi8oEiUaWKnG5ALKnBNypJxj0Szwkb+GX+mqSUx0gBQeiWP8L1Hkyz5
M79xtrncewdZRYtsvWgv5PWt6t3C6jrdq8XmuxVtJZir2UZnik9PqURe+V4x5TAESL2DtVgaH0hQ
7B/7KngH4Xjm8TfR0Bund9176nxkveNHNEAEUi3rXlPVd76yszCHabclFGpUtPaBkpUJeg6oKtJ9
odTr+zsPUHqlHbCaQdop7GC8D3w9AdE/qkS6t8m4NoT3QAhHwPOxZ1d+/57KFtD0cbT0aWclyTyE
bPa+6ctFYloUMNdl/FmNMikxW6G5uqIWLzDQ4uTQyP5n0lRmoIwiheJ9RjCUNnFQXPOyC6DN9EKe
gsMh6ZKiavwCp+HcY+GaiOyYxQcMok4mNDR1Lz+6XtUXbAxmYDU94mw9tIT9yqdnt1PIIJLGORrb
OWNLzyg61M2AnizSQRID4aaD8opBYxBL3XCPRmuARMvkmvgwu+0xZp0vkALzhPbA53wPlE5TIDSy
edvN0c90Po3zDYPBNsLwZSqvPUvzoqxjGo8EEMxWpXF+wQbFppQEUtRJGvDYUxA11Z1/v5R/+w3D
ubG10jPdva2wB0rnU1UM4rDTWLwjzVoqumgSQIetO4TPP6x6kfkDaGZgWTkpm5xEUYSodN9/JVqp
LMz4XPhrA/RTUaOcQBq0wnZGX5qGJjwevnoucCtx5tfVmCKriaiDsQDF46jKhDOtMXanlyizUfmy
8sKDhjizVlQ4IztSha+Je2x56ounrwHWHXtGfJMx7hxGK04K2DtJKMe3+CcMTHZg49UEbNFbJ6V7
AxV2g1W5NVuo7Kbtv3Brw9TQ8TotGLhsaxO2ovNGBfpsO7OvzB/ZawyuuQokhz+waB9WP8iFSEK9
w5NGkDrvnUvgxc5a+T6Gxopk8hZ5m6LcwF2EqOnDnzuXSSmExqHakmQjDJYwHGgrd9vpih/YwJD1
cSosaDU4zPvv7ofCK9zSTgDA1pcDMw+rVCC9slYJ6Mt5XOkCVP9TgtWVUhg/iSa/5KvB/5Mk9c+q
ueMMizwwM+cE7lRRbGkJj1mGOjNFLWgryMVjkUny81ush6mD0Eu4v8bz2gm15o/Tz5ZFT2DPe3m4
nv7YuHdq55283AOkmNjX740JpnHIffoJ5UPSHY5JLWv/veD+3QlPhpnxLxGioS9bNr6AjUfunRls
/IbjVRIvA8TFkB1oltH8oTOaGy49Ch85woqlFJ3qSYkJEOyW4dv+txNKMAs1Kl5VaU0jPNR+qK6y
uI3BOnu3rgqYiLj4VWKxCRelBfkxBk9hk34cwcp19nmKlRu81lnOrcQ7R6c7s1z53Hy2g1xqgz1f
5FQI4/gF3l/exqx/HEyhya6W73zp6DDfdwgyTISEFYk7OCvlsVf5dHNxAGjIeikMLb9Cgs+r4Che
HqBd8KOWoKijfzNFP9pZqTI0BmQ2XuX4wZWGFR3RmyTxQTe6Jo2GAb/+mSwuvscFKfgsPuZnW/aC
/6uN/+dRU6Zs1YMgC6wrSXDeOA5jVBAq2nbqnlPd/PlZj0fME+RET++RenCTrEZobhfMYh8CI8XJ
ljsJkW2zcfzjKvoVDKJm5a/79+G9rxorruz5OsQTnsLjmTAFOQ+1fUm7E333Kz5oSs8FNQVy2mZj
d3ogC9c616DYLIvn1PsDXEyJMSpkUY1JQI3MQCV/054ipgqMIOPP+4FkFaQc6N1UvxH5CnynIPMJ
P6MAxKvlx24pDZqB0/YTsaN3vsvwXUxFwOwLNsKw43bk2sDmwBH1hVn4cX9LCT7N//k6PWNXEra3
IsZFT98abw9G3UlPhP7ax+0m/ayuAWwAAO/CNazivuiGwdbjdNCISPl0zPH8N/abQqSMD7wWDL+e
pnKT2LyNNQphSA6PargEyWIqzA/SkF8Luzl0AflZvyPbGvJNwCeyHXm3inggY0i6ls3g6j9Yy4I4
H87lJ8MZIyWdHD+yavH2SfEXPeXPE4pVWMgEvcWBNzF4vERHpbBCL72BtFw9BaPTpjA9Tg6fa4jz
fRFsBov+wlWyxitEQT8XuuEzROlUQi3wTgLlUtWcHW/SkVVbIH08/jHAQXu0dk8Z1PwMDWQc9KRO
9XoJJghuQSWKodBJgBwQFo485pJQG9k5nZFhGs4vt8pUNyUEn7yumAhbaB0k2KgEkqFeHCr2elRw
UD3/7tkYhmRJUoLS33a3mDBRevtb7p339lroChX16YKo8fChRmy6eOAf1cl70zEahjozcffyxUca
X3tomtxVc759kZEjEIJXTGYf3dbL4CNFOVIqYDbzJV0Y++ftiyynomR9u0wse6PDXOstEmYcHe31
B1mHGfsQdcD+HFohPTac8mYVNf3jvgdNsZsqaW9JRl3wgGWQakR8D+t0MPq44uuQU5Wz7Usi6brq
owpHMpnEfmzLDuO6GGtaBTS2+vxXRDgCsAP5H/S0Xp1R/itBq5SfjiGm0EwglrPrt+/Am43F5eXu
KvbPWxEDKgWdeoOsqDrTp+IaU2ymmEWRo7O9JTx0rvZxmU7I4S2TnoQGH+0w/yMCN5r8dewh2cEI
LhPYCxw3g9cwFLEmUuZi5fqERXnbBLz8nXRVVB/1A31vSDo37evtAic4EIlZCiMEfXk8tFprGRb0
R+tBCEvNB9VWNak5gaykvusZ2IqoPxMUMMelzzOw0FkYqrTDPOFeCXY6CtOYX2gLdBpo7ooUHJnU
hNxeICfuK9QpLsAaoc+SzS0a/MmPutoXL1Pj+XuGo7DoCztgpnqalyuiyWBdTbC2t9tTJLjdLqz0
ipTpamQ3xvRlTbRkInG1sWVVyt+TzpJau2nuoI90OXAzVjMUxk60zmRVxybLsesAuoGzfkDobwQt
KlQmxnOLkkAKLFV96nIQXCNX0S+W84cM/iFlNFALiTe2LXdrJ2PoF1eiyTbLNbCcpWGvInjqgh2y
BrN14iy8yBhYewkg8KiMtvo8IKCGWuxAAcs+V6CdZXuFVbDwjoIKaIM5Fk9k5G4KY5s0j8r4QPGq
ViBpZ+27Cn8aOmi29KpbdgJIo0gNvcEwoeTgtn3SDq00upif7390GTOW2b1F3ii4Gdg45Avp7XxP
0TVCNDOWvlcPpqQiNFYKT1D9q6WmtHbzH85uSehTOthAG8riIztAYQG/YB6sZ6oIGtQxv2vtxQuO
sre5pjubHnqAm42Pgag2LGMnvfmBgzbKEAQV75wM+PCiacrvMrK6AnmgST0O7l6XqOe+bRnhQ7rI
P3BZr2AwCN6mIBjE906NN75k054B4IReCumFQgTl6bhAgtvdCRcMsbrn6FTKerHJxZ9SZZJO/cDE
gwVTcpvHEXGR8XaqhjbQQi9M0HN4F9LJl8qsgdZavyzdquLIPaEg/0glYQTb612i1zAZTnneTC6f
ZhsSvx4c4ZVWXwh8Yp0N+9CxzQJrdwWeidtToIwYqbRPOOC/rFkEMMDUaJ6FVPAMld3xb+WzDpxV
o+k7V5EQqRc42w9r6T9OOlKNCc/zBMjx5Sy+tR5Rbjq/oL9Q5M41ankSgYu23wEZQ7X/HM1kKfzc
o9nTcDEiI/Wkv0LDGkAdQHXIK3WCMZMDdX81/UoNBp/8Z0fR7jmlsvv3+L0mla04kKYKFGSwob2G
bTcatsRBS4BWZrcHvJb+pr9nLqJ7kqVRsUVrw3Eq30MnYyLxS4u+6Y4/5Ci9zjdJo5cejLRykwaH
NpxSy9IDGcN3q0RBQc4EE7qecmE2tunTsmA7RCs10dWbK2k2nFZd8Lk2r5Msj5WZ6W99aDO+1BwO
WmwFDbVDujm3EencM0TMu8CXdJIQoIx/wrG/2wnXfm5u7+in4TUEy4qiL/QRnHULLi+AHZ6uWVcb
p1aozXcsd0RrOaJ6V2GGnPSPxq13klH8AHNz69TVODzrlsu6dsQQL51WxL3fljT3WXrEOdJpfzee
9dSbyg1ulOwiKoTSsDBol7dkZZHSopDxzeE86/+s+KzAw3iAn34dUV/p9s+z1EW/HrhBhYNDSd5L
fkMO34eWEIKwHNo4ILd59IheQYLwTyq4+aWQRkfCHmbgNUzzazX4OZMDB6eQJLytsJd7meLqES4c
C1pmuRc792PngCucsD4DkRv63p2S0G8u9EH3nEqRTJvLPjYw8O3vTT52mDfhkYhMt7D1fwIHD7ww
BoRKyl3EaEVt+UWh+Dhgbx9L99aodEOWPgFuB66N/aSnkOsxqW/kRO+CTLPmTxuJM0X74JH/IoNR
edMAAupCu/dq9CJ8HRc+rGSpIvv6tjoXgL9wVoD4udlQ6mVcdNievH+GL+wmNxdmgSFpLbUH1Y6R
6YYMIFRFLr8LvwxBsTHF397V3sv0zHieTKpGv9wftO9cpAdsezIOBC/3fU/x/dEPFmRA7Qt72a8I
y0fmnxNg2sLUTsroVyiLsuGylHE07S0ZsKY6vPPeFIrFedxX4S3YHB7PSJXzVzXyeQYGcgRLAVSJ
vYrhes3SL50TevYxpKgD+5AdIwcfNy4hbV+T230bpIn6wULXH8YkyTatDMM1Ia5IT7hYTQTDBq7U
s7zkGnzzVc82T9NXbRAVPa1Z9t8yj5E4es0By69chNLkOvztVJk81/zh+DNEZMWk39jXIRPDHlcP
8rxXfSg4629JEt2l/TxyM0E3bI2n2gElc3Sj59NyjZQk4pXkXWICBRq9/BU9Ebvbbr2QePJXZVjM
vAGAIWCglWco89r6AbvjgI+u/bndd5uww/mNgNnEPdrwe2M7GziNJE8OR++vqKOcFVSnoKcc9dX/
sLjD8DTz5OIwO69REgX55iGpZkyMvFN9A7rhdQaE7ub3DkANvkBaeMPceBLgtOcIBi+x+veMCAGj
1xbq6N7jNUPs47fkP/kXuXzS30c5fzXVCXImcFQlCIDQUkxHh+UV7m5oA55PKKRtufUA8HXxtQNw
2U8FwUOR31r/yGbRN75wVeeD3j32now2ziE+VT3Q1YuR9Da5CPrshtoqi94dcyZtYIIouKRcwBrN
lZQjGxqIYugLW+fWN4AVQYqeePQ0rYTXke+s15LrVFsOurSciXzIvPhM0cGoHQM1r3N7aiyK1xTh
M9CrQwMfg3/S6Qzq3KgUSEXbFFoIpwcLnEGRE58JLk7QUEVEjPEuTPS8lJI5uXi/LB8YXNpbgFzn
vJfbNmDuScMb20SyzVLCH9FUb6RkuHUotIctgoIdq7FtkqVQaZtitnCpjcAcmfWwKPdiaVfs4xcM
XckoDhab2UZ+1pc/PEo5FBZLhSgvp0D/YwSFrK9qyAyz/upZ+OK/H8NqFKgOkmUWFxWt55D06IcM
iUZH6uibqd963I1+ZxX+t7s8dwshTVB9J/9qTc4fAB1uhkQluJiFkoyVCKZiy/eJrmZJIOSBqAPf
H2EHrCpOP1nx2CTdHQtf0LXcIkJaqzlBmWoTEwwQIf+8aNyUI72uh9OX/cf3x6305oafnLLnC3iQ
6vaHsBWX3wKoyM6rP91sl4Dsi5Tsiy62xKWhyRdrkxnVMkk28OxbXpjdp0/OIt+skFJw+dsoM81p
ZxgCr31HsMi3YfcqKy5xl14J386Nk4NPF6DZh2/Hv4o6FNA9yndo4TsuylVlIUcQWgWg9G7pij6q
5tcwEsrXsLs5BmJmOsj1LJPsdlMIatQo9+6rBwvs0TdXYhk1qf65mYa6DN/j2B6uYqerDefyTsrF
Zx32jrWG7itUPKCDgpnXvPKaUTiiSDVAO1NRh1si9lYJrijVUNdho0AgmLUTWrIALtbqMDM/xQWy
a4HSMt4kZAYAuiCmiLkkjGO0dvaE0nG9lmIjWoZC4dUX8iUpByUlmjd9fb7EKsgYIf0IXsiPEaCl
c0GRePQohVeaXbxfZ7CFsj8sW6Vqzt0hLrKQCgp2kEl8NQc7KZGUvHj2s6/rz/Pov++N3ttm2xUt
XSRH91un1EbO5sGHYNEbHdyd9vURNy//3WgmPy+py3xmWhgh/VO/3sC0mklgcs1U/1fPpdV08/QD
QXmfNJcAjJgLABLtKtRJ98hWPTgOSUtoDebb8oqmPvLQaVg1IWY5X6fS4t34AGEYjfhxuuMcRyd7
X6j5SYpUOjPjqByz3W5Aah2U6g3VpCGtv11mawK8b/M365cGrly1pkx5gfgDvSIp+oNcQEvS0j9Z
qgECXKhcSr6vFaCHMweSriUboBpkbAwuXtkozWETq551xCVA0PbauyM7k1nZ4PWYToyDdBStgufB
gzT+w+7PHKTpEYBqHtyp+qbRLrOVIEZsuyGbO5p2BrEJPOsHfhd4bHqCvAcKZ7OD49GX0HDRwx7d
vdbX0FowtoFzt0yguB+poDTxipIDxUVAtENiUCbcWxiPa6HtyZ4YHDk6hR4A0tTV/IqrlZXQY6e0
qpcnluuzooxuZveXAPuS2Fn5+PdbDWiMgUoZew3YaSE5fj4RiBeAePn/mlHnDIiL+SZbbV5cKjBR
B3ezmg6p+QkZluW2QNFA2THTfEHRLxja8pNUHN8ULLWpKEI8mB2CZgq5Q9uWckxuyagv4u0VXHzI
KAf7uQLanBmvi9DkDFXCYNREvCUR9+TtxJDK4BFCtQ12cZc+/iqrkGH5YQ1UtSZ+AFsAR0MztMns
F8hHhUZyBS97M1eGgd9o3u60xh76qjXRjGUnmYD/L6vKQSZ1bFUsdnzZPmXld9AU7pPnj0mSW63T
uohIQlNRbkvOtHMOTVc/JpVpiAIQuCVk7lRlvB1GXGi5ti0hZuGBzyu5OZ5JuCLvbD355ZobCcD3
AcZO5LMS+BPHs50wqCkQXpi3+zNoTBRzr/PhOUqkOXpyi48T8B7AUHeNd+/KHSsz7Xs4PTrJD/lw
2pCgAn124F+QqSB4HFV97SkWDD/WVs2wdM9I8TsglDP/wmwbOgBBpBCH47lqB8TH+pUCjHEGeO0Z
VscUSdsfwm/zedjZCW4zkmEbis7X7KgrBY3MNPFgeCaNX+PAa1cYmmEYLncgrWJBned+fUp5Y2AJ
gF4L/ER9TBi3H98WZU8cQBU9m5peg8S31eu/gAKvabSwCvltjVgeJO7mTl8SNWcZQwwGeC4Jc9uU
HRpEZvMvD1+pNXOGr/DTGTQIA7NHVyKkbcItZni84maADynKznUlBO4dkpheoOcjI/q9COzujBE7
i5Nn2DoZzKRBrO7GNY+WMAWBWu5htR3vjOYkfrQPm8FSyclK9cLxWMs+H7sHKIycLZbOl+Yl5CYW
I2lG57+BVs02PSoYSNZy8Yn5msejHeB7w/PHnWTUt0v80xZXLsXiUq9wzGqMWzuZg3H95Ju2RCv9
AyXwc5+KpWivxKkMBVCuE3K9X6adkVWcMDGpIS1UgEXE2BC+TFBJsmKuYPJyCOXhKKjS363+KEhI
Y5qP8TaTxMHYe3pbw1OgDkaiavuuqY+uLbMlW8BGmQ7CXS2YKmK+5VomZ+SVZT7h9IcrxILyKkeK
lPyN2Gp01+qW99lhdwtOjsGCBPYG7J+HtNFsWvK+sivjzLO5XG5a5FfTXJD9YTN2TwO0LCevKXm2
I2Ws0RKRk10UvbkNESAqTdOCckDN7V+z2aHEyczMm4RDU6AxdKoo6hCGC4zVIKXFTQ1jDhzMWj2z
o27WY7KtcJ2t/OxRZIZDq83v/GuPao8y9GNMgRp9nPCmEOWWd31QaDgDsX20S51oJOg3h3mIwO0n
qo3P9skfXMmBdqIVuzFbYEiVqOFmGDnRppxRykpW6sWC0Fmv6WZtSeqBPtJJmEW8pdGtBGA+SLVb
irB35Mf65IWLhGDFm3rutTamv4qeWBs78m7V5AemcOgM+fvs8uSLYXg0E5RzDCFHmjTucj7xmMHU
0szFAWrgwX68K4uCMDrMAF/Ifd4K7lP0J/9eJA0gg//sN6sUMcu+VtRdPiBlgQ7JKlusjwkpwG4Q
tifoGRuKUb9Kt7F85fkfc5OR45FQk755VHP0idPtpcqkYSpQ0FBCWSxnw0WGA3WVAlDkPKbChnv+
ouC30xWV16zNvJ3B9CW8YQhwrXzsnhboUoaVu/xlvxIfk0AuaEik+P660JqM1+1CPPbHYe5lqsVK
FABK1UWHPhhGYv+FRG0XzYG98Rn/i/Fw70K8bUBtwPqrqotCTmQ8z6wSJsZZJbD6SVzmAz5DJzmA
zwvwR7hYXJ8R9bJzudYPcNJuPKgwqLqofNfr78+vSQQIzKywbmuNTNhXDRN930znq/n673CMZzc3
lzdt37rVWUMUF8JykTQ1dAuErdQpjp2uWOs3UOhx6uEq4yG/9kJY/U9spAz6rcuGvSE4wESIxT0N
dZUAkCqwGnxbt3Ch0O8EnFN9UvOHBI7khEISX3gEKr1xDdc4AxD71jA1GpDsNmZXPlx0WLd7Bdvj
30tqQcicD4EvwpetKAxV530mozUPjEYMg5cU2XV4TCyY6O7b74FdLhxWF+EHGbGeLjXN3VINp6jf
wy8+iN8YxKonk7DB+n89DVb9HcfRB4TKtulhJEZaPcE5ff+CBg4hxPNHjwOmH5ulr2qRmx3bbiH3
A/bDRWIzdt4NGklb1Y/3a557g9xLqDP6dPpWVcld1bJyRgrZxv2MXjIdyNw6ha6Bz3E9ZxCry0cr
xJkxwrcIr4/6z0/8spq1HDL9z2qsIYU7hUYQmR5/DTd7ew3xxVtg6QO5IwHK0oIni55su5gHaq1u
GSAZxt03Y5dX+S2//icgrh6u2qtbzHPkF6Gz4yocGVCznNI8POmzy6E0g3Vd3V0vrev/RWLP0rWE
d5QLpGeOqggPrsXF2Z1PoxuZSOV1XW/yfm7goMN5s7ROvLtFliPzs2mPTZQHSzNjiwHe94qoE23C
Src3u9Zb2EpXNCv1EsrEhVxXNgYDTALObHzhwaLnxzD+CKudl66Ro/w7T96CC33F5I4mFtOAizxF
kd7MOIEv3M8GuMIjQfAZNxh3ZD4s5srsOWUQnUeLVRzNf+o+q4Leizc5DxmbByhtvpjT4PwPOsoB
oJYujUaBib8sTu+BaDipzvBlovo5G+5P6BayzJimWpe6JFgIhOnKlRfIYS3Epitq7d6xkVg/GIcu
CwDo2Gw/k3WcSMRFljNVkOWD2QJkHkHpStKFbIIp22NvFY6MTnSsXWpIdYUGmzwd3yLTtZ86uhnd
BnghJELSDrcbbnoJfQUsbKtxB7SZhD8/enDprWPGTMg6j4PUCbRy+fZPIJOSV8cZRx+oCWC1oPea
tE/22lshX2fhlgk/6wfNOpK46vlmeZPZCOylIvn4ybLltMmL9kFc5QvVKyafIfuXrj0YIwY+dd8/
xomsmhwaUJ1QMQOae7Gb+l5oJXYwxdV0yg0L5tlWfgsxpxLcHk1wDHQ7I3DWYXYG8j43EROMT80S
TpxFwMHrfrgIlwO2OjYYB8tBSfnSeFCaT+z8l1WbKVmmwR7/h9KfPtgk0tyV9LKYpkM+CFLVuoY+
vehDPJo2vIFGXgzxpZaJHgcNpLtBFpEoM6dUuMDKleh9RkXK9xZ14rO++f5EjcT+IEy4Cj8ieQ59
TOCdTHww23dN3xdgAKueaPbpumYjkFKfw6caxG9RHCKZ0IMpJbhRhD6xj45RUQ8PN7TgywXVm3z0
Kcxx8kX+q8XRsNXYxdMLaTnjt1w03bD2p8PxD5j6ydYR2Yvc9t3jB78MDtGJdYqETpcICiIavUjK
twvKIlii6xPerw83Qgx8svxdty7K+zM3at4hyqsowh1nW27EmhbyMLXonhZvefHHZFd4VTE3Eeou
sSjcWqf4TSFaYV9X3WA4fd5tiRzWr7nRI2T47FMkl7kCMGtyVNU+XO6e+5ou1MLBj22j/Zr1VLTF
V+jdcFjgoQpsv4wEKA6RKZNnrjddKJUV1qW0+q+j0RNMsGln9pisED24pDuQlJWjVbxv6kzyyzzb
j3o0kapg60KpseXGxKpzX754gjC+N0mFr8xNgqxPhdtjpCYERdYcVADzaT9ycCK67kKKxaCvPhql
A4dA5uSuX+ufOaywyphbc3DJ5RS034wdY0E2Fl6LsuIueNIezZo9gcgkduu28YAqBdW8X93n/V7S
65saQWMj0hM+TK3jVZgwyuu1btCcQT7nNfKnHpYkDl83HZkPWbVN2Wsu39Le0bufMDcQbLu7eCpd
ewPK9pDfboeN8RrSU2ac08cKuohcvjjg0lgw4BaNqd51P2opRrzBcLfbc2U6X+YchWQBDQ2RBUu3
1sCh8Y1oJ7hYCi6o13K1xPtg9/wWrZqL8SeglBRy1XwPGU/wvzzFepr1qGGluHFuG0P8co5MFrr9
m7dq85aPEEkzQ/oPpCPyxmtuBH9dYBZ0xARcgdasVYKTDIcb3GqIH+CH9VTv6Ynz281TzaSdQVDm
d3/zdY8ja2rhdPbExPMye0ORsftKWxYppEUluMQb37YebkpcD8zZaOX3WhSwNQ/PC4fepnT/5RYt
qy4ygQvCXTSYdO0bHcbRUthhdLhIzOGLsnKRveZORrQKbbCtwrViuPYuv2XArEwSt2pCmfZ/qDSm
Xr0WOiTbbJ2iR/SWoAXufwOpgV22aphmzFiKrnKuTpco3055hNsE6SK5BTR0i8bqpi/1a1DgRIxE
VkuMeDqOUTLNnEpgYK2ACoDUEZSwYTG2XAYvhfgnbfzaRD6EhvOTKmio7DnlEOuXHjqhGIWsQbWv
aEiZ6BGy+hPNkEycETj75Uj2gheSKf3mVLWHoQ4NWPE8m1aHTTryIgco5LhGxA8S3d1pgGdbTwzO
jYUJhpOo2+9x71Un8nFTUBmmaaNH/PbpkhlF5o2bOrjz+WH7PnqJKK+ESqep9ZsnY06i5zoZHWjZ
xZ7dUwjIYpPXnVSihVaWgDBmK8w7WYBEd72R7SD+Go21Nz9IOhVYG8s5m6leuWq9I5ZI752tV2F9
psNAZaNM7GRjtxZrTIX8Aq4dmPsAaBNxExr6p0jZJM51pD+cmlKx8InYTDfWGDh1nfJ12oo4gVap
ffbt0Q0WDfdVuIlHyGM9Pm3q9i/DFM9VLCVcmKXGiAu1EKAS4q9jzBg8Jk4mRvmf+nLF81Xbae8q
PpGsdXJIWB2P66LWrOeFBMMXGRpWTeHLw55btT/5S15zViQaVe64uWPT9Eo1ZMmQAYN0nRXLMv1X
NdcxJBQktwQdoHxKyh7qouXondNfQK4d3IDnXYbOhKJkZRX+s/z60E4BLp2fh96ZE0RHXsEhQmEw
/aD6zN5wfx2ZrO7qeZ8XK18ufA18Ji+XAbULCJblFhzDzUQLQgGBAOCS5bMC7/Gtwg3wet5QgpAR
riL37kT/MWAxh+wEV3F0xp/Edw9WUy4Ps/X9yPOI/k3nAlOticlUGz2oqsiiMnjGmTa0beeapWza
Zu9ldjM7wiS4UgfWvcSY0Ga6Sp9WbBSzF5FBxKHoLMxTO5wFh9kjVZjy/IQR0rDkXwfdsg1k6gXR
FDHN+Gr0LPoEqVkSXEKC4IV4uJB6J12m15Bov5p5KjTFdn2Hm7ssBbglG843ZGOQtfDojITNgDT8
Kz99RVaobRuJQsM/x710JUuN0JpxOGkwgUz5LOw8UWnswg9BKS3CR4ETwgDFRELhdVWX9MldGPHm
tY5yaRVFpigMPU9avFxajAMmPgBcAGdT67Fh5H5uBTZOuQu2jRQf6V3bjGqq1nBBDEt+iXg6wC9f
0TNxgkwAb6cQCC9sTrBhk8yS1eucNLGynedrY3RAoqHdO1G7buwNR2yTlmR5JfH0SXZzoJf/ndGv
Q0icfNsuUbvaPE1U8ODkYcpI4d4E7yys6p0q43Gtm4/e2V2QP3gID53q1UfbzI14u7F2mLO+92Sk
kwFzKUwMoDFH+CZfNiDs1+/BwbjH3BxjLVxjDbI9Pqg1+ieFEayqmB6p8JmeBBYDt9u0qmGmMOCX
CiJkxaS15L8Hwc/yjHWc6yO78e0lIvZCfagqBVLN45wWqe/ETXJLeM/EKSc0dhMP+SPyt8J27X3F
0K7WhkuoAToYliP4G0f+zauyJIA441JStGz/M1f1etFNKRpMrpjiDCFgLQW5pUGFko6uvBNjUhb5
mqPSjsGl/84sIUqNxsngzxMg+0LWcgherK0uO1Z2blFPXmn9akob9r0rwE5fIhSwPvrJ1sczDqmK
HZ1BysaB81jaJWpJe0D8QnlXMTH435xs1envqqEVFS+baQXJ8QOPkwBw+Zegd9NidWME3/NLN2U6
IiWlubI1jYSLms5B6D2Uby3hwyrBOww9DpATHX3HRb6UzwXXLrCHK9gr13747VMxNN/di1s0npvy
Stsz7ILopMmfQGfDxmYXn4EA8TDpjsfb6QhTy40vMXjTNqWisy5lmz31oGfbAdi50iWgrFZ/ZMVo
6F9IgoGnrIw1DYfpD7YB0FPykBNAOkYhG5SOILXnnrCsBreC4cRvbcK2s0+/UfHfhW7rIYsfcel+
ISSYiBEP8UAEbzST+oxGk7oUg3CRIsQYzIn0IXbtam5ol2hOOA+k+mfDNzZHjL5QM5L9ByQa22SH
gjAts3A4ZzA5Jns0qHdZhufBRsWU7+eeLRbfq0aIHGgN2kiNQ6ZlPr1gsZ5wg46D25UfsGUuL14t
KzgWylu2zQ0RuNzuisHZicr05Tap3Eale9UB+nlhSVnUe0+z5BWOd7Yv6Jz6hb5CIarZ2Ev8jeb4
SPKTY3NwWGdlrIY+QzMdZT2/f2gvLvTBN5LpCFCXyfks0NkaYVrdSLbrilWi71q8quGZqei7z7Iu
oo94nD0N588lwrR2jdOCRGQy6g44URuDZcqmF3GjKP7abxR+7cwk/6+HKk9PZgHZDItO/kZzLluG
EwrOMJMCv8sWsWaa68DC+PPcj8RruNTtbasrM1mGtlys+9fnRjrrIbW4BZH81TLpor0Cz6h1AcA5
Wu/jF4vQJKbdJvwV+6xafPcXfsLf70Xx6JSmaUGG83sNl5uK/3jbtt2QmY0cXeP5NbCLlJ4/hlm1
+HtLpSRhFZUA6jbEDfBfMYEVCLbmD7Gdne9DQjR4+2xNnof3+7o+5sDLJLK8rwc4ziIW8Jxd1UKc
LqPlpSHdLt+sT7YOUIW8zuCHnOQlC7+xnq7vvXvJPvFb+Zw7ThZI10vBZ3POvsrdOTK3X4Ed/Nw/
C/AoikUu4dVWB6Tqtw+y46ihaH6KjaDTEJvaiWmab9HVRliawY76upfvOSCvQ92wGFy0AFwo6vT+
Q5ZDnTQnye+9Cabm/xI2kP1+2CehbjOJucSgK14NyVYeM3IKDbuRSoiEcd8/WcVn9dYa92PkYSDa
1DJPRHdpw5pRoNM5+QQycJmBfaDhHH3L8NvQVgYDdwdomTZE+agvlDBs8tHejUkgZSIGjGdlDmQX
EcskI9ovrPD7pFTWJMspOG/OXWlYm7Kgpf8Ws3cQRV94u17CmolSuqL8wd70OUyMWr1flPK50Gos
7DsZRYt34b/8DR2HOJyz3ggd0N0/9UHDQS61ZaYGHK0SNfd4l4DfAYDbmoYKJOeaVUF8Aa7uzHkc
bHB7bQX2wAM0EUMyXt4fFUK6vrJ8/r7pvGnvL+dyR/01JlscifjqhLp0Rfy1vSYdhO6mN+lUUGq3
PVt5ggwP8Yd5U5DtScn7FcPIU0hw+apG+qXxMAWGrQ9cYbweIAMQT1Ww4fPOwFZxUFwd+8thiAnF
lqtW49cjT2N2GV+2/pxGbSZtJH7SUZMOuGVI9wHY7sdAJcVBTS+ykb9TFd+/StJK2qg7I4vfzGwg
fEYGAfu2G9SaQhUWV6TVdEsBUTgOALXznh9rYUjLMx6LTsM937WQJO5KFNNZLlkCDzdo2p0URSI4
VoeA6yVhe8qALZdS5ZFvrLHPdHQ+4V5frXyrZV0t+Brv8YsxbRGMidYMw17moDRRKF1F/wT4G6A3
zEIjexXC1H6xxnVAjPof80JEw4yaGGm8fhgKOoS++WLHjxnh9SzbSxRLprBxVF5aXbIruh4knE8r
Tfs1QV3becyaVyjX+bTSDHwMguBLZFuzo5uedOt3ImO/IvzRLTiqwEZ1E2TRGYvpOIaobHcILRjC
n2lYAvAyvwcs/SyKOMlEAqBPfGqsas8qAdaVwwyrMyhP7JEit8HipNSjC19589EhCfzzhGj/6Ni3
iJ5E8oHjkR5tcfk5BLVpBcQmLg8BTRy9BfbQkL6gmGrvDfJDR1yBCCGdYEkvUYIBrWO86Teo3MnW
JaN/P1jloIxpGKvB7zCwqvIntkcFnh3W0ijvhwf3ubP5jBwX1+jO7b8rDKsfhQFu8u8I+UoQ0tyy
pKJqI2oCC95doeYfpkTPqteAygYDYNKo6xBK5A1AR8+hw/Yh15fBIBEzJ+cm4CaDuC7jDS/Nd1Ou
fdGmeSmZWklgTMcbAfVEZwxkLLScKEqD6gqbPey+XwiixA2+LAFOrQB/+akiEkgobNYrbHRVev79
PMivg6x7UPbcdpoSTEWnEq5dYaWI6TJyObGjkC1mePcOyedhOTy2BsFm4LRF+uJ39NB+hKk79Hh8
A1GrJat57KMLnhNwal3yPbadQr8ceo1U2RbdkRpfskQAVoY4VxjRGBLdCtDUZi9/Ga+1TnCpal4V
TsVoYLRsaPXGJtV/7U94zweSHv3FQe98PqnTX+CeQqQu54kKBPFLvJGIOJQj8HuOQmfguvARXpZf
RmOV30S9ue6PRlDrHJpUPbg5syeYAv2wXFis9s+X92fUlcvn3Yk3XwX8B0xIdhWlawaAg05BC90N
F8tT5TKfrFk7ueR9ecah7yJ27UGJCSZfjWYcnnOzVcN05vBd5eJJxNB5JLzp7fP8fROGFv7gU/Q9
TPi29VDE6nk1ewcUR8oLrvHSoLQgosM1HX8zD0GvK5P+xSWnXiftG8/VzOMG9QKbH46ijbyZsKGK
T0VNaNCqtQ1q27YeKR6eyHD5P6MUXwzwiHBOUAuUhqAPaOEOGTkIGhFBYtiNP0/NpRb6xKxfDeYN
tuvLmpaX34iqLmTCSNVkRZVpxrHxvaVkb+sF3c4DgKIMb4obFmyUqK6dXqSPi92XC2I7zVMjC/81
Q5QqhAqE7wvF6DNcH7A2UwZKolOOVpHUEsBN5ySImSWv4qtX47N6eEPAx3r30b1t52jXgJDj8roO
ga/sKjXBSq0H8daum99abZRl7NuprRHQt8ysPAu2TTkPCkxp6tabxaot0Y06nEdxgPgg4JMxRQIL
M5Vpngc7p/i7VEWPoTjccnO/hKYHE+tcdizCNpBwCoNF27BOumXbg8mHI3jQkak7vt+ukm+OkOie
KX/rv7NTAz18zN8ZLWSwScGWVH25T23I7phcNI3ynsmcJq0aL93O7VIpZmRFDuFePXZKxKY2Oi9g
dws0Oh7rt7Zb4oKV5EWW5Y+QMWiGSZJtnl4wYZn7m6bSER0Q5qKyBW/lQ/8/4EzgX9XRY2Wu1IEC
lT3JspG8kfqOyfzDUoAoUSblqCo8uyQArtDcBGDv64+waLaSZXkKxpvPYci31sLlcOSsNkivld7B
LK48r/3vapSIAfFvbmNyeQgthXJWJhAzFUFsFQIgxcLfVtDshh6Pk8BhMRex4Sk1zCrDKC/fYtku
UIc+jTfzvsxfRggklqo+76sIVXuDkWc2a/45pEHVPg49yD5JYurWmBgoppYFIeU2Jmq7Y8PJ+puF
mHF7xUmfQMPeIJ+vZwXiUE7fSKXnnwBKn6Sj1QsBNxVBrpYbGoeb5P9OGKmgBF00DoSLm6UNbF+r
yoXx+g6WXL3bka0kqMDFY9lUXpIlgXEyTL2UlmDlb19JywlBbJZVeYODEaGHuJTVHfcxHsM1U0NP
SeLMSdV5l7+Uk08m8T5NotopiDJGELZjuibI+L36sxQrlV/MlVxoT2YSV1TfIdRR732YHzUxxFNH
qQjoXCopnYs0G55Gx/nudT89HrMT5JYDz16HgVdABoinLUHUjqbjowasn1Ne5IaqwFau3nAaIcuk
e7w8PD05ZW5PJZSg1Ck4Egzp98kENJVGCGJQJWc6h6uzqduRfNJ918lD7/VmRBbJwCtbdRQnM4f8
9dOiYFdYzApqOcEc8j1lEQ7pHlp3az4j7IkdJK3CuP6kt+sBuTAnEfm2SsV4oUiQFNrhwwsNzt2L
9SkJ+l4TbEDdzFw6wIFSS3rZ+4gSb+0TVEVBFQEX/DHFJ90i+2K8z1UKPt0+TtpZH1e1n8DHFFkH
qMoickIcmdxY1a5OrfOZ+V/TzvauUjt2K46fnMVLbZju8/ML4uptVK6wzCAOYT19Vlonii9YSoj9
z+ZhBNGbGrbx3ip1k6SBgo5H6dg5AuBHnbC9PU/fzQ7DQiYfQ4WD66VGR8XcwOODjcy379KqR0GM
JSpOvxZox+J7bHn0fbx5eIUKFHiWADL6472lpFl63RbV7ib2gV/EyNU/1HIG3Nmr9EZTiCo425iQ
OH9VZhHrRhoZkxA9+ha0fx8ETBtI+ZEVilUWSFTjqWuwM2Dlq55zvqh9BHPFNQ7ZHLsRbx+0IUkD
NRuXtcAK0/hr51Fw/2i8z/xgKoX6P38JNAnjATfYwMWhLtUW3Hb8MEjHPE8IbilRxXtDuJMUGTRQ
G4fDIWh35cbaaib8PWTL49RBZabXAz8dojZxQEENLzKQQ8fW0RieuJDNkebkq7Tw1+pc5IlSXYVI
h8TOgS1tTdrJ9g+xb0Nb1w+bafiBGuX03TfoFd6DZuEiuSQiiLgE3MVc9S7fuHeR22nRqrb+djLC
OAZvSzxfLTRLUos6TNJ06HdDwSoXjtuYG8ChaT6+QlB+IGOY9i22MGGkL7U7iNT3O545xOIuA2Eo
f2HlEWYInILq4CN6sVVy249JRHnGfHwP0p8bHy1+kwIcbr+GJ4BpfVF+H1rF1Bdj5AYVcUokuiiJ
uPD59P20f55P6t9ADtUG/TuOnOBrbPKMx4UhLmPuKPAte0bJS/wEeI2dxoQpUpGSPgNMRpmtoiF9
5zDxk5Ta4t8xEJPbQJjA+njTVrMDZBTec0XrtUK1VVje0aBxF/ziUSmISRQfOPG+o0sUWdX16U3M
qenyL+tWzORsKnMW7PHl8MYgJ1aDdAPP6yTBAf/nFet3iue/5OWBsMSCtWbpK+yNqBYzuR//VwhC
LsThYb4Y0W7LSjN9EyBvCnDZUnM3CWX2KhJOGGODoey8Tph4OtkuQ/ctlzBrPrC0u25bpPLOcggb
xEGdVNYh3J/e3l0/xfM5Ql52S2bYHQssME/7HRp+u6veeAagrGjI+H1TR8JcDUblF89nfIs18a1t
WErdMHZJj7xdTM/dwlPuRAyz8BqSwNeoyzr4Lt7dt2dd2lKr1F0fXJk8VsQNi7nTnJANE05Ws7FC
Vpg/DBtXuwdtvp+IOiddMCASbVHP6dyrcgMA4ir0t/WmErRn30VjksnzRntLOVgpBvmxLhj/tvNu
Qm+3IZCjq90c89z91ygGZOHZiNcfX9eSazKOZLQnyPY5QWDtH68ZGmzKgNQy23SJUDmUdGZFdtJE
5Y0zOl8W6BVIQyi27oxSxHvx7NcfivDUqVcrdnQspdQa5MrGFGsGB2VDaule/CJfLwZwwgnQi771
TyOF1vFOWtxVcoz0KfPdNQaE7+eD17MYfS/bgnDdRRtMLmg1syOALYGQA+DQIfz6lyY8nVsk8fRE
3hK5XK78iq/4MscE/yrroJELwwL1isA0FGJkwMNlx3/jtxnWGfsC/PXHkWZn/1OWvpKMHcc5vX/L
ld/f4JVjHbKvv/fbbdooBXrF5qBWU3F4xxVEyeKgM16q+CfqKApoQ2kZZAkb94EQs2XkywOdU1f9
fzpidoHHfKDaCY3DLTDh35gVpYdB9C5os/hwbNK1GbyF+jk5+yijJ+97DY8X0dIx0ZDTvOm8KHGz
nmkNFvlWuSV8bsTkSMk4OtZJp6/7w7PgX6zfg1m0GkQaM43ZgWWKKgK4Jw4AknNC4Ew+fn7XLAXo
BEPThwsxAfXSddaNYl9QaZ5SHCB9M3hxpS/1LYOQx0mpySZmVeSad9ufDN/pu5sIzyMlzBqgaM/+
zZXyHzNVzoySo2gBHCSzAo92JPNpOrKy2Cl9SxVg4w5DqKUsZXWmlOarp8JQvGEyFRApovXmu3Ue
AqEkIzbFRgp8BJ+SIj9U3eIUcFCxxwelRnwH78QV0NINlEq//qfIU9A2xvFScphknYA1vUv9Icj+
JUWZ8Ckj1pMK+pYuT+8VlGUeyIRJjESYPT+z/ZcYBgS8FVXm7umLbmJk6S3ShoVF0M0L6E9elrTU
8hJ4ejSnCCg+Pv7Lw7N9B+xHI8x6cuIKmbscbNeriwbYSdkDkauJS9Y2o0YiS2urLNqBf6JmrCHO
F42kcYQf2R0D+Fu4SY4ue+g+psUE9UUun+UQjXd3Sz0OJxW4oezT/SBWDujNDeE/iYUjbjijQHAa
TRZE7MBv1S7oqr8Xn17S5TC+vOQzTWbe8HSG+cv6RkhPOjeN7FfmJHGUZZBca9FWKTNGllk+FvLe
6HGlNfmITKSj2O9GYHrFxKnDVNkMLDcpTDFdel7Nvw/dcCc5Oyk7lWF1n/HbekSzVxIMa7KIruuC
BKE5QROyz5ssMQOr/A2wG7JKeR+iHH2zON2sabWA5LkUUYaZ3gtFO23LCnUvt32cf4QFCyq6VSx+
G6q7BKtYyvS7oXGPlxVC3cRv0Pz+KilJCfpx/WnA8s5G3SQUSF9QLZJx1ziN/JIfxkqHTiDs2hJd
wDrpcLKBEYa9yKBPAE7y2RiJw1NWZNpDhWxFjXTXpayplqH/7wr/btgfePLKO2MEVuue2x9X34e4
09yku7qNc/ne/Actkxz/0DGqAVmZA7cZ24c5mVo2f9aZNAw5oFtMx59xL9H8YiiMRKt5FZaKM58Z
v8b6z1TE2uTlDYABjANIZYQy5u6HqLrOH3IDlk/X+WyyL9DuFHsLdkSdKjdy7YlCbhc5V0clWBgY
nu9qO/FUzgd+TjLd//gC7Ahn3wwFYWvXzCBnO8SPDQ3FL0wKmflGQFCIGktQklg1EMSTkYId0SoH
0P7aR4+vb8mKe8L7lUyXBbjZJm/qbM7UrXRCUd8YVFjoqRlYdJGJeEKlSy4naj44r0M4y2BsWQCF
UL2QLggzHWY7QzZZl3mRNdvYZfhZ06ZlD8ctEp5fKMLkbdFV5p4CbmbdQ62GWoaUgu20aQCyuFL2
XhjXELAGGkrotIqJN6dy+t+V1FyeTas8DyKg6rxmrfDBStpdgOrl6fyvD8F3w1DbfSPwgLBQduCG
wuLegnk6DxD2XncCZuCAahzGNJCf0VZHFNF8YMKPcp15UqwpNCLMRNf8FbHSRIa7cOp72oOzxz/4
TZEyvwKjK53ubnJGf7nRUNmrd0HhJ+Snqhh224Ev/PmXEtJ36l6j66DNcHSCwvWWlQwg+1NAIRD7
nSMHOZaNZqaMX708ldu6scMrCHrFr7D0XRkwDSDJaK7HS65sWs4xr619VQTSDVJKLlC0FCFYfVG+
+e+EF1anDD2/smPk/PFG8wle+1ell5jR7dReBlCy1AW3Hn1g7JBezQOnng7JkJ/FTZofdCbY/H0B
xK3fk01bsduXGVVWss7JTsURybs98kaZ1kODRsbb/1lKQ6+IYU1qEssm4LRxdLMjsgzxA14al1T3
SfD54g2c2txjX0ickCnDGAxaAHgvKGPTV5RBG8aE4TUJPFjKe8dU1yiH8ycfr4dB34G/d/ntpNqH
9rmmO5bzGSJFdb4yJ+gr0SU9cKCJIehSRKHj+viRIPXNACuWDCKbJjvc7Kdeyyd2Kry/HaNJBSZy
W8tD1A+gyEerUO4DCpDQePOAR8Pb+wM4Ldb3OXv3vqgBiRHOCkL6QEe37RHPfPOnxVN8OIfbpAHd
FiN5noRZh14+cwoD4s1q2wpOg0yvyYAwim6wwy5d//LJKvMtzcWL17Np2J5XRpmFoZOQaY15qy7N
UufjxA/QyrRBeuAnVzRifOPTLwiSOtY3jt78Q0UKf6GJWFY389o0BIVTpXpKQH3U59ndJNFce7tm
o1oWoNeMLeLzjXSKw6CzKmBg6kiYNh0K7a3WR4PeLZuSPpwJ5/kNyz0XWacZ8a1w6K9heLStr0A8
qMc+eCqDsnaDfb00Zz72kAL/6tDEfMCaqmY0n0IuzhsAXKUJqpJjouathTjZqBoqp+GRVqGWhIoW
6zV/2/Du7Hca5du+zunbVHsESsUnMK9nLotp+h0A0ff9w88QANGNZjiPFiTIh7bjlvGBkmwJzAOZ
0tpArkJdc2M43NBJNp/K2awF0/VjfvJMhOff7tE8czHZHennxmRyTVl6MhEDmtoGDtVnrSw3DYmu
gVz258qn8kNL5VzqTZdGC8oOnYQeOHtVYtI8tKKIb4u7DqdnkDy4e+cDPNRC8/adJwbkAox9mRuA
s233mdceVY2SvCK1umGQa1OCN1calaWo327DBa0J+/x+WdVgtD+IThHWKVys2zgpMQU8qQSXtASD
Znj5KeDGYcjDdiiDQvFCWFz/EP8SIMocQdwkbznzXzCHWgl6xfUgniQHhoI/TCwzWZbYvJkens9T
KdSIkvfsWum+lXlchCvDm2wpls18VkCHQZS2VIsXb8WRG+35hSJzi5H9Yt1JPxJfT90wIm2d1ihr
JBMaKlI+xOHAWcTAOq/Q+QfIfLLRfqYubt7v7gbvnAOUJg/REBU2nLoht8QwIK3Kp+DdemU1NBzL
wN3V4b9qkkFQTXS8YVJazS7XJjFFZYSUQqZrcF7gmyzhrv/BsKYdiu1Do6x6gQwYwAnklLhLzCnP
WDhxMGc3WPNV8/MFfrIa76STM1XYRLXO5m6SQZXSMF7iFfZOnatCC5Y/i1ErnqiXwRcTooUQ4qfC
iTp+7FJOYUrmQGQr/gzqycA2JTSyTCfq2Whd8/lwMtI9PotzP0sLDtO6mRxSR39wLQjlishC2fDH
5WdiLBS7QZhcHeSrQT62wi+js0JRdT6gKeYV4xBctnNdaTbvxdD15CCS/WmJ+wmo/a4FvndYUEll
AdejAaQ4AdoKHZS7guUEhc0ZVpbFYFFscPmJ1Se1+EtBzradxgPQBoB9rAXYVsDjLVCSi3/AOQi8
N1+EzWbNCaHtMNzUNx4CLkPiYliJUTSLPzuaH+m3BrsHOrC0I4HX19zV8OLHR5qoqfTFjuzSDMuv
5CB3t3SPwz+RK4fRmHFrWJdtuetMVwlttRgyrXH4EGIesyhp+oDBoIY8FgfLsPAiGr28O5nMP1LR
Ubg6qKEyH/niQPgBsmN59PJo8ZYz/vJqwPGzeTeJYqIfw14cJQRpdefjzbyspFI0XwDSBWK9VYiR
q+egEll8EHuGtMxM53EogxAj231FCqndFjktImGRSJWcY8qy5caTPVvUI68oWOZJqYuUDhNeNlO+
nbAe9848UY3wlD6mVhUsNnsfVeSiE1echqca+wR3f1VItGekQSQ+D+b/OZtaXoH+K0M9uWkH/zB8
e5eJ9mheZWu0EA0+xvfdT72djqsn5W6yu8XRdIP4l1sQ9IaecLVCHOA6/UfD6CFieTgZQnxc3Dgc
TLlAGefZL9AvFvFDa4J5XiE0323h6FH7hRXNuQlwnApM7ctUakiTlHQd26N9ZSHmNxyABQFX1YCF
x8Tdgcces6t4JaqAqh4srieUUTM+Y/asiB3uC+G1A+0vOaCbOPDIVRGE4atACST+peFdE1gXaIKM
EaBvGz4wU742KZ0DlTu9tI/ruiL5d6KbI983ZkvI3MrMm7FkIZ3D1fRZuB+CMRaPsx929x5LbcaD
bXz0sbWvRMLTdR9+S4qTa6W9N+PhKBjxAiQ7gcQdUtSjy5saTrQY9yVsn46gY3CGIH3Fp7GejT9v
CWAW77v/Q4P5PFtMyzKkazoGR/SKJ/9QLXXayfRCmYK80IxJl40PJbYs29CviGampjZs8q43T0Wc
dkzl6R7qX1ktwMZdP3P7CeBsBNyLpBLD551IdOtxs6tCHaMgZBQPgHMcoQyuxfP9EHprruc12aw2
bmkrh1jCoaTPvCHXZWMgHe+xW+1POTb/vZxStG3/ur/GUgfMq90avIg54imInvk/Msbe1swzaov6
5qZjdLD9juBjsJ34KV3qic4anypkmFP9NkTI857EJMp1SstZEGGvG1FvaZ5o8+iSeKhTxFFekhRv
AC2Rm/v4+Ta0NnWKXfxHZBF7C31t+ET8m/zb1F0nu+LIR8GCBacypgnzpn23+wzbyE+eyJJkZumQ
yl2Nf/BhY679pihCrI+jZytJpZ1eCO9OOo6gjK7lsIGKvY87tU2vYHuXrxE4k1rJy3iz1oS6xt8N
hmPGZwcP+ZJvSwn4chS4Syst38uhv7eOOeDTvZSNflzq0ih3mufAuop3m/Yj5y1HeyFMkclMz0Df
u4HsnXY+dyf3Zyu/Tp6nMNAH60TLk/wHSM5s7DHsCNynNG8uQiXT/iKXDL/O0V2brvFuTwksOK40
3y1ln3ZvS49IFz5kHhFrE6mqpBsKOW1nP76e9Wv43/jlrwx3y6gRYpppOMcUcNm0hbLHfvgd1Nc/
udlZNjfhGqedZV9WhLyOz9BQiKq+7wLX2ugDtkogzyQyehqHTBfwjp65kLdGToWG4ZttlWO+QJDw
yik7n1TIDDk1znspeuAj5QIT3FT0Bh/z82e9kJ7YVJYTjW1dc+i0sOEPpQx7Wpo2x0ZQ832/0lsP
b5jRk1ONOEPnVDULKjU9Wqc1QY6vnkl8PjWVLgAuYpMU+0dSA8nn/O0ajBe1Sb0FyONGhECEwTo4
lqcKt+pFIaz3ofC1WibcMGH6StZ7t1Evue6h31lqgQXe2ZqUa2TpVjpi+GgVWZY8HRWxHEi/Eg5H
mk31OK2gQZsOUnPYHifdPDVh6MVdlbb47ugCiUdHK12DFx+Fs1tV5qzIk7EE+MV1D3YGMDpTtCFk
VxGd79AWSgZso+8c3wes1ccyhVsafBu6pnZwwQUcUm3bQ8PYLYBzW16nS3cKkCNlSkSwD4NuIOtd
N71TIFuNUAeCTlRES/vi/dQ2sgc58zd69ebBhJpHDQx/BGCycksT4w7XBQKPRTFJ7I6c+OnPdGuf
ELyFyQEGLKZJ3knruQ6O+xl3oMKPmA0/VYSSAKSIJiTkCUb0ivt8nHXyH7ZCGslwQP1JUheRPR/3
occRj6Uy3bBa2K0hbwjA5hrZfD/4HsgtNI0pN5K7Eyn4TNmhwgCuGmJjAsesmo2mqo7zzeJSm/kG
Noe8q/caDDxUiGZu7k0V1Hnw62PTvT+Zd0hqJnhydCLgvdq6Cogw+dDPsr/KHoBoRw1BK+mGSFMx
UTty1cvcqhCQ2nZDgPa9XowBE9J+uim7sDqrA8s46JgGey7hzLZoFJar3Ac5lTSbf17JJFsaiP11
UQVGP6giXbSQ+0FcLTp930OlL3j9Hk9T2Ir9Tgv2Xdov1wJwoMAeVtRSL2APdy3xx1PBb2k/K7cy
8ZOWCc4Rz32aXhIgHKRrs7dyRQmsv63wrUZxCTRRk0LbvHeUFqNUyqkrCTLe2p99fvkD5NHDvw6T
xmeIjeQIj/cBK0rOSyUkt+OuU095AP3bTwHTgOL6/oyzqvm6F/VpfYUELxtWB1g7rwfuSGX4sFHG
9BXm0kP741JWl4syqGXHrLesiyuoCkuUm95dI/LYw06H/jbtBzXz0b4a8B/QH8VLt0gqu7KNW9Tu
CGDCupDOokMK8LyrARarbsTl8mNczsP0Dtn28A1Ijt4w60HzCYmN5c06BpMepA2alrxRCWMy/HI/
Ey0fM/REZzIKXX93QluEjzoI9YFkiOmyGjp+9Ph1iDoap8LcJV1r+POG7rPsaW0HcQJbv7BRZV2a
VfYyPkgbTdtikXtUh+aSQoU3WyYhbp1RohOGm1lTmiYJFS4jr88isSYQS/7XzK/55vncO5DxKt73
HQFFG2zpv9HGGPBeAu1VnhRhX71T7uWRowfgz+7KsdXpbKHSpgWnWtnzPfDypCigFqD9cs2GK8YQ
crxRgToRmaIzY+HMDhwLG3N8VyVqRZ17baDTlNa5nj9cHvo0eBdYgBfAmUlGbGKLDmoxtULqtM3X
SShz/QY7tY0ng9xXYhNtDcd8bBfw3MLpnOW9+aFme4kv4ro5e+inIGOeWWOofdGdNPTaVSfmYBxj
mXB2SOTlDoygPJ5HWWEBfyqtBW5N5Jwdcd8AyZZSpET3HwqAjfJM4RlEN3CuBaY6uiHfq/i4eao5
IUQujY2X7SIoQYF2YsQoiBLr2EkhkEIMd7TwaP2ecg+C2Hr3vpkwPkCs8dyeFtmf9Mc5DbpoHxTy
EQukhus8TXWvFeljmAD8xOIXi9mj2b42wKoPFW3KvFjCefJx1eG3tDeJ9Ofbg/v133gbrZlDXDiT
BNkBBXp+qhZ3pBjwlD7rR251beMAbCdgnpYs9BVlimMNSKsl+Hc58sTbBOQ/e/HLtD8XOrpFiiPr
mXxWrKIluumMa61cdYce/RDb92Ec+jVwNXbpRgv0Fcp0d2/fEpBUVuAFNpp8z8ztgVeSW77BaV2F
SX8C9d03/x9W6zntpPJXAiaW2zuwPDBRbC1HGXhKSoZrcGoE1DPYENHi17gXMkZ63ZlwyV/dT4IV
oHyZR0e44IYnggfD4DQlw3jh49vYeooKrH0dXS7ygYmAf+b+CqoP0oJBZbJomSjqMNr6DfX4zAN6
1Q63rSXuBviLJllv3c53N33jA40BRRK/pvbfBRNAi6V0RyfWYA4esZiKbedvB04jccHSNaKiHvQN
WwX3kMtwxGwu2mwcx+aNMV47vHqHGrr+dCIpuG3wVrlP9d8D37JJwj06drQFpKqRgAGpRUFaZ4jh
Iyau6p4eGbzpApynAhiMD6tSKdD4IHPgp0Dc42pZVoK4YAs1SJ0QxR7Z8YgCWowJ2wp1+bbDj2pV
BP0FC08+nFsvgsexECl9mj+tP7iWBar5pfJcxAlFA4H1Z2h1XdMVKhuhOLgkLc0EyYu5c0wkrdGX
pcQ6rTEGHgTpFAxgNDAN0g+uNQHH5PWnedd8GRZufKPKCYe0qZgXatcZ4baPXwfQylw9jyYcaq+6
XRB99MjIKsF+ltpL6HWheQpjJR9dELolRVGtb+YAqg8us38/XxKL9I2vbQi5uuasfd0HvOvCMoNp
rcq1ybR3/IlngkgMAbzo7Z3v2ubGER53cJ1+4k4ND8Xf/kFmS3/jX9v7b0J319x2xhirj89lQV7k
XlQ2mSF9qux2r+EKGR4EqJBJM8oPDtBikK9qTov78kVqadtKPg7mcHMg/c+jM8tZ1HasT+ieE4je
Fe8dr9iBu8o7sehbEZD2gJWe9n61n8ciu/WPI1Te/Q1Z/G9fjoYuQcKU8LL9y4331gbzqweWbvyr
eoKPviFgiKN2+/lEpRjCcmDPjeBqwADCqOSXfkuidL/vbtGTqd9JDbuTPjw9fYFyKqcPzBDVBSeW
dgef44kLdK7V/04cu74AJEG83NwxWYK7JlfewXD0ungFMLTrdHrk47FGN43yJ27ShJN33b1Hn/LP
YJ/Zpsdz8ljlt6qZ0H8AQeiFGv/NoCOt0si7wgxgZaVwbmBdFpaqoR8FPEm8rNTG5cdu1R7xRH1c
/ZFOHgGjdLAtiR17THwdP0EJtNczORa8fln8sYRA0e52euMmkCvWRABH7+jETiccETrF0O4d3Lwy
x0NNtg7tiXZKe8PCraIUg9sbj5fYhhcOwXau6aMcUBPBgbUJBYoJOX+0DFRroBpUvc99RtM+R44o
siBeDkzXdJ4bn/Uw3zBxF0YxbdfgXVGtOR9v1hO4bibWiSYqR4HmFLr2dAOuMmobRlzEbU3BEyZx
ZswWNfKSNY2l6bZh40AutBSnqXoHs+iAhBcgdIloYto5TipmWfKL33BHh3jvtdf1GGLAT6dr2VjR
OswJX9lqT8jFRSjMjX1fxTViSmdmycrIMVKMl78C+5aCozJDqEHelsYms8rI74HhuMPwr7/ccvbV
kjem2chztNYovxhCrhc/TZZszlcRLy2wbJxWNuy7tijHIA8v65SF9eDHrq3szpJIgzG7a7BR4IsU
UUDsuBEl0dxosge3t1ogJPdrZOR9wkz6+X3AYDTxZsw+ZeQg/33wkB9S7pBIdxAeiv9+SGpUZthJ
VZRyzwrI2AR71zFfZzlhlyGmnRwVTVe+7ZI9h+mkyT2eeWF0chv1SQx5FbhEkgbr2d+9hHqJ0jkP
00caHqjSk/kvdkIfgx+HswLjC7d/vVqL1sLn9una1zwLGbBTM2JXS5F+yvuslWd5Om7urXxl/4PO
G7vnr/9nkTKnoxp85rDp7m2dUfhGBWr3IzniDF58euHLFtQ8fiSA9yg2ow2XGWDCFLKiP5F4GXbu
6t4NmPuEDhuqICJdeYZUOoBCCfxT3ZrMop/luAHmGAKV/qQ6OPp9T1itUZaVfY13cP6ILyNARKM6
U1ZHD8aWg/wGoyzvFKPHf3HXEIkP1KjPGfacBWBZnCxBid9f5rtSPnMOczfrySyIxny5eKAKpU+d
ZMrnJ4VOzvAZMhfBb3QziKze+18kkCsz9Z3ED4nWcXm+y0QxaJzC6RpKfmls8QyQD2S88PDbPSbV
9m7jznC0UZbDTC7EEdkaAFsNSSd/yLHEf3Srz0Rh8syDLbWgfFZ+Enhh3GyAdJyyHl3BUEW0ye4g
jueoiXd6EEqNJ/+uxPI0X0Zi7ugxYKsf2FxaKg5aO2+lcWjR+pb/HcV5oQ3u8vapgBpHPbHR5az5
bFt+MbvYhh+s9wCcXbRVIJSKoMdlQgZLUidDji1nZhsoHOeYy0fCBrQcu83zzjZOjAf7kL6ophZo
LAIV/BdhfhuaXoqfFoN3lwwgh7Pz07jLABH27teVWoTM9RE55bq/ytJtmplwy3rDFgs0zsUbQlym
u8lWK7zSgFvDtMFGfMgZpwfv02Z+bpMWHphIhElmREJziWVwAmGAjqC0OnfhVV71YZhUq+0GZW61
lm++DvT3X4JySXf5tytTN/mEmRpZ8hCT0u/zmCFfDvNKbYXhluUyRZRAYr4Mv26gMt/6KimYFsTl
RZXf2N02XPC28XbqOTDYEbALlQIFspW2ItZnAjj1xfQ7jOfl12D7Y6t43EAUIKhg8Cz9/eD9yTRR
mlMcwtHp2HXMxHlFth2CXE8bVeu+9UaUU2Oz474n5DWdmxXl3WMvfIbGsbQPJZ0Avkvz+ytfMgyg
LwrXo8MDsfUKyWU3o6hCPfXMEffkBowysiL6aaNIQerCsOtA0mxXlpNDFNBxZgUQjMgvpma+Uj78
x1XBJ1j5j+N7Qf3TmyknAOfUJSzDulN5sX4N27GLj7Pur2qi659GbNXo5kN89eGuifS54TlQQIr/
YTPN6jbzXT/2BnKCViZhuDa5zYyg37eg/GycHKzy807E9ZCaD3mc3Heh/slLzSKWllhs5KnRL8HJ
sU0NIIXl+rfl1rrwIdDz7r0YiwMFseYvWB51niq9A+E0xzr8SojfQycZT9b3SfZeIa3QhJQB4OIX
eDBlw2j+q47WJEMPwzBD/G1x3iJw/4xr3TbDH7E2/WkhuxyzyeGiTTwlQhCAxXsKeFrjKEhuixL2
3oWhDLJsnGMC+InfFrfuBJU+e0kaBbonW3ji9KEjMXo+T1P7X5vcQSZz8llHanyfttBlg+vRIvbE
jX/AVcZOfPQwIthwu0+VKd+XLMCMdEQvblkECSzJHyg5Rkn9CO9eZlUe1s9vt1zdgKPmNtryqspw
RBPF8wzkeJpM0KBZg5FQRX5D7MltiBg2ni5LORVFrHgyoCW1B36uMfFrH1ZqZ/lYuWXr7FlR1aC4
2suDPG8wHm2kNxP9Lgj36L9cHSNn1qd/rcuaOkiGN0OIAwPMUQAb9vqGDnyOAfGl86ZJ8kmMVPPq
x1Jzp9ceDFBaIL75e2d0cwvkMPQtCnRx3Sk1AJdUNtHjKHJD5aFcbAe4Vp/F6lGqmmOcFxoNczNh
oq5rMUkz2YCMBjHv30vFjTQpEsTU4XPstJWLAzdj47fhBFB889LbDLIRO5gWwcvEc4E1LXQnfiXS
K+kEZ7fu2wsNxHSI4AAy6mZqFmJysVBV6QG1BdGoUcRT2eb3MWMfWLIAsz7t0J2VAYIvLNjKWyHS
3uKULQ5/yZjZ0XQslXG6507SMlpsvbmPduypowHBqM4ZBgGVFXGfFprtkeyYnZso5RfY6mKHhLjh
gfCyDIemvgPBCCZ+D2pqRRSaP6uGcyE3C7IZca9R9Y8/HOso2LjJgYntUrk3EOA5AF+eBV6WY+J+
YXrsabLrdwnpApr6edqwkQ0WJwigX44FkWX4dF2fj83Q5pX/op4G9MexSvCABGSa9mYUVm3U6xfT
f0/nP1gMpOGH3OzmEJDRSmZ7xVEuPIYsUepqzoLxNg+T8iPBkWBIVIEX7Er5AkfEHwl4Rq+Z3YBJ
AqJ52tROntl3+eeJuSXyrgYCYv7BpOeGJFhgc/sq75o7FLGqJYpCA3jrjoEV9uV9VHxw9y4Kw5+1
vpZMAenf0G00opltLAkgsxLhvbAhcOkmrxzhMmd4CTVDvY8pTgOMs29+4QSv7jVBOVhR6KyoMKAm
5O+8e3+L6J3FwzPvRz+AD8OkcfOz9LkI2cI/MreIKVVa5kNofplfi8kGFRC7ud+h22EsHWZqeUVQ
WohnKrbtw6tkKfrpEDCXY4VuIS/nyCQw1QBhTKqQDd7ep18mT0C7zHgAtPpiGl22jeucYWwaEfmG
CAw6dlj5KmNet2mk5OvsyO3ZriC21KA4cWtA/9z1ppsmBaWpAvw7uJcpxS/DWHRiy5Yywo51yQxQ
fKFNKTiXwfiZD0r1wB4M+4ifUNNc3Po2qXxKvr5KgEaBUkVjIqYtxDipOW2qHdWiKXp2Duj5uM+G
EuQJOL9netHJKJY9X8GBIvqzcvXjvBlDLx7ajLxqwJE/1uYLSNXBMoaPlqZEeZbj+6SDM+hr08PY
0BrUwBbJxn/mumoc5Iu4/+PPk6E+gCtfvKodAgpxcrgj5dFOAT4nsYD8u/2KmWsEqOn5GmObutCk
1kY7g3w6hcQqHMiLK3Ga6yRkkts8BuES2aseAYcUbsTiueLr8bLcHzqr8RNcRsXc6rqowcO1JEyA
0pzaMNhQVbpE+5MSZBFgi0+Csc0qVYYL4RU1vg47rq7YcrCpheT2+uLNz1PGmqA1EiScFSTciCx4
1YS6HrTS67oSH3PATN3WoF/nwANjtkjNBW4cqlmGUoE+d/tfviJ4TRyJmvJZtq56b+ZPZW/EhkcD
Y6Tr2+U4SNuScgto50Hn0ZHkanC8wqpSul4z5ys6og19HEq1pc4nwk6zynDk/CdelI3azWy/wzN8
WIpLvUW8rGM0eKTjGVPgxjO+S8fI6OjvQNDhoKUbalM+DUEkehD7G1FkSO+Y/NOqcJR6+oJfXo0y
F4rTigMJXhNZbSvULc/5BeOof6tVtsJnKWn0ORlM1f9zs/VN/j4ksqxFf566t8u7oOps4FGWttOM
7VS5+9KG3wCvGAp3CFp51tDUZEgPRVbzyOOv2Llq9DbUwx913VJPKH1ZLSur5YDvj4qKo+s/6lB7
j81oJlxhwDdoyBd+sjON4dWLF59/vMlbf4nN9uAbQUOZ0d7DA/ifOmXtVG+GHTSXxZOd7yjq1dQX
8Xn8TCTt5cUEdhtjVQhj5RlmzPzYf/B/2x5O+fjFGzyLxCFEIf67NVhRMiaj8CHZMoJylqTsyOJH
xcjDC56It6SK5kUanWqd7dAhd0q/LkV2lVX9VBfa4R+IREGyyFrK1hqv645i4NRY582XpqCxl3ri
ibYfauwRNfzDv7oOL/28WPU3TJhWh0G0oKGTkY9FNUOdJrna5IcTOYACRSTLca88W0R2KqpO9fsV
h31ZypR+ksoCam5WP3R7pG9Kn9PO2BUPUhP6iRfE2puXSMkpzGFx7Yn+uYWs2lgkFlbZa0ucY0es
/tucpCccwHY40r6YCPn5Ad64L4vgqfTHcseLfsz45MhEdEE5yEy9zIGTsuxJyDnS/oIckz3xVk+v
ayKU/miSF1wWGBS9EaVprs0pJ3IspPfmD81r8WZlhZ/nht9wPqJnW4ZeQnLI6f503xCwAo/C+U5Z
d2wSGjtemsIwSLw5k+iUk4jqAbg+A6/aLZ3VEJrK6j5zqRAA7PpAkN7zo88hlEbV0FRiXQU1qpZc
WDS+XQVKzDYGupc5hTVuWKUTu3xKw/7TaMtp0MH9NQ38CW+RrZ3TJS0t0h7CrSmykJAwP1ahdMBt
TXxGT9u6TUb06xe7fZLj0+5kpeMHIaRctULK4wgc0sZ7UpGA/gznxZYG5vXiHgZ7D748UjnbUU5E
UMjCyliXX4/1y25vwfJNrTd9EE1hs4AlfVCA80Kv2YV1I87kXhmdoH/GgKrpkNDTm/c612bXe0yv
Q3gszZ53QHOpnVfLid0wpmpBVGBuICplNBXvmOKTsJAUoVAZIesi4IMwWy5uZLGEpTGQMF/Tk2i2
+qK17X0AfrQ9v9XzIkMohxhqyi7xfw77h8DRxWwQzyk2tC+UwS8fG57fxaJMydX/AL156kQHFuOy
ra+yfNtnWecHcyuQ64gYEqsNwBb1gXYMNXYvNhbXzN+lG9CmjiBAS89xqcfDc6t8xKRqo8fCHjqo
avpsko8lN/vxGdQA34ftmheiPK8aAdOF2uKOkZs0H9P6xxSXbEFbZ2X3a/ZmqSKtbuDIQ1SyabZY
RFOFOw0fVQzG4JW3zHTh4uXfUdlIfjIlizxNpuucMzvS5R8BbHGUhGPkPAz+JQMFMUGKyPu7WEVB
w5znUjUnWUh3d4bIMGkwWp1pyYClFg8mcFCWkGT15p8QG4WGk7Wc+0iwGZbuYFJ9S+EjPz8ePtrx
Xxn657r2DG/DQ2PH0bFeX4xX1cVjUzTa6zDxRNUzs94kVU1sCSIEIZs0NfLCd7BV/lRUkk2Ifadu
sAxqDAqEGD4enRZaNY5P3Qqgxu5fqaCSysPSQtIsU2RkzoF64lW6RoQ4Joczrdsdj5iSBCHd43NG
baWUfpUGDQ0SzYgZtga27HNxvCVAS7orHSGSCG3Eg1Jf3lzlZetqGGLg/NTu2t4kpOEd3P3f4bZH
9NmuRCKXu64JauD+w0BHTEAMqfFy7ml77RTOfNKmfC2uigSb0qRQLKa7AeGSlMa9EpOQfXpVYEPb
afzx31A8QVAyO9nGxAVj5GpnAy23ewdPV0GcTmcZRKxr4P//CdPHGXg0HlpN8ebnBol2AND+P9Ee
L5JKA37IOLRyS43r4UUK6wM2ye6SRX0N5OjRqBWY4kBFFpjVwTX33DJv2OY4I5annphlN4Q9ISXJ
vAfOUhGclr7yjx2Fbso502rqxU/UB39IadOLa8DseYGkDpgjlSCfeprshxSSTani67KjecgBMFe0
eE55qimDKsazXlQdw0PNzjP6GEN1zxgAqFAAeJcsnNjRGz67ZsBK480yzVabWF2C39hic6RAOeij
t7Q7gAkM1P2bD8Trzh1l/8eMPfOXUQlC9mBAi8YM0JgnAuSsMWJH15wwXJBOuXEx/WBXJwtPKpS0
L0g7waKqK1cF/GeEL55wd6j3kg0OFSvVEXyaDq0nckdlbFkHEOBEk6xVOA6oNKT/Q+ylmB52AySE
RWrdUkeWCvIua2vQ8sgx+/HyLaB2zpRTxErIy5LAvCYsjv0/8kjOszF1Jfk2jbjeXamdmMDmd1S3
tuwes1zL9oy6EyM3xyUi38lFiwRMhIpaaIfJggTyFD5T5lTyL89bz34I6PTvw41XR8moJSVnwsed
e1tHGj03y88VNVp5+dfrHh/OXeEDf/9lM6Kft0gQsGtsWWyzEIGQxRlC1CVWCk9FdeN21lDadcoi
Kwyt7saKap3dm+EM2waDK6vvxSSjcGjmSzNEH+4EG9w8xgbBW6WVZiZLrjjOwbqIEzMsL6Ii2DVv
738q1E6uM8VgOcY+xmp1/U2h4mplgwN6JXusGV70ACze/P9t8TgJgzm0lEn6/l6iS4d7puewqvSf
xE3JRFVLmpz63sBsF/oc0YQP5xqg+1iVyEtHdsCnxZFLe6wIzQ9PsD4zpUKfISbuv1lFlXLa0hZ1
gNFsnVfd29wjywKUBld5lc1J9A8SiH9SHzlQgwcMt/LpN29R/jukUypVsOOe4m4DY3HXNoNxUeqR
NuZIqSQhZH/8CiFjbJR/mbNLGlJiL+WlrYQ+uZOre7boCO1IF4IKiDHXooTNMtognBbVS+HY+SDL
Fo+XztcaYMTOL6znJWHMnpeST3qRpgcktSeY/SNWK64J+ZLckw7zFR8iDi/CX6DHVkML6+dvDsH4
qHUdy7Woo/5yzw1go6GuR9/voNQzvz0kXOi4KuhOOcyI3MH5IeNeGEgMGzZIQgH/7BZXf+6TR8Hg
e2kfdERGMPj0dQQk+lIQbq3m/T/lt2yY5IrEYujffWVMzqLFp2y9UViMtYe4n03vdIZfW4m0dS41
rq433HTigj38tavnSgs3G2TgwX2tlxbV1fEf6vaVv+kgr6wgQbr4JzrdmYm8yUd32mmG4ra5bhBx
vHJpzSqXgN8avV9z9rLAxIoToJvrCnh7TB1O2rnEM92y+mk9iyWuicEEgM5DX2CbwK6CfybYA3sL
GF53+Y9CE/gVIGQlHWTfY9G/syyYuBBPXC9gx8Irls0CxPB6Ahezc3oib5+O1pb3R7OfWMj/0aEt
xEhMHLSGOVbsUxa5ON9dgla91gZeM22lJjwYX0P2jIcvDhri4XVXOByGA10pGBvHzhkG9cru3V1Q
D+TAqnLTN8hFvf96nv4GTpd+MWCYwgNMBCharH/Y3J9MVd5IrxXl6G5OmJSnUqhzTpC+grf0A8/i
Zte1JU/JNxO/nzjNclxqRuK7JxA3JVocxkW7yadni6eeLcm4LRxhAwoRE+ckbVBd7Gght0pWUXu2
l5kbdE6q6/YAQb5ZGI9WBccl9Td3JkvlDWdk9dj9HQAa0jcdR4qDowoTXHovlbNA09p5TDRY+YN+
Dv/xkRVXLEVBPk12n6FXIXJQ+F4nY2xe2Qgin8LlGZW6Ar139C25WUFiQw9vFEU6ORqKPa00wxCk
hhqNivzgRLLtrsHvflvK+F4hp+uShUHHzS3+cuR0bsZGgE27uzVZTNLNyEN6G4ZZJnFotW22LwDZ
jdOQIWIBh+4J7XSHUodY4mxyS51gbR9lvXDz1aUU7g72krrdX4E2WWEpZUtdL3tKgJQeShyEoBUN
4cxy6uaTKSR8VyAR65lVf2HXVtxn3AnlKBxw62PHsDJztWrWUap3v/im0PD+Z9PEGHu661EybLxV
esCviU5d819y9pNqxtGde9wk/DjwTQyAxxeNQiDUPOzydERf6BObGqrj7Z2TYIlpzvzmVqFP5W0R
CIjY/UqnhiMuVsPMuHWHLM+rA6l446KfawrQ6+UJjapia0+3lrU6jSp+nAWf0p+mZQ14sMborZOF
xbi5KClezdnUM4X40iPLZmpOzgGMXkqempkBwJ4EQl23KWPY1UKrn0LiH76pa/7mC9Uorh2voYWz
qLPtgbZyyxyaywdwsItfb8qtUDpJvXxMu4hal1dyGdcMNRshcw7Ma2xaqWyO8XEGKPZKuEnQJQpY
S9JTOlyaudWSqNkY/CPy3NGKb0ayqi065y6fssiuzS1zM+WfiEMRR5Srx/OO0bV2xhLBqotGxx65
bLXwgfT7KDY6bWoivGONVTMhO2tmfl+IF/hY0M1fZJmsmefDgDN7BRttalcbNuQDML8vh8BYHBJN
P7beIzc/hd7ux9K+5kQJNYKn4D7JE4wJ13BWlvsnHClnJRi5ZV8k2mJ5b4/irh//AetPqzOkgcmM
ZQXZchspCh+dZnCtUnLcPziJLAJN/A3AoY5faUZY2z276suIDI5IV3OCTvaEoFO6mXKHUbBfwdVA
t5M5R0LViEzDTL9mN3fsK1Il6Rfu/gfZZh1iAqn1H8Rg9o6j21Gq8wyYhSXW3Oyj3WigK9tBtFtD
//W2wb6uy7daza2HDLxK2wq/lDqbmqafL5xqCC2scMrHi/GAdOAo3C22NV6gRc6G5sGW4kzV9DDp
KJtlxXdbcHvX3YkWYfjCQ7AY4wrsZzvkz/zYEN6rs2kX8qFBqwn9uR0VHBwJJT/Ric55tYdTbVDL
qNJ/sqJAP4Oq4gqLeWMbfHJss9/UNdTkb/TGw9PvEfrMvHWwIODq4vTMlCGeLN0vKo1qMmK2Y0r9
M94wfhdPfxXaAFlCMnmqEsugmVYJlnTRk7pcwfyOYlxDj6tq/MzcEhLZluyVzQ/63Yp8ljHppoZj
BOcHcNgHwa9IPMU1nKR8jHG16mWUY+DvSMo+bgLF48W19T41nTybB9VT5owSe51fV6sNkaL8iuSQ
74BBg+dY+cKrNibfEb5q3vIDWL2as8kDk1Yx8VRKxQZWuFqoHLLpxJWldxwE7L3Ms+NtqwQdSDl9
mW1ce0RmQpphD2QRIGusLp9EHhcOz5kEqUkE76hJHyKYpmptq1KGX1YYfXAKzVC/DleBGtTMxKVn
41yAvR7z8V0hKiAbMMUzYOBwH/XoJMG0ItEd+CleLxIXmVfFtDJswiovgb+Tqd96ZGet73KCMr/a
zgFJrRDm7OE55kJYErQSYNZB+2iqiucfgAG4o1jzlfNHWVrN74nZDOLnOiCHMcDKi3rTtH6R6f9/
8/MjP/BJBt3Goe350XH6cAXI1vsYPrY7MJ9SD40FchTxnQD/ixmQZwix+vldwXyDU3qe3YehXvqR
K6KzGbnsc+SDmW4o4hFZgW9DNh68S6d3CK1nh/4KMufLgtqGGyofajBPGAPcRheQb015mewafLGR
ugqeMEWDdOYsHscTOCldACocZFDUPyHWwX7G5D9S89bHDPNWmOqX473ilkwX4GVPb5pa4u5X05hz
xP22ZfRiJo/ta77hSmaqQfIrk419lPi1PzD4igthaD9A0/q4sVDZi6k/56o5K6ReoKQc4CRdAcCC
K+lToRl8Pcqz2D78kmq/FeDYgR/NNwiWXwHK6Pm9pLZNz4sVg0HfLddu4FgOcQ8h+vlMqRa+lpre
YSM8NBEq5tl1XeEfhXlWYBDh23tYxyLUU8pVnUBVGiEflKQa7E38sSq2smzsEkI3nFf0lsjFhx7q
pckxGRaE+Za8Q8dz5to/I6RPy0m2kHXjz5RtgCaiyVVzS2vrFxmDWzfO303HuYZkck2ZADb9wXL5
8Q7CYrhauryMpDca8fvZ6a8U/B9GBghIRmleQSdVJ6mQlKfa0v2LN6KwFJdqN/AOU9rkYoZEgx2R
Rc9MoeBYa2SnmqpB5/Ph2Zz5VW7Clk8lfIHqs+sOZlLHVFQ9H2zddNsncRZW3U+BkgqOpFjW5tz9
SjAGi4xnhgzS2jltBOES2QQ38caJhoZq/vz9XVKUEoIh7z5eHfC1bg2DBo4MJKFBtRsv1B7Os/sr
WGFxIAof0ZYDEG2KUwVYAukCpDlvgePaxIRvDJd8H1C4hNhpXjtrcllBln9rXLz0tSYdzGiw+jXk
kRViAGSMOVN2hHGxbSje/ljroP3lJdZV6qMqP7sVszs5rw/iPB0Gvst3mSRm833ahdNkspbYphPq
aqIyI/em/S9z2ozfjCpXVCv2Tnpi+s2w9nO7y4CqzzcmsPF86+i7i+aTHKuWLuUtiQ5m0akE7D1e
jNs1+pHETUM401WbH+DTYI/15OhpJo8mLnIBRLp0GHhu56VwYCjc3GNSp0/k2nJzdBBEk4ABht58
sXlvgLD296lDBzLDVYGTswkeTRqIl4+ZmBLLa2gRBtTXv7Qt0raBAg0IEwlHZMt1MKFK9muh6a9c
Y2MHvYmAEDugHvMkKKP4+Axc61eoJMsHOEJV06CcoItFxI9aXXPgbsY+MXgZWwmD/9dAGsn+HnEl
MQV9MZS13BKwEgSJ5Nc4UYcQ+0cYUQBmZt9P2hdAPv2TE7ao/6QDaxG+x4w+IQ+n8Cw6mZ/nFUtc
7EJ+0BcqtsToXMEinw5taeS2hDHOtiKfONyHHP6I4zj0r/cSODfp2dKMfgrT2g9MEgn7CmR3AyFF
RaQ97hg1eUmeDOvcgYZG0fhZpC2LK7ygMvP1XFTDsiO7RWNpm3VQ617SU/II9f1LIUrindTyQa9K
d6yRAIZy8C2tVJPXTAflkyfnIj8q3Ms0GUgbuKg2HtoDl2HmNl//5rtpx9f2Q/Im2SJexYBkxe7M
wh2DgpGOaW+zUr8uqrjEBf4ZeM26LVMAft8SQ5Osn4L/b16Nn6f4BgVkZzLZ+Y3cmhFB2Ywn+Xgl
RMJ1GYNpvWR/kev8tQ8d2WzmXw/LgDbZUeOiqESrKzVKtqjGwjjU30dfO2B5BB7h8bNS8F8t/dOy
yNAh7W3N1eka6p8VW5bfLtVnq49s+GUA8gvy+LDd9cz2nuB2NEqV3sYKn3R9isTen7rFk0kAwj0H
dRz0VFo9g/RyolOem3uJoT9Nim/N2PW2s1pUrarZI4DjMCja60rq4/Kc+9vYX+BIV079yJ//4sQE
c+aOiFqkPecOhP7e25MyKGFSHuKqmmqWIUPV6qvWlZWpV7mr49ptBF4eY8Lo8pYCUmfGFEznN1sh
S4xRh3zydSRhiXCA4Jv5kI1v4wLY0+weWVRMtv9TWZEj96w0JPfQD64tbgR697SXpwsDg+044MGM
j8Udcjf6DccOsR9hHKLA0YHfdymkmCX01SJZUOZtzTQsegWf0UUPMhsxQVAlZo8dtFWxlcnt04F8
aNc4O+KcIBm/H03990L88wJNDOx9blNfyWmCPzcpeW6efiTIe5MDyaQ0nsl2ZMVJwg/4Eqgiek3W
SqzkKxmVetIydVh8oSsInpjY3Aibl9yBpEkHk7isaw/LlwSQ2/cmLTyBt/4gfkF4kX3FU1HGoLxG
SWa8/E9/6KSZk7kFgXpNnzaIDpFd1otoc82xOanR4VMehk9HPGbEayp8W2BRFq1RPR7vjo529k5+
PYas0eSPjG4LeVOi6A4URGxSib4FZGhrNHl2P68bMLH2tIzKWfwG4yYIjQBJWLmdo4fO/o7qsPi7
lBxyXZ6k6Vi9mBLg+NP3/o15NzVZKvV7XL/LoVrL5NPCpunRfzU7lqO+CQE0xc3+6d75EmHdImvV
tj7hvPn/5v0p9/bnOdh4llJEjCdS9tToB45BKoaQk70fMj2/vsDjzD2gOcIfZX7d91coaufgADe6
vy87WcRXvEtCbuu30smUaN5XXuSS1nA1uOWT1TcagPwwB52yiGJGS3uA6tSWdlTp3aJRMK+2sqj4
4IHtFRhYTK8lLi+p8W+/sAvrVLi/PWa1LLhtfP/9TugOFfLSDDKi0pqKSnnzuGACCgELsoiuyZD7
TyYmb7RmVIxngySynL+NUn46D9U4jEoWza/NYd0fP5Bu9MlCQpiBpC0lguZmZO7GvhU+6GP0Iaap
vaa6ymxcz7sWh1mJ9rp4qZr93YhACVvFK8tdhVD4rQnMUFrX2AYkWAY+gLwsdYTI0QcL5wrqxiXR
oLpb38qs0q74PEicCLS2Sqd+YIlo8IwOHurIwQgTZO0v6AkXWbfK/UjKWJv/ylbFTj9hDDGp7BZ2
/CZwzd4Avf83HvqJsbRgOSTtJ8whyP8lHd9tT5Q+BmE+7t/Sc7SE2z+iYkuSUjg//QtXn5C1iVaH
iyEhoVdr0jeZ0xox2B5UrON3fDjcl1XKQv8RA+s3t8H1tHej5elIeOInhHgXnGS+98stAVJl55J3
OnHWO/r/i3P6F5Uk4bkGfs06JF+Ej04E7r9LfLMv8OurGwwZp/3eN6ly54Fua7Bv9mTPchObMnQK
Cz+3niu6h0qeSjlW5GPGrTA6mONTw9DYTgY/Cip+OU8wzG1ZeUjdV+SwOn3kw9nxT2736PiICNM7
cp5AEFatxlZbWPMzKAlzAQUKGOg9xplLDd/v+Gcpy7jVPMehu+t9lfjFbXGY3XxZ+QgVIz/T5Fav
/6nk+CjvN0o9vgd/0SISuq8gw7o/nwdt69B/lXyNdffBFgbNb+ewLMtOoqu7RnLv88vV3lkfcjGU
n/+dlRK29ScGcIyaai3tyr31sTcTtOwv9R/c1Z+84Vwv5HOH3PYFOBznZBf7dfx0oUHfOQaOyVCk
PL7wj5Qz5fJC36+eLVaOxGx78sAFrS/D5PP9awn9DzvEyP6GIg31ja1ZcFzsaOanJbYlPe6IaPIR
4gaokVy7eq0n+wo6r0vYP/ySt11U0clTSdvGqtH33DczeE20FZFXxBC3lN1RMA9PJOxI9IUGWxQ7
k6pJx7jvfUQaDDq05Nj4IPnVY2EYIQT84gSqp0/8CfMuKgctk2fh37JI+bkiiaQ/GW6WE7CyZRHi
+gR0dv8PGVVMF0Uw9d7DtupSOO5IQ1YGmtwSGFOlag4+ut3/wdGrPA3ONlgVdE3mbV70l2B1BEzA
LVzsLvZX/qUUHR3sfMGV+/uhvezY1ez5GK1s7WKY9P4gM6PlSXpaLwDAXnkgjgkstML7UhBDxct5
C6xdz+GtV93sdLbUDUkKYrVFmFBweC10M1SKOiLbBGDM+iQ2k/A2VzPTfyUdXxVUnm8x7mHRfXm/
oI2te4y4rqIC1Vzp2FJhdixdJw1aZY0oL7d78fw9zVEy3S0JiR11z9BGIOxy5TSORlp6ujhZTKai
hWV7GRmDU34k1IWLMvxgLQsW68BfFk/mGL9CbodSsYptjvmH2urL77eQput8SNyao7JpysmkF+88
OyLxxOnN8BNIsQdaaNplCxGbQfGn9OL3Igq0jN5Rp8zOh/CyY15ZApPIZaRD7ox/dZ3EHWip/2EO
6NCFEdXP/NvA9kdJxA12s77oP0gp4zCybbhI6QqzhPWjPMJ8Gdl8caadBP8r1vHYvRbPjm6KbO6H
WdJtdEZezSso5E/E1WjOwQ5hC3PBm0Hb3XIVTgb6ZL2i+Ab48HRzxX09yu19p898sfhsaolYkXY2
M5a00XxX/0M/Y2G+PZiNDhXst2GxVuGon/EFae9oiA1NZL9VWBAEudtoTfVT1pj+B3mJYz8t2mnK
neqBokhPDxd3KFb6DrNf/Qwn9nPVgWVjesZLTw/ESrN6qZNzIseVjQVsLrhwR/ArU376KY2zqOCN
Cjd1OzTNACKxm09s8RU2Frc22iJDYD+YPmTedf8ldhyNWE8VqHo/DEc5sXkEUG3SK0XhSjPWRKI3
TJb23AHaB3sJu42ebvvO6v0ZdE2tkSizyy5LUPyY7RbBwysnk7icqpJHg8zUhIxydfUiO1aXJCiI
j/Vz6U/WUhbqT977HAHcjZeT52NfYXYFtke97cYGnv+WjXZR8Vp9WhzoTB7Aeah4ANUGhaF9PXse
l+TflQONMwXrnq+0MoVe1ux5FhFT13JFwaiqHfRoCnHNIFZiX6+KjewCbpDug+6018QEGEpXs9Ec
YsyT8RJ7dl+li2UdF7E3cxaxc/UgEyVfxEng67ZHNnpjpPUQpcaZ+7rp+QpirA+MGWY9sP08pKwO
BvEt8/EhGYNeLiQyU/YxHA/f+6IMXciEN3dVziTur2/SC3LnDVuyit+ApAHfIbfO8p6xw+jwWLw6
5S48o/RT3QulW0VqKKYsGc/vlqBAKaw85WNFaK4Nuny+69iGmsVWz+uVkooEavr3QNtjhqDKxOXI
x/Ej8M5dor3H84OtVth2QlYPJQYQTkH1buL+zexoDFvbkkK9m8bnSS3S092fON5dxYv4YTOK4MAm
Xq0u9lsq0ODqF/5ZR5hk5mCndL6bVB4hykVoX3zGcHgIdJY8VX3k2VjFts1VtG3+/msrQoJQJ/Z7
AeaRLuEZWmlbv3YMmhiHhPNI21GgC+nMI7QzRRfXEapE6sw8DSDq1MRw4RgMdIuNBeZFCctZwq5A
TaLOIs00+RW/ZN7qnxgFYCA6gthAOqo/fgKDnI+INp5YNeuFLEf8OZ7iFcCIiDrI2uJEEs/4U7Q8
b24ut5LywRPBFiV0/P0QE8+Dsm+sib9hzdZWl0XcPczDJa81qaDFY4z76xkBEORJ7EztpQD8i0Ti
0wxSRjJ73d23q/1qIfhND7XzNFHwt41iWTPyGbr+g8qrEQOIVmNCYtcFjwZ0R/EeglIICd/lPHkv
JXJylksmfyxmwr0rXE5V1dIpsaAboQsil7kDAZgvnXHsvD6u54UnTsVzWWtX8q04bVCGNNHuPOLZ
sZ5KBxL7e1fDYIw89O7REtf6FUsk8llA24848AWAbMTS48cESKrc2m/p8hcwDj/h3249QPd3AzHZ
Au3Q/Poh7FPjbqCAVuySpRt8yvYipJhlRWCit4QUDqlJh9pql+Sj+cfchNVWlw5gA9fmV99Z1dV3
YmiYnJGJ/vWmw2y/2IYY/mjfY1w76/qMbT9o7WTurP0D+PQ7HfpkUssz/RPrvujmAGtKnAz7ZTOf
iJu5a3UYAe7a+i2MlX2gYWvlFsNsHl0Y4+s7GqhHD15V6bYARPsumC/7cw9WDphqBTTTx/zwQWZD
z4ZnBsl8Nl0kWrpMgu7UORzah+zI95/tFjX49CJMs6JnzfR7xrW9Ld4lb08C48Dwsf/EexQoxZr0
ELSP0CG/F6P+sRf3cvivzPatJ3LwW1zLGm4z/hKZx81SoIYcAP4oG1mX5URHLm+T91AtV+zwWB3a
CnQKrPkhXvfYtfoffu8TR/v20Vy+xApyzjOHOm0VQFyjoVnvn+OhMVS5z7nsMbIHa9DiST4E6WUr
kT+ylouaVysawT/myQBgdlSSpVi+EuDQWl8WjhzOp/NS6kameLgUNFCS63227REtXcam4FQEfQyS
1v5EWIGu2xvxu0DRLn6nuMIFVzfw5qTO2h8T21hR9RnrYSGsh0E4XHcr1ELNi8vtKx+fojnSC6Ys
6eYysM4Bb5gxkrO9MmTepUcqceq2W9tviFEwLbAoP3jK5B1UKI4loABw+txO23Y0leKZogd+AKte
gF4Up7+sx0rW0R0A9RcB0uiRFvLnfxemoMMEzLOTEJOmbXfBxA0W8CQkP4zmZwbOdqd+wM2pdsv5
hOdCx92YIXh+DdSnxjE8EKgybYvnDTZ8Vy912LyaN6cXrH2tAqUW6j4/sFpaAB3meDvIo/0BdBAk
BMZat0qPA+De9DjtWH4CPZs/Ab/l2iZ0SKszAjMNbX90/Rw03qGJXdjo9iQKKYaUHOI0U5r6pMlp
ex2JSca7MDE0zxxWxnDEabd1wdFIWN/VTUp1ZDiOPEcY6lnvQjcDpTux/QOgoBBT7yl2XQ19nmcS
U8R/I5Mxm3RL2Ai0UopRJCNWuO7oZmYY1EV8C5d0Ef7KvfIKDgcc9n+VG4yUT7MfLHC8EzWEGGCi
XLJP2MKNatlzf0QAmMg0EbyFiq7Z9JZeFpn8+CKyyjkrZP+IqO2+UyXGut3f8QDW+yGArORKrz+N
SdQfLyDBhVgBCd0xF+m5c5gn2KNpT51S07h5C4k94npCsXGgHIPyZYpLBtGaI9MeMYUVUN6xb6wX
j6Q0sjJ40YOanwDngnEl/L42CmZn8r4Y4x+ckjqLdcvrxDV2WTSAKiKkrl3KNC7IkoFKkkz2lCCi
ptig7RO0axu1qIAlX7I/7vFXshq/sZa9iFVWb8elI5B4RRr6GesbR4aSqfzbPwDNgRUXNC6FLRJH
vCIFyOBUoLm0VbPeQthD/DX3BydGUrv21UaOrd3R1Rp50NBP00VhNruv8NJIolbtzm8bxOv2ftWp
39WLef6VqknUJ9OmWppQn2UgAD3ZE4igrwS1fnpYnJNKDj6U7gi0eZlsFikMD6sjmmwXN414MnM2
/pe6BYDGaZ5sQPtUbVDr/7N3/xBbOiT1sgzQUI9xBS8Jo8SMCgnsRVzf6A2z4qwIT+WUEbgyGhcX
cueT55TVfQ4627J9xNav3vSDo3NAPlDyT5mPaNTXQ4hYlLDkQ/dAMwXn18iLNdov4eMaT2Qb/Qxr
1XBXWO6Os+b8A+bC+4r800UGkaMSzlgNBbnX6lerKQNrEMi66Nqa4LK7FqllPT4FmSyOXtWJfZMT
BJDmUoRvllE74PjE4FVdpf0MA8v2CE4lZeV3CbwjN02aY4hCTlWd3wlAmC1/NixQbds9+qmyCjSX
hjZDcqNafJdEDqt6gBvVT0n0utwWGuzuZDi8OhsUvPgb0WG/1CBtHVxX8cQ61OsshVo4qTCPZnpe
kCO8utTeWE6kYxyb7S2u/Zr0pHKgSvf1DKeaYc5fXPwdqFcsCS0R7CSvSzekO4g88PGy/W3Elohp
G0YhJv8/KeoY/axAtblX8pBE+h3z6Nxxx6oII7qkg0huikAzfKjt3kUQCae5R0GMBi/5rQWZfhoA
VIAZxNljPnV9+0FJ4uMHCkNdWwmU2hADBaoG1bjnLNNr6NSqn9XQgcdue0NeWasewoj1kxXUG5uY
NMNumZrp+oroIWS/87X5jqjKVuTxbEY71GMX1rWo+4h6toZ3wpXCgiCAGNhCE2FPtMYqzCqQ0ohk
BRb9qD3j6L/ar23j8kNEw03qQ8WHSbVUajSKMiTk7hZkxaLtezV/JcuXcYbZiLmCXRKjH7Bsv4S4
wA2X1rJ81+PhiJlPrMYTVvl/KFizis9xCAUOXUNlBWla1iqDpFn4XFIjdmWFCVJj1VhJkxHzOnBG
gKC7ImRdQZWTE67NZQEhErd8R6Qp2JDrndOJagCZrPaIEQ9lkWGEAUI5Mu6RezBNMW7yubuFwz4Y
nUT82f+Ulw4tDL+Bgj1W36ueN9SWXQqJadbVbclD1hqUFPdTCbrI07OsU0HjMtuBjiP759o+Sd95
kquHfaSlaHJmJqZ+fVxMrKE5oQu/hAfjl8DPElNnIlpTWVulOtjtrxzKE38Er4qOy9rFD1LCWfb7
EpTI/J1vHLKNgDmpBpY5Gs+1zmKZo95xENoQCnVrpZpP60uCc9HX5uZmeIZP0XWNN7b0TLKWFP8W
gWk27J46J4nR6ggVDG8trYQjYMjXxxJBT1rtuijBeYNYaNqHNuVLhc1zZ+sfYOBKFDK4QOvszLkA
JNm/DwKItyRPW3a1trC/EnzxVpacxb0XDU03vMS1Xb4HQNNKSX4pWTBEfua6+w9smq2hexDVuarF
khqoGQ+nkQXtdpDvOJXJ18ZLuKbb1eTcciTJJOcaY1GUK0lkmHY4EpR1Gz+TD21bsnCLqYc0Mbse
oVNzd4hO45JYYZ5CSpHGS1NF1zwd03mNIhve8w1xHOTUJ1eXbgQAHiJve93o2LNa8OAEsa9FXax/
OrwrT5rn3i+frXPeFJjVXxXh6aJ/bJesWwMUbiRkksozl+D48sOnh+0m0cb5giPOICdSi7yl1TBX
SaBcf8kDuu8jecpLYOk0ou/sN4uxzprXYaFaJB/mF/7mCJIEoaBWCb/dOB9vErhmzVU6akaBzGxA
cHgPoDmpL5WGwTVtpYh6emj6SLZKMWHw44IC72WorRkvwpuwJo3g6dCXhtDVuH225cIn+xxGwykQ
or8HTkjJjK6/KVRqGEd0BatnswgbicyLlcEOMdL4n9UqDGlatt9DJgSGusANVd0aK+i+ABwH+6h2
sTsOWCloyy8322qmaEFeof5iJDXoTGKRC2QGbvftwbjjFPag9Wso3FhpdmTCub4HPt0TBvRu84Hc
Pgnd4SZ3Hi6JJhAM5Z2wImIRcImXiv2Js/d8sR4S3l2hXv1/Z6o1pEW38a9m7XV208sPXJ869bRO
ENU2hm5FgNDEpm3sRWpz9ZO5QaVgyNQcxodjkXdvbl0WwBEVKCi/VfzLi9W8XGYnNEGNxgQPftN1
/T+NRKMXGXYqHv67medC43ggiMbAR95Ug16sziF/Bo99VpSC3J9y80zt6I3kNZgFJHu+ulAem68M
Ofn3466bRPMVz7PHryHNKIel4UUQuYOyMjP3TcGiv/1Yj4B0QOI4Xd0AO0YIsDs80uzES3Sz9uuW
fceNnmPNFIRdYrPIYy5wKVW3klqJyeLhmN4Sij39suPoargMwG9MLXm16RAEYSsUtJVURKizcR8v
mLTMxSsry4k3M2Pxo9aCkUc7wfKVKvtl/VAUiRqsPd1f7qLY91cqDgl+922BbbmWH4IV+/wdxFTs
dGRRoVijBAxdD+qm6gRy8lD0B4+dVyq1ZQNFjI4ViZEchDaL1D+yrao7tWBkKqoeZKAmxzKD9mIb
/MmPxYrX4dpIosOoSlFaWqx69/1wqfCPFHchAUMC3isym4U7s32SQet4mzq/Dis5Xr6kZdDB0pyj
29R/QxQzShGF1YX7kllkaVhIUSs1Kk2AwC3e/etI/dZxwWt63//b8uvDH6zoxex4ldkbu+4lN0F6
m5SGGZiOB38ngUvzwnRWTt6NXlAWs9V9u3VT8Zm03DNPi1hfZNYYOEt6lKww6JF2p3XIn+M0SBLG
Rw8knvXbpsQCFm0F7vNkyo1dnzq7PJqYmfadjGw55AgT9n61G2YE+vGQVgKAW0uHlnujymm+Cdwq
R7AEAbU0tLjmvOv3s/E9hwMCjTW5WPmFTHU2UAcjRaS2U21GOaYkkWR86mk16DkzGxBBis938UiJ
48OpS/ik4n+t6XAgcnpCnZWRIuvsueBecXKiFX+z5Q2xsYdi1ktDoZqal4EQnAuSrvjjpE72R1jW
BRqR2L6MzGL45xKQqu2mb83iYv8q5jbuSr1pR71H+n9PKVXxui9PcZA/kguNvZ9jz9aC4WQlOngU
Jt+iBud5DcB7xvL+CpRcP8jzRVj/RMe3iOx//x5E7wKq9rltfd1Mr1foKyKDZDHk9iATOq+jGaVz
8b4iP3ryxfgcD+tIc0dEwhSLsgk/DwXwrDSyKTCp8lijtGpDjTTMzMvF6H+nvEuhwUw953g4kYuB
HejREb8JM3sqlsj1tSCt47NueOr/H06wVuDNajndjy0XGHaqQri589NeInJESTjgmmWwawM5+ICH
3XPSrLOLpHZaT2BBszmQpIu2tTyUCTJKGPr99u+4ijXqJSYAKcCR1DCPYId2JCISI7YTYJy/zw/s
COJHWzIkyU3SMTepqKMbFvkjuOB7GGJHdGIu1UCOgAdDuiRRtc1R6fWDRuVDNBtn1Cem5F3u6ZXV
RlnuDMuUCXlDtcrBx2P/yi/Xkzj7KstCuumg0hIPHWqPIa1PsEb2WYwlX45xZOE9wRhkXo9JpKvP
1XP5L8q0YBqkFkeKOCJwl+lQFXiv58aLR8Vxy/YUb9gq0aLkOhlUAP9U+v1CiP4SyewC0vkwbuz+
G1vlE+UfU4aZHIvYTF7gzyiz/q9m4beanvhBdDYWAry5wYZCvjT3DlqkNKYXGEAH/g/HUrqJnLFQ
XmGpyHcbsCIfBtcJyxSRRtkM26fhXICajpvAn+XbOB/TBDmdJRF0UiBjl8C3cQvhNz3WjwNOkyvp
dsSwQ6H9J6lh3yE8ukreH0CttT1OuGOXc6PMTWNNOwdWrAyLeqIhoC3QHVRybqIzbtfhL/FNQ+z6
IHEqX9tj2QB3Mxh0g0lDloh40esj7F4MuUzwn6XW1sxjVTJHlqhy+cbv7mK01GMx6c/LC0A5gH9r
wwi2LiDRgPhhbLlZxYK0cfegrgucF3OKTW6aButaw6yrSUDHGOB1M30Dv24nlp4cDE80gTg9KpYV
D5SeE15Iwo2GtS/EWmt9z+8BMY5JBCzNTjl/Zarxpnimmt6V7pGZtkr/K1cOQkPCZ2nRKyGbTvCe
2YiE1xSXNIO3JJCDqzntws6fPim6l8g/LZqP+UzF9SXndqrC4O79B6lQtJCw74B6zdiJm3+yykGs
Qg2/nUdLxTqDmFkw28/J4zBTOT9kiJ8/NEqZAxN9Xo4F8kUQCIu9C+8PKFBjvugDiHJ+Rn25+WJ7
WDrv7CCY/Pb7zNnt93/N/0yhs17Oy00961gfFKu5lRaGzXWXgXey8wlSn5KK/u80uoffkyG4uMBF
LsBhLIarWlwZhhYgBE8n6Gz4N8SydL4Ja4gYPv15a3pGBgf57V3xZi7xCFLlPeTmmGLpqAKvdyzs
rA4Jip3rivsIwpPX6xn9w7FsA2Udh0uMHBa1XjKPcEBXDAk8rMf1iV+ObhbTY42wQvioA6nlTuOf
Z+gHgi42rNDSfIWvhFKl7qO5EVJmkV/6d6Phqxl8d5wlZrpDLgqRurxC0EEIbxSMHhYeIj/qUV2b
G3MIpsrGinByq+WIFAxaTGGZjNg3umYL4lADMaoYbsiIXu5eH6VkG5oN/99vNsGMH1fnNWTRbm5h
txF1SQXk/EH2UQFLkEROGppTNnpjant9bw3yPxoWQkRpYBBFjmXmb/8uZvDYO8RPCZhlS9BqCJgg
LjERN7H8AolJj4U03zRLyTa8hJOcmTUH6QGzqubYnOpiRrgDLDDXBVXP1Doogt/hjco4zRopzUDl
nQdIBZoCDzk0JjWcakT8ylQuPtES/5ml9gRz8Y1OBK6fXsgwrM5d5zsdUI89YRDWx+MOYuDooeaQ
/HiBNqeOIx+ni7wUtl6XiVl3e1p8JAqT7rt859W6jr+Bdh+ygRPoyTvuH5X6cizWYTOoMalmNkYt
32LdnUv2WlRhoVnROej7ykubR7pYLVA31qoFO0Oy28DUUqdPyxx4uHH/LEW07pgYFx5doDlDVknt
8DR5BGvRqaVk9bhWHZtyruL0nbrN7PZyaiwhdPev73ndBrQ3I/6e1swGLsDXfJ1aYynVdjEWnra/
b6X+R8/UUjBwg1X55/quRmBnnS/BrvMVngj79OkPmOKF4eFZIKLOCHzFt7sTzapecdJz9eBHfMal
laJmGenevPfyHoWr3lbHhUHPhujmWGy1lzuIoJV5zcXhLFD9ZWc5+NFukCZlyl4QLVats/3LJxgw
kM/Y4+Lncmln/qliRBFy9AxmSh3pAUs8gTkn2l2HyZ8IwobXevP6QrOglyRsAxP05kcE53BUj45X
iRxE+XMFk12/MnZqxctmMeJwMy0A1jGvXklWyEL7G6OBv6ux4ZjOsOKteGB90dPKWVCZbjeRNkqZ
x7wq4P8VI+Hr2dbmJAYV6zBwnRx1JsmKvmk5W9vbCNWAPbvAOlP3EVCgxaco2YekW7/A4uGAhIW+
pn9RGWTzsltR+ZaKtjgQOXZiuB3LnwF2CzJa3FGnmjEBoy0JaiDjzJf3lJjZrIQbJiLGJ1LDutBM
XHuXAobM+ju20YtOX8lAHo+Emv6cIZlZCXQ8o6wEFlmjgtCnU03LoYAtoCV+N3GDXdQgvS0EFruB
WIkyNfGrn83Znsu3Hu6GWhFFla4A4b3tF6mmrn1vpJKLQuaH/VKd/EQRXodCVe5mBi5Z4ONnMV47
qiHN/ThiTCBVjiavGlTSDGSVzGIJpg1VjItHUsWYSZoaaSzRHZedH2gv3esVXe0Bl3YNyEkb1oRK
yiw85nXESqu2nBWnElzyV072XUhaS66UKNaSHwRVdOhtK+kwmvtWXMgiBpqR+Tw38TQts1N9rmQn
mlEFoQYYh+OkEWjvUDJUGYAeWSbX0sM26GngN8NdFzdy3yQWzqSdl0lP61bn1jclr6OAJrwf5Ulm
rXQyDsObSAElsK3rZAkv60uikR+Gnu2jAzuCjS1JI/DJYCLYzEbhWbc9aqFyMXVIzcjg6XhnT4ar
b1GLUtxGHuuED/zQbfZGv0SUIbriS7Y517Ypb6AmbnDKo6nbgApIJcqbY5Qz54EWUffd0qPSQDNj
dDlvfbEwh+t83yQ845o+Pkj9hHZIvS8COFvsOyPkl3QlAfoL3Z7exrAUo0paVKQL8tbPysB965zX
DZBr0JVLhL3os/Nwri70dj3FMtM2WKM7h1ltQRKYLSRdctYytaaiZnNoU21cFG/X4+qqq2+b5/Ul
Ku9AGPQ13OqhWtJGmVgMSyPdiPO4s04IShd0TuNlutu04fk+30b+i9nNRvpLNVDBb74T2jH/Pq7N
ri1rP0wIq4ybtWwbXBnWwk14a4Vsj4WqrWqIVAjenBOTADbISt1s1qqMkFEtjz3aOgacqmNxV++N
2GP694JjSYAp23lRHK34tr/LDZRv/KGJcaSGIekkVimFkRkxsHYnc0M8wsII6wjnEDZngXadafh2
rjrExQBOQllzWXtPP8e9YVhQrCOysyQjelE4moTRCvRgPRqNZv5S5cbLQ5nMjIpkaohp95rXmdBY
wkqVOkAJA5H8xB1G/vgyZKQqeFpoKpBCGagJjCPSD2d1zOk/h2Iwen4MRXcBWIef1ciiNS0PaNpE
+g1IKa0nW4x6WNRjg8q7OtCnwuV0PnPPbZLlxcuZiLeh65kwhXX7VdWlQSlhohzKIVGqJ6Sa/bN9
x9hhDMXMbKbZvUWq9eyDaE6BzmONUScYwBB1f+GcPr1BoxTNf9sXJJHU+tMFRleNoPO5BAlLcQw4
e+Z2QpEOIRehADBJ2qcusq5r1i9KxQN7Hkyc5FeGZp90LIg9Ni9Un+EYXqNdR34lIudIM2CaFvPr
1G6Ldy0F6W+Q5cFiu1C05ZzfS/WKZO0x5Fp3JnWqfC38vUcrlbN1zCzh5eHtYGDtssqauSmE8QiV
QcP1sU5BtDTCdaEF26Bovt4G0ygKVw63S3WmeFl/Rq1waQKpzaZ2TSUH9f7UHMy1SS8Jabf9BSru
Qig0nE6XDybgnOoabnrdRFLOEe4I6dJg8uPTjpPuQ4qzdCvAq+K1GXmY0kU8QiF+YxzRvX5LUW7V
WHwxucdnXWFkq6Q3ccARNSu0gKX/TrQVKlEAtsNWfrcGKd6dcfVtc0LL+2aZ0xsvqzZ+LMubsLFO
8S5K1g9VQK+AvKaIu4nkzOq8c1O38lPtxcUxuL3gm1Mi9iOSfUGT2WWGY4itppaoLWCvtpgfDH2b
Pga8bhv9mI3Xt/Z/MQvmcJQDH0IHsViNiiGsNKtiEQmFCJjTRA+OG7jUtM7ilBvF3G5DKGOp0JWK
Yke7sbtw6XvtSy1qTyLk3LnEAXoesr/z/w5wF9QfbEzEUZIfSG9UnNwrdGHOuGehQQLve6noqyS1
ADBgMeDEuryrEwhrVR5UPRUAvhMl6G+qWm194lIOuvfUhJrMMTqc8NR4kM5QStgLowpm/3EVxDf0
UhUYG5GgmBTJi9NCa+gMN+fKJpbuODVfEDpGjcyvxWXpVzo7VkvyOXP68wgphn6Sok1O19eDYADy
JbK1qPEqP5pkzznBluB1bJrDkuA7nDlq6AEF5NSv4d3cq4p1mZgy/FvxswF98xiRFSESzz1YznvO
4va5Q/gBC4lbzt1kizsAmdUlNOXg7ckDMHxekvVg+qI+6tKT9oO5UAZREnm1YN2TB9Vlezc8y0iV
dSkuvmCjKnTd1dQyeCfozBboLx9vmx45d/l1kF+riAb8YeU3ZeRp/s8MoxsImJjAtnG4hZqbCJmT
A2W5tX9ce3t1uUHAurQUrj2USwjYFcnPuI3gAc/1atRjG0lilQiU40JUtTO1E7pQ+kiV670jZFeS
+NuUXdQTNggi1x0PV/bJfMQjwRR+B7KO2oeWztGvZRXz7EX+4e/7LZTPDe3zqvj7iAtNLDiTKgCj
EfojuRrTFMSNWdmvEyRdUSl9tAsq7NNisT9YM15/iPr1/9r8R60S1laiY958uGNu8I2iASEA37ik
ehxRI90gNZ8zK2DeDuaPVMV/Ah/7KwmDRtxA+bdIxHlW6eDarW3hEma51f5WisyfyDbJQ+QPPY6e
0tBhcLHmhGfUSGBCWsgjj/Mkd7FVuKEjlb4MBcl3LFyMrvcl0ThhBuEQWzC0F0fMh0Tajhb2zzwl
TJ8WEpPuNxYQiRuUEEcBeT0aKH02biHqCn02di3d3E3C0m/Cfftm+5pX99G7vO+SRgi7zBZD4XjE
mc3pTDo8EcxBGiAa8Ib5CJlFvjEWVOZjsrek5RnPmTAF4g46Bcz/BMNHsqL9rGEKdg/90tzWA9tU
/gRFscfj7DlvrDoXek3ELrcbIkGEuPMpToPBF23YzWjRk0s64SFV0vMySpouLdQdPItvJl6rByTJ
O4ZbEvsDr+6AKVTrK56XT4ukVzbHadJTRR/Vy5qKN9+eUzqebqts7vT+2aIQ4zQ4PFKg6Suu7PMY
39cuasISSCIdOyabP9BS9Cf6nP7dRF1TFI1M8+tNyQkvyCFKp0t+2Axm2CrKCgra1CzTD06trlqa
lKUmsTL2knp+C0udRnh3UQ6yYxXtpgicRjCQpNZf8wyWyerQb7b/VMDPImobT9YTs6VvQ888/EiO
cT7PRer0/fc6p356FQ38aOWXV7w0goLuCjUf2EerS1luWknVsvGQ5XbF3KDsoPXW6kPgiNFf47oz
jVOip9zMAlmF9DXqkjlJW1lsmgT8QNAeBvV8w4WqmxS04hMSoQkTX7YJJxShlYKBOVN4HH3uR7mF
azWPKyXgIvGK6/d70sUN6a3IH1sB5pwQEikZE9Oc3Xzubvglmjtf9q6lrvHVC08lPS+Z6PBq9sME
BLMn7TyrR93//WPnWNK0vbZe49mjxtUqShpyvDPGOC5UzyrAmph7mdh7XjvTYfSzvbWrkLBLkDAs
hagV0FmCKkGo7Vzg2D+ALBmTwYQXuzUjLakIGMDUGNR9l/qO4wNOtlA4naI0GHHHjLwbN7UGkOWm
zdnpF8UY0YMo6NkhOW9zfMygNlTOSDhdh4xXxKpIp79urp7rJYFQpTpPIbhPpKNBILnw+IJCRoev
hkzi+GY3rlPSMUNScDZiRghbejlfdbaVUwOmdRuEggu0q+qcilDVy+7GrWRTCudF2I16r4iUUTeC
aqmyLAcMO2ZYqt5tPNpFIVMs+oidSHBWmS2lPvoIRfnoMnDagUufRp1ttHKTVJOOetbmODwtV2af
Lt924NtbFUuorNXGFvwfpgI2NOzVmcqj+eKIn5j8y73hEY88JJfGN6zmaoH+nsR5t1ycig7lYuWc
FntarClcpeToY5EelQ7k5g1LwXuIPwSFlDjWKIQ3SVCV1tJyDftL1ZFz14EZ7+/K8BEXE70322K3
RzixzWGVPJ5JfqAmDdty1Ru/2UxOBmHV4NlGKau8HFgLS2EJRUlt51LF2ApgGy1d4HKWl7RJ/LRo
eaSlxEOl/rPUk0JkxItbmBwCpT4YPUUCCIA/uoMK2ECRBa+eR8rhKYU7USW6cHdlFHxJyy7X42aa
Dz95LZp3NWqx5qfMUi6HpERM0zc4Fpx03Vqq2/a8S33TtM1RrD4Z6ZebxP8RAp+KFelwkxP+8Wfb
c0RAPuBbC49OxyssBxR0LYNUvzl/ABq66aqWYYVt5Bm8kcH9nTsDg799Uj9tXg5IMSRdPCYYB0iG
YIEXH4MG6YetegCAUZnT7Ms66TatyzpXAbNz7+MQq2Caslk597r8wnwktuaO+IWM1rJNo6DRpRra
Hjblw8Z5tLhYILDMZt6JPcBvNvCsYSH6CShVA57iRxXWsA+wu5K6KKBODLxZXoMZKDd5mKr97U34
s+9cqhbpFJpBio+iBI58cOUbr4ouZZrsb8z9pGKpJffvx0s9Esi2HB9F7XHmxrPSK/VpbHIN5ySW
V0N6UaXbmZt7gESnY/ejwXBN+YVpGp/0fVnaIzFULBa0w82XnddsnmB4doP77+E+/05lIPyrCk9u
aottS6awW1HBfwYbriUEJyNPHzk/pee2pKrQQ2JSN7Evfez9b/z5jKYTlyGgA1Dy/2jHRaaVCGhs
i8HkmnrdFLDRvW37etgO4dOZlzFQatCZ3DaPMZS2PbUxXmQJsq3WlgJbyBnp5DdkOcds4DC6qgw6
MRs9fv76s/DSlbW8mlNdsaRSe55I9QkTMRp7SF/IxM9jXMrcp6VRlaje2Etn3uo+DIoLM3jM9egt
qv5eoDBagkcTuSuoe+720t1IBVOZJtie19AmQrGzvI++1UMMFoSKGN+/Tj7rwx/D5/6Pnbm3yU6h
FiJ5/AACiPolWg3Q2yBf1r6ChUv8dXSge3awE8sdnNxGa1U2yV21xc5r0ZUklZ0hZ1Gd30FJVpAb
UQLda4wN3vlAqCDxP5BbEsI4nde+BI/PoDrFPanu24IG3pNUIFjt9Y77fhR3bwE6GLzVXtDKq5NF
3jT158QhDNrbn2NknqhNkseih6rL++Z8rmxhq8hvBO5xGzjmVyPfRuo+nxSy/yuzJCOc9K73o4Ck
S2ExM5irZMYIf/KBOJFprDPoVbl6/GGKN9owSSBV6fnYeDLGGiGXvl7tYS5JEYFzz+JD8W8WxcmW
aQX7qRxUii1Uy/d0z+whKNNFGzs/VQ2s6WBgB7QKXXt+8xFf9kYwihjE1C6wqPv5LHVF1OATIGba
S+5ghThZgw9notWzgWL+Kl5cFxFAdiV8vKZJhqlEy4dNTXeBY8iKzqCPzSWVB+/wiPqRAawEYh+j
bry2EVH4TSGLWi3u08uNDwMmasJf1lWKgkrfGLBRHIPaGZmQ+RBQeGk4IomKzqW36dZiCJ5isdiv
1dwC55J5a3g5RgdGPQ+Y7dwRCCeG9HkBpWjdV88qT0KHxqwYKXBFQQvj58V0PzfMHJf5kJKmRnNj
yNIso5k8FB+gv7dJFbEggajH8EZH1uLlJD3pdNuBr3OEELDBZMSAjP8U/EWXAYD+vDQPkvp48DBR
+SZ1pFMgWG/48a1cGKyTC06jidvRGT9jErmxL6oO6EsN3KcSFMQqUMSAI6AroKj1XIP9A0Bv52jZ
20IbWBNk1u5iB/Yr7l3/UuWOILpDAIqcsirIXFAkDbwhjVzCdqBVODGJpfK1k6j3k3uYbK+OrsOz
T8P9yYUTJXgMNM1fp1RZI1hFIw/eRCaz5UgCGPCP0qhsOXeOn7TgUyQNgmMjMuDxsaVaY3OOvgCC
Xbph2OADRO4Z9HHrBbpmFUFvs99aN3mQCTN6A/1HTZbYB6BiSqMT939W2QB7F1gi+W5/p1e4cvLj
BD98N/ihB2xZ2A5/mPeV0J79Zdv5iWHSRtClbIW71IUGMX/15Vw1owXk0TcX3eQDvKy8+oXOXtOF
PajkBHS0vZ98v+qi2W8LwyDIPgRu5Hx52GlCWM5DL/h15idw9yVO/vWU//KsTGyPn5UWIW1chadg
93y9NktuqWHYTc6Lj2xDZh3em15Re+Z3wGckdl0UCZoI/GpRWMnoMKFkzSav1aL7dgLOkjob6vVq
TIWCFD0KNI2yxl8itePYFD7/ArJbvGWM4+v3AU4suGRS7FwPNOFMc2YZhgO/H1vVKJXFS0XalUrV
MPfGvhYZ4m4dbQrOvCM7QfmolIeFu54SunnMjtpQbCER3lwIRKdPU9eO5CtDqT7WCM2Tl5F93KCA
h40Mxvf7pQo7f+/bHRXH5ToyuuFq8+SWZkjlC+ka2YHjzCCwCSedubn0T+Mt5hDJk+wbdfULQZp7
lH3bLb+4DtI9g+q7hR4DNiNI50vsBzyOeTsNZRq3aBi0z4epUekuFw1/O1DpKeZyOEfkL35gYFxU
JMw1x0/jXXrp2jYfzq/avrErPlcG7h8hEchasTpaTNBRStQlY74zyDIkqrXGTuCDFUpCEqdyuThi
4VK3yGxItJsGrdrQ9F14CnCDyY/Cef9exauz04mNzKhsVEjNeLvkVQnNtbBJOCVeMkZHX0NjpKNQ
ZDeVuq63rqTJWWdHajzLPlxLbL70PPifi4g9t6jNQ2qL9PNNX65TEqKCD5BRfnppMXc1ty7rq0HK
x6SxgBfHlOvs91vGBFXrWmhxZHoUyqOWURbhOgJtfGRrb3CSEAeaKE62bim6ZoHshoWadLmG0J08
W4jT+iOxM5t2UHYyY+/q0jGO/jhNfB/QS5gtRdS8hGs23Fq+NIPtCeZhanRHP6AHy20nNYshLjuh
MhO/9iq5bylquo6YbC2Ux1vdyABPomntzIlDQJTnVetRonDNClXY7kb0KXDIpDUGIaZshSAB8hxV
IqQWpSTgDXpanaKcvS+M9gNe97zE21erT3CTDnPog5bEWIdbamOOQW61CrE2VQC2j9T9uLbKmrQZ
b8w1mjDhbqGHzAIVgng+fjPIpUX6okI6knjr6NHBbFzvbYi9LEiRMnFgAnwynd4D9auO2RK+Fi0f
xAtaqizPvRB/G4yToxd5aUrbzQdVmwPuA5lTxHVsHM1qDRppmIt4R39jY7qK6ZYmLrZzPfbexmeS
sr8gBgcSMraZCED+jfjCPhDrOVprS53U+wWBRU1Y3ca//X8VvLxNnHjhO1pyuWwbJefE3oOJS+ZO
UmCfyGkLBoI+P3QKxeV9ro5G5hpCSod0cQznr/FE2PgQmpqvGvf2xWay1NtFHG/BvevxUNbhe0MS
u5Ujni0tmOaleYA77dk7FHDFAEY1LD4FzMolpBVTwv0eitUdBxhfJgBefYRFjHxH3Hcg5mleB7Mz
Clxnv3zZenpPFxTQh5LS9HG920YOON7UHwAc9zkn4WW/4tcPE6I+XzaCDpRNjFOHhCDzov61tk9n
Vn5ehkRkX+PXeFnT6kL37g3VdQS3nM326QoJs9gh4whL8v8fOUJTS9vhkZKo3DPwLl64DEAl+TAK
p7+mJmFEUkZK81qR2Of/e3cKyBtNcaOBJhzEDFlXe6dF18aM31VJyf6MVD3gAxq1slt6lpnJ7wQK
yT86pNORwb8AkPb8dDQlRTNzKXM00BCOKJgD81okAYsgBQWmvURJXsr4bMJMGXx3VZsUh0PqsX0Z
lOP+CXh17dKbVsqqubt8QxNADIffewiJtIZkEiveKDQ7XyMdk9rUMBCNwt6kET/aCWM8pDw+5265
qnBI7CqkMba58IfTNsXm+QwOlaHIvyhlCUd+lCeKen2h9OzQ55NOpL86iMpDtjWFe9E0XfPzvivp
k2mn4i6biAVxikZDEJhjGbB3yA02SRBSEtPU1Rq2OKJ1TXHdWN/5MW3C98nFLByU9onGBBiAvO8w
Twl4YwKZkfOsYuqwRnCOmu+ajl8lktU85sMGLW6zTexeKhr2HT0xOeAw0kQcNRlY0Ia5RruOzZ5P
RKt7PV4DgpjL7jwaLyuGCGkMv447wEPzLWlLoeNGcstPoJwUY5niqB/eJhP4Wc+QZXWImNFI131q
BqFC50ouo7dtlQiSMLChGxeNCvdmwwNouurmuJiJ/DKewElCbTgMxt9+10glujYLIwu6JOVMlK6k
0/YfIs5BYEaysuex7W074xvhej8jKvK0usPeWIPwU5mcRpBg3ymWF24lgCnlYdygOhs8tcEJDNN7
Fr3xcoy/4HnXRLam7+BhJ2A0HuH6/1AbdbnpzbCvVLMvnODw5giR29xQpSlKT1SpsgjxCGGboE88
ciaV4IADpGH8TY9bOw5854TbjYM//iM10uzMBHdwtTf5SztBRZJAny7rjqX4zxjok6zGY6gOuMTW
TfZOMLv7pou4bmTS5XBwE4dYQgl7eTUGSFrWEbAvR9KwVKYboaWDObNFjx3MnwisXsLGUizxymo/
QNKvjVircPW+xR74s9ywpGIvNAEpO2NT4BRxWf/j8flPnBeaNkYC/Y1v18iJwIEbPwvMHnMozAsQ
B4VL3VPpd2hvFrjxbMhQKsg6RoFbjp5JzE3ottwP24nkNo5c1Fun5cY9yK6/YgWUqL4DobJtQxln
+nfXMhSV4K4+egHAiKzmr6dVVk8Opc1bIOzQdVJnE4z7SBBWKTAVVl2tqo8grIbV1Va2SxCYq35C
qCmalpTIuTEpsMVSDZ1KCkBWTiV+XEYionlPs/ZC/z6NNfcDAfbhyyOeZzLRUUpu7hUN4buaMxIV
D1Mt2QyWAlRP1hUrbp94i5JZS5k6RMs4HfCkvKPlYzzngd4FAZ57RXhHJ+2FXsg63/i/rlwnRMJL
SzyUtpQ7bAMDtl1wgKatkYCxr7KHIoR6Po0tl5bewbtOfpbTv4vCuUMmvkf/7aWAGEgoJQ2umX9g
lq0DdPPzVFg0CCTHq5t4qAH9e/w7/eM+7vl8FDpycDUYtmtu+xrz9wD29Sc1CygAe1bnGh5bQdd6
9NUnSNFlhGX4nbeREB3nnAHN7VQwr07pKTmQ0Cbtj3l98BxBkZzOsMbQnRINsz4Ky367ggwZP8PA
d1wWijot8QFSnd8Zi7uCRg1TbFnLQ/Ecxz+lrGPVElkHXIzGcm2T372Bzr1sF2XgoNvJprx7hDLn
mxIUwuqbi2piCBmKrdpXJ81uB36pB0z4e/8FOdb7d4ijmCIlt7ny27Z1pHtharGAaWwAK2zEmmF4
1C8Om3XBFb/XHwJ6kJm7f3xEQKNijS7aCeb2u+FLmcAnv91ZOUYmJq+ZkWIk76aX9ztJIEXA+G82
YgTJwjR5DhV0RfMRDarZOM30laGpc90Bhsa9Wz1j/cK8+Dyqv/67JBF5i318IS9QfzJsw+PpzZNn
dy8ypA5+7ORHZG68G/442iGyKMTyMKeiYjwVpdL/Bfm6O0KTCB3Hy+3z6XoyRKZMJ9gdfSVtfgfb
s7c87ozhxYN90p6p6SzL4pNp6pOAAEKI4iLlpoNKOUjuEiyL8j9sMBCMX86ntOZJdMz7QZhRNJtk
CfbFC26irGYHziVL1rcuhtyxtiKWO5488LWY4UOgl08IQL2M5XR7AtX2XHqvcxL/KCZQU5mJU6Uv
a+urIzmik6grpFlLvT2Yy2Se7VFNW0IqkI31EC3ln6eq55cf/9RByk78TVlkuqDADcLEopcz4AM2
utSrCksjO3YVhK5B/trTgvyz0mgh/yzj2Z4smv9Ao7GlVs/gjsqQE8oqD2Z6doCJpvKCjARaB187
gGYai+pYy6s1gDLTK3OGUonKXNNz2YoCDNAC3e8HNRONxVyA/nS83dGjfO2Nh8UmWGLtsAFb2VJs
MfjccU+AVARHZZN3kI0dTkSPhLbg9DnDLRjesq3JH4Z6XJ5Ns6xW3bN8xlXAwGehV6bXP6aUi3ii
8L+lm1oghUOwaMoZrREPBSvtRNCUzaBD1hvps+WDwcxW/5eU3sfc/g3AzXyyIqAxwGklAqA2DPqi
i2B7Ob3w2XOoSh8E8D1jiSF/MDMRDgKnOMsNFZkZcGrmRFodrte1w0b0Ku6yuNkaw0awA1JNiZFZ
ddsz+OVdynSbGnkd+AwXMkU6OVwcBS3Pt6KwDegOOtQ8IRC1w5j6IzYlWJMWADoqQCWaeqlFl8yG
x4OXG4BdNv5G5Soxg4z0WLdOS2jmEy0Q6Ht/1S4+PRzJkcA3g1zYqWZlZmAbW55mgKIFYTx6ynpq
gDNUwB+yWa0G+e850tGQNyXC/9lUD+NNpMruFgwiuZaDcEbcixqkSrdOy7eOuVYtXopsBlFKzawq
hcYpPDa9fPBB2AY7bNkVrwsRjbWqzzZDeY0AAtmG3Yk64Ha5qDOzdxpcBBm3n1d0gwKBiIpZNl79
LCcJUtVk6tk7nqPffzKglahPI4bbPGStm3UMiaMdXpzVmaeCL6pNwEmSocfjkNHvPy1uj4OI7URH
aPSduzut678QGVfuAISmFy/wDpfKaP3LOG6uYwITJVXWdCArM/rrZcBuUftV+5/QdMGKVmjd5zzM
rjWHnxNqyV/mBztRujTebzLBz5qX6VqCXMrqXoZWrxToBq2qo6yFW0y0gdayoIJbj8Crdi8HnJwQ
86RHGFkEY5CZDS538IduR4jLizmsYFSIfIwPUbuGRGwwSiq6pRud9f25DB98UdHbMe/yPtSswLam
H41J6xJNYKVcPOsgoWq2i1ToTA20rBl4Ed/ovcLQ+Ll31Jv9nYauq9JOkfYSZz53q70CIpA9Yyif
gJDPKCJC2WPh3CfVbQt6tYIxbIzTc+/3lOU3Ya3Av3FAx7d82rlPUSJoiyRfh7JB3hRKqKrrIcwE
8jNHsB7j+lIxBBW5QrT1g+NMayyrN3ZAW4QC2SgpGeMKcGZ0BR4gZqm1rtEhrzecXWYBoUFUpzrf
eDJdCAA9wCDcxiku1+qs/X3xO/bMbmXjjgdXsk6iGKv45vgAWqv5Pl5FxbNfw0Pe5ZUHkIyvkb3W
Pn8DDvjP1SHQG8WqKYVGqS7gnE7GmDJUbrHKrCLwJ9CEveSXjX/nwZ2dcTPzM0+Tuz5BRX8GFdBJ
E5eZ7+ZGSkVrfLCHjqCTOyJcMGiawTt3pZWYWuSn8w6MEq72jI/8hNV7xbqvwPTj+tLZYiVwd8Ta
cAc6lic5oyYE5ANfZxjrfI9LApI9ax7gJMAzJAAoK7yZo8N94HdnocR57epAXWlbQNReIWHsCH/T
QfODpXeKllMqDc6xw1tDp1s9D3eqC/gHmyG8UxJt0uYqSQN8vKc8mL13GmyM+ZC6/U7KBjEVlm8Q
OaBltnJGQnQodrVs2r96cxmSWgGWH11+DUCo6xF+yEMg2zaG+p9OqYI6miDCfdCdpnZb2Ctzoa5/
rurkokMJ2UDL1EMkoOf2MyQ/Uf3KIFa285tP8l1dHNrTMux11AGsWaBZO5Ph4GT8ZKjdXUHcgkDF
qWhMX8bqZvah0fiNypwnn4VmXk0avNQLZ2Fvmj84d9qXNjnn8hgULBJ54bzJY3vaiHd80CfpEnqu
cnVChQPdJW2o2fLsV7D0YgGSE7QgWVKq+cQTblUbA/Ptqr+ZJdLi0i0sKSAb6qSbAoK1PyUniejn
Vc2jdeFYG0V0B99ISNfPDlbQsMNj0vRFDJDcaH7aTFdmFtTWXeWtdjLapIegZV3jnMsnMwBtHDWR
W3VHQJZMIHpwiMjx0Ld27vCYVMChmRaX9pKNpJsl7ZcJ2hmg/nGipbxkAP2cBBKbpW2D2JdPeTIF
IUYYcygSKvLCga4xF5F5eMJGv1MmNJNGZ6RYfFLIjY4UBeZA8hodAKLr/pim0oKOFJrvW5fghBZr
C0wBaTg9sBI2Da0mgd8aOkGyH3+87vqIzKhKGG7IoI6jXpZeXMhcIBeCadkbVhtYbe5IzwGzzX/M
ibbl919pewVwbn5Ao43cztwMPM4cE1PZfSLT4Wk2j6X4vSRztj3rRJDibYgOci4jtD+ycY41o+Ka
EgzPwXVLYrGagxiIDixwAApN0Bu1r1RuZ8Xx4rlDIXMwO8yB0WNry16fE3bKP8KRogQf8651enwG
eJ4hco6kwsaAso7J0ywptICefWlV5g6hw8aX0swAwrgLZioe1zmYZ9XPseDBzywiVUOZYWxDbCkq
U9cUrvyQjlwXUfZh+NfFIT8wrVwBwwL0OPKoElmAVA1Lsv3uE8P3VpjwpwATSDfNhelJlN2DBvgE
aHBqOtUQyDRLe4dcnvw4opLS3xt1+a/y6o6JoE1waRWJd4KU5fRzH11D3XTuEgysRBDGUH+GIq7V
JivZvK9jr2hSOkuEiyTtSpTAAP9HG6nbyANzptZC1GI04i/X1LnXOLbiO75zb983Xy+QFaBlVBW9
F0s3/nF8IikDi1TB/rz4z77keqr5poV2jUYJrnVxSlzdghteyph0a1o+Hoc7FhCFiwZDCSH0EvZR
G7YzYU7ARacktLwx/61hOxsF6e59cn5L4FhauL8gV5mkti2uGRJxlEvnyoVGNUHx1jxrBERCegRA
tDEypgFXMFdswxZaaY09cLAxNCahLAsTWMKYOXaF2Li9EFVLikwve8gl5V0n6etL5+YjCixr4xWK
c0weXO7bmce6MUuwm85CPrxrqYtQbzul312F2AhHW481Ilez042MAPtEzIb+fNRNZoQmQuhbjLbR
oUX+XfQsQt2RQid7TY2ad5t5J/VSnr2+hO1qosGeyACrc7vhzcO1jKVP5PoRAl9/+TW9SLEmcvvT
ciM+4FQdfIc/hCfvSElwqN5mn0vV29M/2Z4yYS/q9EDDyTx9AD3LPoAVIdEvnfEMm3LTpu/gWclf
Kn9mwvzBvJKsYcf8folOyuldasU/CahqMYW8lVDqhInoMNqvmqQrTTDQRh6ecY0B44SxFfhG+0uC
9FTuDkl4K8TYF+nraGrC1XPxlmlvOly8zAuMYNcTFn4pDl0JtW38tWrPIzsYRUNT+oqgjV6fRqtX
ScJjujzU+oYMH53vsQmnz/OPFc3nfOeot/KbF94yvsB34nVyiwtn41IojgNdwX9/wGPNC4ok9hY/
jWeHY1rc1vXYY+eTZe9Zu/fTKVeC+Ykfx55SnDzSvQdSmaQqkevtn/lvhmXKxE6oo5LqvbuQ2FyY
D+wo8mH7+umldLF+mE3KCL/A0OKt/XMvc0Xu7c/+utsTlE45wvDGx05a8w0zzV7FyjKhbeTlGzTe
mFinXvZMrjasQZthkU4vcO6SjjDGkbVW2HY8BBaYbJrmUB9nZDtTwPssSYD4tBqdW94dkhHdaDX5
eR1cE4vH2MlCMe1RsJwWbLBJBtQmTVrYrtVCjdIZMV1qLzykFOrhoOpxFc68XMMajoxmcZ35lmUA
TM8JUM56ZXLh3T3uDGQoxe1JWm3c4GCO0GWic2XWhz7/FIO6LzI1ntpbzxyQWzBAohQNNWnw2TIO
QRFNcjr/kWwWHwIMC15cTnzHWdjIc6V8AdjV7ar8XsArwLvxVXuVnkQLsytU63Xq1SSgI4w2H+m/
JrB31mF12cmMABZ62a+MjVCaj/H7t6C0JNYnmvn40HlpMw3tbMln0vcNI1pzkpVFER+7wOFIySzv
Q6ECmXCcbKGPEuU263oUsR/S5Wo3PEJ/VBVJMfsjvKsCzpMY2zrzjkyOXxZraaeOer7bqAN7gdFa
oHB5BN4hdqx4qYLGrrgrAFa1O4eCYPoTsSyh900jP7eGnKhtv7vqLmpg52CpcE9hhUdfJcGYUgaG
zriTTmcoOLFaVV1izwF7jCg269xTDT3SkfbYfsMVxzkNBMI/tNhUAE/k59bOWH/qV1HORq3JDGmo
ttPmALbfQwzLFkAjP+WgENmZT4EyjpUTp1vyjhj7GIA3mSry0V46r7vTP4nO+S5zeOnyVBTXPSRn
CRUzmCK0rl8iPZ2bat5U6CksR7/WjdsCinlVxTCALPIiOBqlpU+0QnNB2ZPdrmteW+lU7RfTfkOX
9jH68HCGbCF7YcdL7jbpEH1/yPdcW44reCk6hrh6WSSanofBwm9H3bFJSSM1zGZU3kWu/foJKo/q
q7bZDisoUHla1CGXyP+Ce5EzYqjzWFOMnNI8iFoDOkyAQnxMrUl6kzXW8VfKz0bouW9OkmWvSqho
RD22R37S2YWSmTIVRBvPZDKMLllAJc8R6GTzDcBjRV6kquAvM4gSnMgNyITLWkmC1oUXZdv+7qcQ
ZN7P39184A+YtTe+HH/vq0dkF2JPOyNThdZYoensvt5KaI+Frfe6caMWnkbgv4ZCJFwo3Pus+8pX
zmr0xMYqdNUTIHqusiuRNC2+fKZ0XDpyr0I5X5pdof2v9jTKFYMW51LP7it6y5GSOlgR3KamdWBG
TOm5CzzozQ8XdgOiO8CXUb4h5wQJalD/x83T5sEnnTiE0zJz3mLHpAmn5LH3HhaARxjcGlPSoeXA
XyDZ4hXsqCNKVfmriUJmEYp1AgrBSXiZNJMqFQ2Vefm/O4guOu1KKTnLOpr21UeY1aJCS3udpjDO
M0agSs6e4T1PEAcvXyt6q04Qqx7o7OM8ONKMN4HOgozHSRHwgUgCLm61/2xCsya3Aklw89EIRUyv
SQkXTCRJ0XYUTk65wkftJ3Q4movgwhJrVam/oqQs6mv2hRIYwOOzCK7qc9kzrEsYAmJS8lSNV87/
E4I9lCOYz2dstxapilC0UPMci1lO2blZmI1DkrZ36AZWHhT0HH7El44yXxyraxJO5hZtpzAz0YsB
7iEoGq1X3Nkr3nKJOGcr40TtRkVsDtfq85roI8JUeLnpewE3vEfdpqAaVdrUCmWDSnChfuzYaOuJ
QVxYmsPqygLchf+RK8eexYSqwQHb90lyS+mzh/soLKmPzyFLZVdNtRaT0ewb2bDeu09ec05n7BH3
4A3PqJVcflLYV47MJO4i7axlOGMoA5CjERtwhJRabk6ahJTm9jM25KNJP/LPMfgaOHZJm1T44d1w
8ANr+gOplmBvyUUVgMa7Ap0QEW56dnnrBxCkzB05CkhMa305fIrE7ZcdxFCjE5uNWH6c4DnmV3O0
Nhg1kUHXVVDdkzty4C1/GIn5EDOzTNVJGRQODqrXG5PpcLQEwxmpRyF3FcUP5Voa7GlyNQkXcvBY
OIuEjhq2B6gJMFJqIQI73ackF5o5rxmHE2Ecmc1duTzgAwrEDuI/JG8VsPF1H4hAw4q9WDxgBmiB
PePqmwom0VzNHdIRU9eTsVkkvpy4c9r2PA7b79YzDjAY0/h/KOHxEjqIJAnuslU0Jmrri7yl5gaG
6YDS0uplM47fBilcEDKa0fStxbA9YPbZRacdzImPBl3VIU9R3BCmI3lGo3eCWv6iw/+M8rN+DocP
MU1ghCQhAsdOk8xIrvHQRyrih0L4WlZPe/G5dtZLFGxSkVBd+TlnBMG0X495QQZYpoJAW1hb/Nuc
3cV2fQ1VT88ZtSaT7Gdq9ML1Y3uW3o5uf/asnzntwby0Sn+YbTV/8WgmtfNGiaKAn9Fx6z3IAh7Q
ePdyBrIFGAmZmvR/CiiJPVr4Bi7pUQCVhmG2eTIsDutqe1VohRFr3adjPj6IsGq6GixDep8z6x1M
fFNKcN8sM3IKIn02Y0HaE1wWQ1iTX+TlXwlGdAIDTfqMp7xfMvnasy4ofgW9tttLwg6D4AudDw4h
eOWn5QxVlgLE4w+lkqYPxfLSeqBpVzmGhBYfwdunjIilNY7NXAnisJZYIQYY5BxjRUheDJApQ4B/
Xib5ndr20MXmtNBJgqwz7LjNmFlPDSrO7kc/UIJU1LY7azgKMx04+nVTadC+dz9IsK2oNVTrSkvo
EqLUgmMa3GPUY0XbJbYx0iEd4cD9Q1+/P7Ms+2vBCSEG4iVQ5lWRGGL/iwCvKzVOqA28dcVNxFUA
H989EH3HYVS5/pi7EgUW4BtIT4TmL8XqWGNPisYygqDiR16R6yDlEvp+JPOh0KF2FujlREecNdMQ
ONVFOwU6uG61dR8Uc1wptsmjOv/ja0U23Mh/9nvyCHCUdeLp99AXkEvwnZMOun7r7W97iNGmr83f
MPt5ivGHPRG+BzR5v4WAFuccd3oHgh2rDpEkDplAoctRKwIp78cb2LnP0an2vI09PrtmE3v0th81
ZwmUzzjZsEr6a79JwA8gNn4PHQdnDHyOWRfh9DPpjiiYaxDQ+AN6x/a5qbdByWJStgdRN1vwQ8Ap
BkDOpZPQ1li8gLp8bcZ4wiNkxHXRNsOHaBz3/vdtxKSLMrZrD0l6/clqIviraDppxHCaKCP0N+q+
A+oia0m4MAZW3nkjTLqMxRzjERwHmQh9PtBue17HdBIryyrZLwhOxMoqeUVMEmGq7WsiuQR0aqEx
YF22sy3nDaJOGZWqg6vuf+mFu9cBQmaI2EFOp9FcPKGcQ40SOWfsfVVNASDKuOkgFTpJZCh29G07
0ZP53VmyDW405JVwGpHEx2/Iqoco6hAQ1UpcdPlExLL8tvbzo3dZcseobSWJXO21YalPEI4JwCpc
sgF0smOkTHYsZdeOxDaXgZc3PZA+AKt+9wpEoF2491tSxvfpm03FldX3kWWhev66ghqdQsIdclFH
rLywKCVOGYHTyv7eLcn1W7yDJh11Y3bBTiWTEaqp3i4jQtQ2Z7SLd+ZkVK6Qv4vNW4wFQ0HMzVEA
XTHqvlZ/YgQ1Ez6TWZrANIewlR164J5mBDaJXEqY/dWZT55P+KF7Y0xsYBFZt6ATcVFBX3xkiNzj
7CjLcXwXCS9Fd/SUcXF9S77/mDHsiU0Jknfx3YsdaT2QZqzCkOPVbbxgNoVrH6nRgJYZdvqCGICm
aa6OY3gM4CNEZXOJiL48E4p8Ovr7K1KSKErLlTgoe3eNyL7UbYZm7N2e4uaxaxVrG8EkT2XuYfeE
9LHMlv5jQv7wqHJlixBXx4U2p6ZPwAILriceT9GsVoGf7q6S55PsOugPUlqc1NQ6JGYV4JQcejEj
7QM+7RqXqrbUwTE2y/E5Nk7EFAdu2mSeL7ui2hZoiUKYumfkPtIYksz+yPUfxZGt4XdgRpwRwJxN
mZm+Jk8Uuvz63hxH+P30PL/tklhZjwVfXxAqZYWxIAN5nAGySJxucKqkeRVsNRyOazDeysutiiKI
9fskuvi08Fyeu8v6PxkXgka886sNSZY1RonX7oJVXFGqFhulC6ahhs64hu9iJejdJdjTAywkXiWx
+JOXSTA/iIRJwnKsTCcpongZvPUfhF2aZAzjIz+urCYOfJL9humW2GrHhBotWpDPeEkDtugf32VN
DKGmVG2Gaqii85VQNI6v1JuG7Dxt2eCxqhjDioLqY8wjxb6RYhDAcezpPzLWKMUfqDuEXkCrhIBT
tcwC/HcrC9efJgqwCtMhkMaRg46DUwz0YfRGIHHqns0yoa9tAHA0wC1/NAoxBTSZNmqme5OWvxX6
oUvfH+vdkDWtu8NBR3PFS+nC60IIphm80T6b1XIn37+cNIGJ9lye0M0ovj2iqLtXJQPv+JxvWaVM
nSuGWykBmA4E66VHuAPB3NWc5rBjVZNnI9Kb6AdoNpZ+B5d4/2V5OBXUUUPTy8IdqXpoPtghgUMO
b+w8xO5d6IxFUVpHbM81JueWH6Td58MY3eV2vji+8UYtP/QkzrfThVxdzWSE2gHVFPGtCoUW94mO
6g1HwlmpOpczaeHy6svD9WWVIMarmPWPQ6OCEFmnPEi5J90lbHcJnTB6WC+CRstB1s2E+YbY+Bkf
0UPZ+71rqXaYjTr/oCn+E4m07W+pxTpQ/kbeGzwb6r3K9DYagb4R8FN6dOfHa9oc+wm8I911qph0
yRkZn68tdXCyn3wAoDliA209nrr9kJuKGhruuGot1GjOQMjQd6xCMF1HJrjtuc9vHyncnzobOkYq
bPQAJJJzqjd5x3ru2I9IRLAL2MXNizKzFrRTDCBXo8R2xJXssBy6377uWNV1vnpBK0ftjbrNj5zJ
acyD1iNH+iWjAPX8mXr7LvLeeuPVfjL2AX8vPnDUgYPXsuIn1vFZFvqRzXQTcFc9WtPozEqv9GJR
xATNJcDzGHiEeCkw7/UhLgGFW57eE1IEna18hoSxp/pQT3qIaajqBe/89b8WDEWqlQqiAHhDZr24
SYQacPbzIhvmTsqZvoP3Krq8XhJgdJ9dxlIUUWw8Nx5gYp9OmswcupbNqxZsnpo0UNnAh/MfGp6c
N7PCd00xLovTJEge3r88e3dEE8em8GU2xZKroABXyHQiy6skjMCiK3CfBGMAQ2nHO3eVJ53YdS+t
7DZPzSi+iluK1Wd5bhvUZOQCJyT+mR95nuVD+NTDuzpIVJJmkmJP3tv9Fep/jVRX0juP7nDMckFv
ZifPUlOb6txVhqMdo3dSzawfmO10Y7AbYPAN6BuzmCUol57faQDi7jAJ0AC1kaWNmU6KxLu3LEDI
vK7za8dnuS5qkj0QbCerVbG4cu7IMVZMQfitRItDrvDhFNo73F7knstxG2aQP3u0IRSM8tz9fAWp
7IbRW9XKUkAyuENilfP4ZzHVqvf5ZDt+DTCU8MPHyTFY9yTv/oeBpjphSxm6UsGrmF4N102fiS4J
v1tcgiahx8RgpSG9iBFCQDwRqO0qyLm/1eVg6hyme+yYEqBW4OylykTR1x+i7AVMLlyx0F/z0yHG
yRisZOXxBTVJJ29HO6RlezTKROvMNaUzsyAV/9johge7ssA+AMKDa8kAQjUMAiD7ixsAzhb4b9Nf
Ick2k8Ial1TfD/0lPEyqgKtT4MHFqWxusuJn0rXPNyShD/VrX+Yn49SVyQtq96/0R6zwkLog2O/y
qgWCR8mdMSrgG1nVVM35diRijHp52WBwGjkvGwmyo0xFhyCnzRcLCHDPvr4RFgj4ghbibic1Uxoo
98AyJKF6COaTAXKonOyJZsbdbaRB8FMaL75YFul2qQBQdJdGWAU4yKbND6VSHmkzkbAxe2w9Slev
jS0rPtXGsHVAlCO33Ch8L8DVmRwOl90+U5W+4mf41edYTQwOf9HCVA2mt3V/a9q1p+/5O47LMB+l
C2RJnxyJsdxvkJ0MgeOVTbHFRJvU7eIzOL+JLGw1z4tMOk+beZTwGenql8vNc5ashAiyWUIIHAzB
1rMOPeIWwehx8fjUR4A2CaYbHbiAjKOvk8UjH4UJ6j0cU7AFG+Ha96sTThDYBZ0d1IoOUIF7KQoj
GDr9HEmfh+IyAerYuILg4ctXU3OU+fr5s107ZPdU0y1VI81F9c8meBZ5RQePGt4zjHhU/WBMX8PD
vXC65PVEQXutaa25sk30ZbwBY+9B32XOTUbLva7yXk6dKUEMETlM4rtTABq3W7PX8IP5z/WEsv0s
edOi8hJNaF9md+J1d8JQtEvMXCqGUZfTsv28lWKfCV9ierKPRq9Ryaq6r63RxFNu4LL7/yoXhIHo
SOYVNmgueQHCaYYV9kO7HvO7Z5zePeVX4aotcufAMg5leSwa1DP50u/OTbcFQ4OnLFN1D0/CGQh5
dYyH2aam1OSDuCOTr2TfuKDkn3eeRYSvzJ+Kfooiqph0EjFoLpmJJ+mwTw3elH9GqxorUlUY7Mse
IG+Dy13dASEPiKjgH9qrBj273a4o/yMEjKYfSjFlr7MK0OpF6vRhxtBGA0MoqriUKyHsnuL6nE3M
BbISdGGRuFMAaCNoENVYMalvsK/Sl51ggX7/HR/5xoiIv/G3ByLfVhturptrrHg21fA8yEANmhHY
d/APghRgEdDyQplcDPMg0jyrprZCGNrbnpR3CEEZngRV2UhGL481QAXv8ZD1c+uhLEO16Wy5AIDM
y8vQurXXqq4oK6suLrjXYQTra9INziKm8IJnCcXZyTVbuUqcrcVj3vqGJgInSgcpWkCYRXXzeomj
jJtWrtrivtrD3AEVlk24DZBcxOxVRmdE2T5i97AibcBS4GcpaAclJNZDicfmJZKEFCtAYsHDY2k9
/HwazmvgY56Le3ckWR1j3ML43g3EdGVTX+ao2vWFCElWJgkdzyoIjOrGxNMJ7udHYnlBHJOG/I8u
krfCXp66T2Mb6xj4SUXTDK4RUNdliodi0KgJOUdtCTtrZC4j4UTo2mcO48KrV6HvNYgNj1dfx0FR
IX6puz1IVLkxRGK8jdGdNWfLhGs68pPYTlYPaD3wK1t7A1QT6LPPD7WflLjGa6GXuQ3DtYS4onjq
kfFBWJmpP4QF9oUBiIc0kMggvhbOCQrGOS0TrQafGAv+Qt7roJw3cvFDrOM0GDhcoCvtSnCK0rhj
uFcTGSCps2fG7btP0kxdbKMHsU4WS2qVnHQ7/Frwj65dYbyT0KFciucbWg1MbMWTdPmZR/6uuHds
vANMhnv6RtBQdDWn/g30wb7qLA6p/hpWJNCE4WREJU4KQFKqdbaXCZyFy0I6DPjOic7rAv82dDgd
apwkQEkgMzI0K9SLeH3YlOKZNKWmmJytYmPoGWNwbj6KlRfNlrERSlI3A3PfHGMxfe8wxF6esokJ
odBSQcw3WStYJsLaK/Jb4Wr8wAVpK0C5zE8SSjPLYHsg+GRSxzQVTaArK7dyu58tDugUDkTSlgpt
d/koQL0CKEL8XerYVT/BQ1mNN7qPRule5NFGy8FC5PvvQFDXusNy0M0i0BdQDiU6QIzuV9KoYOGi
rK7BXhEIDCYcGJdvHp6yFUSU+yyfkACDC1J11jHtZFVnCXzLeNYxQFYcF5riVHaF6TnAQdAw+DQU
D47YcuncKRCUllnMzO36ee6lxZilemYheuVfgzW2ckaurLO1891yxMviIXAgmw7APdx/xzvlgXJO
o3FiQccNmfuNhFd8H2bkzXQ5chmu5hpmki5IaBGvdc2offEqiWCAonNu8xvmWWAzcME1uHWS9do/
lvZ4IMkV5tZal5IfQOmeIaMxwPIQvggP6BLnlNROcRfeLmXqM8DTXEv4fhCCu1e8x9FrCQmf7L3o
+qFc3PD4hF8uMtN4wCpzerV+8lTHq0Hg2PBfcXSR+C0AJKjs/6abJpcGlhD0sz5+exuGR82nZ8xE
hP0JQjEKkuBVYvxAUjOnCho0hom+hfh3F7iwYMlAgx7HCSiNFoe9cFyuodpX03Xq6yabZNSRCPoM
olgMZuzP/ofWJlilZ3/mVP9ihrTXG9wLeToydwzx/szOS2uoY2NYQhCO3D+N9dutOyav2NABcUO8
+56JD1iPMkJBrWSAaRgQnWSrxhnCXneBTFT8P4QvKQKDMt5YPUsMqWNAhsbLYUyYsGX5Rr1JRIal
Lx2wv4BWXWrybsGYmQbZbjZrqX0UjLidIg/MCGPOkuQ/lmD+ApVmguhGIYmzs6faRfJywnvDfFFM
Vx2ECuSXZrlvg5n5TpqOmyvptcrYSzI3bmVyFO3NSj1cVdRD2t8iwM5QXZGxKS36m8vi8UvOUvOi
LsUAEb6P4WoZwbS6ZUaN1PeXFui4I/V4JOmIeSNi59iE8ueteTFYDZ9jLqoPBZviOv+FYOfIY1YV
iHGD8Urz3Rm0hJ2nMluONp9P2x/e7Zao2ZVnqa5XDsNTTNX/T5fXixv+BSaJCo0M7WyDV0CNwuU9
lPSSWpVUphRllzHmWRJjJtDMkowcDFqH3bcnXcKmR5/1KryfY4k/aHx63/JR4zDmcWKAk7hE+Yft
kBRk590H5DY2kjUjDDykwT2iPLuTe6Hm53DXFtg2fG6P32MiMT0UpaX07LP6X2ibg+Ge2JD7kjyt
ukw8IVV5Wm17kwx+hr9dOTgoAzzpz7Vc7pR1vV7S7re6dd+K3xVLYYaAijAyR7LxYU+4egUyu8nK
OAisc8Sj4OLTp7Hzj/sbmLSQqHFbzDkU0UzdkCYNBOdS0STuUM3Det8CUa7PNTMTvhePZVpWEF1m
9cWHcqTci9iOzyWWA5ce1xayt2/xTpQJBI2DfGb1bkn4UYyb+x+jcW8DZKW9Vw5aj63krWqP81Kn
JM3zmsAIXqEhhGgYLN4JrXAWUKmqpRx2vfjXMqN9xdiwusCDQvqdtYA3zFtCDyLVQqf7OqS8rngh
GJC3BAPrlWeiRJH6UCr9kDuew8yCCkVdMAwooJV8JB+sezEw0wCVW03J6078h7yDWhVi3rfb+T26
9Ex4g4y25TUiswxVugAui52CLxOjM2cMyCU6iPhQDF6OCGeTEUh+oKVbmnN9Cqqym7gvpuoumEKF
2RyQ3aI1u0SAMFnlWsesgoGxJEzFMoW6nYRiIhVNCAzODHdFZwY3VQEUbWXAjFMGXr4NZl36FxI+
ZU7nelBMqWSbxSCMlfAZyBwRWGrdC6K/V/b/G6OJKV7ZbRExSVvFZzFkMe7tee6LaXNZ52lse/uq
d9kzCPyPvmJcJKNh+wfGKDFJDgJH6eGNNh96UIFpNTUpjNGtVnVhwXHmPApa8yM9JcYqnJAtpQYr
E+lkwqerqfyfVcvIQdRkuMhGKM4Cu8Qxkd9sTz5GTMv9YzfSc1m2LT/M1GehJdOKPc1/4vKIHVtN
wRxWOGC6FMV1Sv0DodtpMs3Ich0r7baVRgsuFM97HH/hDyatMSzR+JzxwrtQoZaIgQr15F16YHCo
GrofDRl40hr9o3HTfSeGhhVF4pbAqGUc3DdT0MY6z9YUgQ4o3AH799f2lgRDstP9vfO0aGN/L2MQ
BjNQSGhpn0lsbQOY5VrBCeaZNNoWaE5IvaFrV0mJ/0tub3zE0YQW4mC03JyQQaG2J8fs4wzPIFOc
GsZDHq3i9Xqkqtgd3Pvi/gJWqIpb8gS5baIbkPLXsnSVKM9Rh65KOrXjwu8+7cqf6Ihl20jQ8Xq1
Ay4rG8ehBGlYrNfu9V9oG8s7l+pNs9eq5wkja82Uwo8ubjbrQIwOOznNfh8ABQfVNsCLhkySndsI
JimeWVoKTL+r+1ughkvpJd9+uwhWwsIwcvKpDWeeH4cB4inVRdx/2MBt8aA8IlJNrBoOGC913GXC
KBEmSYAhokaUYiPS9FqhvwKjnUVB/chfznf23RS3798lBuHpBtqXrkamS1EawyoJy8UjXNWn2I2M
LGfLTSraSabSdGRaSpOGmBkVZcLdzgBdcmKZ9oIrpbsxA1JkS61U1go5x65de4iEPv7uXGKlE/Fr
DSRtECM2Y0cpRk8MVR8bw1dcy8yb0FnSDeutSgkXrOCHZv0xM0mNCUdQLFplmHkfzWb2dbWSzsDH
4oi+mBCQNQvnZV6V0mc+HY2pXEnSckaoLVhUscDo77SZOlMceGyTCFoK5NVQyFD7UG0t+4hzABNM
aBNEYRnnR1Mgy8N6+o5JwcUBZ9N+uAqapPiJAzooialVBNrfQMXh7c5zgHalTebMUbmZsHp29C+y
PTUJj4uiy49KtU0+uPH9UpwbxDGvLwFwlkuzDT5V8HISMQeS8psBTpwe1aOOZYsh/7gm4DGEZrVa
4C5PwsH74XHJy+IJD2UpjiFSA8A4o0buDEminMW8vKc2IhlZv4cQWlDkcDy+n8QCUufvVynLhb0A
h8lBN0jMesNbw47aJ3+U/pIeExo2+mby/LjiiYvahfVPUbex9Wo95sYKK5Q79AeFMPIGWFmcBVOc
2hh6XC170t74yRxX3cGnxn1JW6M6d+xnkm5hh0O+TFpnVSjCClyDyLnPz8qnIuiKCIG5IeTt/OZp
FMJzVBSaCBf+zulILvLSm0bDLwwT5YLPuCJ29Vr5zXoUpt+17BTox/2vruabVxSTQrbmy+tYB8E+
EHOapsgfZiJz2UZDhIUazPDk8HU79atjvdb8pGa56lSTNOijhJ4We4jB8mvlepCDKKtkLz0IgOXm
y9rD4aVkvN3RzP+kMMXz2GmAvirOjBIJXosXB7/1b1dz+Zta3idamWa2nKry8ZsZmMlbVSUKMS2E
UDj8g0Y6O7OWw2Q4O7hkb+w2GSpiRTefnrTLunx8NXQzdYLyd4IW+Qf/gb9LChPWoGGK3Vtqyg9C
sOy53HwKcVAhCj8WXSfVj2R4tOe3h1oTnCIbvTT4NStj8ubbYY1bqxJfwPJTTx2H4DvxnpF6OSQc
uVBYzRSQH/zh9oUd2D8s/Wbz15AUg5WGZTwTGxxOT/Dm0F/VEqbx4S4Rgdz7Wv+tIn15WSEYP/t5
pCML735squz7IdWLYezsz4vJznW4UD4JZ6K/nQ/K3SfaGXAelhtpedjZa+ebRZdVlMTpgFEGHtDW
jxrk7Mu89wbpKCW4ngdffWlGEMark5ra/oso3ZudBa9FOCNlVQtQuyuZJVqdr6JDBS20xOdbQBVv
5HZnnkAvjBzTCGbV+W4GK7ACrVPel4ky3QPV8X8vJHhBRoP8Y0rolNFeFA9OwX58dcU6GPhj6EMX
5lrE//rC/jElhQtrgaDYWVKhqaQm7WNu+4y76L7PVla54P5HRe61vY1LhXLJC1XVpv5qWcmQhvgy
1x5SgFWxdm4Itln0r/aefUHDqD7byUXZeK5ksrkwh642qJPzqwLT0EKWkVUzi69yBZ5o3bX6fejr
95Wn5cZFnB7yLmOnZNOf7YuBy3/uFEEIjGkxCrf2nBEkJ9wkI5AZ3/pFNfORUxAzn6jjdBObUTDO
BywE5o6zyZ5tUq4Np8EdKx/P9Pje3D0e3YXdxJFnYNkzgfi7inKazpszRAarucV/XvnxmXXNF/XA
mpBfX3wvFnSUI23BWubWJNvaQ75u2mHXkCLXjlHzKbLwNEzU5BO/fmM/lw6cQpiIfJkrl7oyKxdf
4lvZdbgBDxOEEsftzNt95W2ZYRxQFYyzzl87xOIVnYSfDirwVyJ9XiqOoxpqpt4lcY8PWU+aqZ1z
l37ywamGIr3oXBlmDlMrpcOXslVw4GNH/3O67LjFkAfpud5bptDZ+Cf+pJUFPA6D1XGkJWhYqbzN
VBUJQJCQJbSUYl6OpknuDwaeEHvs0WUBgRARr68vZEI9tiiVvpgSpw2juJaeuDHmed2zS1z+Wink
A+FjvvVBZnRz+lSqgW8yBqyJDFtcluLTs0y1gWaiIeJhKnDJtdhZwulUxqXsa6F8nyK2boZAu5uf
Q6g8lj6R1J7ddYARIk3iMFdO1rnWCJt4+dxlZXT7yRNWc8vKeOM9gZtRjnzK4iDKIk9AnxKr2ytQ
vQ7twC2ndkeC9sAlo+chQfuZO0gaf3wWCyYRBdYshoF1H1uEmQ1Q3Ur/AUrJfiCio/9Bdy6KGz07
ofXe5Tr2x87sZXQcwOiebqtK3cwOFBK3u3Ow8apebVUvSUrver45nvqYNzmGaREPrcfGaDCE2AR8
vf1ZhmoyFKUYrpFhIyKmmaH7lTURSzqSRCGE16NG41FKgwqjUBlGB8CuLpFyAPFi703zaBROTghP
7H4s9NRTEAP8FcjP9qU9V2pNw+R/d+9EMhtbfdkPWQ0feFpSGxC3mnWILbXeFj34yPMsjQ8j4wDP
OA6/svh05eFnXYObNPPzVvumcL0tlIaBTt6VKi9h631zh3SvbCuGR/xLY+K9IKCcfLP0nPM1Nppu
fDwtmaqa7bB9BBu5fQow2/8yrbqS7IgNDyjlKKp1W7IHrG/bPAdryseIfFd7J2/U5bnPpSS2N7Rg
cVcMc3hOvuLA/PuBRvnRwCnm0L4B3jlNLr2VMtszJH8anYc1IjaaZhDVHhEA40yBEJNNxzWbexyz
fw2sF2FNAHhsohmwQ+GM0vttjcY0Cdz4DfgGg8maChJ8sNU8JvZQtdX182CEcmvZOO78T5nxfi/h
nfxr3otL3/HUsOYMzeUoAPbPZi/koem+XKJWQUEyE0ojqaS2P7gmHSr5fg7xEtyezdxqOkfbO8Eh
WpFPC2esjyzCxy8HmdgBmEDHhq2fF/SJ52IVGN0elFeUlBRMtWBJ8RoHgjWfhNZOeWjKiPX/Ubn3
CdyuLj6cDK2QK635ztCRA2Kpffopcj4Z2jDk1Pt90v+NlrmgzlHERNoCZUDg56NBNZiSwrEHu1wh
zY2m9vIP7+kWpjHZgFTPeb2Ah6oF8erXA31fZ26dDupIjo+NyRLHYU4RIqpncoda3dj9w9jpChZP
Y7UhUn3tvegGr4D69Szjj2GOokxPCUgOKL1Q2EbDP9CTD4UFDaiLxIPu14YtKxRmmZsIUW75MUbS
1Xsd3XasAIrTd7YTL+w208femSd6QieeH6UvgxZU7dzgunYNJv8xqtPVuza0QPzGktPAV+a40Vel
NkiRVMlWxd3XIBdJMUBk2oCYDQc3PdYBgEb3seHDGhrhhtosfS8LkdCvU1GtrcVS9IaqZz3FhDzP
8ZIzreGygK89/TRR0omHLlXk8/pe4JZRDwYWHPTuziTBhyYHdioFLMsDjdP+fMf/wCJL5RIok8Cx
j48wef3CYgwrCA3T2JQlmqIwExj9McBA3lR0jefh+Kw/qe6B/5EZ39xWYojLlcHPRh+NQqiww4jC
oHq0FOL0Lv2ntI2PiT7qZyDbjtrAn1DwkUjW9lKexamrKZWX3aVSHwQ1c852cpgyOkp3LobUpa1E
wMilIMjPJlJlBpggtZOZn4TVcF4FC5WXVS6ZtMCFCzxIPa0gvVzsY8ep5j5GBcnhWLXTOBN2SuCj
DV0asX5t7KeBnLZzlbDP/kmcg/0cemKwtcZTxwzdGcyYyLEbzd3APouurnxvsABfe2c4kM3/WnEr
IbRTEvzWEkARHp14BhnIzRPY/AGaHanJiP+LvOxeA9u97PHHEdiNM99riCNOYg49tRXnEQbZvA3Y
VavRh2rcxppA0FtIx0g5X8pipCEx6wezNa+6W3BFuwKCqOZTThV8vzdd0FRqgmWqbvfrB1oZ83hO
1Ioj1dwFkrAdxuL6L+3n/t+qlvF3P1miQtPV/To+GWWV3cIAKb5OZNY5njiPfx4rvSn/pFzaIUhS
uY4RTddKuyP0jzG+X4JP9EdZXnELT6WEQd0kt/skkqfRMW/q6uoBVK5NOF74nemr6HBaaPPcin6G
+RD5k2FWHc7+XsR6E5sYmun3aUGoB2kJFoSW42kVvYH994h9lCa742xRTtwv9rMSW+cUJLA9/BEz
5rQx5oEZAkWznFNzv2M67MPuIvdOBsyIARG/s4mPiZiVPEiDn34XkKrP+mQZu38SfoaC1jW/K6Lc
oYvedLVRMHhAyBm5DdcJ+0IgFppoZXOHPhVffCL1TO/INHrqJutxNZJQ9js/RTMdRbIsloGtKQpS
mRTsFWa/BLHipTpYb1T6pjThuOst/Li5dlAX2svW67nbA9BcmHYlii2TjtQSYHei7HSAQ2nHyBum
S1DTziQJ3sWgTMfRArFBKD2KuyFdPzQTaTiyIkfZ2967IKXOWi3/G8jlwcKsATchd29K7CwYtpd3
LYwo/FXa6ENK8jqZkZ6RbR7lxjfKbHuGylyT440S7FkLCLvLm/74a+ZIyIW+ymQYqu1yktKqO2uN
NVYxo71X4IYW4ceious9ijDygjdZSNCC+BWVmqFpseKGiPR3YWiBSSavP3EAlM/knwI9PNzkwWfh
8b1SSNv3C9HURuIDHVV8BIFrPi2fEDQpTzpKZcl4SLrEentsRC+YYI592Liyqm6ls+YOr6PdxmzB
XtTuo5ufIs4rnWJ9RtZ2Rk9z/XuA7abJd5vdJ1PsY7rq7ZS85aRshUPWGPvZG6Cw0GlO88M8/6d9
qAzQVGlhU85LIiyuIaxcrF0zH+ujeJy8jF6fcMpoMdYfvdZ6dYiW8QW9aqe1/yqg3T+K3pbV+Xw6
s2guBNsg6bINkP6HqDUNCCEZAfniAhhlr5vWcQn64ek2wvohffudLCUx9JRhkjM7MJGYJq7Q++dI
TJUGEwgqRIS8BflKy16WDZpYe9T0QjzGJb0PbmxM/VTr2FiPBVxYHNpL6z4lZEIiPKD6HNscP1wO
KzRJeED9QK7TXgepAc3Xp79dk/gmWscChh+avCJSnW9ABUiBYnuMOTUeGoj7j8pERi/PYqxVKCQF
paNSrUyTNsxlsqfnIQDrYoi02hwnZ6uJIRiR/CMcj5TYPKCxvmH/n7jpMZxUsi2sZRIwGK/uRYJp
TgJ1POYfQZtkNEoKS5ApctwQdfdom6TgBrjUEainGMmhzJp0OiVIW9z5U0jiHR2M0EN7UbjsNR5P
82xHScLsIuHCqIrNOBSbWJc/mHZ8JolQ3KKneGD7EmlLwVqVanC+RXkiOxYIJwnGvPnYBn3OLNdG
AaL/ri6NsMaeezSCSV+jf/HD8kh+VMfn/Zu4lVVIQAhGYOMhtaYa/t49/hCLHD6eOfqcawMEaTVQ
aUXPkIFk+SVSm1xRsj9Q6WfYNOOKBrAWgPbGoYqTdtqU65mFyDTmjL5/qjiNNiM8azEzLbKp6hFp
KY/+78ha/jd571TJlVZaSbNSUvNh5Ka3yIXBvl3NcGkoXoXlLpakCxJU6r3OnTNcLkBbsmJ+Pdim
yxqFbr2L7l4d2xWYavzTcp3b0n3FYDQfjSes1GxRUunFslKXvDUSz0WvGA1uSnFMb4szD57fkS2c
Kh2PQZ8Pa73vnNmcQipz0Db2V41Khi2Ct7jCosjS9m2kCe36JJkA/ln1AHqcoTwRIsBQy2GPLx+g
sNrLNxFhJ4Vn3zWT7B0HoEXXwldFpmfefUZ+qde5sxbHiVPr5eA1Gsxjic+iYcMipra949OOZp6K
tMZolJLVgL5RSABMyZql5G+a1S8rJMBDhpoc156031V5Uus6C3k3CboRr1zx3tamwgZ9IdU73USL
pPtRXPA0BHNx8gya/mDVYgCa+ssWTyc54vwA0rDlkhqOj5t2ttG0PLCFSdUYjAkR+a2c8IBPZ2fL
jDt//NqCOks+htsypDkKH2iaPQqDVjgt/nKVlebxv+9Ox+0+YjQi0nJxGLB0Zl4a57oOGE1nEucm
S4I1sEsLdmKqOhxmmBXzDDjzvpNm4C5Fpw9mJLiKQoClXsLgNy+M7nueeL/AJpkrfpcj/eAlb6Bt
JtuKKI+Oxgb9IIntf2mi48kFlVqAi2yShTCfw4ZlRSAd0+23CKzquV2KAWFdeh97gKcNeTzW63rv
E8BenjlbNEzBtrdp5I5053b+Xl8hbfMJtyiJsJ7Yt1wLwbJF0rW+FEjkNTmPgaKxOw805Trpclyp
8tR06O+2bbgiMO/4EXzENnUggdLRYUyKO+LsZ1Yqq5oCNM8cmHnIZtC+sEqm8hwA7eUOb88s1zxM
fyXzCV+28pdjSPtlI9mgBzhgLhOnOO4Dxx07lNhMvTrQG+biOIFyyRTK9lOY1wpLjZA6qakxYbnU
F9OqLoU7ZIsMlA6u9zbETtguVvL9Hh0P6PQMCL7zXZKLCMbcY4jn9v47epiJEimc0CG9OMEoBOpo
ehEAa4YmTMuGVNm+7tfW0j5IW9lEkUH/ydLEsE6eBPqaPps2+LEdLFec0NMOp4e/DKnPhuikCuts
z4ZVTu6JqnMprp3yupSIA4s9hauNjbINONlFVhDtWCTi8Mf85yCllP1LonjuC4ATZnjeDRHu5AQV
bOlJy2ptJ3Fjk4lr0RNgdcRD3EqZIdCMY70ykurkCvdT2M1neMKukXqa4lcASvoWuU4XhwTPlh2s
+FrTu1+lYw2G5EiQJQncvKjTNOsIdBupnNULTGtIn6ygzAolnnjqKA15vInP7UuSd3bFNk9klSeP
sKJOHCP+FgJAZsyeQ7OSQ1UU2W9RysNmnypLPy4J+NckyNHnwOrsfmRHUklK3T2bXcSNeFtF9NYd
W3p8DX7NlYvHdzpyMpUZCr+JSCwtAhwA5C+RhBioPVITLmBdlXtRPSirSZD7Puh4TPfTTDHo6mjz
VFcTSHYq4EtxSOX8wmvDJZYkf11Kc8S1M2Uy3V1RLoida9nY+O6dwEszaDpW7oi13MYevM7EqPtd
0gohblYMbllyhztdlO7bS4G9dxmmlgZd34JPJPU6tOTzIoVZkGNLj9odtvx8Fl1fOKRRhBnCU4nv
zS8itijazlNfpfO7IxyYGXZqQ0DMnAe9mDSI18cZklyht6VbQb8db/G6ngv6Iu8xhD2Y66bdd+w9
u9Yd+2/ZAnQRowOgJ5tDVHfiM/aJCg9iD+1PPUpDOQOZq+V6b8Up05BKGXIsbiVcWaY3pTmLFTxD
+inG9WWorxFhgu6T12uk06oFO+lsjeDBczS+hUSWM1PXBcEjV6nfHt77Hu8fyMTmo5c19vYI36F0
Bz8+UQybYmooCR7SD2iQSPBTa5nbRfuwFr8THSJLSd0J2ml2gThOfrjtUjhi67cRqmN5I6M9e/oi
iN/UuvLZSoUemZ3fwuvUlgKAHxQ3hXj+ZCGBPnkw9O5f7mX7QRaUFJtIfEcSg49WMpk8hxqhzuIM
CrSfXk2Osjltabfu6sHxWC6PYYkqz68oZlWxoHczVJ2DkhHk08TgGVBeJX62RReMHIWU/HqtkaOX
nhan+elBKdU8BXphR1efwqggbUtmFzMPqDP9xDfb5gBt2/0mFiXQHHO1oIHytUZukuHVhAz83gGs
+jw9UnE0MuP4wCMpg7huXLk4xW1iIAoEeZt75qoorhh/4P1ebYWEtiHbs/JaXqoNZLmBIk7Gvvuk
L3oewJnOCVQt1WUtCOBOGUqY013PmdGuOD6QjLgwiQo7A6opnN1QLfPCQQF+xtstsj/d3pM0aFT+
G0e2qHOQFGT1DcLmZRSKMRgBWtM5fkiO2AI2ZdUBY624Ew8eridv1yeDO/mX8q1bbvrY2tG6YhYI
TcwPkT6MH/HyiJPC2/CKiMbTYqEdOotGoGGMSBZKrMHq6021veNa+1IdAAu3nR3I0iDY3vU9QKwM
tRJ2jyBo2FDQ64JyWHplfIA4jd5uyk17Y28UmiTC3ynfGlQJp9MKLBRZBtGiWLXhzYfbHEaxrUSu
uM0eOvjCO1pBAHOsVN6uCP5vUXNdPySbB32XBweiUJPdBT+K3OxxeemWiiPPZvWOBqaJclcO/dTO
Hofd5+Cn/Z+gEtrWGTHhtI96uOSOB/u8KpV5aXKopnIvDIJG+nrDNYnz2d9P0JgIOrvjPB2iIktI
B01rOSutICveu/52z9lPDwm07ns1Q7a02wOagjAQaTeRH8KhekPXHHQf/u7EM5DS6uz2JWsnecpP
7QqUGdIq7WOoHST9qTohW4ItxwlC72GEPFnSQ9MHnYjGrT9bXOmDqNl4ADWEe87Pk6volHuahiOO
WakwqZ53wE50yC9YE4bQ+fKbNoGWB1pcU55g/ND9zsSNzTROdnU69dxEeyAGOxWpJkYcITb+cCO7
7ZblFCjK7Mbm/dRFe2ipT9hnRj5hibgAD2Sllj1+Exwci2sZdmvrhKx28lNPFPRWzfP3z5ov0VJy
oWBRe3KNZhRsQ815GFxRjxthxzbteykHKJBo7dREOv60DKlmhn98evKc4BFAAR3QSqPLczDrWT+Z
OqTXsdq162GvOi/XLjAUDpN7u7U5m4H7TLPt5R6y5kcLxYZipt0V31xSOScGTBty/T4Rz5Eyiq3H
L/8LJ5ESgnq8Sk1jHDCXmMldSkgieNf1VPjddOTOD7QzaEfwLG6nAlWPX77StF3DPPtrWD4hPuBQ
PdqJJiTnqU+WU5RTU7cXEPFY4v37KaGY+1yQDzNRDZeyIq5h4I4Qhj/VQxLO58O52Gy1QVfMJnEo
B9iIbMU5YiTCBXDudwvABUX/4vGMvB3f92/PrRk0WHwsLYoIqs4BylD0ej2NTN4H66sXnQBuj3jw
//AdGMcxZFlE7SyeCsrLlndbYjvpk36oOVtzkSf4owUyoOgA2LDsVMY7KwLlHW7LdBT7H50n/cpk
27i+JxS01wQkFv451gtmuKome9HzDPCC2iUH+niDBkjPeVTVKj2PncPPvv2KH7Tg5HKGxbDRHm1S
vtF2eLmKDgClHfJM7/1KVmBcfx2QzeIGiJg42pE6E/K4ybxnQKmn9cU3b0fhGhW5Z9XThIVqsLhW
0ura/xG9iM+j26/b1Mg33wosSHiskw1XvQwUVfgcozu+J4IrjnrR3rvsAHI7zmuwWVjfJkEVJS19
WyySBeqXgCdwYIymL6mUzRn/AkvMNwbugemR25j6e04oGSaCf1DmV7rzSKgdrh6+Z6YgfVYCadVH
ppolAwGaWziuI5ugB5pZ1joQpQWytE+yX9P61ZfV5lEWqaHr0fn4ouoz7OJbxeamgiejCfo4nD6u
2EkvJB9tDX3lcoL1HZOUEr8nCqNov2KNtzMZVbTJ3iVjcDq1EfXxwOJrcvpwBiuYCvhCEGHRAQsK
pMyQWCShmZP8wC7mX8i8PojnH94bwQlZZuPLpmJ0/tWKmE4g+knDG9L3AneEWyaFGBdlh3T/OFRz
Uz+bXiSxbGdROBlNL6ot2BidMOzXIDt8q3GjY/VitQQk6PkEuiqeZuXTQRt8bUjLSjn8qQ8XScFE
DsmnzWgRdLDA+UjCNZVvUjeoczRqVXDyjvwCsdg9kDaojoA2vbFqJIAnX7iCVxFkQ0vOeq1QW1L1
9LpXa+S7ffx1XC4+DdfOae8OY8BOr6RJPJp9xRdFWDE0d2vUQ1b5xwB1z5eId9/FO6faaNGNgpPQ
mX+GO5ZzPthQBZs3Q2KN/e+8HKIk9IL9uIGoiBuYprNR8OfclVUQYrl41C/Sp6qH9YRKthoVp+x1
nbKdcGE93guLxmlVnlEzQQ3EVkroeUDrQQW6G3dQpqn2Y/BPK0Vq9VHlIzYMpfy/dar1lOS0+h4Z
ydAovd3ms9nIXo7DjvdFHgdjIOJprsTLlmeIZ9w+uFUjaM/1Vcv7CAMQQSFF4TxapYXnQqW57RL7
LPI9SdtxsIptiuoL95cm2j503gtSueVkgtTLoWvUGUQq+ucdnczThFlJcsaN+UhGNRtCdnksoea9
KbDzOFG88/LCEdRjxQGhbV+rwlxAw9tzurei+TAIQsIR6HTe6XT4hDgBe4aNnuD/w/8JIdY+7FOH
kEtx9i4QQhpATJjn1464CI+ABs8cfNf9OZzuCznLAwMR/teqD3M/p8YwLV5kipRC9ggGkf9QksIA
s3QRRYMTxUIKDPmhfqXmgGf+QoNz/kTxZf0rYDY3WINQKERoSo8FLVAs/SP6otXfJWi4PQrHLohX
p4txwkRhMZUk/NpY45KnL7NQpefnaJcTwpbybCO4/8L4r60MUbXN9g+qCTkP4ysyanMxVScezl9n
/Gp8Jl1PJ99Kln3/BpZwUUsNeES4514Ac/evU22d/mIxuOMEhvxW+Y45zDtxNECwK+HMxbzY/MON
iTi4evVeoiSiVmzvUcNxweFrxzOaPhOnJvVkHm9BquTvCTPiDH7FDnXvT8g2p5bAvIDxJhvkxDIq
b/dtupEgGvdztKPd3qj+d91UV/tCiqbJ/eRM37h+hxhc/HnNlXb1j0cQOTh7Wz8tK8qoFwm5/EMl
Un4v6ZBHDJZSgF41vhqv8cYJl9+m8qx0Db5doTpkbxpCqccOFxbY0ZofM+fDjGXcDuZWoxqxamS7
st9YxneORCLfzX6kEc/SrFgjhbWNvH7egkpE2wCWUm+IhFYAEEkxO1kLDth7LtQJReFuRVCI0TMO
gQ2Nfl4gRTjHt81rpYt+nXPvX6601w/QkQG0tsCZ2pJfNNfWCNQbGzlQQunDMyjEoLDzdcg9eJ0V
rX5j+fcRsvtV8yFFtVPYuEda65SNdGv6egTVVQG1Rf1nPO3EfGr9tXZyMJONGyUcyHqauWkIcTrp
VEUL4tiB5vzcqcrJo2IoX1zccFs58bkxSdIM1panwhB+yPhm7tskIVWSKJ9SQtRetUtn5TwQjvXj
yUjCw2p0TUUC13jhJYd3Lx7mOIb1cMWyzlHDQIrouYtINoTA8ylA3TwefOC8runy8JRX+H35NEoP
xyeJ9YTr7Ngpf6KUolGBe1JJOsrXfnYwPgB5hR7h/tZhsi6hjktffBUPTyppWsS+vqM1jvxLRKDE
OywTHVeGmMV8YpMt8iexHD3XYP5lhGqqto17uGLSQftsggT+KTUlotmq7LJlDWUQjUHVoHHLJHI1
LtNr9/8Z1an9611X2rLWZvkIyEv/eNnhRlaxjfWlyJQ32HUx41SthwoWn8VJMsigdFnIALgSTtof
xUbtyP3wchtR9KkpXEC1sISro966AYgWzYZxh0sgzvIQXs5dVSY3MIE5WnMOGkvwCxTmJJRRQYKu
pYzGmdrxwXM1e0foOMqzeaH/CF9su5cIilOE1GHGv9JQYXkmEA38RiuGTv6fjP3FVZbLfE818QeC
f1yq18vc+svLiYZrzEGoKJod7XL2S8cbfQ8JGzYRFcjCur9bMM/GoY9nitVKLxwSZaii+Rj7JdCV
D346KuiMSU8275zAlvC3VoGbxQl5DeEc2F6LZBsGL2pL2lH+k8sa/Lm7SuuV3gNnO68PhmM+bnas
ntmRpl0e1xBhmFG+UPorlZrtcKEwdWWzp03neVG7PC8V4Ugd5QOk2WlSh/hpG7t7xgI1H9GYlK1h
KuKaQmjy8TXaPYSRwzeZij9K1vzP91QiO5oVio9OwKeww5rCmcSCDNf8UYYQuBCDOxPpFWaSBIbQ
VxlbsdD8AElshaSEVy82GWZyl965EN2WgK/KmL7EIyOgWZV8Ywv2j0tGimdDKPWeWn62OErtvroJ
ER+O4Cj4Gf9ypgTiyT73A6bkvfITOCqqXBjJTWcQDIt3Iqu0v7Ks8gCmC4H9XjMqWtEYYmACOOvI
uR5avgzSPUdMSasc1eBWlgw0tM8ODpPUA3WNXgrSaq5APcRmuSWpmL7UqiiXBzDGD2dj4AcrktQc
4d9ZeYY9h61Bfrk2DJfTKJDREKg8ODWEyWNHacPzv3AqTVckW9aCOFgHGnSDX9UhggqeKn/ZBal8
kR6NGICtu0pO78HxGgC0VfR7gP8xOteX1w+j+ufVyeOasI7iaT5pf9v3TvB8jGkLjpI10IgBbH4c
uhV+dpIq0/NemofV1km58ezWTeJKegGmIrQeFS3v/o4IaS4WaHixDzFwXjW2xLl0H3Ba/dga67v5
UPyNioLjOls2a5yk9F3BCEoKuNNDxkiPQ+GNI09p6BlFEwKiTMCwpwG+7lwa8HWPlswMdpYsF8Po
bISO58c7sYlDucPIXrEAeG+jhzDZqSUIsiCO4JBT0lvUvcdAM3wzFNg4SoGv1aMi6Phn0wHBEJlW
MwXQ6NXXy5W7MwRO85YG/ixiEXzmrdNKvNsp0bBtFb90RZqLgE0ZBaWJw+ol1u+XayxxKrLt4H2k
e3Tw3EAYAF0Q8lDAh11xYoN/9TsGEd/JP5vHXuKdtLoOHnhaikgm4QdMabMH+9FRMLUh3fvK48zY
PyEJZ4uDB55VvLCVt5nsYb4knjIXHu6Rj6vlIenxQA15QqBq07w6OTPGkMv+4PUmX/RyIZXq1A+p
P29bEwWRaXxX108ktRy7wQP/1KWmxufwtaAmnlPbPpXKNJiWpXYWvpcnc3+9sOWv0hc59CcMWEAw
LSMDU0YZ4AgDNlQPPclFeRlbGZsgK8HHluAQTK30qbXzn+BjfF66ccHHI4OxQd9EINR3Y8knj2Rl
ffE9kg7NOfGIZIK+Mas3LkMZvzJIraiOUebw8hcyRvB3AVH/XHVus2CJWzP83/k33BkG/cUqfPzb
VyqXLyLPeTcUOSDIgyhCtQXzucD/8Ec/RmRD4VD3Eg0dt1YUVNtU86qrvnbtvrmn0EXF1Ik4u9tF
hme6dqUFFf98iAz8ArY9i0h9uxyYEhJqkXYgNqQkzzkCu8OlgMuLvZsvgyQOF4tb6EOqNn93+zOV
wYT2AFbMp6LB31i7wLuee6lHVem0s4AXUyGblRwqUV12RgAle02jtf/71QcctkGIDyoK6rs3xW9R
a0CsVCJene0twvW3ZH+FTo8DePsXROUakhtbDNZQjgzPiaNt7S85/PsmHqqXL8Ca4ZPvuiwAx8P7
4TXqrp5FsIM6yOtFkYItVh/0x1OG33lgEYbuu1Q3dcnpI3etAi1A0lHHyNWqflV37qpbO/XUHTX7
PrMQebtguMtyXlVi8rjL/hrBzHHXZpKZ2xe5z25V6RdVAhBfClonniOHcrXWspC5pXhVTJ3ooL4s
QcHRS4/4r82KNhKWB4RrMJsh5Y8HN3cEwORFjkL+eagNbChOtsiNOyBB/sEDSuNqc0dzPBXXRgKM
ukxn5fFJpQjfVV9ThOb6EzZgpAFYlETj4TtHmbK/TQdGYOgKPw+/O7vR240Qns2S/dZGlyAp3Yfv
8l9Jcq3I+yp9zcevjOeOgVJ+x2puog5FsK7HJP2Sa0DxnVnIE+dKMCx6iMbYou6eX2eupY0+dX8s
68t8tsf35wqdTTKip5bzXu5BBfrtuYTIXEL0cIxi6wVJoy+gsk3CN5HZIcM+jrbbAJfD2gvX8D33
aorW8mkqHPA4sKInB+uix8RN6TWD5Lp/t8M9KXjDp0X3ehN2RhR0Lq6t6Unx/ZpOYO+Ogilo/u9H
sb0zYOhcbRB1A/VnYkwZwOt+o13C0IkVxF2MZCLRre0JS67M9dR9bNpWGILO2XuA2czU+Q1l8RIB
Qe4oQQspM3+lSOQLD1zf0OR8gXCQ6HcABADU7mkvBZrzTXVnWykF72HOzKHpcEuvWwStXAG3VWsC
LVMyu6lh28uIKllHQd//Lf/q95Rg78izU+lTHsIF9lxZZOqqX+faF4AE0UJDwsyW6CtninCO0Hx0
uhqIAABmNOipYLv31tkH+fE2Jzv/+3zJzO9CyPGd2ep2cC6KswALHtXfCB1hBqEj6EOQQwIm3af1
irP8540dzvxJOv/QyxST6HEdL/3ByV+CQEj+/c8YvzDNrXnlHRaY4jOqrUc3XXqhWx5AULQrORFI
AKOAsnCds7mtlCNjhmC7f66+P9T1QsXRDxHG5TZCPmZho4QmuEEqPYho2APrTyaCnriLLz2lWIHR
WnvGwtZQWeXtyVDw+OlsyXpHKAA0UgzbVUWlrkcZGzK7Cdod7B+weyq8U0ixmUhm0mp5skN3BVJr
teTQc96EQ3k2X4HMny4oTGFvIesG357h6oCGFO7xEyvgRM93vTzgvgQqmjPidfgJxiEhOOVf6Z7Z
a3U5pSWheTmhB7zln/efhHP3Qk2YNLuWo5kWJMnAB336Jn0U3QczFfbBrHwHCEt9uS98tLogsyW2
RflHBssSLSwcPn+pZpZh5iw0srfD3edxISEXIVnn1bLhrIeP8Zq3qz7a8NospDhkMOxE6FB6fMwh
sSC3DHPM920MLuxuh8SK7FC4MLk0LZpPNVYJrtpj3cZM+R4IV1jHFHW6b/MEQ8Hso7C0tpnHuL7a
XSYViOSt079iddszXJV764R0TfbuZiTKj5OMk5rQldvabUyPA01p5hKbeTGwwUnWEz/uAsyZ4o5c
02Ktsf5IwNlX8oXJF76326uXi6aOyS4J37PB1oW+wq9IfIdeSfmWfOT+ldh9nE79jdtMij/NRqBy
SPOJncLzEUWPr5czNZf0vjHzdQW2vJrILHq8rgXSYuFOWeQINBCyjsiRtrzFY2hM+ZHuzrBnaW5E
x+p8F2Sm1kLfSKrFx/w+YoFHZlnPdocwmtW2x9PSEVgjlrSaZZCdQ373Z+4EjWI1mSBcQ/HLTtcr
zX6ibYEjBAfWZlMuvcGX0epn1RLUAp9BYkW9/VNK57EGcljZTZ1SIRZp5q4D/VfzIpRnThzVDG1j
mz20Zu2acXl4M+szX7/ByOiNxiknoOBmSkFtZOidVkEgDHPMlscpj4WyGEti6/5AVIkKCMHxddgY
sOcGmco79bHKfeeQVKqurPg+bS8MaDE5C+VvsFK916rVAc0l0TqC5awWciXPuuHbPxPF++vxSmLA
BppgPoeYRGJDc+mtSDNw09iWD6fARN04wGWCBdFAY1aXl0U9TFsyChKY+QDbcZ/pTTfMKwJ8dxWC
Ygym7lS2jeVEkifCkkmc69s03yIrMVG0jwI7Azt8bG/TT+8EiGn9wXH4Gcw3sdkO+oIxJwIM8cr4
nz65fZePi5N5FuiM7VrUKkiSuX+MlmvhcesgE3V4A8E1W71VAQRxZ2rS8xveLf+T6IDY/XiNNuMf
87Jpdtnn4rLREXGAoy4Py4kk9djdr2nsUXMZ5Ofc2ShP4ODyNcXGoN67TXdjpUG5CWuw7IFtHhqq
jaesjnTKAJ1sks89IzTTyi46dLIy+SrK93yjjwwVLyDpaLjHGI5H5I9lPYQeogJsDRVskDEcXEsy
5DYE9yFhb2NsR1QCVxFkiUB5U7I3JmiRnxoTw0XKI+UK7xbILHFQ6d/YQbnmgnNMFsVw0Ybq8mrF
+/JptxvP461GYw5nTM6EUf46VmHW7FZXnYuEyUVKxwsNPO6LlYkSmP12bs0PvSd2FYTIiMooyFw8
8VxZj5kjdZ5d8JrfUAwdPmfvi7b0H1hSA3HlbJJSKMxFXNGaqJPrbOgLsYs+X/L96h1OD0QJiQPF
a9LKHO3KQUZ7GgMoscoLj5KjCqwAW+Q55On3tF2qGmxpDVVdo55WHdvjjpfYBI1g6jHXfvHrquW4
HWebR5gpmDBXMGgsSI9Wa6r/zOdWkrIitpQaV8lr/crTBL9QmK3ETpUBHM6p/RrPQrTJtCZZD5Mc
12aSxYPfSI0iW0SdQwHBWthI9VpdTO0tTjbMMZ3uuzTL3M2G1ett1dxv+PzPkdmhQ/805yr2Uo4L
/RvrAdvQHX6iXli8Rui+oE9P2mlvYitt+JiccuDluzaiuqjksBffHGloAkny7OyjFvdHaHyjxiKp
Bd7k829elOMolMqER3s4PCqRqbjgPpLJjLsDzCQFEu36hwAVKN32Evw7w4ytnNibCrhrq9XfLc3t
UF0LKdRSVnmk0UZmAWnylyfcdi1yv1vzg47IpE97pDlD1+SacYApfeZb0JrJyPy0NkconvMckbqL
A6mqBzOgFsNWwt+bXLMWIzgSoSTDNi3biBddJ5dXIPrp4iD9ANCAJDSjUSsV/n6oEjYojix7tj6y
K/it7X/UOBQgNWdhEKBvb4DC0h3zC0uJJ7IB7S6eahOZVInd8TXWwMiT/xhSyR7IqLqQMOjkC76R
YIANGMpksn1CxCqDnCWKbIbIBDjFtBR3ED0gES1ZYOxiQ0dRA8/xlqMWWa1H9pXVh1de/GjEAS9q
dh6wXxw1sFwJCb774XI5z74QN/4SJBkHjaBStpxwq1eKIB96xmc0VmLkDN7/n+TxD3xpi6HvB8Gj
iOYKyj3ES8N8FPz82YPvztrzM7QWKkbSNNHN/L5bGFabPjzwuoMQ962Q7qIrdXovlBMLdScytQYU
kI4AntAjRmDDIfwgZTeh9orqUF3i9Xb1Py3zX4b8wxMv4pBJMOAxhcCOWYIJy+iMtJSMrfbRghp8
MlwpJIsGTeQr67TgzpE48ZVD92dBvn2krBcHi+O7XeRIWS1CvxyKl6A5YDmAX009SACRkbxaO4zn
VlhWaekIu3KYHgGDKrDAMb4IuqzkTe7wAT4rowAbSfRoWPTq6rPTBZ3gtVf5d4m8DE2a1QxaOiYw
POEQVnmRd+CbqSKVzgIEss9T6NCqMZYZXAgdvWJj1q1vcdCOXUDZqUdbyyT4l0SRQrxIO0v3ixLJ
j7RB4xCuP5et4K2rHi3MWTltH/NnZxSRLGDgKtoaoG5dsJN7BNXp59d+5a9kWoDPRPu/WCvUgI1p
Iljrqp+q6s2Rya/i2DVHKkKfupN0+2G61AkS3tiXtB3+AVvjl0INzKpEXYm6+vRR0kZMIvvYxjqD
4nr98X+3xTLKjkK/gX9qQp/k86qa8Jx7LzdcqdOwY9WpMr28CPwztKx0OIHSfYoj66SaeQYzqkod
vR0Us0yBNP5dVH4Y5CdUrDfVYey5Axwtukg0+ksCD79iXlFl6Z8gv/xgHc5/Dy7PoTZSDmiqr67p
dAtPKZnqJov9+EVvS4p1CPuYNvZiVDe9OoHbfqxaUCRyKpx9u9KA5SlKdFt/5572+XTShS/abQu0
gbKq0EZXE/7slEkpN0haQPJO+3lgajY0zOq8613+Jes4rgdH7MKI9nJp5iHJoY2aF5+QGHeJGbKR
YX+CBppsRR024qmtJCRjIe4zox9AjY1mVg/ClQBYy7I86lHG+2eqCmCwtTY379aVcXyQfzJNOc6P
4LxE+uFw0yJ/pNKmn6vH7mMZXGLKrP19EG2dMHbmHOTLf9bihFuUsnMyvqSmp8Js+ocsP+xFwzkd
PqNEBhmhDZJlqQk+WiYhRda1QTGUnOIoiq9n5AQn80UoabZ7eHF1XpAHsbpnGbL8aYLMCJotNTcj
0f2kibnAO20Ry0Iv1/BmGyR++2AKFm5XV5HsvT70SZqyn6BN+qDzmH7gwAj4XVrNckvUzT9rHO2p
iJmRQX1ZDko3wSpXQovtkII9WajWIYvzwqCorYhdYowczGIYcy318Qd8q0VlV66648XBw8+5Oxqo
ORzCIzdtyglnnpzBn8qXbzVBg8ftqbEUvuS15W4uEFxm6SwEuoqcnqh2v6+T21koC1zLbuIi5rN/
ZbztxMBQEP9pj7OrNnmyBmUSulrxPNy3iSUQLR5axZmuoo2N1a5HDzBk2loGgYUNgtFdGH+bAVqm
WMXTLclUh3bkPXWd/weZ9goiJtT21Ic8lff6R1hRNNumRZFtqJkRGTdCoHHdDYn7DV4Py+G0QjUv
sBfabcAg52H5b5yaDCodV8i6jRh4Rabqrp0pwbzHtx33Ce1BbpmmzL8k8PPvpEmMTbS+o+JJmRyq
FAfdqRw5g8aUIzn/zsbzE0lbtq9eZZGvPt16qI/UmAI0Oj7viFWPpgTaIzmE3J5c5iS98pp8w/E4
aDW8y22/8vq/kv+G/9IohfW+gPeytLwz8ddy3/9BaO2uOqfimeokukrcGDJLk5rY6lLW3WFIZ5IY
8o5XbMJoUfvzUoOJRsnB0OTUYmcT7OJFmqexXLuc265SIt5xODpnDq5ghhBMTmKw4kjpiUMHrnnY
5VM1BvuDPsCy8E0ViUbHmsfkPF2dKM+K+zTLGBonAGyOlElXp1T/X9zbwZuUNIPBPycMg+8HBvH+
zClKxGjqKIoT5QOPrIykd9ksUQDCV/6AHU4eVZ0AgNG0WHs1x0wcBvY6ziPKWyuyKlcg4csM7wKZ
O7pNXd5BSwyFzQkusi+c932F8aESGeTcnhvzEo/Se/HZbdtToikezoJULpVZVwuY7nHDyy7vJ75E
XDaPb0rdPUdZljSs1aaEwvnkuHNZK3bTIRudnGmmk8CgaFCNQIm24gCLNUdhTMyXzVhmzs/2F5Ml
+CkAM+LY1B03QP1EfkM3Mr0FrMl0G/4N+QiBBmWKhgNFqjN8YYnArtpENm9egZOcMhbMwAZxXCoM
7yfWwHCtM4t6rHjRK4B5RSbbrWOlxseTbI7Fgbev8HW5mLLIR2nxAfbWgmvjCrJyxf9DvDRiZSlb
TVjc3HuWFuA73Sw/Hmxlddbk3loO1ONU4yT8pQ4PNbRtRMZRsnk3Qo6ueAGIB79lGbT5CSc95x2H
uxk//7uupx3F1uULXmN4Dp/qcbmOrbTvSPITGmhKNLixDz743HV/HPLtScCB9UVkl8hLjSzRtF+y
jlavt99sl+uwQgthbcckKw9YbuyBgYThzFByKNcfDBDdsmLcZ6UUgQmaX6a4CJs+VfiDm/bFAcwF
h0Q/EG3fb8Q22XWmxwTxkUX2MZDgox8auPlfhiZ4CQYI9dth50fIaAosF3q0OADagcIXPKn5YzPT
Na0b5tJK5epapJN1eAXVCk9r4U9f2FbnfNU1V4xY8pvMzJP/Qi48VVhyPfkTxuHPJJrZh2ZLCTMH
/XHc1JTppU5cRV7f8qCpOvNt3Nb6o/srp2DkLSPQbFP27qL31Y7cuiST6+cWf7cZVIuQCFiPXo+U
Dek1kED5jWTydwYFRzawclHo9kpfgZcS0O7vMH69dI3BsG9r67vmEsf9XSmU91lRore7PyUJ1Cye
yjE9NwVr9lwrZbTBrrsYH6PcXUb9Ue8ieS0XpeYfgASS12T14XhT+mzVTxRlqub9zSrw304ehsNX
dPVy+mhxRzlkH6I8OZHCa+z8pyxQLj5wJPxkGpmDnrGSwFWHN6Gy1v0xdWiPhCDRW+aFufxvoY/R
gXujTnQD0j829dLOfsRu3O4JBOWLdZ9SzXWCUcOMnw5dRfQYUIjpFMg6GFjdwSJJKStuPA2ETWSe
LnGjsLboPz4CHgtY5dAfp3jgDH9OgENHBnDQ4aP25VzpQSW4bXuhMRF07xB76gI9nCaP8JxsQ6oW
se+zWN04+QEC1cs0bPVeQ1ExBcQa3FZCWcJuVTZhU1DJpqlYfTkBV8V9HfdtDzV+zlO3D1eWFXrV
2d6r1fGVryl2hEwNZ2rnmpr+Hhd1NksLuSN/jbz5f787g2lNiqL2zfhElQJJlvkjQ05YGjMrbo7j
reqI37W1dAYtxlIaUPnQMyOBkjbZSpU0aqWJLsXK1SgAbM+/wvPBLBNfiQ/EaHO0JV6Dma/eVV3+
3ujow4MEI303rf+FnKzpTbJRknroDGIHK36NilATy4G1252GRl4jVwZ4TIaaqlL2yDmG5dzg5yyA
zUQslRE7TidA/a2kn0TCXyuxKU5wwdRLBGIigR/lIdw6KQOelTx+nucCf7nR3Cv0b88DyNuPpaOk
l+e9TXY+Sd1Hd8PydtMwakHoQBh5Wt0DxGpJR3zOCOnYzNPcMOTZ7cYTSjOHh8OAdjwTJz4Abulm
m1hBinu19alzpdH729yc+13BlR7v4AurG7ASm/Qje9GoXQyzvO3V+mYlcVD1TuVj4N/111puU2GQ
bXhKmG0zGjW7aRZooWSUAyOwMNINotJrUYoy8/S5PcrD/7ydO82qvukMoyfcJsZ8a1GOHB0Tf4UU
VsjvwyzZYSTSQXHWCLC1I/bLCRBtEN8lrlfZiVAEpmIjTHZKUtf+FI7ezSP3RsV9lqzXZ+BSQ/Hy
hhEqV9ZgxyNSgCeORPDBk4LehkZcxjdtkYIsxf5rBYHXh6l9sUmzU/SaiFDHhX6n1MsPocKIrIT/
y9eCzUcX8nK3uYkNfildR738Z7Y3kucI7IyRICNb7jedci7PCtLgeQ6iBDC8zAiqAB91poZX3mRS
bpDhyRZnhEc8fPl3vjoXByaWdcar7bU3i5VU7Y0de+7YCkqwBSwGQcrueTyfi5s22fXb0J9Zq9Ia
LeKkwQU2xz046Jnzai6dUDxMau8fliMy0XgThYy4gN86RocIoLhAMjqzUn0xRmT8+LfqsyF+29UY
ZYddUIQ9nxasRAjFlDNg8KJshhOPda884M57PyYJALqTW3d9C73nGlpEKWdQ/fWr2sxiRZLantyY
QeAPOYQaxp6PKozzUjgM3sROPXtTKpwxvOtAO13xEFnHmxEgi98aCybwyXBxeXDdz/q93cgtHSax
O39FZwvFxLaqXDcPSIIHsNgvDXzaJI3FgUFK/qg/ZD+iqrgZ1w47HM1t++64aOGe9xjWBzcAr3a3
2Bso0MlJyBmLhcM7z8NgwhYYyhJEZDeIyQ9wuIzyYDPh/bObr/VmZBhJ4cKusO7OKp6MOFgbfE87
Fevid3KLemGGteYhiNik1BddAn6kkD/HLKVN9U7NC+uAV+H9477enCniZzOMiJ+C41FPW02v/7gw
616RccYgHHwax+b24/FQ48vx97gsD3gCSWt475s0kcK1OA+8fXaRTLC+kREnu+Qshpd2A7Xbsywn
JTuw5MA1GUkpNZuza4+pr3m5+fYRHpET96GJjx/10GISmzquduSgkBIeSDsrl5bICcYQ482FQ3l0
ZwjwO4qt96EAHgNheXohwn81OQO7lNChQWd8p1SPYjvvL8EJmtnmalQ3Nks+tLo2um2dsr3uH2XN
+bgm+KdEnLHvZFQLEluFX0PVteQsDA2SAadHOSufGqXZSQtoyjUXljOBYweS9yhNgCkHZbgOmy5B
nca5+fkbmnWJyypOiWUqxmO89APwcEAB2uczpdv0EQW4hVHzfpptek4cv2mfLCc4L/vGSlQ/rPYh
xaL9+HkE5tRGGN2HoK28a0InAXe8vhvCdHJpNBUW1Mdyx0tiAvQEQuNvEsId51XJ3aX4qK9pQP6+
Cb4b3oWq88T0HZqcNziLKfDEm3eLVk8vzM74UeN9rM13z6TeE4/AYovXiC/hi0toACB1pq2twoni
BUfYbwsqi2WMGoG4Xraua0tTf1h7gN/5009nTqllhmo9t5vaF12WtHWyBkiV4XUl3jP9NFwfxNlR
aQLbpUysp5dpzTnUL9PCiAuqH0kS6Iz2/4J1aLty3EKjxq2lEZOm5B0O78lBpGLRYp/n/a6DoEEv
y9uR1k/SIcf0/c8TI7tNmSOfPgNsbmRPBd8dOZzrMquThn/UupNgZBlyLCfEglmnWg4WgQnFC4DK
mfSiMWt6KZh2fN9YZU2IdDUlREmk6lLibQABkV20COCaid/JgI1MxmV6kgUdoKlPO+sCftA05qQH
Bu4e9kbRoAldgQyGHilIQnESWZMJFqKhViVRX8BEvcmCNQle27nNjVdgMHgbCCOg++b5Nb6uL4On
/ifm6OgFCSQ9UC4YHVJsbfx5LSRerPxcRuk7hBuJHs9NOvp6U4RHLOhozBDMlRVnmvNpj+5+bj6b
A3eignFfLyvU5w5EBy10ZzxzGikXSoEkjnsxN5X+0DG4NYHqP4gBmyZkyX+iETmCIe32cBgBJnuJ
7ak6H1hkOUIQg0TLUifcfBxETPzy4gNqWbV7lZ6wUHfY7gAiQGQ8TH4O8D6tI+MPVx7rMvCTfqsi
Kc47OorrTvGFhJiyflRKBchB/zkza9DP4MXN1pDr+RoLRc1clof7FEwZmIx4zA66GAwMoN63BQjD
xBuHtJA0J8+4aRbTKdVzcMWus4z8JZSN6pWoMdjZEpcUCtS6FkFsAIS/G5ivLLdhJSz2u2ez54g3
vzYfaKXJb3zmesBmpJLyAFYMLZY1qJ1wQsGoFXFJbwLZofo1TTGnc9gwgJJAhxzJEBkzjuLQmy2Y
AmgxD6ta70pYDrYY1gHr8Zu+0BhplN1wMtyKzTiuSiqW9Ab8jhb9zWDxO8YWVdtzGxgtJoFYcYnh
LDDFIDxoK8yenWVZtbEZ2OCQgsAdyI30mkm12E26QKCYJ4mRZ6K4X6SDeIzrAsI6m4V2B1Nah/cR
weSt3uJq3CnePRbxI6NFGuVZ6ildioPKLwqe2pCX+Xzwh1bXSxz5zU/ZGE8MqmUa2kl/JCuchlVK
FoFdY9IZSD5FgQ6CTW8carKICDBBrQcTndS75rL138WmgRAWUW4akCfL6f4B9Y0+amUvtfSfHAML
6f96xphv/PMgB+fkPMsd2/pExP9VYk+sTxjpirI/xNaOLwfKdYUZT46CeHXQU0IF0XgLKeGd5O4O
qsifV6euJ6jHXgtvJ/y13qORoryV5uuGVBlT3MVBcD2p9JDzu8megA449gjN5+YsjzH5JPAKcGNp
Y8rY43J3FYk8pHMfSYUmOTvTsAhTi5nfqmeN/aF5EEm/BsxA9NwXNsd35NKk9DcGcVmCVbgRl8xa
lZ1UYgh1o2zflzPZK1LxDk8T7f0VsmzIZRwuh+MToFAwhbzgHlpteYmDYlN1AaUvP70D8xz8TKkz
KlKoFnvB1G7ArRIeW/JtY9xSwNr0o6eVGzPb5VQ12AplUR8wcJZWk2ez7zEbB/73DFKt9OxO2a0z
nHamgU2+aKC8iDe+WizElLVRrpO3vZv073Cw/haNsnorzlhI751lDfqXSA4xPseqZsiE8hEYvs9w
n6la8BlmfEC4E88qdmLP+zxjEdYXxWRPOUtDsSd2+YcgZXGwCNjRfN8H+RrZ/g1ckiZcTvPhA9k7
338pCLWSCulC99BcxqsysRFEt/LZ7LAAP/rmaPgXX/s1/xhSgFewiKodAlGGWmz4+JCL6UvcPB+J
idde0yL4mEghV956PgS4tl23I0RFFptcISGBjw1abwcOT+Nf6psB7BlzDFXyvU4hyRHJALcwYtPr
S4QYqmkFOyCTG8L31+pikDsdbFV1t7dyUOCxbm1BOKI+e7UBMlrGzQohZucPURd3X+k8ez76iW8e
FfnpDEzXIRfNqKMX6w6NdCHygYc9ERnNQEwNHZKE0hT+axBeSafsuBXJxPJtph552G9xJc2zGUeI
bW79P80YR80AjQYrYhZWGO8HnpvF0fsK2hAPWoMDzYO89bYankV6HaShlvY4h4dVGgyJITgs2Kqq
7v+9uaDhexgxqCZSebwxql2bL2f14+sKCQP8Y36X/N7OT7egHQOWAEJ9GvIX+XyeO0iGqGtbtrPX
XWKvYo4s1HUBnN4r8jPEaNvaZ3ODD5qowbkQVmVsFJtwJWSonC3i935zjLp44lOt4k1MHlKtgL+A
SjLPpu72XVln1MAXw5p1y5NmeICRwY/p2DS9lq7YvffBU/5MeWFrkeha+ewqdr+mnuVp77lzBshS
SlpcpbOvnPx4cYjO3QoAeYbvwXjmnAi/KLmcK449Zd5l0d7P4c9L/ZuKohkyLnw8P+5LJADqYX8H
NY4/5miORrn6IYMacO/7Ndj6lgRrwB1ez9OR4SrbwdBWUGBTCVNVvYnClm/IntOLrTmJZOu5BwYS
MqdMktr1x/DPW/AFQNhKpJydsebR9UKIE7DfZEF+2B4LJPvtXJT2z6DUs13qTlpHihVrF4jND189
wbfGQ4fSpNqEJhT/qfVyqu1KnPbkpWwWJ9t1AZ+l7vV1GdULiveScFlywvFzIe9JY1R7iu5zSci6
Tf3acOEOH1xmz2DW1fyYVRZqGrXVYKDRVDAaprvWfh9ZoGbDXO6NKOGFja1VUVhBb2yxXgYwSvaX
b+vTj3Fc1ekOf5PZJPol1pJjfKQxqWnkP0P7DCnTiRCvT8BtIm/vUbuUfmS31blWmzmcgpoJpOM/
LxGn3g85xZunSLrfKfefa9P3O/0Z85cATg7t56GotmrvrdATMJfk5LZCt/+9tVIwxrqFD/hMKNIM
S4OuRAPG9OXBZL5twAEvU/RKoG2CjXL9HSYzvGk+rpmGMZgLWFdK/mstmqwBxbQGhns0zV4WEZBz
0ETPeJ76z2CP6lB7tOMcRURgSwWrRu5Uu7MTdD4BHOXbXvxXVwpehlZkQKVJT4GAF1W7u3+FDh/V
iGV3mPH2F2bMVKsecvqHA8nVg6MDokZskufmRXe2laym/tkRqstgY8c1JIZnHSCFSXt56RTADypS
vRYCxo9Qb22SeQSr4njnz0aWj7gJVHTI6lZqjl80ibPF6AF1BenEWM8sJr522k4NKpbfMWKWx0ff
6NXVJQrRlSYU5qKBrtE82j0SaKeawbTZ3NerT2/r45drZ1MarGvfWO8L1rTr7A3ejTXaPDamrr5Z
lLCoaDMO+Sf/MhIhthP05j1PfbqSPKYe5syaGSgOgLw+SFWnRbuuwzfLnwCxDiwWx9Q9C1jN4OF1
s6sa3fiqvwsIRHA5p2pBfJ227Ic1c5IlADqitstKR1hpLK433HSj97j8aXWfZuPsdnmeemMGTZoT
HsOPNITPEm1ijQGXe04D0U4ECWvMP5V1HfROgL3TfOFDfToSt9jv/JXbaStW+kju6kVi8uoKDzrW
5Ff+ZakwJMzWuGLB0miwkX1Wx2PpjeZakZhdOkZECVbk3tnJ0Z8lXsz3fmxz8lWD8Oa/b28q9x/K
D6mdCIUx0eM3/xOmGktuYOXjaV8kTwPE+2JMQD7QZZd6ZHQgyW/lJf+WCyPQiGNTjjdYTmoV/zY9
QUqCl/5lxRJVXcqRS4pP/JJlbn1866oZ7nzNcP1Dyd4zcFeMGM4V0gxF+xESbEJHdct+EbZ62HSd
ZFRiWoQX/8r7+pYF9Q5pH6TnXQDzkBk7KqaZz3vWXe4+5HrtOktKcfjDDvqTGP8bgRpAjbIH/naP
H3ToHaSsDVrbIg1zgpxkztQ/edQAG+HALBMLEvY/5OO+CC9jGBk0W2sD9QANgjHKizFMZT9714E/
qoSVa0+owXiXS74Q84xzxy3QgcmqydUo+1E6gLmNwjsACeEudo+nty3+tclvs/Gh0I20LfnUdcng
UTuD53qInUenBupUMCbFCht8qqve616bO+thNRi+PTjEuFyF7vGVTtqQOpG0o56tGnFnN2pXb7Xw
P5LnwvJm4aK7hF4TOiJoOEn/RxCoBmuUYR3hGIbvqMmAjJkCSX3VJz0YDD0128A0sFwVXeSN2f3B
Ptc+O3IUUq1y0Rs7T25gq+UpmB/qoSqeRQ10E36CDYTOyErWNRx1iInnTgYFn05uJOnmGWOHqByD
QBconMl5nFsrbhpnTpMjOimDyDR/Dd+kdiLmf3spN4k0s4S9qrLU6i9gUUurFD7bFsjKAdE7Xlau
t5xGGtNKFjAIO8ij4eahoUq+chnmVI05EmZmoEA8QPZfIaoOCEkLqDpPpL8fmL2aSCrr2a0EmSDn
p3Wmc2h2vOm3173QL6qUw9VOxu/LWRX17jTT4Sjprayxm8wsMGs2x+igPSiaqNV2YT4fxFbsqkcy
fsooAn2zv1ti7BuseeBcxjF9+ZHFj/ky9nFF7vHsQwgTJcI3vl4KgRskWt/BH5Sw2b+LDr+n+tPu
jRCssBnzbo+pg67XIEooQK0/ZSFc9IXaORGW/j6URaC/0xLdddjECngmksFrZndCqDIpCgNDd1D7
0+3OZX4GlHtJ/0MUMjFM//pKGXhCd4hdjLSEbL94+w0wf6in65TpP5iruvPM6wmtsihupSOIlqZr
NLBeLG/Ff7QxX+jdgpm4VyoeYsqDmzLwS+SqezSptIk8rhjhRyIIlFhsV5UvVA8+8bkNeTGSSgBz
vDQ4Mk2JovbQwwLAMQ1y/aaGEn9yAy/L42RLywtOSpvxK275z0xS79DhmYJCcCLnWYvAaawNQpYj
fl4vpn360QF7arfAv2/YNeqbOfD5KM7qf/x/pxWW99GpcYWGRNW4l2yYWTWWSp+114BOuvoGO6J6
p9KJ0YWNgmFI921quRrXM7PMmD0HNurID8G3Kfa94eUoqGi8tUNe5OOzJewO7Che7WIAyGn5XUTc
Kt/RD8519OEeu8s6r4/7QhtzJEL+kor1JBPmOB1XEYKiG9gMTGwVvFUJc0ijXtyG0qLqxq8kUUW0
v4wqM39OnKTG1hgCsy8S7L95jlJFDuAfA9ssoTvVDkOCz/m4Q8qfAemuFRWxlbu0VR5MnHCAlLxV
t3Dm6Va+NGq+zYvArT2rxrWabjZSPADOuXrebQEpRGEeg0CCtIFYt+Xax3ZYyL0zO0jOeDvC+vcU
U0FUO2gQ8j7Q4/o66vd6glcaMJAbp0wrTkOQRlPuplFPKFAPH/QVMrd7o4ecCsMKZKsbuliKCckE
PEkgE62LDgJB1hUEdWXeXuO6tbmuh35lipywbzwVhQpeeZE9hhspQ6a/itcHOLZPercmc2GSoiHQ
c2ptKpJfgYADmAdw7orsrgZwftFBCfpXsS1+y7JdUfxnoSl9l4dyYGeGZ0zjPvLYanus8s51b/jd
Cq8gBR8dJhZ4I9tPgeWYD0gTQEKxMEGfmIURoebUA1gME6b8PTYFahVwEZ4cPLXdCFkTY9TCuIN2
siGNot27zLU1jgffJbQBz3gwjt3eA6lEyFsmMFN0aJtflJzN5HPBQxPSPtoPgcsr3Z6zvbBOwhDX
CEwnBSmx/AHesTf8HcktDql6e48rbVdz00BCd511Et9afr2poWVCMT0Hc6UDnIaQsRpJ3iXzXO3R
tAkpMfDeO95uc0nR0YJzCvG4PIkF2gLztUwCBL2Pzk8NDjBEFDqWK5kKLm+ePQ07lmdR0x4Q1Xd/
fowkkO1Lc67OXBqghTOYkuwRa9Lv+0Nt+ZnR+wEX9yMOmc2NdfEOM/nlfUOT9wY6vzlgcahhIGdD
XLN8qMqwIJAf+QV50ZCZ0sexxQu1WXlF7e+lxUYUG84rsLwQ8eM9OP23sRkMS6R5l62zPfMBySIN
Mlo4hntsVFcqPJ9ADBcOUIhOTQONeAdVB77Sbj+GlY2xOvcF6CqbccYbX6fQjDR/lPpQve20ok8Q
yofhptAqJIxogwbu/jlDo8izQjFM4gLJME3J/5YKeIDdFFHHgPTCD7tC1K+QPZRbJZiKLzIaNqzs
mPNTutFw9MYx/MjItg6GOVS/NpfvHsD1GAGXR+Wfy3qlB60Nkreokso/EUZLLRiH/zWxjZx8RhD2
rW9k+Kv6IN7+qyEBe6LCfYdbrAMfha6cqI9XPqlnHIWZg1B0hGDC9YNzKBXXRQLucgKbuv5KwxHX
cRVp7V2tHvJ5HTPsyKivPFjJjOwibYadftoZfOOoyWmYbwuqw315peGBFIMuqxUuRGPZ7cCoMY2J
WRWV/vCapGqXyQcBE5h4dpODVEGwqSqNZt53sf2gpwh+0mHUB7431AAcNreOgIgHkufB91sQ7VBm
sunULZpa5fGh/3qZqMp9TFtstcKU7DdidPnCW4k1os74lnNlDcelmqRNPl+cIeRlMZjDOH+0LiDd
BTWZIx8klIw28X0dzCHzuzsGnc9EAjYhL/WtPL7odt6i/Xaa9MDE1F66I+oLDaAFLfqzzWkVlLMq
NYvQsZpLj2nmCP2QAgFXYnpVZyhlF362tkzjZzNGnOzDEP3NhjfsXpoqsvIpzuyJyjRlP8yDRkEc
vk3aR9dhgxJzFxuGMvvKRNHyEeJaDOJ1tFvThdrripSb6sYiHzXwZkgOymNgT3zaItKrJtGdfstO
/P8mV4VejHGJ6Jj6SwRYJAnw+bubhw/OiW5xi7vdAw4Dyz8Z+BaHzBB9Psu1FrSZhHRbBpNNXAkf
gkaMZTgesP/bs+AQB4tIxzjUs5UK5f+5x1mku/BGt3Z93YEfSUk8uRO9Nc4ljR2Xf3fdTKytRDp8
wuy915zfPOVBxNRD3lCktMxdMjRnpzEsPKCLiKSZQRI+GjpCjXJvHZyrtJDnH+OS/uDWAvsuqTEl
ZZ9TTBVkBqkLZ3i6mwBuF1iKTQmT6MPt1jFSNQOJyUClrNnq7w0AVyZ3CAHzS3Ysi1zMbu5reElk
L5L3icqneoMLSz1ZfzbbRzQg+k+i12T7UTJ3kYwBs/NftHtpFseVNpDGHjqE+BBU8vyOIxWr7U2G
0KHVFJ1lpz/8B0W8tusg/X5rC/fZrspXrA7a4pP25tJhZyDFF+xc/ndbdZYcMtp0/nQGP8Zqb39q
I8raArYblFFi+5loP+6HzKNiX9bsD1qgKQ7wtoYPYR14SCzAYKkBjB86w9YtrpQkFbHMPxwOKpo7
RxWWCIXTU8t7tWZgoy4aelGLA83IUtzRaj+7rMNp60gBDDxHBI4dFVv1x8lviAI/CHuQhMWHUNY/
02FaQXOLyLPXqOtMfhxwlVTT7fgnH9PtjLuixrujMQNNDk+r8vJz4GkSC1qdWl3/9daHHmHc1wYy
Q3iJGYJxju8joBnfwYtsBTiZbw169hV8iYZ7B37PjOCzhuYU8CkSXx2qJCWpt2nwnfPk1h66cLkF
gNTpWOpe0jlUAx5LjDyhpPyuVWI+HwrZ8dbVkQ7BuCaDgp/ctfmoZhtM4wMKLmQDRWRAFS5qB9DY
D5NZqxgbUXPMJtQVYIX7ClxU4rgqnI4veZM4XuyX+xRHnh8jizoWTG0miZozag3S5l5/k3dLgOVl
+WaNuR9j/7JOQRt/OJPzpCyyooz7zJ0vYUBB8lbEE8nXJdYHhSp4eVKNiExYDLlipNEBuYqwiGjX
evoAlj7OjFKLWt2y0bvfM8OfDjSptsQJqYhObXFvBcD3xSkOLOD2lShILCcAMcqybjlX3OHBUW9m
bhQ/Czh0r7cL1Lq9PdqC+bYobDGTnGq4tXliRdF/R9kSS9/4ZBZt1KO1PA0HIaX5afNPSh4yH4Eo
LwIygiM89G4MdGdjaPQEyMdipK2Nd5vgjcaNVOQbSHkSrXvnGvAG37iclu/3w1ACbgKsue1/F7mr
Amvq8fTVgLORrAog9i56XVBwNtpW5tq7B8BAr4BomVwJdLiu9ri2pq9gPN2XLynwkHy2lzDgFYXJ
3yiyVrsaNQQ6e3vuBHpjDJcoMnlDsAQhWd0A9QQCbgJYsbniKYQ+jCgIQ/lzCIac0CKUYX0TSq80
QN1p1/T1NlH5MSdbSykOBzupNE/X8n5z+uyk4/hRBK+GmRnFKBTazF0e1HQHW67pxzH5nHhRMd1e
FPmo07Jy3X6JOQUVxcpS5Z0ePNGtZmlcFJ0JDyLeJjQLwJNTJFf3ZZUvGw04uKzGdep2JanrYU1f
WrxEfNVvuzsaywkSSZWc9zbSprYLGMblvdzwQJ1FBaxjbf7EnhHQSM5qqIj65PXSL3G6D8zyoIs/
RrIkwWQjgjffrD7O95YDj+z8h/2i0Oyfy6u6UFCwSbWJy1khKp5j/KXaeqr+oW0O6Ifr1pqHKUBh
RhK/cOpFww8s6hOm1SYh/rT/rg5M+T/XHERMLX1V+QlmZ+eZMLhM4KNUTmA6w0zNLuE3pW2MXkRE
5Zi3YAwmzUd0dGDYKbJNJEa0rKK4yi5OEmgY7Aqd6HUb1XZnhdX34N68hlzLHoJsmlXfNQcjOfvY
jbYZY4voxV5uVBfwcDTG34nkysRR71yCHvpRA3NOanRx424FJPGiXq3fMhf8ntETTr/Wxj5i5Grb
6FeNQAyXgdVFAJiAwqh5T/wdp4ogrjM2Hp1+++IfZVJnlIjP5gc2LrSWoYc1YGcrZnKwru13rBNX
3v9Befyats0pPLqFqDtdAKlFdWHIzSnglx0ZZh6MQTa+RkTbEA2jG3/RfotkohVbJK0OFLwBc2vu
zDzqS6nbzXwbZVMZ6vMaa3WDJGjAbFZD0JGeo7x41wAw6IpypV1Xk9+p9dCXOXRDXpuTf9BxUl7M
R5lWjtFuCkp8BuygRKRCgoIzE5WE00Vf2CTd1dNTLYodI542v1vrb02SpX2kQuOuTBW9OpV5i8YW
MOqlZ9PyEXOQz2VFz4S6woLxGf5l7KR8/SsyickoyfsqZik2h3IwuWUW0rSwA43EKs2H0oBxRRsW
3PAsaFcHuRVzIamzaraIiepNw1JL52Y+BA4+75JT+ccbJnuy6O5MRYQQNXDnhLXO1dAcju9qTszn
UZ0zNTWVU2IY8Gk5BDEv0Kd692GnNDRl+GhJuJeTkILZj0cJ079nVFI0VRVyKtspY+m61wl1u53V
SEcCh6aU5PA9YKad1wi3YyHXlkir9QNBOkoaMXf8N2RIRVEOS4gGuJherR9gpHf3YUzu7oB2L+pn
Q01rPHCh6NyiLIwwkny6CdNn1ETa8vDxSMJ9sw3cRt07dCxdJdY7eDsKIYlAWMhSPyo4RPnsuCn4
ytTxYd4O3Y/n/l0UVzbn0/RpzmSPfkDiduMnu17j/tZd1NY94yD9rnp8eUoHAift8ZwBLwRafokC
VV7O1ZIB1fIJsZ1A2jmM/RNev1yBgW0DKc0lZVRoj4fVzrquyy9/1iZF4SsjGg1vGMoY2NurzSgt
dnYdanoc/CVGnUg/qV9JNxLoc2nS6P+md5R7LSU26+f8JBfqnHCikvmryZLA2LQM7VnDGrxmtXk5
jUVn3tWJUEXk1fwREvQGeH9UJ9mUPT4DvI238/T/fJMr8om1BLiABqUKeIcoXqwMY0Qv1PQKTU4i
VdaGNvkL8DUC0M6hRPgbLJmxSFzoPX90AD7nsVr7x57gyC6uvQ1zmxF5ck2Tqzxr4SIZ1NOh4wfB
NDrVkesm8R/HqURkBk/ekunuSLHRAST+A1w7R2JMtxZJkqVCRI6OYjQEM9kEGHHZkhE1MpGmKoOX
nbh+9UvUZ3o4eMVr5mjfqNDh7tU3OzXlN0tHTELhteKxwDAL6AxnZbg+o0qP509RRFfLWTyouxhG
RWK7F2O5i5f2ub+hEauIsQdO2mSnOTYHGMnrOijyE3NsOnn7LhRHIyks9WD7srXUg2OfvOoPtPv3
yTTbz10xbAhaZZ3GorqsW5C0o93PsTM+s2Pbprio5UN0QNbXbBTU7pj698gHjsp25SF1F51iabHp
ut/9H8taBn2zifhSThzNnFoQsbaRQvmRzy5iqtSYheBa4zrQwXDrTozJjzrLSKXpr37w0XpUJIoL
jyUl2p13UgQnbiu6QBHfjg2JFyYWpVvW7udOm7WxyVAr8VZu46Qdf2zIAo4BBlsOS/Ytoc6MYD9R
oMgxWyebAM+dswRLrJayaLjtFv7oOeI1b619O04VX1FsZvnTxs/WvuT146XhRVV4sMI8FhmaJnr/
SWlDxxf90u0T9etQhP2/JACADqdECS3yUp+QzqSAk6j/VNlj5ZCvS0HQloxE86RfkvrNwOBuRatu
Sgpe/f6vbtzvkHyvx1i4f1wG0hJOT7kuhMAIN3Km/J3uB1ycpwVrU2aXTuVbOPueOJBqYxeI5AZ8
+S9Vfgs7hxCNo7Qs4DYLo4oT8p5OT204PDA/slZUChEfWuFNe5uIlhYlTLxY7C4rG069GlR+tmbd
OP3/3HBSAKOe8GXRu3b/E9RftXhK6/3WJa8lKdyCKepXXMiR51xbp9kPRXTm+Ih1MiVn+j1rBjZ+
5KYJwdpTqQbBGjfC4TjVqM+iczUdxBpDeLCmqiDgqXYPLLmIqRM7YENB9EG5HNSZRCZfs0B28vjn
6egKaFi98rfvlfIxPh77jtsm0WWMwrl6fU7jnj3crtLkI7MAwoTkWZT8Rk1Cy0FheGnicKFBvXNj
qTRZdUO8+vKss+4D3hSK0OG5I2sql05+SBVMWYIOoz9LkpCLPKUxzHQhd0Y1k5ZCaGYx7xjHqWuN
Ts6wk+bQHZA4I2z5uViDs6bzBzf3/3uCVqf0P+6c/hWStgj3LowzgHNGvy9vJbx9GLM8ouHaHyXn
DtYAo+F/10kkCnLSjluLa5Yu2Ch5Rf2CzLo8D92j2G7lOnKKGbkPuK8gri61vlz9+h0jfcLbVPLJ
ZGY1I0IU061VmOF78RmHLjhs/pozKAee79RFGF6aw7XuXuSa54MWqPOLOZbQqVEoBMUnHJeg8rlJ
hI91S9wyMuKOCjMGHsdT4K98TmQjwZRpBRMMxXrdw13KWInasrtkjIEq3+5vt0YMCC0YGMb2JqI+
NDHBWs0WA2XT9F/qQ56U/FwAiByvg90qCa6qI4VeBuiv5ZcgUKK+Ox0uowErbrkYuhpIAaKcnd6S
kI7NEVeI/ogY/RQ326IyciHmuasM3Z+iQZiQcfzhtr5XVGHLSeXoeWO0vpZQPRF5U5aXuolOUDj2
2ev7siul9sWu7BWkLhb9dVrDTSSVs/9q8HzqmmyAntkNEI+PUVWpbtt6b9hQzFgU4xmzjG4UvOKR
bY+sWfpiqGplQ5eMca5Q013TH4ldVwK+5IfkhOijVsQ6oCn3q6luiLnyclSSM8vf/9VPm/1xqUHf
XFLJmVbRFoBI1r6DCrV4/j4dQyjiuedkeNP48tlU9xT/VcpE9+yVvc/OlpG4ZGpncSle4Er5dyOv
gYJBeUYz5hDKzCyc7xDENIZwWl7SJp5YwmthLzj7GbGx7wCT6Pfrccw5+otYpLxDivz5Y2BYIrG+
44S3a5ybD0lMbzaaBMpFMRdFLAhUa3qhyYy6c9r65FHe7mXAPxb23fPrlIWdgLQZCrnqKMD4eA8C
XOsfchn9kmMMceEB6OmmSHnnIUllMwjyxneOy76xr2eFzS7aUNS3sCNMHF33o3/ksOOpXfu7ZTmT
amvJoa4kiukdHYvY6Y2ZQHeJV7cAs35uMgRmf4NvgtsjFOIaFdjFliEZPAeE2JYdPAz7UKnhjWTo
02iMliQTvjoI5fSvbSYJ/gpyWh/a2hllBdn2UE0nSe5k1QKGFW0ZiCA5KxwNaYaKVorgkiIB/RXQ
9C9tw7X2o7AX8JwjQRPb+hJr8CKEX4SEVueWugeyWsz04nah2L/FoW7K51QW34RnY9PMG4vn1fAR
RbIPkZgPKXqopjN0YvyUl6quLiQTvRc8BQWwy7AlvKYfP8NqfKM1B+CRcnG+U3PtjeRemFnRemKA
nzXBSWOa7BqddF5ZwYbJIHN4B7ErFU+RKjODm79yfK/6892AHiGwIgQMDSLdD1n+iKwEvPf+sqvV
AiLIkn80+WHmwqeE8txooj4Hz1QuZuLMW4WRisXW0MuWPE5cv0A93C4p/KtE4zaqxSyk9PWH6q56
WIf/HcgClYSrotmJFX2UgXSWqTU3+pdSKpHbR3F1Il0bK9MEofPzYTxVatD7RO0jyOzi9TyiTxhs
ChQlmjr2KMFqYcb3zligvAXXTMXhkuDJ53E4sZObFNRk3mR0I8Kq6L30JAqJjGuk1N6F6+49Gyzs
0Tfx/G9UaShS5WnVm2EWDKI/r/Pfu/EXPXHZRBRGEK1+b8LKQHXXRqwpCq0f2VDE9VAQ99wThDWK
yOvI8BOD6fYqTlUkdSEDb+1p/S0Sl/XyXiz5IZYEtY67SIkgdNkN544CCEB3xv9Elt/KtlhZKvqn
TZld4wlddxgfJ9lPW6t3aX2XMpzDpss8bPU52VwDUpFOtUlRuzLCLhipiLajLC17UT6glA4PfRSO
pjqyl4Y6HSgkGzzjItg5UlKSsfzgcJ++leOvJTuSVCziZxhjirp0qltQuu6n7Ksir38tqJJDnamw
xdsTWJSUFHRddDrQM7NNhtiV89YtFH5Oq0NWt/6dXHYyAJDW6IyLe4+1BT1I5EmWnZMuvPRUSlgg
DkPp+6bMK9TKwRa+b2qXU02G9+b2k+hUR1qhoyicGBtRfneHtCi8AeIjqvqYQnmEDe0E/7v8eEL5
J0sTGa5Kclw/N+6dWddciwdiTi8vQTwcJri1dWcov99mt8Y5GeUNvOrfQbeUyuB9C/kUwTKXukrH
9iXRkQcjmz8pgAxrv1jFNFqQT7C+jEemFsV2F8BaaAcunHHFrllQaIWTyWPDngEB9rnYuaS97cSB
dHvZlEIOFbX9RcmVucQbWGou5aNGG0YLpz7Xfs9JVsyyxH6qj/yxsnCXdzPd1YI5uEBBomw2Q7EJ
RskoRkpo1O9Rh2BXSCGlpgxQ339sd0GoeYxkM7MBe3uAxjGE7s19c8f4vBavsbc8lZwl9x7N1xg7
nCaQGcWJoty1hBtzyeMkcwQDRfikhjey81D3r40ABcpOJ8UefLbzNaTIDd5Y4pPOfiTTA+tQgAKk
+SZbD3+M+F1SFNobVI3JPhJLec++ndsXBTZKlAQmPYxfH1jd8zN1/w0czqcEGm/ngNzWcF++PyRs
mBpWox4mOYCyGIJXoYfF8Z1pKoGYFeK/T8Bbv84/xPUR8mDhlngYMrdHELV605UQbDrtlSGVsQz7
7hwc6G/WOxip5zSJsOu9M9aTz+s/tAwMk1SNemxPIQ6GY6Nz3QiUyZKQUzvqQpkMSGidM4S0nBZu
As7/L7mao2jEVTq8AnXMY3JaKs+3dQMrDtsFDo+2zybVObNNF+HC/tcjPRl0jjk+7coRcCrSWMaV
g0/WymbVgD/SCAXDZds12YXlHRSfWSO+LrAVFCuW8eQf27fpwGKPanZZwcwJS56XdNQOmyxnvqNM
+tXneJZcCmZyMy3eIMtsTDIlOU/SZ9v0rl7hXrO3ZUyruJ/IDdtD6SXc7rYbNbFaQGGhsLnruIDI
av4BD0L4L2+9VnylsVboOStO/GhTh9Zelt2Fd1VdXhShBEb+ItjVRhPtsPkImw9CchBsYrZL42Po
EjsilrjwxcgnZEDyfOF3KYjb+sHbhLBiLJO6Zrz9nSat792yWJ7zsiRgsoCMkTZL9bODctxCHDVE
rZWCkAmp03aZl/vyQ6KQGuSkCiX1gNmrFoxG6e6w3XwYJGcXeW0zItOI6qDCMgqR5GlApIryVKkk
erq+g4pqG8uw1qy4+/SN6bOr+FEhTwOb7rQdgAPcQck5f3vKsg0dwhQ6606uuMMFB7I5PeyC9+V3
wA7qYJs0hfSzZX2nHi88gmHBo/R9hNYCZ8NqTfipn5LMmPBD/n3YfwfctVmAP9zNFiKkOOjUxucl
lRMtlc0FPY2RtlRhFeHwEegtbiF8FGzqUPeP0uHfGIDwpEDeTfyCLD/T65R7konF0OzF2x1Zw4oj
z3QkOc3eOqh0CPN8kmd1WIdIt78RdAGYHk2CCilXzAms2JAUcHlgPVgFxMOz9xZJkmITJ38qB2vc
xytfWE1CeWmrlw+l7IGOz8B4ih5g8USLE5zDL864CIuVx0cGCPsTnP2TAriUST2JcD12mclBKgfs
kh1lv+OvMXwsTFw2QK4CoLxaBtI0RNgvN0esAzjT6dcsmYl69YFW8j3BpyXNik2/sUaIjfsKWbDy
zFF1bCfmWY4xDw7aQ+bq35BXgMBO4LddvKEfxdwoEQCEkNCaUltrBqelKw39bmXSJPU4EqQ9cSol
7EVm4bACz2RUvoQcujKD9DjZEY5tppvCqb2QJUAZ56ORv+Lw80KzsY+BC72IudTTHWIGe0b/STfU
B3ZutjGHfjOzeUJJ/nwCGevqtB9uiu7J+fMw7u2Uj5Z0UwcTeQcFlp9Ey7cnU/x3npZkYKU4XZHH
9mpgqq1SCN9Ikb+NrOhh+Btmstz3+ud6p38Wvbfcgr8brJaqQmfexH2AED7M7aqjGo+pD7/73WXQ
3oAu0prwtT5/rlOD6Gbkhs3oPJUlQkx0FelF2Tmwq4voWxyY94DAw6XRZpoMyr9vFDqU9b/abww4
J6JEIbG+cFDEzeTOxQ7dQpST+nifC9ihdWgzdFoMmqhnPTSkPfOj1LBCyg0UuNJrXwtOVAIFZPPM
Kq1k5wiPscJN5etJzsuvHxpyzG+KQK3nyddGavNCZkks2pkTSOUjN3FA7KESoJH4YOw/uMTw5HPm
G2/7f+AXN09KYwKPbiz0YOnaW96EB9St7yqIxLmEqfTz+zGBI9WSdmbi4VXVA3Mkx9LcyqqPgqC+
y5HaVyQR6kyxdjNLH4SfdW2ws6bJ87EA1641EqbaGZTwkjpiARrRfPuDUy4VKhxbPoLpCuBJ57Ow
4zYodVKS3/8J9pkXpIqf04Eit3ENKIfjZotTAKZri36DR9rksjWKnVcuTn5dTx3cOMl98+78xmwX
qxA7pa2uYV+3f+GMWWb76yAOc0cQd6OstJO/ZD7Im4SIoZ/UzFqXlktqjqPvQVkior6hkrBRmLe9
QF60Yuc0Vm13n3ig7FIdtDasBEp36sGb5TOkM3kyVjmZWaRCMevas71OvLiW9rKhdWfBON+Fh/6H
vNNPHWCTdCuW7R/N+MqJK8RYM3sHR7XhRuBEhgGpSPEkioir3QwmeKC1SUpxog/ugaHWw2vPvvvB
/oP1BQZCdWHhhAFXO6REj8GSs/l42AI1oUL0183unbdirQTbRFEz6OK7TZekCn+AQHAlHkBVx6wd
1S7WQBOy3Ew6gcl1q4KxMe16tuWtu6cFFbfkSSPY7+ulKLXoCWEW8L8ipM+1yrvfpL/3kZIPlWyc
D7+3kPbI11V0nifiOOBlmN356DjCWv2E5lhSySJHK/lKDfmYqhBiKkaR2nPlhBcjbv0JaVVH2Rhq
XQobKHVbDqKU9TRKQpKHsYhqS9OKfd9PVNgAjZrEL1xNgfIWesSauEVkdD+fF+E0TLZd+lzF+VWZ
1W3ymIAowe9Fd1yrc05S0oXSSOhP/DDF4EUPMNBKM1VDCHkdLRBLoYLHKykjU5qGp8PnAVE9wlo3
FQ9JxDDnXrx2GUNLJ27D1s1VfYwqdBFcUjrEWjiYjhKOCIJIwCQLeK2zEnK98pXTNDyCAQmbrx1C
PNYrqNGrCYqi53uRZMenD53s43nrBy/9Q+W7p28K/rN/I0ctUY4toMiyq5U2rBVicSBCeaHW5HWp
8abBG+5FWmmDDflnESsHh5cGr7BKjix3LJI1jTp8iOb9qbCVN4FEjywdWc2fPnrE4vG0DaXJQXmF
TqXFiBLsW+Bug/JSoWz7RhfwWQHlpOJUddE3wOtEwQnDvQbF919MqDXdAIPR+8hJfrOPVbeDa75R
yYDUpr67eZ5ysnNtt7uxMxt1v7/dOMysNhuAIBgDYUHY9QpjHe4HAraj4gopcTd7wo49G8O2OA8b
fJIZRK2QDd8NqioMArrJ2UevzIwo8IfxGlZSkYWYjyuQjCJaXCfjVbiS9muK1s7CEFfGIoq7wIUc
308PW04sM/ETo/mRZncPnJvZ0SO6Lh+JYEy1ZcoQ3Ms+O4ickM/y/sazCmQl2C+0zS/X8ZEcsZHO
0WTVMTznLuYlYTooDMMMNlp9SVXf3Nhrx1H0BvG/MyRGdoUxyHaOW2wLKGHpbnLJTeXi0lko+6U1
6v1j87I1p+npPQGl5+DBDNzCC5fUzAglx7z82XpGZEcH8QoYqDUjFrgqB5hnYJaruRO8/JYbQeob
Rp/Pyc2vJMzu1KUVMHggl1ikAdUd+6EgPVCbkwIJ/wXazovN80GawjD/XVCgyqOsjMThZMjCF3ST
txl3g0fe94C0VKqmjONrnAZb8apGtN/XKC6VOYsxmmhhPuKMoOAKXfgookHzQQ4kWq+KsA7qYXam
g5nH6e9pbk3pxKgkYiI+ZI5Ax/ZV503NlrjRABMX7PJ+da1Jic/utXONsASFabMOZiPpdu6Tvrh0
cggA8lKCB+qxBk41u8n/Qu3TcvyCAE41jnUIdhsKBNUlRPOd0hDOiM4HC885/mfAdfRzcBj17d+l
erHQeGxF6keBtulqoUMiviqe89NZ8vtEoWEFrF6exiMqzbkzv1tGf6VmrzFLIviLSO3aTscLEeZZ
6aWVmLjR7lYRNRNcFq/b3NAdqQSYV4sLHBskd/mVONRwO8BKKxmvMc/v4WRWT/d3NHvhs+gGl7OU
12Nsw0kcWFij6v2CXIrJEDXD9nluc0+qCQIueWx/CZQOv+K8w+SRgUvf6yeRFIqlzteD1TT/F2QT
wTGH3dhL7+aVfoGUo4tJSA3kyjkBWhU79FPhSfxwbKp0YQL8VsCOOTtF063TX15Wk6BrJOaMIDDY
2u0SyfeR/41GR5ULU0ILGppVuoekG+qN1MhfLyKCuUatEbjWBzPNwdtfNpJ383t9G4xVJsc+jWYU
Qbhq/MdK7yPskdT+ofkE+XxZD1R0/S2ZCyzVhpRukEJJzRg3M8XqgxSW5aItoZlwQP/abkhNSMI+
Vyhaa8xZXRX+2QMfXnbcSx7QR2dfnSsqwWtAzbzRifK62A6nLMvxBhZAkyPVnYAbvd71nkCTHR5a
tVz9wwcAzThp99vXiWgF2FpkWnuaV3wf0eFGc/Tk7dVG17Ab/w98W/UPplfh6RJInIIunbtpHH2T
Gxx5r9YYsXA/OtB1JiIu+ZiJh0QQgUEggoX66IOeZS7mTKCpjbBA2TE7++vxWv+eY6wfsGeQqxDh
0B4T4/kqupEe1Ei8r783QQWbwejcjBy+4xs5KbpBtPEnFhyN85fNHagtN4wBeoQ7K12lmiuxc/Ss
r/3IuYewk3TlD1ekBqSxBBsrLySSmGfalOFmzPFRxk8INA8vmSOROLgtkX+Q90cYQBJUIoqA2vo8
+IHJe/W+pIDqbCyrSbSd2CIrSCsge7j1EFGVjT0eLlKYnE3qv6BXpQDzGFUuBH2vPFTrEsFNFhJf
ZduSBFuTQZOutNmI36ZpxOUO5u5a+3vFnongD853hf7NFys3SSBgiTtBWNyMBYBZANqbqRM4JqgI
D+XLMd10oDznc8cDNVtiTPAO0Tx83xquth4ueDJnmikN99H4CQxdFc3oEVmqqws8O8rt09YJVqAx
Op1nsQatZQmk0wt28EmHE/QVGc2xzCrT1vLIslVz2FKw/o8HDCnlOZRd2SuoYETLuG4kp9jQ+prD
icGp96eg4mNH8S8nUWgUs+BwE8hbNyAipCGib2Kw8uNExpLXMB8mICQpHgP2nsrqFj6bnITdQbXr
OlK+4Du/HsyYr8/Xo826mwox98d7vVDao6DBNFncIKqb6pyKMURPUnrj68AaPY9Z7tkUsQFf2ziC
APjX5loECadz1LahKfuYdjeJm4xuuAQu9YprDdqHG62qrwUVtitPUli6xFwS+AUuW7FzcKxgTUx1
XyE5slA4K1NXwWsBC4T3CaWMMvhNDLKv3R1yLiLZ9JcZPUTFrNaTh9scxHL5U3+G/H5WzzpMv15g
5evs4nlZ1Wpm/YhnuQFrLxzEZSMuKbLMU/OmAdpIbFjGuXdVVgj6r5uMR+gsv/RwNuWTe3BDrPxl
V619ZVLaUOHY24rxL8ngkn53pH0gopsU2bkitzkHjBKeIjNGVA/kEyLzdqqIhOif9/gahStoSdf/
HvAPFg4Tc+V9jRBOLPNYMeX8DPEInLMy4gEXE67/Tr6silROsydF0LcuAEnCgXHbJ/NlE1QnnIJs
d64A9Z6b1Pnz4HrAKFwbbMRwaTDmtPEREhEpVtOgHsAYPaO0cgD4pQgpJGNX8SOYs1YLsc/RAHI+
90ETI41o7dhMSPyGJCaNrU7DbkCU3yZqkUSAv489uFqRbzlPqPJzt15puVAUP6zwDVfukf525teF
iddejq4mpMyEcQpqxxwY3wKegB4+MhNUgq5m6/bIa3SRhIHKNr3Dy7mrhAwF0cGQnKX29pVBvW1R
pFosevor7wKFdXknJy4NiX//6tbU9k1/5rrjnMiDjkJQspanVAFXQWRzp9arm/KGYd6QfF5rd4Zw
tNBe3YIyRqSAXx/AQ3wYt2jwfW5NdtDr83uVZRP/2N3fYY+LAgC9NpcLQ4toF5J1MenN+E/FdH+6
DBcbErR7l/0NQXiKKPmpIXdYyD2pNg32yrcom7C3xlAkDnuYBpnrsL1MiBJFgFm2X5U/ibOFicUf
jmMbqB/b9qK5n17aGnJmZNlt3Ezc+VleMSt/R3zktw0rj5BxSaG99qs7h/e94pAbfNerL81B4VrO
jcjOrV594wxQPxtx6fZjxnQFlWoDVoNOyZclySQAceWfwK1ww8fvBJjqb5UOv7wVW/3SOJREDsQw
Xw2/DUdEz5/TDZezniAzV5jX9FOcjjo6EUF1/w/GBFT71Q+9nKdajGV+rqo9m8myhFz6jXFNrtJd
+BiEnkZerCHo6JQkpd1Y7bs0aJYNKH3+UJxVjgBC2IfhqHPMFbD11vIUT0Oy0dn4nQlRhVQ2T9YB
c+axCwgWxK4UzMgGTsfua9+Ywx1+kGD7cAHv2it9cywg86CMu/Wx/AE1AdxBAknFex0XKnVE7G13
DCYuyOsSl5nV0Mtj13MPeq1ejqlHnA4eAOJJFcCoDy3qMAmn50H2EY+ScVn/yKvYBdtzbyGtT1Og
nTR/5Bmcw04uAwhuSZZQaCSuSrkDtdmflEzwX2s7J9jTooI2Re2Zc0jNFpMiDlnUbxONW5F7oUjC
HLgKxMtxwNEMl2ipr8oJZAcVMKafo7LabACkuMiYMqdizvPD97lKqmKa7tVUdariF9oX6GxMl9Ni
tLsgs3XjcANPJ0LcfDNry/XD3KHBtpm2Gp1EERfNqOYVaFhR1vb3Vwuhb4zzzpuzIRxliqyAhi9n
4UL4xZ+WwjJ1k8YRiliBF4JvTfj44VbUA8rZGxr2MMARIwlyAu8469z0pnUThJdhdOhEw5dh1gaz
72XjVnuad1lyBx4vgBriThTGfUUOs3kQ77CGVmSMTyTewHHyVQ2lv76qQeqMEXDRAt+jBHnci8T0
su+doBofVpZ/WSiqWUdG0angbt03Szm8cApUZzaAYN3fFXHOfTFK5JTL0zwMNgMs8xYM6viYd6Rc
rW61Fu1BzYmH1kPm/5byFvp5pPcs/Ux+RR/rn61f1WVzmXLWIKa/PpVvh1lX/IoKKaZWWAVWkdUr
Gncrcp2jCcXlKUxIdp4VQA+8+kLsyxJAKYIQXyAQ/ni6jw+Fp/+bUVzHUuwXhw2Z85Q9+pBvHWuW
uFKhMTNSI/garpsu97QjG9egiCtB4si7FuUM+9fu55wlcIi0Qub+i+k92z/7yDYQqG3AOL/0gM3U
/uNFHviEKUT143tkKM8rPwdH3pdkV1tCh2f/t/JhL7ND4D0gsEiTovSWmEn2M6UbWQfEwvZg3Pp1
E8K6+eobWdi3qveA+UzMgzmb+fchpvTaWZZELeiDH+7UpZEQz54VPge5geVJaaMB3SB+NacAQaAm
U2eNHpgzDYOHEK3qWV6z+92xNW8XaSIZJ3QpxLtOzofhYmx70BFwhI2JCn+yYQESv2lfa484C835
KUmYbufXXdX4gRjdP2Lo5FsKiRjQuuLiFdEo66OmSpK7PfaXPPOG3uSOzpJ5DBcS+uEHAadgHsVo
VG71oq5ap2G9xL+FpLaG5agXdXUySJK3ryvNa+HLrva8rvLk+Xqe3RgF6N6YcMR7fklJpPABX4hR
3FywiNUDOyyLn3KEQ8TLUwiTUOCrAu2srskQ+iI06f3fyA+Byepvfcnrbwb+WfReszeiWjNTfCFa
oxajEpbwzSP04v6Bno8QDsG3xv4E1FEXJE87pIOlXBrsEkjAXRAI+5ZXhsMS+KVuNYB1WU1a4GhJ
LiVE7rH6mCM4ZPnuW06xrVjkPG74gZIXWEefW+12xn0oElakUazOhov/ZwJqqERx/o92mVEqJHB9
qi1KCOvSzl74Fv5yOhIip+Wd8LgQCW2xiH2br93LT/8HvUl/aZ7TrpIdBj8+FjFK1JA/gk5n1zPt
JktsdF6utc3S8bt8U2OB0FPe6iWfEs/lIa+MrFUNP1iz8lqlcvmb8G+h763D21tT3+ZzLjbjRI1r
TsOyqwWUgDsJe3tsLsRpxpC8CWpBWq4VcoP+lqCY9dAeiYN5g7bPt9OhknehLqkUWckqK4kuZSrH
EwffLUc2wHKFNCu0lWNUXvjc1W1vl+/XhoRZXbO8H3zuth1Smspel60XrPWRIvXp7EkFgC14dc/2
O8tH0lNAtgrD84zHllIkApoOARQ2rMxyPLjBJIQ0Dppuv90CTjc+/kOzMcgo8DY50Nw1nu1Js8lw
hFcOOkbzK33svYstOwMQpsUZZKaLBdjXSxmjIz7hFypM5APfVOJvA8lqzVpl0fnztS2Ohkj1Njru
H44Lfmyz6jV4en1hntnrkImUrzw51jMpevQJ+Fgm1qYv6b8tS04ytYLYPsI+8+NhORzjGApJQt+H
6KngDhcakiUCHzB/7MLqFaOSntaZl1Yc/pYqcrfwpOrqMRUDxBlJBY7iE/Toa7GNV0BSJ/V4O240
95/JKHd7TJZqnKO2+7PzyNfayPCuO00slsK04iGIR8o92x02lPxColu79Tdi3sj14TGf9kDjjmQJ
yVit5lebPsYryKOIsfdDiCfzHXHTQP44o6LNA4MnQDoCt+c9Pfj6FGIc5BkCUNCuidhWNJkezKED
9yi0EcnYqV99b3Kx55WIJ8FULxM/lwWzWInB2pnBrNQgh44IX8ipaZTricH6ZkOjjmfyA4IxVf+6
KW3cvh6eqCrimBNFhbhsvSpZkoF+KE2/pcSvem+chGdI0oZAcyOKjZkfc4gd76xICycmfVbyu6Ul
S87FfUauEw1L35bxhdoTMR7l7CKH79E3DokZEORy//vf4hrjuQFCA4FNA+BnfTT5yfdOrG3+Cdf+
hqUgL+C02uO+PR08GfkLFNq3PfdTZzIagAqub/ry2ZVMZ7gM0EEfiemtKlAM7jPHSdmBVDPTsKle
YaZErD0I/h9W9ua/jRJQVLnW4bCrO1B8cSQn45ElRUsoqDk2PXMlqWj7RkWVwL5ICyptcOgJDhwn
dNx5M7xrNPG8ODHGZmAwUqpmN5lAVZ18zY51IBG+oTsWcVwQSBsc3JJuLRsh4xQQ+HW9RA8dHR07
fWXNOyZ2vDWPh4QXwbtojE+Pg3SZuu0JayGPgnkK4D5KinWHimkZ/jZz8+bEzkCoaR/1S7j1wKPO
3CpowMEsM0BmJs1WtycPwctrVTBIAq8nmvW5O9hHZYl2hRXEcDbx6T9HtSq2KqCDi6aNviaTjbkC
GYUyAm4xr4ZHIalTEaUQoDUhcnfhjVv68Y7Od71FN//JlXy3DihTwcZ+9KqcbKiuO0SLKQI8h5CI
xNo94jh0cImc4Ywyxk0qiwodUdK+2MvFnwTc5bF4jZ6sNED50OR4WvI6/o0LJ7LSlddTJjqOnW2z
JJvVh4CFNIHp1hn8Rj9mc5+AUAjSbX8MURitGe0vSoLhLdasBRmo5hOl0Lg02p+L3bFTWDDPCp6p
wD73KUTFpZPFA8WU+q9Fb2BGJonB7V/Zvr1z3iyR5sQw7ctIw04CFu3PsSs94MnWDzh/sBI5zZqm
Z/wP5m4jua4rBZCdDeiA7mVQR29T1EvciW2uCrW1QFf4I4DsDYYLWSRcxPUL9pjsG4iEw5xvR42S
jCLztusJWY0Z0/7b4tG5OVmqFlZjb8E23yJEaUzkZ1u6wjzrEVyEVU0QkTCM0dxzarX1LO2coGck
IHknXzl/EmtPmkiay2cysvYBvo5kb7Jlc3QzvtKC2s8fElWR9loX4NauyJkaV/j1gTzWH+hd9t5N
hhmfOQlmDUxj8qzX2Sl8znV7qzd+pT8Wb6xdAAnFz1RiYa9Df4lUv9ZM4PsmTUzAIgVfGLNSBWP6
TrGDuVMm0q7BzB1IqMKUAYv1HeF+9NJegYYjmpIBADYK2rZcHoUSroO5yQU99YOt778bCakCBoTX
IgJk/C1DKWLJlQ0m6K+PT9C9fXDp4ofTDlkxCWCyMbTtwY/sjVM3jPxlveqJmYXGsLUZKLkkuwGF
2BQtMb0g1IopsACtQgLub519aVbIhUgGgFUD0IVGHqjIAEh1Yu5/8uhIhYPzJ1UAAKeW3zUloJcD
x1DULxmO7fNw7HP8zW87eaQJEG0SEP+Nv9WI78XyGLg7JG+Li4CFmyKg48KzlSi5wXNcHoMwdGni
yoVm7hKoxQ0tlSPruvUX9q6+Q/X+rt50GuRvzWZwuFqTiBbWTa7rNEer5nH+MNekSWtY4XbihNNh
yg0vkrh2XHZ5pkdjKlS1r2k5LPc7NEm2O+S3A1ok7EI3j7GGFchT/P3eH9K4RJeInTeQ7RYtRdFF
EkigX0xehcUOtJ0yYHxE5Ygu02L1xraikUlcEIVKeQhtdesAU1QY0TrjWdvo2DP8lCGenztvOIpf
PkyvLP65JqeUG/Zz+zCKfAo+BuJHBOroCjwjQR/bnf++aOB757QksIyscR3WWnS5ULNdijayJ+kf
3DmaH8qiFPBw8Klf04w5E+8zgBDRiX+ZYeMkqzjpm1MqPsQ01IyNIE2T2AHs8ZWqbcm+vfvG5hlw
fumOEDoz1X4qlvF605JfrS7x68ssBIcbUahT6fC3BAZVt0rthld7SWTbkN6+AqefGb1B8NtQUPqJ
JnKnuEzT4lwX18tdotyBZjjc3UPh/RM55dJQ8VAVJ/meCmUYeJCQSs3rqFBNGa9UY91lltASAX7T
veihN9NWgnXQCH1j2GCO81at/doE4dBqUL8X/GFAbtC0WObb3/RksRKk1jPt7XfOXmdZr9zfDCTQ
RBdmqFmzfd1GBZBW5gIPhdHyIdqCM2VF5PTvKiKsNotpZY/mZiooRkjt6LneJ+GeZlJK25vSY7/b
+4009fzeI7/MiEwBDBLO9SFePGhzA9nW/iOy/byJd6p41fpKk1epy4W1p2Rlco1ifTQtfG102NZq
VvBA5/3tToBRpaxvOh4Su4PsetKSUt7ePILAOi125469dc0Nty6EX0KIABAmZTkmCoYTjqDEUZba
g87WV4SIfELMfRD/Z9p9HcPeJN+1onRoh53Z7+NNBA5qTywr0r/7P/AhBW9e4JjJQqisAzdTKt/1
Ikv+EoCoAB6Ynuy146E6XaNYie4nlzFtd+Exofn3KUDKU9AQ50qM9ob8kon78D1dSOVEZq5eVPtT
B6vetKIRF4JMjDsthCaUcI8FsAoTh+vJTvz+3HuralcP6A4m3Jit2tHhe+XGdr2rh8N3IQws+gkz
tFPyT4RyQNcHg0D11FadBPQBGBXnVEllunsZHxJvX6wGCi1yB2BKGJJxTlRGdI3XUdbJnnOuEFUA
66JR9I98m71NwvqhgsAELHoy9h/tq67Dl99I8NmIlqeCF/Ic+GOqcsq8vjxckbLIuhjYhDpj/E7d
QZsLpP70b34V6AoNLWsD7MGU4lUu/VObAarlLcpkp4RO5unCLMbH6ZJC/nK307D5Ei147J67NDze
dtTm4GkHmRXNbrb8GMq+ylWVcVwUboKrnfVO6nw6+YCO4kE1T5owERe9qgnaqGOrY0Gw/tjU67Pd
4lPoDW+mqSYPhX0rABN9ljfX6u53CW71/O7D5DkWPRSYo05RYo0yKQxXAnvgHkeFMWFwt3Ptg43V
ojbtzBqxTxfU5Fu9/BOP+kYw/31AhZ/MKC1hqHeSfUrHjROllW1f8Whsj5FKBeFRoRCumkgyKkhO
CcwAfVTdi1Kapya7nTMPgo0Igh+xwzOHy1La08DHXJV+mIcks32iy3ntU59tfmciB1cpDUlmcCIC
oBDIvWHpOsa16qnRlobF68gZ0AyW6n/5omjawU68AV0VgEfTeoQee0c3ufhwbOX9uIod83HYzeHu
PNSsXlszbGXM5C4NMar8lOhT7MYXUWAM8lN4wlysmVwRfzgFB7pFTJnh+E7xeE/Hh5bfRW2bNfTt
3hQWiwcpjCoGLWWLK2w9Ylp0KElsIrTiWkYDlGZLj2Uu0DYZqWQiBzI6K/WfmMJp8XlRMkUOfExz
r6bNPT+3wLP690NLzh3osbSql9bm1a1xWk2EXQZzktfaBwyr7LgMBiP07yW+LA96COHFw72Jq5AF
lXMXpm8uH05/I2OrUXipCqnqSEdkQ/BL7qwqdYqlBPPyMFzO55mAZhYZkFZwyly7GcN/Kjr6WL7A
lVOTLvS/qGbhv6w3kU1WZgBdhlXu7HDMZBLFpEXRQBGCSLikA+7OtZhIKx5p1LrCBsBy6NFqkK9t
6b0zpV4Y2yFEOg3twKBJza692BYbkvBufUk0tCrDdk7wqPXERAOYMkGNQJAuYlweoL+qYQsvTHN2
lsuroWiQoXlyE2ZT4KEtF8jDlCj1sy5urfwRDw5udt5r17Kme44WfbWWlUBwrHSCwShrkV7DGFlK
406No/MOTB3rsDkTSsj42RvSWef0f5jVure+GAbPHcl3Yi7SDfiLJGsk9WovSJonnW6mXISKR1Gk
hY41pJSN7CARGc+LS5mXNijm2AOt6i6eL9K9/xpDbxdZH5kxpmH8hN2VbL0H8CSU/jBaUKL6Zl0R
dnWYhTr0zjsiOSr40yW/p1uMDIPDp/WnhWuSV/I3jKUg9KVWQL4dEgOgrA8pKLexRKP43CVB/X3M
I8Z6oU2f0CN4WRyZQDOPimP4ViqxmPzvq8ylKVzmtkFYXA3qkpvWsW3YNahx+Q30aWD+9jAZ9H8W
E6pLpFsuEJYwDH4NUWAfx20YLD83RbAwP86buWEHGgTHt5Yb2GTFOzcxx6XnvCO8HwEWH4DmiUyU
wGhm4CBa2UiL7By0dTF9doCjHdGhRa0fXscwvON5IcdqtQc9yvVXL1XdxSHNdPCHct2rTz6wNoKZ
FFfMv/uhsfbNS3+hHh5HyCqxplFHaZ+OxAVBHlNTh0OOx9p6iueX8QHGhPBhNLXLERCmb+nggFv0
3PWHN2ISiLbi7ANROI3Q0GA5hMiVuCpyVMiqFGeD87S/kms9GinNmfnpzSP41oGnOMTShOQfSzlz
B2eYyHsW+MVDVdisDKHsyGaJ6dH4wSOvKQAiXhS4KswQawuTsvsaf2KPWXexCzyWXR/tr+goo2aB
22NO2zPY+MIa4RxXlNHqAOLdks2oAPcgyAsuAloEU0VFCenGkoFPI9cNyJB0DXuYzpObLNQkCG5V
GQPk2RrvFyLf2j1bT/QeDWELZHI2x23V2W8WEbcvEQV+uAXVOLeYfpb08qZLz4kS75KgGACX+clT
yyAc9pYU1jtH5wxlrM4MuOttbICxqKYTBdQ/MDkNqmAFqTNKfHNjBY181BJ5sXmK8eqP3uBD8Jj2
L5keL3DEyF5iPYiNqOlMoT57rQLCdQyyGrrPi9wtRer3403fzuyHaS4RPAtxsoiv2gbCNNtc8Oiv
c9Jzd5C5E3l6Z5gCdQG1KpYGrgO/t7FKMwboGLqroQX/4fP7fedxKtSl7KCmDdSfbS/H1Ysq4E4t
A1nzLJFbUWuU9owFHimnDIqpyD5AkwLrVUgb8j5BkUh0MZRxp4+zv31EFitVLIceOYzsQqoGpyI8
0GdcOb6UU8L3jE/hqybErLm/WmFWpMMMyEd9Sxra8SK8xU1ggEEN4p4ttD61zkWxUD/38ZPp0rRx
D4XdRRPKvpEUCdE3PfwYZTx6dtV+cAHgV1uTHQ/CK3Hgic2riAaQF7MI5TukwLsINXSfqA7DU7B/
E0kSH/l9G9vbcL2FUljcWv98yH3bV8u1js5Y6XgIjkcZys2mSo3IOwLTBj5JphBARJf9uxaX0qi6
XgpsT6os0oUWI6fLs+kyT6yoekrk2wZoVyyoDSfdoxl41WoRmkGV/6aoOSMTF+nsYsp07/4nwWVG
kRY+OTQE/hiCcj8ybtqNd8KKXOQsw9Js0UGRZa/jcncZUhEZA7UI+SQLZyLiHSW526NGjudbpSM0
6anRM5g7iGGpQxPvudWMJOLzWX0zQCdw7gO4l+AymjYFHMj9X4Dcba+v78qh/TTVzrNSRmOS/HDQ
Abj81gbFLk2Q57bFunqWUz7rxyzEMkniI6nU4IQ4/fUfTfdj2MNmWPfK5bWGIJRbM3Qjag2WMuUf
U/3uRZYvGi5Vg97+tDwMpWHl+plRfqA6ETqBUET+T/YVnf0gY0XslzyWqbrR5uuJGmaCN4WYp7gl
7b7POEJago8E3JGMOMIioFC7B14UEk8jp9a6PjONaxwoJ2jnfHD9m7W4K4xN1GVXQxaUpf5xBG3u
TDq4tFdH3FE4pN+mtAo7pmMQGPW0c6KY1v2pzdaKWVJ7HFe7PQLGEK0x6tYW7DGpogr99Do0O7jG
hTDs5+phtZOmK3VvWbzD4VTC1TMaZxY3e6hF2zT6bsff9PlPm0bPrbSO4vWhRy0d6Y2EOnJOhPvN
lj/U5ikXYzBg6A7AtsXpV+17X6l/2pY0ANLw//ja201QQYHR+yDXxdpMElPPy5EgVru7gOMkhSW2
51TJ9qyCZupMGQgGJfCmF+OgTSwsKc7FJ7bX4gPyOTVok8m7iAZtxqeoylHEYClEJAT0csVnIlI+
KzBnnWlynrYrK9D1+fBNFqZi6NCC4/XUOBjhWNwcdCWPTqmAyQGlWWYVYR/pWkjid7qkwGsPGxJC
2RE8cyGBnOO3keq1qfxtxCeR99Kt0N3ylbE9u8SyfrvilXkFwKsT63mS0eVfWIyUs+C8sHcpQRpl
VI3V7/zEUEKIRt3PtKb/wJyzBxRlpS+6Ryog0kmaCKdtih0gxNrF5gqRRSUrsE8jm7pEZ1NfMXQg
lSBRPp7mBZ1FI6ck6xXH4fwc9i2WkDXileadLFte+HbQAqxggfIN991E9FtrP8ef1o2b8aShIgm4
TTsJ9lMLiGBujH2ggQC1nmzZH4U18JNvFnO5TJhjNgrAViIl/Ldho1J/+imBLDAMWVSFsxVwsLcW
kH4H7GD0Thl48fP0+/UcgtkYuIVMp6PbXJqjmDMEtx4e5SWRAwoLCD6xW6QfhdgWyJFar+JjU8re
+i6e45EIYL1vd8MkM7qMPS9LprGwtAjGQ4yS5Q69c1XZs6FxMulHXGHE3/Io32WUbgBlZ1HJfzfZ
nyQvaJoLn820OCKuO90DKtvIDTR29Kies5rJW7GSN2mOwd5kL9REm+H/AC6XjdRqLN8cbYPOBp1z
6ExdL1ywsm1j5RO3pZN5cw/Orm6YTkphMy4W7+KK8lLjsue3vgmBqo1vzj1arCdjseAp5UAbEwaK
8JUYqoKlee5DheO9vFa5oc4Mnmr87MWTDidmBIw8ZeQvYLC9eP9193GQ1GxRJ9S+0V6WSKKTweWZ
K47yoZxNK8r8bDBGLYxe5f19bkLSA9TClDwCefKnCVcbkOsDZrxUfguvDD34VnrbaovwevYRTRNY
Z0pZwQOOlIVLdrdPVavr9h6PeU4n4Wy9XpA1YEWJNqIbZXSLYI35vsjMFL0Vx3hThbdxMp5kVVIz
b023fm5H/of2Eo33MqJdfvRMbB2EreGRuumWT8GXzTATFCQ/gqacmtolfbz2B7N6UxLWcg/3p4Os
sACoa8z/Tm606ZLojf1imJifnA+hym9Mo+cwlfWAdCijQow2vj6iwHre0FBXNawDmkmwEMeupYkH
CTAq2xDDZ/FEBd5cT87lR+QRiz227cmt/cOOG3o37k8Zayrr472HS52S7iI+N/CMTiFSlbCbj4OF
/Arjp6XLhhUN89ekVJbGREOKQczhTo2bS8wiWG2JiyRa4+AP7DE8A4yNY6FrmTBOpgBCNDK1q/F0
516JeDgtqksIKs3TvJ6g1nzvtqWKgFXtlxPpqLan2WD3Rto8/2zqp1u/xH6aZTMbcOYMp4A7I0BT
3RJUSfiuTSoGLQZ8M8ONwNmmC42Apcbsel9EjtL5X779twynDmZ/BLnuGWre18K7vlvAJCb0TYN2
Wyxm7DNpE7TZUDfh8XyWj0OdogYu461C0xG4z2tTvw/v8l1nc+mmkz88xF+/J91EKG4+hwmDRnzH
P+Q3FErA6W0AWXufyc/jRfZrW4qhC8fqlUg+N9ddMH2fe5k9lWHO/wja60D6zHTjXR8TXo6dLxl9
zNrZc3zH4nZw83DL5/jIk4X0JnF/NtezOewYfV7a58PV70StVTRdJyLGaX1BsStH2QHnBDw5fuu2
I0tlKocCNYvqirK4CQf9DSysEOrGeilD63j9n2puPbJwb+f1FKN2ac456S4VUg/M+jSza9Y1WXfJ
hZ1jKOTTTmOFjyVyUokMMUzzPotnpPmjGqrBFknEDuVnVDYU2NCieoWbQvSVHrisvh+gteY/LsuH
ZBjeoAE9F9+aX3dnBzSn1YQa40gGXwYASEPz/r1ZzWkQh3g/OfD0MLUte3TcE+xsB1SbP7yaQETn
kAIjudv7sJRHmX+f3/YlNl6ONaKrmRcn1SeuU0dEmm7OnRkeJozLbFuT5ynGEPtYxSDbJNxKvkn2
3SqZxek+CIRkoB+CK3Ez90Hz18ND4cJDE7em6qlJXkZPwbQFbzXNFR7pvjVeqmBkJ1PjeqYxGDQg
YhhFqX3XjbfdiutvNRqz4oX86e7U5uuvmjhC4GNc9j2HXqqbsJfKVTkPTLeguD3bMU+NTlihPBrU
AshayU2L5VIQhpyO3Tm4LsX18wX46rW3p6nhUs/YIWZoO0njY9hweVg3Nhb6mnY2vdDJf1iyYC5i
+frMp6VLezwjktU95SdJ7LOfSaV1muVhxlgWxqTBQlxf8rIs8GwLudoStnIH+mt+L969sNjSFNcP
i/aWFwjfuhlGD8Xr74bPEUDY2L0SpqkQoZKSman23lxKzHtyz1aP3FfKFxkFakWjMhNYr92+RWBX
UR7RYeZCQk/HJPcSavx9GI1ewap3uB8dQ9LV9+PPkwQDZmur1CVSp7+DkqFua+JrOi3LXOomX1Zz
kMbV7gUH+7Ozd4hFbxiAaj+3X6ENVBfxP0L81/niZP9oMGbVSanqL5GCcVbN8twHkNYvXyWZlhWw
K5j6Ftmv+ogs9djre/aPpcVHGPPCxEOEgRRr6fk9cYa7L0518FT+2WpRwsm6t+aJiKUAS0rHeLCT
cxvWYMwf/erFxIBHd8Mq4rW9MRUxs8r5D/oEB0e2ZgSl8rcckwspcAFApYbgPFqbWdWIyMR44E8m
pxeJGkcwt/FlXEn+SLvQjiuAVhL9UJwA5OPwpLp+JRdwEXroOdFR5R6KKWW44TcVIS9gSrnTjq35
DyHhk6jafFD1ECnJX76/shTcrs5POP0C9svSl1umwYBlCkNqMo1vK2tL8AmA2KKlCw6gqMV5fy5M
m4sdp42Wj72ptMHGXK+sNwDfQTycPu80ZFUffneo93DvqBpVnQirPJj/b++qA6xnw0z3BlZdLx/j
qPjTIsh6d5P7iZvNkolkoZ/y8I/+Pv8eNyF4kKtS3m3On0D9aSXT02IgOIZ7+WP9pnRCQRX48xFb
2b4DkJjg2PvAPajEOw5y53qDHFC2wn0KhsXcmdLoCb0fOv/ZjnOgNpLN/XlYMuDYIP92G8oMWykD
KvpcWqVZ7IclxwbXa3SkUGEQvk590OVBKogeVjjmig9zKc3C8ACyz+Nm23cPJxI+iqS/AkIfvS1Z
ql1x325eIGH9z1TZ0vqKkzAYs1A3530MwJrIu8AFRkqqAYaMPAzx0KK/vQabyIDfYm88kKEeyo+1
PReajR7iVNStyc3lspBPrzk/SE8VTeErpO4dCgFWmNtCjGCsY+ouGNpxW2drRi16JbNoZZ2hFi/1
5P7sd5djWsha2UsxlFOFEXGmP2cr3UB5eCMl6WA8pCqglQwv7YOApGnpTCY6r7uoJyuYpuu1sHI8
zoLQSMytyNPYW+iylfiRUF0uTOpg3tg3Z0xLccSKq9RBN3cjkdu1UgoVDmEFI4oHaIEPxka4Oyzp
gTag916iMGz92zLea8kKNx1xW25auelxTGFw97CyKwYcX3N37Zp/ln+n1HFCKcxgQOv8nad7r8xF
rqVr/pUy2tLFg9U+RVSDbBaRUmGm+5jMlVF+w8VkoU4pg15CiTvDmYu4A3xrOy+iXTcTCSZ9Sx96
n01rvf4ba7kxL4EUNwHsDaT/LnMdBaYYWwq32XXo4rcQpJC6ZAphoUzziireN+XdjdjPXqJph14Q
5jl+sJLcMENA4AlKAE4LGKnFG4rgYKWMHvSunT+87mgkB2oRw7eONtXvsqbiPVooHDk3U3rITXyr
kSvCyl0zdpziev7wTKjVzTXNTT0CXKVPtrqx8G5MXHxSzAtbCuenccf6vhU3znscnMi3KI5B9hoF
+21sERs3Ta1iAh6UuJl+iVKBhK0MhA/zX+/doxk8+8WEYwouQnmSCas0y5tITrUoUleZRgJpD7ls
23gJK83E+RHiRphN1r26rK3wSjhm/I36bQpAfgQRSOBnmI6JPTaCdU+vursjpQeyGDsIKAZI6NRJ
N/I/bF6orEVDp7OamQjSOmxthf71WKJcdha3bNbW7FwQzTLls9Ylxwjh5E01Fq7Va+j5laAyP51L
YpfowfwqrBx0378XfUXHsHOBuzzY22nhz/Mj0wf4/hazEO+QT33qPEYucpdDtaSFLsPvWBcDw5ns
gJtXZPnVfPDn4v8diDG4W8REwXzYbweCCtYxjWQ5f98wdNYj9LGA89oz14yxt+4oGHD2+IvSEexj
+bKnvS/NrLoQ0ugsImVMnNgQ75mgxLbSU/6Nnpd92cVD5ECw1SaJy8URJKTeCvSpMoo91bcWxNxv
o8DQVdirM0ahsDBGnWWbetzWdeMH6DV+HKdOIxyevALWlS5mja0x5FZIP3jwUpKzQpKXxg61Hhwe
C61VKZxSosM485tRjWbSJTySNrQiw4+dPUGbcyL2FgeuZ3x6hy9h1C4pXSq/MnxUwiMYCLVLcWkY
O00ISqLcyaVcW5GWpdybS3VmXhwaxOLUf7kjbd6fNrcgrMz2Zcgmw+4oCO+UDPoCleJhvUrGlygm
dp70l3pdy526/2Lp8MvS6TqymzG4vb+UB9y4+qJE1SQBHjxGrY8sBA7jtjUJKsNyq/Emi/BWZU7+
GekBZAsB6b2wPqq5bkNt36dZa6rWGwD+9T13BFyGnd5tV9FQC7/+i9k5062DIh7v3yFyf7XP59Ro
tlisUGyj5K9CPi0ocr0TKiSHoZ6mvOy7pZPbZZG8TqF2Fn7Of8HBjQUkoT88tBnMLYZE+by9GG+7
DEfpMHuHCea3R1Fk9c4L+7nsD+1JbphFs7uZKvDcdO2T830o7t0erDnEfk0Zi9pI/lZG9EjH6WOH
XRURGNRIJO683P2xbog4J7rY2hf/iV9GGEAoYmPEAK/7udjuN4+0sCFo3M3ozBeIXuBrPcQx03Bo
wMLdyI3rKQAc2VuK4/xXMkAn6BChfHZWbLmJ2p96EvjOhSpcz+3k6sdT0LzOGJf5cu1pU8ECawMK
M91VtWrTMLuZJ8SnU9pfy6/YYDokfOKaWRxJgIWfppqSEps2+MMa74c984ym2F7Q0jXJyJED0Gls
Po2i1SMrHAQ8Gc1mRsugF60ydAMfPYxTx44TkfInm7uBBNxRVE+AbNdTpUaMDp+3IzfUSj2w4CJN
OAnzBrQjle9MrrwzPgchBJyTo4b2lXmdSSfCU/mMz/WNTv1yMsGILiYKzvm3cEvS3Cn44/GdAZxr
esdC/8OFFm5ppF2STCGTfWLdiGSqp530yTEc3HCMDU7B7wr4qasrrEnx4eWWzAK89J/AjeapnNU8
ozD7PjEvYGCj0ELOLz8pS0dx9UwDF3pZahgm9JnejWJoHoL5UGLZKpWpRBkk6Er1Ng+miG7qCtJM
PShP/icY2aV7g70GSSnQ3teWIfjioyRpGltkafc2YG0zJjVrTpEqatSlnbN9wpbjEWl3lhBRlBJb
qIwKVP8VNXVuiHvQc5L3+nlu3i1eqhjSbY/DFlA9q85U50Mh3X+3XWWl7mC8flunxxbz9w2ZgDG+
eCWnHIdtoxJWTN69CByLgjBz9XG4HRfc0K1csS/0AXB+EzKKmeZgR4OzA9e6eSaaYcy4DjqC7G3g
Udado6hC0wRreKmSjxssnsuTsQEDT7cH48NfmrqqXsVjbzzny66uRtxbAoJhN65gJnB9umUUL8T1
boF6nws/11GBhKMVBP8Ab/5LEMi+uVOpL2BILhi8NBqDRQQHLVewcT7FBlOEhgLkIXL2OEfX+A1Z
2u6ReF/NtKIHEnf3yq5ZqM+SiNCZg0Ow88r29Ula1O/cIzlQxEvV2sbuyxJ3i2xBOawb4rQeLdss
tszOPUvdHl+oLDFZwbs/hZMv0JUQFg8Pz9MOVprHLV9B1r14Ydm2qDNLfLx3VmzIxQRWk1vbCoiU
Si4cF/kKdxlL2t64WilZauIj1s5PCifmjDALohICFOOj4p61FA9bQtcjuLrHsRWJMvE8jNEY0eFS
XLU/GITVmdo+0FPCM07p0K51D0YO8RhxHauGegmSIWt6uyaP5CBqUaovM6turaoLcTqZ4EN29l4c
wWyeP6P+bZfZEnvQGUdAl9fdBaAhk9GS9Bfba19qa/JVzeT/VSScoZFL5n11YgdHp7q+PI20AJJG
IROdrHAxe8/WcQL/0Ap/xx901bHqd2eSog97yBtkUW8Bicm2yGH322U1coH94g1fniyVMFXvRN2L
Bl8oAUBnw0MN1YCC+88c1Z5RlDcShQqsHXcBF547o4r6248cMpefGBf0nfXhslLBJ7PgOFNT8NLb
QlHCSkJ/1YiPmoxPCPZf1E+ftTzfVTRcvHffxuFsM07Wb1zIUIi7beiPUh/5XriOCWgV5tQe/RUe
pS8GWTEfsjmR3w1JUdkXALmQ4Cimj2sQdygKK7wsnPAXqWM8qTkXAPUw6fKMcS4FG43ym/ttGp3h
iBQutWHChyPFLqLIUy6D8mQ0Hlh9sRt4g9Rq2WqnjhrmDg0Wgyn4K0xYQQ5MB5Bx3mtyw13YUHpz
nSkx3ipW1vBt8SVywFUVmZ13Gqq3xAehdM3c1LTR1dKqgB0qtyok3zp/bo8KS0QAY5YtF0P6fdGl
JrFqHHBvuwphnlrNyz2cPItt3ioQfYSr/B2EXlgncc4Nutvsc43JivVPKdMBhu3hSIQn82GQCe3S
1X/rRQ8xdET4+YJ/SnrwP+2axFPJXqwlwcqRv70BfkSlLjiRlB1ta0/QENc3dbThZ4zuLYqV9DLj
66EE5w8uPSMv7fMT9n7a7X36m6/ne4dvYEWtfXP2qCklsMqykQAh1jGAuVDL+ZRANzpFNubxi1SM
i3QC9BdH3yNDB99lVbnFMBAMU3hAWQ3Xm90Fngalub7oboDlUpBOOnBMJ9zCqSC+2F+DYHz2VJ3I
8aixxIPV9lQSZB4gt5g+C65EN2Z9d2G/o7+N6RVDhoOtpQkz9xY4scpq0GE1SXZEPSoNmALM7Twc
bmW11PT03TB2Yv0OT0e8DyljUOOdd9aoypbId0fpxqm+NS4/1EoKEMd5wq7v/+tEcCefRBV/uumz
jqdWoRAv95Doo/o0h8DJN7QVJq6IfBI4YgJo4/aVGCzc5k5hgf2wnZHL8SiMXN+aSHHbCEpfB0td
r9jctUH4ZhKww9C1ycK3Lo5Cg/M686+ze3ntrJLaVsv/LWLMsWqv3r2I5nIkP4PiwvfHIyA0JDAH
SQ/e0POXGL+GC/EJQ1Yo99Z/zsu9zBr9Pzp6HRmYt/8d4vR+No8LhMX5kMtErP6EaCBLL+ztkzFG
UR7J7i5Tz+61pM2/8bIwwotUya3Q6ejnVog7cy1wYl5AmUZGViYm088lcmDFLupTdJ6Q+4UbauQl
TMzeHt0kKvGIS04690NKumsZsNhLVSO9uQw4R8qS0wEO0k3/434iELE6LPpPUMZqTl8FdT4xrAcq
OrMOUja/dzrxX6SVMLb/QPikzDIe10gLiuvpyA4p/hSshfaXpR5rG6MLM688JTTNNY/6eT+naClY
BnDETCK5b76upiYSebMQy0fr+YvnvQjqNcGftlifkA7C65zhRY0bBV0hErxrhjudR8tdLX1x5/KS
o81f/my4KhHGs6EEJFh06MqwmudEUf76voLUlumplLHDTbcp4qSCkjDo0n1A/wacDuJHHSmQfcDw
7JB+YT/u25sZaR70PUHejBJqhGQCe3TWZc0z107E1SSUzWJDAOeoSpcF9ydJdK5vMgiXmM3QTUjT
dTAOoQC1g5Zh+/KZhMrqj7Fl0NNmyUGFIfV7G7KgOY0o7oWiG4npjsZ7ELhGNQU9uN4RDPtGIeUH
l/RgI1e3DLftWgMhwVXA9erJEMy7LKn986D7eJ2/RcpOHZ+ayvMESZsliM02tcP35HsYszuM3dqm
yqYlRRz9CuYR3fc01WX6iI/+qJpradewzSMVZ757E6jJ6UUhCb25LxS7I1WMLat6fbKiE8hm1Qw1
sKu74a7HzPSHqcZpeLtdqWulYvui0KrVYR60a/W5VVHOaGyiavb5nBFIsNj5gv4q2uEnwchaRlX9
J8G6x0t0B2dlGNgmbFzazCzwkFK6fINYpCiQQ+NSlqmC1Yi8XYstu3khGk9+fSCa7f1fhi9eLPz4
M9abwewVQaC2o6XoM0IcVgtnXBtmV+/I6FGM0LCNnFDS8ZbGIqLt/MyGd/RKusCAFVuyABPjPaLX
sTkbPR46hql8ImWK4iKt26wOia8tuHuI6WyK/XW/SG6Uzzl6FOwxYAnKxQzArBd7YMXVY+LfLuDb
UzJRk2U6IF0YkOQlneufxGO59JE3jbFgiKVUOCWi30VVjPJop/pw2NCRMm+sRLEPaYJSB+6zwuBn
bUc3Llg6sc+Kw702Lrn8Q81jNqMnLlwTbyyciWCbKtjf3/n6d5TCDltn/GYf+6TnXdeyNaoaM+He
CLTPs+KQgoPx5sELfbtYU3umPEKTcgMLF9OTAv4MXdkVOWx5R6gncZkUjc5KGXgSYLSxcFtihCiw
Jr1LhWhgl8/E61fQ53fFVazUsxhk5p7OK1oX2vkmDT2qK9+qv1ORr+oVvAIVcEH4DlGnVV6qwrZF
moQNjtNJaKJQAPMUI+BDf2jB5DEBpMzfts+XvvOqS689UTYU7dGCt5I3KLsUg6MyTiR0Ypd9g+aD
IJLcB59j5HchANQ35sbuEp9kslUWfT+QHjLB7h5umA4XRDAvbaRf0zdfLcZtxyQgbOjZIw+shAKN
iVxuhJscfmseiAKtxYWkOM7t6lfoMluqvR5rBSPUIlDFfUymPUKzd+nlXmZ3sdG1ZSrmGCID9a/g
EmeKz+bTnsTivSFvO51+aeMc35Yg9mYHKSswe5NPStRXXRUeb5I5+AYoL7FO7yzIdtdbd+kEY/vy
dsqr1iXTAzpZq2SGdujhf6YXertahH+yvr2SITiO/oY82hS6NlCXP/eURkLgV6P+kbaZIi5m0Jt7
bR21vM9VH14OCgjXt+fyk3ec90BRzxoDWlrCrEMLo6Zl+XED1CMULLmoAwDMbTurzqFxAg4v0olO
aMtIsYu3iA3AI4uf+QWRqUN+HALwtEwJooKBYj/drEOsD3unLySOpUgD6rel/HTnnj6tDYC3ma2C
slL5PGkpVffzRV5u1ADmKjGNWi9l2uU3nmYWL3XvWqKz6DfBukJVf0w7yBBOkkk0Anw5XdGykWAg
B8Sa7xr3rOBtOFCrZ9myZQYPm7GuSgHC9BylSNeII43vevtc45SgSYJXX3XQkw4vp3CMMNKYL7Hk
4WlpUQXyh2YOEQZfU+q+hhvG+hHeGTSxBRclZx+yOG0hBjhZ3+YNb0FuJhgePccDtpUrlnyKrdaj
2HYbhGNhnh+Q3hjO6zyGRKYwNslI6p7k9IjfdUpNebJnGed6muJX82dgfCSFQ5vD1/eAaWxWpCa3
9QtJ0Kj1GFjsxu8kkISUy+NtOJpuKzc9wuSrdk/KgRzI2QSSSiDUV6V837U07QzmAaeDoyUBr2uM
wXu0044HFB+PeUUTUz/PyntbfP/NGkShxfSkI4hCPBzH/T/tiC8sbj8hUNeRXGdZXXrTeJ5QwT7G
wImBSWm9nLVuAIvopkvnEFPdyMYCE4Aog7mDDJRdlyAEMcHVMquiw79BxdwiNKEzd4/hua5ZvxE5
x611XRpPi1CWPM6WD7C+3NK/H7h+TYMpPgnZj0JzmIkkbqLwijWnowcOKKOtWUKRE8H8BZL86hxt
tTjT2zimmyXVRtPnyfO+qQmCA90+HLq1h1mu5n2Te6dtcGHFTASiDrxYpcAPq48Hbknlnq0mEtt8
b3R+i/GIE6bRjjDIrzoPNtbZ2bOnkDzkJ4WaSSkJyTzRwwonUCWnsBDqO1uheHtpKmBkeM7Ta2mk
fLq7bOqWPX4DHr0eewhGfKe7AeRj73jdGT3wWQp2j3/Zza+GpnDEn/iIN6UocDdZ0baM2ZqSEO/4
HIoUZ6naYL9Wht5VSnbQSBZ/l1uOG/vQNsfQuONq1PAsbuIq0n0V5xnGpqIg3sF1T6jgRS5uovlF
dBiMBvUgwEJnak0U5P37PHZ74zI8HOoEWXqJ3VvHMzQcaZrH54OzfWS5zHHExV8/3prRHIt/4z1Z
NAfJgZm5iwh16l99tYlkMFVykQjsG7TZxsDUR62709Ci/7JTDjKh8fDMiL34R7DDiy5wIuXd5YdI
zMevn1lJCCugHXJRzLi4fnf8wlcZedFFvJN4Tm34uDBzclcIda4gTBVrmK0XyNo/nakdGp930E0X
sOJNN6oNVJ76HfIzBF3op8n6/P3Ui96GEIqa79pAsup58nGeLAjIkH7mJ+m8SkAqWNVaY8qj9sB6
qKXTo4puPXCDH3/sxVCRwxv7jFAybMAIb0JGmyS7KDphnTCoVqxF2OQcMeTrMB8/AZPJtr3aj/Cl
W8b6Lljm9DIW2XTjSNO8FvVXoMwqNbQbr9RAG+r7tp5dtIcW+C+uTfOHsKFd49P78cgaUBrN1tpt
M/dN4wZ03M1tDgRl5wJkeHaJn/OgnqMGDKp3IdUbTf1miubsc9jP/edcfyZ3yUWyVTacJ3sG6syv
xgK6l59N3/bP+SEXXgiVKm5URV1XoG4MosT+FByekqPhjLw+9sL3SJihaRezH0q1U/Y0k4AkawIo
HuPPZ7XZbpxy4L3V3+H4jQysbdk05tiUvILwZeBu3fnLNT0P+D5yZVc4QSsjmQygKu19h1u0b8lA
iPl1uo/sypu6fQjfOOQfVa5dpl+I2gYDWxIVssS2inZFtZDAO8da2oLMy+rWrGA/wqK20gI6Y5V2
McGpKcUHLVk0gExSLlEKAbVsPnqqGlD0h+j/vFxjZhuVs3xkthUtITiMgwGOo+BZ3I79kt27IqsK
OD+u/z5URIvK+mJphVsBecZx+zxLzQ2H9AD2uN4oCWZrgXjTZe/qifwxRkKkSl6bIyyv3fuofQ0N
L+X46Kb70Rlj4a12SiLDeloQSj8oLomJbQChxqTK94yH9IfH4GPxgy1wyoQFLSLamvypuuEmu+5a
t+kbuuuzSb2qOyCCiktoMiR7dBOhT7WeVd/pxCTknTWjcP0JgxGD752Xod8H8DSWVHlvX1b79w+p
QVbP603WIe8tzDEfdaInFsgDjBnzVXwRy5vhREX3hCIp/io1lbtI2dEO3LyEZuj1iEfOR/1EFWqR
qFxzostfxVVlpV+qAQtYIYL5Kk6TrNXdS9aPjhw/y4cir4ohw2TwCyvjt6lKnDVMAuWMBv1vLFsv
dvuZ8EF5LwBhpJ5pR3Xo3YNvd3pyT+bPNLEVstUkJFm84pZc8HxS416Ug7RDXslEVy9KvUnU/F9P
0DnH+xSCrmUgL2QYM3QI22DmLb8sSnh1te1CPXc5c5JqZ/ncbO/MeKY+WsqzHRUTuugMot4eeQqf
hJa+3mhBKhCE7M7XFua62hebsHW1TUFGCnhZvKVALureRr0VVdf003pb+glfjJvYjESGj/FqQr+f
ardnANpsf4Vs/q8MjuU1QurZVE2ILCXcUlZXYWVbPCwkVA1L1iUa05tTvgJu3/zsA2Rp7Xaqv1G3
No0Lsdtha/oSTlH4iCy8U353BQoYGAYwFkYUdw2WIBXjXXj3Y4rDJwYER/4uw9L1g13Vcvurs1U5
uRYt9aC5KjazYb1yghWaJa+U03rGCMQZIv/JVH1pLEJbgn9kfZMTfLXThdmHSX9eQOUSwObMJCyf
FaMm6icixG2N+xOBjgHvV7WIBdprsJNzkmRVeVhyHttt7OPpScpXwBUjPyOKiR/fNxK+OF6wHl49
jMNmz1cSLH7w/WPHi5Q1lQSVv/uHtiiJV4YmtZLykOuvR2rdG9J7BuOYxi7OqBfjxLpOde0WgXUZ
s6nCn3YQE6Gds82nn7WN2Y8jOrgVh90Lx/FDq+WDMKjQ5yIulQSD7jPufysKebe7H4n9Qv0Z4zsw
2NvgcXnEeCKC6qsq6jWAOxFJtdq4Yqw2XMz+GJVO1RSg6Gllv/W7ksVMqr1POI00Fr2Ypohr8dVD
oMh2TF+p+yv8uJcp5ryPnJo56YIqELvmHjUJFlFUT8nx1Woh+CUDNDTzd907ET1FI9XUs9BiMVfK
NZcu2K5SsIQ9DBLG5ULG9Asx+S3YbnJLq52ClNQwoPeHA7nVocosvx8bZVIrQq+dY0P1ko/SCsS9
knJ4novasZ0V8H1t2M+gK8a03BKfo9RxmlxVC+IhJJeG82zp2cLGWwgRsQzPx3BSOMfq+PmSkUut
FQll1KpRva+I2Qu20fLkUEuzTB46Jz9Y0u/Uo8rlf+FoN4cqlcvekSTvKP/z8J95u73wbKhu/XLM
DemYeEaOiHk0ySi5LKV9DTsrrb8o+bfBQxiGVt+b3rDbDXNPjiyQvSIP+apbhzgJrvwEw9foGPHD
ITHCi3gGLl+w2YuqN639fw3ddCwGYt4kU41Oxrc7dQ05pjsxYAJf/+rl404f4Jc1pNWC6eZFBRNL
LZ0/c5XhbE8UP8LbTbZNXV3WaMUtNSy+3M0zZHz5XnxWi9URPZWytW+NEtgQVIZerEuJeWSacdG0
hYyYG0ea5vKLsljjIHCxIpivaLteELJqw1cEAt6Z7qWV0GL7JRRCedzJ+BrD1X4qEs+5w2dAIj5i
4/cvMYuy4JBJHTu3nOZdw2IErKgbSqnxaVx660o9KNH23UQ7hCEr69k12aFOP8MX+Ipp0h6Q1Zx1
/vR6+DmeXooeYT/l9dYtP/3y4ucVCk7v0VNuxSyrftsVfsOkMUztE0wDrd8hHElZM8uP2mGqsZnf
m0ss8nKwShsurd6UcHx5PnHTmpjK+qg7jgAVMbQZMjAycM0WyN0rUAG1y+0l/350OJhBV6GNXvUi
ZhuOPPIw+vjn6Bk4qOnYYzLOHGc7TWWfzzByDklGzWPgFNsSg/S5eW070AifVVL5PZq5RQlrzR5t
/iYLQ6o++Sidb6nFWChTqF03LBQ0mFDeT/pgoRElwfGlmGXORCKQgiF1WikFYpyeqrIwypUJ4Ol0
WHjUACnc95mZOW/YgBYwan32wx6uuvFUMrwYq9E6E6oU6kwLewT4TcLvVySfttPBP45BR4AVdaKX
g5anOSEAzXQ0LEXqYpUAqLRKW+sszYF81xvG8QzhL6QonJ633zh8cxstwXWvGj97WbvWYpPkDiE3
sR8aycAVj5cLulSm+sA5utxDGydMuas+/ulIc8XpLBnyyuvvgyvIgX32Efwsh+6OgJQJGo6E0FEK
c22oZHKhGKuu1JnB78mFdZCogldNz9o5xP7IIkYWprcQCmwrjeXejkMMQfQv8gXG8QQFCUKb8cTF
RipyUZz9YabKc6o/bdODMbQREL7oGURD0gyztfj0xcBCuHtn5VdNnZEJxkQP4D9GUaPZNu+DcLxg
aO2LUMPgzM6l/Mq8kiN66FZz4xzE+XIKcceBRh/c3PUl+e1cNJdSSHAjKlnPoffbBUzqBpb+CIK3
d2emSAGQ5VnKNwVaY6Ixyc+PDm3zq9tHgTa7pN1/Ws5jBerZlVyZodcPZmhSizlZzJYOI2y6Sd5x
eCqPW51GV0pfoxGl6MrvyhntORDTn74VcnhkmbhQwxEAzSqQbpuf24phQXVvGitDXz4AsNrE4vSb
10URhVg+X+Czj1n1olXxDrWyF0Cm8fWgAq0VUafForZmYNJ0u5Qe4F3vaJlNCYSQg/ghH3OnNx/R
za5Jbmsd9GwOedNg6CWh0ps+FCMtbY1oQzNkqTRXWKJVOzmPf4PrjRnLN/jzgBZbq5fbRoYRjk5W
jxvCBy+NG0vBRkC9d3ObtlwVkmMupQ0O3ufSQNRpF0Gun8YEhTyGAfGiYATcjvUYWjksJL1NKKvK
8+MC5hTIFqjH8+3MXTsZ2YGSL4K69SvbCsV7bI6qc58JA1NkLkA19yP7ROZCFdaiOpXScWUMv1KU
F4YXMo485xl+JC5ExkPz3FHk/o0CnfINVmWmmgoAm7sFzG09yNIl4X5F04yQGV55GxuEENh49rb+
vltpP89ZbDHq1Rgbm0VgapMXQRZFDWGeZny0OBlrpmi19v+qyGyvvkA+7pY8nAILyEY/mb0mplrU
ulHBmTcniWQt583BVmaRYs5iRNnYCpcshNXlJSn9La+UZ/Ya8Nv2kxSuhV2hubbV87n26DMjycmg
6O0p0R4v/oYi2ZCFcV78RLz1DrT+mmYbRq3F97WH0/x6jMzGLvbl9ZDCrcHqeLlxoxMcZ4T5mNtD
7hmhCgRNJ2K1n4LJhLYV8s53qxkaxo1LRUpWOb0LDV9X9PADFY95wL8XE6pB1k+IBGe0TQnH3hie
WYXnXv52olEb3fBxibVobsb6H79lwKnseUPXIuJgGPxUMXfGkNAWjMNYiHDYhxoM3qcEea5rgDur
qgRiWU4iIRu4dEsYY8aieSNuMerIaaEizW6KP7LZfB8ezEdL4okDkCdj5x2yrefkibsFXPIw3BOg
TkFNqmmsQy4W+xnY7RBBc24MLbQIPSpPLa8+Ye8R2gFilI2w3bRLo9RNQ3bMP3sPE+P8LL7bHO58
YnBzKYJzk8R/N521dfjI+7/Csw5/jqgK1rs/NEE2W2HyAukQiqxl5WWyOqGVqEBH2QSybaH6V88U
6UcjCyvln7S5LfQX7ZdQMchLo/UQ0EXVaNR03eGh4CgOlqOQFr2LnqLhq8JMibdDw7IVvSHzbFpy
iC9E7NqZ8IvA1P4z6NbQGRHgsNaB1D5kqweceiAW63IwxG0MKEwNFCZ5X3AsmokQs45g0Cnfiupj
tMLPn5QUVRDP2auPMtfpoPWL4nJDZDW60MX9tJEw2kHgb9U/3WkBRnCy4UGo2BrKdU42mqR1uPVi
rax8EB1vpxusoZMLzeJXRoT7TJo+RAXLVCOQim1TZZcPu1GbedBizPoVVpJQyMB0Tmf5Vsb6j4cL
AK2jpvLCBC8VSzwAZ8I7FVLNUdKcw0Rjtt3tdNCOt5m85dg0O4fHOKd6BPlvKXDsCBbAsCB+bK2Y
wBHujr+N6i+FQDOhi/t19s2Xhpst5PQ/fEB0REDkeSJR1sXjN7HWIh7XhCloHOBamoVbP8RcBH0S
3ZFuebq3q72uvarpqtiy9dg/9kZ2T6nX0zY7z764Mf3rAONpyn05Hac/eUlzUQB7pdko9VYpHHZ9
Q1SvhszutYknbDCRSPvycGZD+/SDTiJjn1p9KCRo6mN90KIsLg0tza/Ut17/oEDD03yR12G9RzfZ
Wirq6hcTO2HM37n/a4YGPDJ/o4dju54QkBq/GwCksAxcTHHvPiBPi7wB3DcjLcoJDzgljE8crHuD
qYcUcXchreTILxMgQYwrH/D2VMOmhBrt3cBHfMSTtAAbsOr1L0STPYAbOW0XRleliOcsFOAppLzt
qPS67LKf5wz4HWxctaPo2mhZk+x/GAJZ0u3eCRpA0CwQK5RxJTL/RhzB/7G/eEKOlYg/EEiQRsVD
fLxWvZWf4fIO4mZ0l5OgCj0aQf1Jqj037DRAy3nO6XTpxSLMvYB82Ii/R5LqtVu0d7kj6bHxAokM
C6SFaaAlcuHQK7l4R5ms3GQxNH51JbTHX8PLaVC+/J8i949Nl6nprPJCTHaKAUHAjkjeYEsTnHJq
V8JOTn6WAB/DejJq2hj7JrQ5r7fO+t/PkXU+Z3Yc+W0qcLvF0bL7Rk9QOFuLlDqIUSqmpuXhCMps
xEFgy/aDFCBs5oYorkeirLjiLhN0UaapYJ+Jh5s4IlWbvT/n/u33m/PAZi534Gwsjuz4NRdAVaO5
QSbpcbCM2dvhSRKF7j72Aq5HU87CbP8TLh8am8+cS3d3DcPFfakoPGGW0PPHFULSqBYxW5Fem+v6
kvwVciXvBbSXAmzSVHZ5Rzy2weNOxD2LsgLQPj2yqV91FlH3zfRFvRv93Y9byqOJ6/UhaQb33Kf+
aP1ifPnTWADGOhb/EM4zBx8hdAeBbkmGSoHO0sBoN8CXOzddwc/Kp94tDRfUIlEsh5NryAhPfM9E
z1mBTUQ79eFir8Bpn59T1C/IWJxRv2DXdXuBpWmll40uSuTLDntCeUWV0IijdgOXCc3NJG2VdiR8
2/EQ5L4OClmyiDXvKd+jQH0r3Ub+WAV6xIdtfLAk8yJhnkmm53yBdbJyk0/Z1yjDnA7wqjIZqlUE
KCe+e6wb5Al6iJ0+q8IZasQUI2mRstHa4GiZWMyU3ZEtk0m6vPEsBJDbGjaajoJDEAoML41mt16s
zX6Ez3WP4887amJBVmBrTnJ7anOML+ZLZXSRjmqB15R3AuPcXV0FhczViOe5K5oKGAoSpyfE2omq
Uo7sGuFLtE6X/CB3+QNjrtgsYY1VnbI0uHVT4VqQEZhD59OtJp2YFZEXI4zMWtzRkm15jrqe2T5X
Ul1Pekn8tehOCw9zfyFE2Z5fr8D4p3QocygJ22AjNCRd0eFJGU0+HogAFw7BkelLazWWUBcCj4s+
MQk2Dzht8x9/7IS0NggV3CayZTE3YE1QoQw6G7uegczY4OTYW4JE/Er3ztoKu/p39RoSi8ZGW23z
CF9rLRjZTodOrgEDKm2lsm1++ESVJP0k9Jq5gxIJzOQDFRN1PCwMdqnowIjHo9ABTBkIlLXy7jBH
0qDf3OsUdj2CuLE+G/q4mEvKP65muqEjU/rP21qgQ6Iu2NXOHqdqtXJfPkDjuI0CG/t8o9VfImlE
D06hQ6G+yBTGss9jcNgfun/B2NSUmXtYzlXI3sqUuHZnLQxCoqmkjd0J6LqXznISF7qBdkPXyUGF
tQ3cPtihUeXaxiG4I3AXniUQ4r4tQ7yMXR7oags6ep7I9YO9w5InSKSUAuZgL9hjjz40XUQqf9ZG
iLGwet1h080N2oCleXMeamiAcTlphoBCa8fs3lWCDv3z439de942YhzXSjIgQ5ZI5qbBrzq6kK3A
lXLygFTskHc2mEh7nxhA4GGD9lRIPgaAsJOCsHXhTflvab7X2IsEm5xGKRCLnmQ1c7ChMYRDyhEX
2DVb/NtKZuvXwQIbVkOL8YHBwHIjYp6vC+gd3O3T3xDxMNZvLi8jEUMSsaPTAHyPOKyDWdwTYmK5
77YfbPRIc9eCDaExvfMISobLujVBtLqV/3gV+2+H32jGlz8NPHfErvL72v9Yx4gdEGZ0DYckjvpT
a5XzJqUv10+mQLh8WyLvuIM35rbd+hVYC9pYXbpFsqxAyX99IvRkmkUy2JTi8SxEue7+ygEiyUR9
s9+q/m/QizVQgFO56oZvfXqDfxDQKVpHiiNErALanx/t8bOGUWHUHw+oa7VEmGZSQZKgBvCB9eh+
omKBgesGisTri2q6rOKerAnTQAnMKjpy22jnJ98pA9T653GindORe4MbRkBI/niRP+ouOGs9vAvh
RrkztWPy74GPkFgIhwWGE9cEBcDmDMWkCB3wWACxMgLUFG8KD5E1vaKkPhcN1aCRb8P/KSebUKOT
Hbmrh6/J0FmgaMzeD61/4/Ny6bavTW8zdsJHSOj3aNe8GgGsJV4Aapc2iaKbdRk21xciSC2y+t8Q
8mJd66Z7S29XKMKIz9NjI5oaSksQsQMiAWagBuyRQYBh/twWoYm8Ysm0KgIhhkcLcHDhcH0bYqE+
PYHJM/ImypOmDGqH3100PB1EA0Ni7KuNpBuMBLJJbUePRUty/sd9ulXis/RKUVBBrSr7fOg9d7Yl
kG76Mb0ca7vwYZgF7BMr24yq7O3Mlc4LTlUOzxZAz7HEwhV8/wfitZUJmKZJjuVZ1g0M1WgZ/kyx
ng1evFbMEufbHFVgWiCajwbSFg/etN/AjzpcFPZ1GXP7mVY6TLoS3W3akB7X0sSsYKK5rdTSif8T
fO7fsTkZ7tYy23heBGX1QrrAVi9oZ83zX6a9LzDHesqYRzYZHw7eAX41TTFiDdaeQMI3B/Ds5GhN
5qlL0/aQuEugRQXN5ukTLbWPzu9nTBM2LZ6KFicwx8NyXqeqaTefq0XqvSZjXgPD04L7X66eUOzl
HxCJc9BRhqHS0ZHc0DHffpiU61hIKXRXh2hOEFrWkY7/NRvplJlA8+UmFfHX3nHrUcMfpZX1XrAV
8t+/8yNUSnar5z6loZwmy/+7B5q5TXH3Nmvi54LJDIcvF9MMfQ43JWlLbRndd54FCCBjDYzGoNh4
phi/9glsg2PQI/ffJcPLcSQ8tlEVEzWNF7elQjkSVK7rwT/tv21wwTuKydpIKFou2DhTmMxGqt0O
ZITBfvPy06fdxIIp6FtOFkWEjs5UhByIlO57YxqrcUcXZRZcfhpjBb9aAuiJGQE3ftFyQf14b6Nq
p0k++BV6a+/Dgwh8YLiW4j8rfzE5pUX0PxDNml8K3ABiL1RDNP4rkF89BP9CfOzi9nUrVm2eo69H
qiXbvlTrzM2zKKEUVUD4lWkdAR5DnErn1oaYSTFUnG2uutYJ25vvZ5P3/5gseNvsj1H16h9chLRn
pEdNll7w1eckZeX5yZDXCO3MCQwjaPEgoyLrQ9IG4aArwLCXCai6NplF9EAmXaFZSfrUsHiJkrSv
LIWmLM8qn2U8oNryxe0EeCG58yfahlkN1AUKXjZ7Npe3+v2TqamVA/f9R2ZvRmb6jPanvttooH1Y
lRe/EE/O+NDPFg53SkTn4vYLzEDeihWfc4g+ps9AiBWKcVLz3WdxHmzoYIwa0GUHjpO6xxh2yruq
VMiq36mvTI0RRGFNpQXJOaKOHmaWryav3Z9qanhqPlzPLftu2JPkjcz/f9p7Dm4PPIivl8op2cx0
iqg3wqvKMKCF0kg5uySqcEJHuYHJ+gJ+ssA+LNeJHcrDmA5d+llFzEobp967zTS8Hgw1z9CXZpAA
a7MFCCMq80HbRMvzz6PBIr/KoC8uRegReAqpylsEeiA1frUZp1bGTkQaFC7en1LkgTL7hy+ee/pr
fuIx25PUY2/ypqjvLbWilBPpweJHAyFUA9G5npvqj8n/AGi5JpbGfpyNgVD06XpmADwxk/hw477R
Hn2d4tdfMX18DwKnLySnvFAlxSSDg73DzfMRCvIzSxTjoquvyTvkOm/q39hcQTa2a1wW4M6vP8Fe
h6r6U/R0E42zh9ffwwpthN9gxslnLUsT+OvI7ffkcob7g3OWA9rD0AYPmdRUAxe/9kN0VBh4TvaV
h/oA0HyY/Bas8Q9udhUbyKV4PHHVndv9YJD4cJWUQNd0SmgofKmwAWG0DJMLOe9RAiOkpHFPhqVn
9dXSn+6K3wYh3xuOQhJyMNJKDBZ6zhVi/elDo+g44yRZ60IrfPxyCMdtrkxSNdi83F/6UnYVQuaA
sa+ClDmaEmutLegK4dAyug62MrdPb2uaiRZmdOeIYHi5eZdBHBxRPONk2QhZBeRaY41SpicUTBzJ
zKfFNalOpMJoKT5eDM7Pi+UVaLaIbb/l++bNtUgUDlFVT/iwzP9tQ/BX6zKmObIbQ4k2WzDW7aau
JP9VJItjvX1sIKodXtXaL2xp6yCwnbetgDkRBJMFnPPH5bKYnATvt6EgQT9kBsPqewFTCAtlZ7Jl
BgYJppbh4pEv0f0QB8wFwZY5vWaGvDrE35BfwVuhndpkC7v9YzXg7PmEZJKGxxIxK68V/GzcXFXh
xYJy3AkPFF1XMU+GBFTEF5aNMhQtwPELGiURzGbpqkvF4+DW5r9RiaCD0LueQvJtJA/I1vwBc2bo
gSjmUDyWqb4pzibT3cRKyAfJDkV54dUWra72Y4+XyoFzNXlYM7JRkIMt9O8QsWsmgJfFtEz427iM
mZubpHWr/Z5lpG85z2rIPKawoPcQfGfymPi2Uj7uWssZpKehVXJMvE1dKCp6YgOeaCu/yoKcSSlI
BfzbBdoqwM5BO406LGMcdKiJbBFqvYI6hml5JFx0vOdBgC+8GpiVs5m5JZSDhyxLds+83rfjfP6b
Hu1O2UbY6c2uuPkD7UmNMALatfTm6b5oqkVEZpMSWtgpNiHfQmvbTatUBfwcTlBWBiPSUG5oSwJY
wSL7ZKjRwKlmXw0DQeK6BG9GimpJWnJsg339epmioSR3nuoqzBwR94+//SO0/l9BNHSxxjDdxl0v
RrVkcUxfvnWRlD/+0ef/Hzx5b8j4YmJhrP8HTHXHIiaMg16yXOiAaujKBSn3FdElLBHxEzFB7pcH
aoO4qUHmG4zPjn1yCYfXf/XkejP6/5E2t7ye/RNxlWFgqWD708PXRtQ5bT26JiV+Hew/xn17ktjw
Inh7OoZuWPkugO3F88x1FZtosMB4mzJiLsX1NWLzOyDKr/SGGZnSYWjn0feuR+xac/hkYtcC64aG
FSvnUG3/PK2yph7XqsqqIA4Htt0JUMNwmxhv1PuMLSZDuwUBQud9qZvm6Y9V483nTjPxfQWfcBgB
eZ/K3Dv6bjlTrmb6N1r5vSxloZH0Q3noHDekANMy2nvgBoMbKC17DppMNIyPC4155ABIsW7q4hv3
4yjh1NGWlpu4chIv57u7MKzEhwxSs4rq3x5ZKQrf/yaSzjNbfHDF50kigvDSGvmr9niLqu/dBeha
LYxFaPE7skaplPCHiag7DVYckc/5wSBnSKvAZxrQy1Xe6Ux+77K2r1pjr7GIE77FJVo6MS3U7GiI
ZYCb1y3+IB8zxp9bw9bYTrtNc8tpu/JbNAtJASdjW4PcHBTI0MqObsmXoOARp9Jw4qV09LshWzQV
ancxi6v4ZG5hzqbZ4JoACIt9eDuOceWPcOH96LhRFv3h1OfKImuybsKg6S6HJSgBEvOFAFcrdxDD
WXT2gDfowF0JOK9hGkglaxBo1HtdH5C+sy0dMHvuQr3gbnsWHD3EheC+avmadtX6HNpMn9rZxNkQ
9Uw+ixqhJ2qTY9qhUzKGu88ztQXo7/uIBvJqEb3DCZik2Vqb5kXXT++3Q2vSs0mDB+xCNr1X5a7P
+A8Bl+ydQQ05maj3gZgk9MUN439vrcFZ9TP7iNcXM5O3eA3ws+nU9JDJBxZTxUHLbKEdPwoxZu4Z
guQAhU3zNZdP1Nt0EYfwKAGTkLJorpZI391goL0CK/uRq2Vm/kny6FR4qaOJfEHLsZTdK951raGr
eQNM4X+henyX5RNjhWyMkgWuZkQxb5a5q868yMzXO1iCM8ThAy6jYXi6uJhgSDF3bCKelrOVwsBK
AwnoYc/tsF6TcQcITTU+/wYmojl9l2ZBRYzuWR7oOTNo8LXdKqkoGYOJ5wZecrzL2wHJ8jB6E0P6
xcpixxHsoFeWxDen5gPjM/5OmTTu79+MM1jSC850ZldjbOZ9AQBK3UWK0onk3ASxncHIsfg/0dZe
PMsfAdfOVkcgw6OTVmF7BqAQSvYFavi//8BxkY66xo5UM5Vm4J8ra1mMTejNoQ9iJB0G/NCdkwGb
ruUOAJtMfe9sbVwEGB9MKP2JIR2ROQVWc07XNrepkHHlykTVsowy/dOhlQQXVAqSogCl0W24f2c3
BAyxDWcQkpO3+PTDl0f0SQrRGWVC3SWD82wk8IR77y6inojB6sOfc1wKoxdW/7INCtSSakiNRf5o
WxzdmV7KbGhh91VnsICgKyi64zfUGmMu7veI2qwlS+Vn5p1EYUaTycOYPcwuz8yTNz+anqxyReVO
7It0I12jzSi34hADkCQyZ1l2M+Z/jC/gllw/C1MX/WK0au6MwP7XWerhj13iZb3yFK4XGNpwlQK/
/3R14bycYFVUZVb8s7eFI5ulfSJS+KJiRRH/0yS5UpAcWn+qLhvB2Rlf9Xq3QLku0sWvZQ39UWS7
PPYwAZUtA+cqxXziQcuj1/mQWDuquA/9gJNBJr56d6NdMaaczNT6mhFq59joFnO8+F+n58X4OVvk
Y807NlsPOJBSfvNf9+zBsRt8bGko2DjWqxNJLpp14lu6jUMW7UWq4sNCsVsAyOOLYaEg1bpk8mQA
hzEhWb+5LGhg5Na+wIx6OGV1tnpl0/PnBNLXMqd2jzWYjairfDyDamriHrxraGRfIqSKTrlpsjII
befc2YXjNy2w3KqCkOuzaz7PD8l923uvcLU2UJqvBdZJzLujWsC1StDCchDPfK3SK9gQ4NxqyaUf
eX2LZDygBHZUb+38kEILN+NAuRENPJiJ4I6ARn3PN3Lsy0p9LvG8ji0us4TeW3BGOSK3eW3G6wJy
d+6ewdPh1yYE2ybuX4YlasAlE7tLoZFw28q/ufDfseIn1tPySgKzl4z9Lgum00ozQ4QnowYtcMJA
r/JT2eZnpADLfsYjP/zsZ/3SvPhUJ22JQ5bOEpTFCabBLWyfiuWoH/QMcdsOkxOYGun5yX0+ozJS
RLVAiCSUd8iQRmzpihzBOfas+Y+VFJLxa2jcgmX7b88bPdVtySEuKThXlZE9W4prF8qnxWl3rBrm
sY+oLntMpHESrVBenBWfH3gEf08CA1zkkscRn9u7/cuRnY5QLA2RzAZujjz6w5IWNQfk66La0I0o
Y7oKjEAOWlrmKhQmisRZfHSsRLbMrtauX8gq65/yovBytP4g3mN5wGzVDQRWDSBFRS2hCtcwout4
7QfVZhQVpjCkSa6rx4Kg/mqYLB1FSQ8wdPla1PLJdC6t1JWHQJJURpeHOf1EzbjQEX0hfTqAxACL
80WMYn0HHgbDpdbx0OHJsjkWsRSlzTU/gT3NlB6LoXI3pTO+Xr8jvuC6g+WCoB/PwobL0aXASKxq
DwOBPP697ftwugAZpEw2qvqe0FLu3TgOALMfCd/q3hp5iRzyZbLmeKSDxv6HdKLpm3tzjy3T/c5T
/uFES7PErlbku81s/5l8+yKQ/lqZD+eKNaeLniwrbUFr8TjTvsZElxJX9mDvrbPxS0V0GqWNe7/q
bWbVT0NBJh9JeGB8D07QLrB5udRoquh4y+2U4QoDM0DwCiz0WpeGl3ZVJuQIZz0NCV1yoA8AfBL7
+F9G/KVlGEzgviCFdvT86upQa56J5/WTOT51n4A5SxtAxaob258gSZiXVOhuRBHI8XWDgDRWlime
QPk7rAyZWHiLz/SUUrwdEiofpytj0leYYUnXyMEfu8G2iN1Dx9RmpaQHTqCDWm20PSFYpGdjsc2T
2R2Dz0fZJZx+G3vrbDiH5TxwFjSqeJkPJxPxG9Z6lQNKvkk09oPf/jfvT9HDBf3nm1vwK1WtWlnE
A3EPoqfQ6Gw0l4OwH7UV4k5OVzVjQ2rSKDBY+EU0te20oU4ECAXzNHKnJH37W1S1A2A2GknfxrTv
seU2xkdK1sZnTB5QZEA7eJTrdzKz88Qn0Qys1XwUWuGWxaT/p5WuTG8WytGMp4ph97dSJ9GSrM1Y
KgH9yQbjRS2YQ1AU07RpU0LrfueLspUqaNe56bR4rslWdUebjnQEuN7jFjFvz5IrsOEeg4+kK3zj
d2B5mxce7gVg+25N2SkRwsPRnnxTo95syD3lOm/suEe8YfxyyEPXjc/GREPkf35SFrMZ4D6tHaWn
gpFjmC8KNygHpJUacwmkrQ2tHvpvQYDezMCjmoqaDNrIdcDEULnqi/liptaITi9lyMQAgOlUS0VZ
ShMrgO5xX1k6om6wrAYWYedieO9+cvDfpAGnTk5Orh0gBuY2CA/cKRQqsbffc8lPjyLIDbrO4ZSg
hNuFxnhvedkW8ivP9oXc0SpdsXuY6A1WVEf3APyJoiyyLSRhGSlJo+i9NalEGTaCDhDkoiUsECVo
fl7hzZf8QHhr1H5praS+ikxoBA2Ig4E2U3VgS0LkthyLH/r5xsiY+wbM3iDbtbk+iFoTVOf4+wTk
n3rZR0RHIuYWuhSBcCWaPEvS7LDpDbDrugpL2LQTDAnaRGZHFrAV+0hatqENRbK+hCXrnpq6COnm
hibVRwiFC4TP9yHIMLxu6KMCoM5WIWX7eKahGx5qbIkN4pEyMse0N7qnelGE4i//0D0JfrziDcvx
9sXpXo8YJBMKyHP5h2FKWLoZ8bCZnWICFST+xlB3KjtcGIhfNVmPI1OiWH4ea4Y6Le/h+gi3BE+t
JviwrQUxgt0s3YzY1YG2TCcxMRwnnlMAS9SBYfwi2zzLZ9Gx5mwelketVLho5HdyaBAYxgOmlURl
wMy3d4QJbhitn5+VtFqxi39JyA2Tt0fUhRbGWoZ8XmIPLHCnA8ptnOFdVR9ezkuLN5hi9v+T7Rzw
/PJZjKMwocXxvtF/08OrI8XX5DT5QMeJtQd0fC5bJSWn1t8GdQoIP9Yref1SnW+YO7AXvKbnMA6q
tmRxrOzZgaOsbHbI1HWCq1YYfeqNGV4gBdns4FlDJkVcmDRZhhrIDY7UL4htVnGFVUckyfI3Q3i3
DBKHaXB4A8Y0t2XfcNgwy2QZnemzc0YJHtaewdRpCTCKsuELiIWHDINC4SVLCVgzOkRrCeQztJHf
vfPF77sY0+XA8rXKRo8ekYuaerSBk1PEOcmb2Xza3dsSibmzmu97QrM/HG0saD5UuEv8c1dDghnY
BQT5V+hD3Klw3uUyI3EBAjVUM/gS1ZqfkTt6/ULMYj+rW1InSxWMrKylD+LfIMrKqJk18bJOU+X2
QculmZT5+1tMcMrAbyQ3ARfN+Jqhf+3f3YpSAhPAGmZvJHWRNMtH6cSSC0OvCkg/Nggidbw/U+rL
RdNMBW1Oj6PGQihXy3QnB4rsmYvtgI6ScBSR2NUKy0BLagL2dDo61QvZpS2wG8Xa33hRit4y45Ab
vcvWLvWCOlEUdIckjXpUaP3xgq9xzl5/A970GVva/etgqziNb67Y5uxRSQnO7pHA5Ur1iea0MirY
2w5rphHaUXr8F5oG6vQNJWn56S81TF8FoX8Hp/g563fmhfTYxFgevXdZ1WhrNDOa2BKRK313azeY
gFsHT+ux8h+qXzPsf5tMnBovwHabbeupL4BzSFX9RnpuPMfd0w5Ay+docD63hBAwxt0StIh9xBJY
fIdq40zSTsA3a6bNKcXnBkbpTYHdEiPbdpMREHdPDCwKY8D5dX8x4aItX7SW9jx3snn63EJ6vrOH
h/cVwBcQoA+fTZf7nEGFQ+AXImgn4NdmuX1otLcvEbMGKBfEql4pmrsz/FFh1nCetwvwYBdfz8mT
Pfkhk11o+aFAdHe/A8VJZvTkuuJQgaAI9EMbu5Pf1v58S8tUNSDZfkVF1QKI5UIiElPBYDdVtzD8
tejMlzIBRQbuonslgRFX9nAoUUGpkrP2pkHMjMPwqTAlIg/ySNvqJkg+sXr3RlqGs1Wgbqb9sKik
s+u63eXeZAE26WwYEhH1oML/pJSTbffWUrQ3ifanDArxqtJ5DS3qSRTivnsnOIT/vpOtenXa9Qkp
qmnV7NUZXtHzjOEU1Ij/QlmxnrCcJzq/UBEgLkUNa+rdGR5M4JwlGKhNmgA56bCqCQdWJE7JW1Wn
Ob39l06OWDhia4+WVYKohDy9wiIgZNCnYnywUGeRBIae2xq+zFaCH6tWUgIDDvE4snFOYenJV69M
QVsDWubGEf7byCSvE0RbCR9K2osgbEbltRF4A/21yngTNqmGb/ZAFrXKXEypoNqOniGsMslO73u4
q/0zUik0h6aAGNAv2l/iIqmXUu57EdvKxh5WE/Mh+R48vh5Td8CUWA3QBXINLDWZgxzCCxD4xH4z
C6qAMoIr8T9Ij0HOu3h6nFyUgANnelCjGsvViM49GGJBCTxF0ukT27A5nOPmkrZy8eQoF7p+ByCs
LOGVq63eWumXN6D+9MoNWmX+epii/BhtPxuXh6zlcmn/bWpX9Xv3pYMgrVelaVZZU2H8MYx47Le4
jFNG8omDN9DC8A8XYD5qxhAt1umO7lg1KvDDYk5hiip2c94lzQdph61Lt5q87R8KPjPnLRsHX89S
HAVCpB1LY1LF1hLIFC281hzymBiM4s6iFAIFHaWHYEKs0LtZNvTLpwDo/vZUl1zCs+0YM0XRB2xx
mi2hPh2wfjUtaF/C6ttWVEwQX91QAUXtfZJANZtJa8OUtciTv9EqgjD7SfYvVtxQw5EWWZEZ8UfN
dai5qvI+B461jjOuYD/Gb6eLmm1yVnXExuqphf2DATxPQ159SvuiNlNVNyzE6sF537ihMHcOKL7Q
Utvh1Qlc5sPM9uQ2Nd6ksLI78XNLsM7bN41ZK0vdwTy0mNvjep7/mRImvrcFd4qMw2Y9w4fYk89d
Svi5//X73OB4Kji10ifjZ4hWzs1C/hcNAgGC4K8hg7XyORk9pCdi4NHI+2f25Xg0AZ0R2Fu3J3EL
Ug+bWYxaJGkGBfmOHITBGBq5v62QdfXvnAmquHnF9qM9XuC5h1au97VbAU3UyQ5hdBKA/osCIhXL
sB0WDlt3LhaDgEKcFkW1+zSxPKEQYEERo5uDt1llRpJfULIuechnCWJVWvGCwopMu8cqLfoBXC3C
8azwe/UMbaim81LN6ti7EU/fEevADb7QF+faEQhdtSoh4ETDSvSjilLbGGv3jLBWofY4kPHBIrWM
k+wJq0ePai8DLuhMrrLTssvVxd3weJuwHANghue6bJDhbZrc2hwERCewoZLmmQ+fsmy1okEqX5WS
On20OyvjwfMAKwQrXfgIMNn30rCQlUnjCNsfz2zFOdOr51KXoZ6alpVYceGzxwQqsILgMR3o72Um
/F9m7l6ziuC3INt7wuhucs3UIG8QDfhlkjcqk5+nSTazXY20E7/RfJBiKj1VOb+qHDuDoryif8nH
0orqfRMV6/BLU0bLwXPcdQyPpDf47UY8xBdvGDr9OSmX69dj+zK2zKh2yP9RCq0rCergwCx/MJrf
SN4sbxLsjngmpslGsQZNgGHZ+aI3fl/bYDLb8cSbe2+WJ9pieW4/QRyFH3jkxZ2AULcDbjh5a1z9
w3ddP0p9RkEfGbn8feZnfGe4iNyE4RnhbsNOWqID8Y9bqTHQo74I5V3G+88xYFZJpo1+DRzupcOY
SeA+ktFhL3T07Bktmi13hDKKaK8eIx++R8DbhPODYvPtXuasyEk/rKzbibZM1L6Qud6WhEQY2fKT
mVwwvToByUXHNgQvY2hxpJ4awayJ0Lq5y5Z3gNJ1FUIWQ76toBm/gliTKy3ndpVB6lkShXExBHf3
4uxXW/weYfngWvY8kYtRCSKuqH/LcO43vR8sdUZ2H1Dl9ArcDSrQVq7H4zFBQHWZiyGAtyqLY4wC
ORnwbVxkLmLe2rJM3FLZMkFhqELievhMzajKq2RIvPi9OZwMi2295mOVv9/SeX2DXv/fOc1wNmSU
ppKLijOJK3aKaEfIUTMFt9fhWWP+hbJ1l8u4854unGAFc6ibvEOUra2FjVFeRqj7LCMrSvcEGzbN
mrad45YQ+fzhRfL3ZlNPOIwvBugyL6keGxiPz7m+XQmPSj0zJ6jS46Kbl3oQprIfKAD73vTqdhuz
JD0o0BDEU69IMR3LfcDutcAweMI/f4tvBWB38TThREsnivqS/GvegyJEyDBOSQSBQzyfwHfKGJk1
LaDu9IHT4XnwPLsnJhqjZJNcegUbI4clhOyCPWr22tvFahx8mFutLAqKN9UnO/oyLeTHLy5tqDZB
UVrz7pgjw2KYP4zKNfXfi6C3VrZuZh/Sl3rI5eDuP96sBeIZg5p4v8vCfCYPAh7tFSXrXkheyWtU
e9CCT6SJbudhXh0qzAXUG6sRpXbIYo5PChdk8Nr9zKCEoqgczqqiCTLS7mpjvvxb5E25ut6q9DuH
9cGPV4EwXN6G+KYtoSJfuS4rXYECxHC7y6QsqLTSwcHGyZ4hGH1QFDmU6XS6QUB8d/eauQ9/6HMx
YNvz7anP8BNAftAM72QN1ULgZddKHHs53FKi5+9N1Y932Nu8feXQoQGuURwYmKRBOSb9BoPcUM/U
zVNyXHhEOFu9GO5rTprgcHTBUpcM7APRLTR68JtlwY/GLE3nE7dRn72mACzdWmUTP0KROW3IgryW
JFZqiiq0KxRZJmFjNuz0GvawDwkjkPHXv1cogkNmMmhf6yP6ocEiM2/k1r5uBSV7HoSGMq8fWOMs
fmV0KDpIZOLogD0CF7EeZ6HzZUf1KKZCsiUee775Sa1vaU103+vfYlzoVU+geiksNtY1Uis6IsbA
zbimV9BFWrngUU7ueg57qx3umhWpMHq2VhJIQd4PzjYzt7+NpwnIrr8RxtdGsVKHRjXxgt9NFNK/
yBxIy8GzupoFhBizHi2ri2TIkZQ914RRD0lkUPygkn7Hfg2COqMhlM2JqST3WdLMDxJ5cCwZTP/N
UGMG93KRKj2QOmRJxZ6/GvEeL4OszTUjWJ+5Dim0dB+IkJ2AU7BWOgNUH86GIT0yP7LluNmMVJLN
EQDIzhDKS8Q+r8G8Fe6Zb42Z6dwnUMW3V7ik1VAqQrdFClyJAWEOcfnh1GceKn/4X1i+bwqFTt++
uRWHVLhOh4j+ogTmUHk16cwd3L/FtxB8ejn6ZpLgx+e3OHYTE1jppWPq8vh8zEdzpP4wp8kZwZ+T
89GbiEoUcxZ65LmoKl0zjnpXOrFCyEY1wEXK54xscY9RmXNm0VGOh3bShB8k9QUj3YVWuUdEGXX3
w5eo1MQFnbulyYdCH+DXiWMVqU2A5p+agu6x5hjtBdMb+hMbTvd4txeetiP5dG86zdEgUqkkmKlS
Ww3ccc9Xfp3iiOCn2511h6O5Ub2oWKyU/wpjLe0WPl3w/cLmmo0EBIA7luvYrJ+RL2rhmcLJYjwO
kjJvyrTkCXS3gkDdF2KwSokD2yMjrmhPGHWJyqsay0SJks17H4Mq69Et1xOkI7i01Ra1Wpomj22b
x5teOskSjUVDT46/GYVbd9qgM4T6XzdZPslk01kirXCvHaiOI2OL8Mhc9h3F8BBVGH/msZAxPhxw
1oy4z6SDmw2LpzsEX/s5FQLNd/q1o0ZNc7E6FOuEyDKWjybnAmqKG4bP++Qx82bQn23sTaMKtlks
lH6dxwLyr2ihq7BEnMz+kgg+RogeWf1L+tvY0odtsqcXN1gXO6kgfTxzm4vZtv1aP1kRITUV1REB
kuuzfwbljOVMKFMZXPgOguT5F4nRWNDsySeygcmdBQLfk+GqXpOIatZiCzJwBUiWjWZ03sswAfUH
nJgGQa4oPm55tfi5V2iLvKW/T/evTOv79P5t5OFSM44cfe3lJQGdcUJE3SQTRoAplhUTRDfeF5kc
+zJfyeFNUyjS9m59xGLmgaRmbE2KgiTaNspKp2JnAQWR50x+e1U4Ur+DXnZI6ao5/nYS3gnBP6Hk
7geIYQYgE3CscRs/sZHvbRXCeIXlT5cWYZS6OmiEpCWTsUSH+sGpu9Yx7uRCUyQ75QM2J3UaS03H
OT120ZPuY1Mo6PnVGPL0e7m82Gsdhrrs0l4U6OlCkh2zPKRr6KVulDsKHkdgo/rIJf0zVJKIy8vI
tgabqF6xAtkJaJQxIVvcOa+jhfguopmPuUUB6aBOBYSOCsKIscsNmNH3MEXLmvGUzKWTMYiewoIk
7ILOzkwqJpdkv21DXMtQV39K8lM+VLy+oU14dGeHIr9vXcn6hmuYZCP88sI4y2Rw3BWxGMM/lrFa
OWklfL5nShxVZX3fBpdjcPSAc9bxnDp+jmTlyIbG6/FvXYR4iFFufz9Sf7aab3GZalRx1ACilsNS
c9Axwg+taHi044PyaTBzjfnUomY2fYwx23RqPtUqtcAXqfS8Af5/aCHWRrb/mzZeFmFrz1OC3Q2C
gtDUtAMSV57h0Y0QZB5YlC4eQlPXQZ9EKjXsuRWYZwvIhJNb3Glol60bH3TnVgyn3ymyrCidpA+2
Bfyzk+6PO4x+TKtst6mtP/wQlMk4s5cKzsjgz4IeJOdOXIDNAJAHy0Zrt72l5jyqUc92uQf5bNeo
05BWQkB2tXo07B2pEPE5C0+04nSwbq4T77shA03lfWXdQO7uModviTi82iA3f5T5DEI+mJIO5N7U
2BsJuN8bZkfWHbiGlXQAF7u8H9FGk8OxfH0D7iIsLQRlCrhQAt4ICEeIEi464Ju8q46vApaP5KyD
+Yug0c8a+SAMI8sYbFIFcCa2TldJidqw3k+jbyl8SAZyJzZyioA5+D62GyTSlMXhFBvC9aXuSXdF
iyntTrhxsICSshnzkFcWl5rs9wTrDCvh+996sePPLPCSEPi83g8ddjzBvnMFsaz/NG6GvzJjL7US
CNtOgvxOAwsvcX4rlxwGsC32Gllg+9fXvc2Doysep/HwZ9VpagiC8xSNHGW1RPmLL/Fb0Yr1Bk5B
6jQx9Fxp7q3oxRp/+qCzeLi+fw5tDK3jnAMMzw/3hIZo3BPNHYTItpM41cd2AErD9kxuWMvL9VHA
L9UdycI2Hg92dTq5dUo0N9tRXTBmv2Jl7HieAJ/VzqwC/LCFbGPFWANl/XAR2ppl2Qzds5i0BgjH
R6r1TY76dk11iS121MyzIcjb+jKEdNEYcVlr0ARjujt75EqTJEo+Xsj8BaNwBKYoHyAChyHlCsgn
nHZyigZMAu9Y8YbtNEzb6AZ7CAHP9o00y+4r4xcjHnyzCFxX+hUO+nfvndoaBkLeLoyCqY0nI4jk
Ct3GLJnQFjdcCiOBzneuwtzmkecN8brCQ9api6lZPHlSfi+1XIwggoMCEM54c/KIgsQA7+f9kNVQ
nQmOU2oGhvZBgr/602JUEQ72t68SbO0lprNFyVvgAeInZWZE8V13/nm+U2OYIzzq+0NakjNbolS/
NIHWgslvC6bj2frnzrwxEgbaNlGbE7U8bdukPil1TAFmWhOxUzWAo5jHn9KFAaKnvCIA/SuufN7e
sD4VrhoHae+v7tIVLPqBQvd2+ezb5xfV4qgjhAjbqeF77MObPx2NRGy9UMcCXGBqlswgj2rKQfQL
1+uzwXUelYx8eR3I9ffAh7u2zHLDgMASHkxzymwFF6/BLDSSMtc6b64NuohIe29C1LmQXqxxOwZ3
lhD+9xg7HBDXgnMYG4ii/JG+DW6ldAWuZACl0s1BC3X/EAglX4ioPWHnu/ueWrELsyo/uSUCBKix
Ev5Lbfz3aXETCiKs2xJVctw/ETPcX3qRDuomnNTdsgqFj14gTj0mkBCV623aCHm7ZkeERwC4WucF
PNVgS9Mp+BAQWIEyV/aGubZaX8rGOea5Z6+SA0eerNmDUJ1nr/GzSiBC39ULKWNA/UG+q35UCyso
0vnHds2YkgNkr1c89lodTEBMGG54AqcJVPRtwMoWpYhUwtazFzvr5WNcUzAlEE3BE9nOw8ikephE
5g+vkbppDsIPrVnrDpguJwJeoMh/Qi/KrQF/3jfGEygwysqBY4IPpoI02UnMbLHTEyrzLUCNHo5/
EETEDJSZf//IX2VaNBahhf3te7ehwadMzoqvncHelofRzzyQiKSMqtdBt77GrZZLKuEj4FUGApxc
k4knGjeRTSC+yRsoiA2/50iozteossNS9XP9esSiS2c5o+XUBoPJc+vOpwfviahJhsAVuUfUG0AI
h8xaQJqZGgG6Ybbezk1LguaylEi8W5tqY3evenbKR0NNceVEQQP0+zgbCyVTWmcgvw+7VPcELnPb
gv/fxEquA0xYPRb6U+PGMhjnIhWDsVIJGJC8DISfOe/rbYSSpv7mEmB5PlEsFeUQBXYH+cZFZs9F
Ymsuqrfkli+ONRhLlIb/BZKQ+djTBIvP3bHz9oAxavr7aXAHttWZcKyQy6jPd5w63kjdskoLYXOx
PsrDK5wpcqTG7kP/hKvqZatZNn7tZf6qbjZgx+i1XwuPyd9noJxxX/9zbt5j8CIBCThgTwWxmSx7
G8g5OOJi1A0DZrsBY2fBgsTD4GGF+GIbHYeRZitquKdsbfmNpEnrj3aZHDHkrKdCf/sCY7xshjNo
YZ436w/aBpsrWzYb2rTGYNqZ3EhROr5H65LJCvcQgoez6NXRiwXzhJwn0uJDtsf6Og1YgGaS9Wg2
vLkHy5iCzhinN2PAet1iFgnMrR2uKr0Tuh1HF1oGpgC52pkukozc3IF6KjpzcQ92lOvNaO503UFb
iRO8hADO65eX8OStW64UAJGybJWQZ7twm8OIsoYcCzix8L+o1iPD4s1Hr9vOhq+ZGFlS/HmPZU2X
YMaFWj5nUDI/a6oLU5SZ5hdLwMJeFQe/Cc6ypHwsD8uptiuOtJlYZOoR9zUZi/vcqpu7e0aS9yjh
HBjlz8yG5daSxKGdC3lSDd8oCBzTKwGx6+QQoBYD/oyHcm2VfqnrE05CW4AQxTWsxV6Vhu03AIjL
YKaMKwePIVLc21pG9360VI+uZZT/MC6Nj7ggZXL6iQKKuGd76DqOTUG3mS58AQt7bLStXm5cpahg
LcKkgv5NNjy8Zg2j/zpNhK6gwGz+cvE507CRQhakXc5G48UJw3V0wS9yCqtjRmdZHtRAbjAIVgbl
U+RWnn3Ai0rAvrKwZG/f5nMDlBQtlzEomfLAoRuBPTBlYfPYG/QlwTCxUuQP17bC45LW3Pi6GkQu
qkRtUBt/BfHwcb41OfSFUIJIHIm4Rr/1+VdxXAkTAqC+Z0XWa9k6Qq0pDf0TZEekUf3YXRKt7rE9
YCO2d/zt6nCytj4MuXCDzMXLy+GwMw1LQDLrJeilD0fwiHRaYaaoMZS5sy2EkFu92DYUbdydSnQ4
0k1ymDDf5ZccXtC2tjmsj4Dqw9sRsPaTNgxbe2SUsZ9uW3EJCjG4ytGzFnsfIyIrPyVPDplE+mmc
VqpU/RcQ9GL8K9l6uw4Dk6aqfkRvZAdtuyTlvdigsdQHyXMz9etOiHIKO9wo0fSM6P0yYg4vrzya
7SXF4rn0QdigfDkmids8PEkrk96RXOUPbysBi28AEJMoPNo06TBpgxUQS6Qbw0oWXCkiqlLiHUlR
zB+Xe0myKDdSBXp5L9QkcZtZq3AdfwWbXeIwVXbkLHDcKv8HMrrho6RchBWva3oVXbULUyY22aT1
KeWVxdaghwdfBmMaOkRf7KQexMFFD3Ppp5DAk472Mn/1XjIyyEQWoWZaIABamCkjgtLmIIiLgIJn
Z9P/Mq9HbAWuWqYAU9q90ODwUEjeYJEwvskTLY3LmshYYLc8AmHHSxq8plenZDUIt01iC3DWSF1s
ugnBxLLBII0zMnIYeJtWQIZZyCwZxNS65ic0IvFweKHraXXOdNg3PAM80Sgc+kraSb40Xjgu5NcE
p7hAqDvApmSFAMlowvkJm/skEHjgPetN+qSt+gydTPe7eSFgvs51W+24GKxnfDTdckSoQ0ZszWV4
hCD2eodtiEXB5wii5e1WWCntxFbG54hR2O5Uou/iW13Jtag9uD7PdziFxA9A+qR0DufLHn02oS3q
5Gf/zWf+m5BuJqHOGqinfx/Gg9ouwGrPG0aEcNQJ7/ObiVeOH2btIlCNeUPe0dLCBllbqvwANrBx
ufEeaoQOlbQ8iy9aLKe0K5XE+60E7F6rM77a/NWDckO+AgTPTNRD/g2IUffagT+F2kQoH9ir1V+4
rCyyy+3CvNiBpT6EF0CNVorSnsj6OxqBXSeBb4R05/XK6r26X+LHg6/6YgwTmiHnN5vjESJpYBkO
S8X5R1+i8jGfy0n2o5NQNS/66AceM0kye7npQz5YTEVvcHFiGZJ25qXfzFFi+4yPA2X1Vaaase5D
NL5Rrci4oEFb7VqsRQGRGSjxCaaSkJ9MA21fE7adYVYSol+/loFsnBWCJL3+LA0frv1R8uWO7t7Y
jfvqLUbKXZE6KKqbjzPP88/fLOuemhguBtx7eGFIVuMiLA/kEim6vUmCywtMbXNRBJik3ljM1zcg
0+9ToVvcn+2btcxZV+E8/aoeBU/01XJLTtA50SW5AnZWoDYJ3jw47ThOWsOedxfMSHwXCQTy5Aip
23j6jSDuC0CXk4BIKAa+iDlwJFFwcBeY68jSUuhlE4xrU0vR5c0E37XTLrP5GNchVOacZVbaJp/a
Wr7lV8A1ZzK5+ew5BZrddrQXxNfD6kNcduk+mx3fBpQdApht4nySKhvr0m9o2DBa8lHCkf+jsePX
CXHcV4asKR7+JFgqr5hQE6jDsFPcAEcl/n5N7IZXMDLgQvUkntB6t4CDVWfzBjqzB0T/HrZ6ZhbT
OrHQXeWNCwfIbENeiXQoaYfwJbTSiZP8wUZflBfejZn4+YiOUEZJDX7DB74FCEP6jKByUDeIwZYN
iVekJpOye+BASFOeK9NZhVyS9Jis5/trG/jJniTlmSJn0Q9vCVNd8/JixbW5zYBul48ePAFjD9qC
oCI5CLASxXXeimuO7LsJrVQHWN/gb1Dm2Xueh0Nm5+cemLgDs/pkYvBwZkiWxVo1vnfvwaIO1FJg
Uxt2hYf1WXSND6E235UMyuxzn3T8Qf4OXXcdkM/C2GCY9wEXo2Cc9hSoNPtzwdYkFOX8vzs78igf
tFLLgMsrl1Hs0Vjc/Sznv92hOF9Mr5rwKyEsdwDsNo/um5wAtRNDKek2axr49hx50CN5mys5+ZwK
hDI431a+ivA6okCxMZh6AJUY1CUshnobozQpO8Hi/l4+96n5K0evH64Az0wmRKUHNtJnlUYH53am
coZD2YvJuaKXP7kP4wmLaD0o0Tx6xTW23DiHMPTGNePdCt1rbNDI6z4+PuuUsE0/GeNmY9CoRh89
WxQHXwHpmwS2ooEBoR0VxSUeCzYkuId4SlXHIOU/9i2UfbfNLGiQAIBIBpcwvxi3NGDQDyXM1ojp
O/BVif2EIbY2dCuF5buzZDpkAMLigLkE+76YxCwNn54EIEcKrqjhjgcIOghVDeTd26tSTFWbgDlX
o761JPHPwiH2ZpCHiUkBTARNKxLJEFIOU8lFYDKZis4m+/c6SbVDeo6x+IT6qT/3wubog1UdkJXi
8dleT9tC69N8/sy134WpEKrmADF8A4KIcK4RgWGdqGmmcpk+bMroMcs9h1GWP3hwuCMzAr59V5bE
fYubCkkt/kp+mVpWaMj9OoXGDMbxktmbhhn4FObHzXNCxwYPMvZFqRGOKUg7RQSqazu3tkVOCgrO
Wq871N4KUCjPhX5svg+VFRCRh0EgzmmOQ09zZ766fxHEMYWft8FCiMunSQ50f42Tx2OrpfLTYw4V
Vc9/It5XXWcoaJeeFUA3XrnPDbgZpOm83xmCxn6mxCIhbY43PbZxtec+kyVDhID+fSAt8AHaqzz1
m6zmCY2eKE4ZnzgPJR+VdqBLmZ0F7OlnNdyY4juN8WRvUnPlin+rjb64KuxZdKz5O87S2Rr8Ff40
xSdoBgVSjWIHhLkty4tCl1c6ASlPGv+J/4sWnJWN3GtCrz8DQqzuIUFBr+tGGHsThU5mPPC+CSAu
6J2vS6aimlAqisAPAvIlrPesYQ69JAzU8gIxzztzsPjHCNedo0BWmy56OQOlYBx2zNL4rjVzIeg2
scax8yfFRAMc/ouyJVglEiKqU/rp+8EvWrjRx9yZ23o1pjQeQ+sPrX1zh+uNjnbdhGuWNvCwnOuT
FxhakD0duA5FrXTLF725l50No7W76ivtPHHSCfhtZKre6B9+D05TLmngOYqDOP018xrNAE5hjAfr
l4xdH3u+85GElpgGWfaVSFXDjwVirqNvJx+k1MmzYjfVsf/bYte0PL5yvATlGhRT9X9le6XvjzVl
603pORlAHKfHw3y7ZsKN9yynaFrkrg9Sfk26i2o8MYhPTovhi2Ra6fJ1ysXglY/17fCt5wjuCcdV
DzxRWANY3voqnRWqO9gIV4LWQkcQRC8wA5Ebj380lYAD/bsXf23Fvjt2slUNB2Zc1DM0ihVw0d2p
HmJ5wZvqJeBHej6N78ByGOHyWh+xWWK+lHSsqYpc8kLzfvpsYVmQiVNzGNA3Q+aGk60Y/pqfgA/N
Ofljvyn/qkmybqNSCuR6uIx738uNVaJzicPWCfJIm1DmPhlKOkMreL5b4OH4ZnSRTWh+7aDTmg0u
61061txsVW5jkI7af9xMf4HLDHUbSqniaWxPAjmksTA7N4cxzmN+CkQdgbndmTH3WTEA9QrmfnOx
ptFOvDaeFhekigNjqxQwWY6Q6DMUekedDLVgAxN256FKHIAxFdH/RImWn10pwRNGwVSbRYh17Feh
gEnQBe6HO5Ddia0nV2V2dFwjvvlj3lfW/JWOulPi1MBcQTWH95V4HrW6Mptj1AA9A+IeU+VjOLp8
PxhrlSaF4zQi11jRzwipJoiKRkkdTQIOQyBN36gkmm3MNXqjMM1KJA+KHk5PrRq0CXnYOIxW2A1L
W8WkLQM5NhmPSETDXigvgSe2wjK/0iHSBhZM/p6wVxMBkm3CwrpIXAn492g8mZNPMv/VDt6H8j+B
vA57qyQuXA6bwMDLlXBPrDlZuvwIQinXtJTRyyP00hwTfqUMUJNm36LzJ1rjuGN1uOVP2bLUgFF8
+s031I+c1cDxjHv1KwyLrMRSXUTnUWjkFq943owcYr6gZYSnawQR922QoIk0mR6oWIdHsJYMN8sG
M4CFzKEuPt40VRi6eyLh9RAT4+qT9N9kNynVgvWxvl62SWOxL1SYhla6mGIRuHMNL/FllXFx8EeW
amvHJkxVFqoKoyJOHmOwVKTHnk8NeAEAOTcMruZCg7GSjjqLysYyVBrGCGVZjSI0hAWjxPyFNdMt
dk6ST0OGfPg5JGIuISkroRp6p16p0jueBQcVFuTf3LF505bAqIdmztfgqHXGNT/1xu5At97QGHlG
tvuNCGE6yzmXjuNnb+gEK/W+wWION6BfOtMrYA7YPQe8/+vIVjcl1Bv3/FVEG37ujv0dExrxPqFI
KNPYXrkVn0gg+YApXIR5xx3FZwcWTJsowYMsnqY1VZoEr35T26zFNs+dkizVywdhyPOqJSLa/TKG
O4xMiga50DeufyskHvx+mhIs5nYu4fHEmoTwKsuEqLj1P+gi+ZNH+eGuMj/Pw2h0yk5xYMSo4MZS
wwRQmGei0YPeyViNyhz+xQ6XEetIoU8HQWzgkjlU4cGdKogc7PlbkREPKBYmqHiKely4iPkIH2Dl
PwO/dFbtw+MKE04ZSEvGu6z78GdeM8YukxrGqkKhcDnczr7lSQVwXQpBc0adlkcrKLr27PQQv/eN
QVMhK8hptR2PH2rbsmNxI9uS8n6V9WGdWaUpkWS1cSp/Nnvb55rt6ixH2h64FYZJiQD7R6ie7bJT
0L6xcVAUQctXpBbLLtyW/ba9Pf2fX2eMuBAF6/bh39EgU+QMMwl2oykQvAZ94zlB/7fmsn8HgDqu
lfCAHEP7h4nWUUaWmjarMwWumaSOaHZkangovHWqmAu+einJp7j4JV1YQHBsHbz6mTdy4w0P67M0
jNKEZaZduGXlO5+Sck13AVhZ8z1oZMm51mqLr5EemZCuP0RaQ2kTg8gsDi/643D75Rn2YcqHMYUt
DjvakA8DM08umKXfshDF48BkmmspipDQ/i8aK8CaCNx9ylqFF2jiM3RUz1Yz+YtrhdJ7h9nf1Anu
hSssgx/dAIL4/uWmZJG9L8/h5LtLylljfk0vzIP/+M86AzsIgIAnbMDR4u8XFYWam2sok3bS0iHK
JNP2wAO3jjZLflCoBIjjoRo0F241tMkpiCl91ZDVqZ7gnAj599ikrQNL5aBTbmoxNHbPY2Ai1D9+
aTCyRx+m+XcY10M0hgAZOehC5wIYwYUBPQ97Fd5oYOa0pJfiFywQY1wQeOom2tfi+B0rBQb6zNrD
I2GN/aS9p7PS9KaKshYmcT18fzLl+QZX7333ldpDQR7luZ8vrJm6nongCBquuXRCwZPmQDKXUMRc
Ezd57Bt7E+tFxiL1crRbqAU6x1jm178Q3NO5hGQ0xkUkGB4BzE5N5PbITCRzZTvB52rh9S/vid47
QH2/jrxi0znJPjmHax3zT3kADaJWQi5QkyJh5KQyPh1OOUntjkSelso/5O0pUoi3LAuAUWRsWk6F
hkI1t8oPlwp9EYAtBa8TgSTiujGgWWa79vlLC6nuSb0oC1QSvMWXTTHWrs6wW7Ay7IuCXtMUVymg
TUqQ3TQk1UMCRaLwpZR74u++Bkihdo1XmG481IaS9IbWpSPM5eJgfk2NxYOOayZvBxDhe63ii6Q3
G7xOj7HntHyMayeFekRU/9Z3sZXyfGBU0HhVp8KIJKOXfpMZmTDYFwSHArCM358OMqWOfinLRXDL
oSQOXjxQZWbDCfW00Jm7Ir91Ofw/HvHVb/w484a7YXrYjRPHDKoH3NprjDJBkwoBSJjCOhid94xv
5cptHMhyt+Zup573a7J4POMpwHK9GE4fNgHgxNrWvHOjChy+nf/sBM8vpXQVg0oC79zCZwc0W+Wp
3Bzy2UKoZzbkAhVMKQ7bTRfGIcP4GA0N+wmISe8XrNvs05TEUCEMfvmxJlyq95LAGvnmm4np33Ju
ujtPkz+TzDVGuiafgDWgFS9hmHWmSzwvqoLWKn4QklSAEcV2Zh4ktVDRWHF6/kRwAk6t1K0LFM98
H/+pYJWf3p16mnaYejXKNtuETgou36of0HJNxd6LeTbL3PwSa2dUfS2iLQaZYZF9snsIjC8pZVY8
dTmJvdBLMwUr8bwMzsLwT/1Rj9n2r80SRQNmtW/50vX1QSys1y7GAwy7JrkKa6eBBLjRG6DH+uwP
XN3fF1367Jge12l1ku4NNiN1eDIjV1T9/q9aT2n6BfVZILFaF2aZZGwSj87nVdlolOsPmYYAGy2T
3HKVFmQJrSUXWg4+opgT5+eB5MQt1W8T/Alt6a4Mvf5Hni4BOehpqM3ySq3yuwAlz2FQn03gQZGw
CGcveycORMlNJpGS1uHIJdF82Ejbnrwe01aVJOzSRHoyhemUlWJabFblYucpg0yH70SxZaquLCgz
fehfrNg7RxhRg5xX60rS4Tx1PrPlOJ4nkEB/DcR03XLWefr85VFI8uE+kUnWI8xLkk0EEtm2R7WO
vHTJd59xm1b5XC5aZ4uBn+EayVJDx/4C165x5+nTgV894U9+swucEs+XNP5AfCjy1Epl8ebq7DYD
XElof8hBLSIu4bCbZFpZok4+TaGZadnU1aFQDIpuHnv4OnnxlfzjhFY6rfkVvZuDQX6+0Q+Od05L
m0+Vhf/Skuo+klYDQNnhyaN2GIp+ve6r/SuGy8IEgR4DKvXhZJhkliIK6eVpSyr1G/NVoI2Dkx/o
wj3Ibm687irb8ll47Gdy2T70i5Yb8hoPFrtYoFg/vGfavLl6tSKvX5yn/Zr/mpT4+sxZuUHaS9QD
4idHcKFsNuWhDciAQr18iiXIp+eT3RQx3TsDLg3+6czhrWc+dgrnSZjeTj8N2d0dl0brQQrKX36k
ts2kbzQQZ/gNaJL+ZA1B6l16m41xW4qH6FBK/kaxVJyhJSEMQiRZwgLG6PffXDmodkJHQvdV95P9
b+SdSfVF46oRQqn1WarPmArIn0NNZVvc2Ldvu/XOgwuK84/+mIlTITZ8xTA0MFUJjtTBBS6Ue0wN
HM+99KGfduxtpcaFW8ZDpHI9v4XpONQpaNx3VPdgRM6tBg+CQNV2mC/72wP35fSild1j7wgv9gpT
cRyyBytjh/f/UoyY7SOBa46yvm8QKMtkWkeGjUpupNd5pGOmJ9OtxNoc/Px6ZP0XlSZ4bm+SFuNX
3ysXArBB5ljmzmeJp0mpvUMGZivqBild2YP5sFOq5LN1JfTjFyaaCb5i6W76AsKZ7IbCh5ywjvxq
qVCG9aGpMXj7abYOP/haLlzdg1O11RAomU87hIJHao7GqMyrIeqnu0SeGzeRGht5KALJFIuz8wwJ
YvM79mu4n2wg/AjsWXvLapo+CSkZbJgx8zLAzix2w+Be3GUZeFhshMa8HFhovch1MXSh4KJ18QrE
BEKeUxLm2En2f5HRjTY5+FrR2vpDVorfx7hUhKDiLG+ugHEb49I5NP/A2zFYgbhG8pGJ2aHVtmh2
LJJbZCfNd26hHirbwX1HGboABU08VA2QgoRHnQyeyskfUIQiwFaRoCZoHDphFyARX3bmAGDaqquS
ifuiKLHoAHeJL6rBc2+V5JPs04pVPluNKVg8yKh17Tna+WDw/J4tmVF/ti74napyboW640pniV1g
r9T/HuWd6qEVGwvv7haiJVRtFt881YWGZY2Mb4trLnqnEIlfMXywA0I3Q8H4O/l034oaskNpi8BS
/AIZ9SQuK+l9+VJwJgqY23mrZwjkZuTnCk/HYw1rFhaK/H6Yx2IhBlDVJGDMeATAxyF0qamTx/ww
fNOxXpTKDFZbEoslRD1b2gSVnB8hmWVwEmawGVw+jxOFGBE1YkaRHwgbthl6EvUs2Z5qKGKvwTnx
kMmJS0Bu7FgR+ZTEUd2zAc8MFNfB4vfKWa4+rwdjnHYwFdHayel3UEg5hI4f8NM0liMNDxQ5/BdE
1ziFoonHR+ZWvHjIxdY5lfWx6UQ36PrlxWactF22y2vauXDtuS6mDLHzYnFlaqLUJxXhhJITmTNK
lWTLrR6XoV3Yk0VFQ8Y4lrl445GVi9Huk0pCkLLnvwiTOhwK/F80TO9fzfxMVfYY0yFaeMj0bV8Q
/QzViS5MhBi0KIr+NZXss+lEWO5lPVjq8GrAioN+uHeWPCD4Chq1vCZLAN5/X5B6qy9nsRfe9y8G
pXnekRQGbL3nq8RZViQpmleR6LNfg6nCfXhUX2NHqN22A7DbXsxG9pDn1qg/NXYRupDvZ8RZjMzA
VHiQ+xsDroyqIY9rVGWSby9wK8Lj4aJ8iNGSq9H+HrTMjI2AvfufyS2pYwh2LZ0zmq5CNt+FOdTj
kTpsonfWGfjmVLBDlcnc9gmKST7f48wJHF9JLuPyrcGkWJARvzU6VJROwCzqCoBtWwc9n9KWXjJp
lh4X0wq+X4hmQLDYIlAmi+FBIOZsELwiClQvGIg2lwqZZDYLfsK3v/I06CfpLW9qAc84UpWg8Z8L
I7ew2Wp1tDGdfa3emcf8kZSUoSsOCZYYved0tnQtFyj23l8pKFFpMejhnzd8vm3hHqS6JN+etmI+
b7TZhupKEer3U0Ke/I7KdhObVYQ7xuZP1B0NV04a5jYvYM09K6T9EvIFFXYOe82Pt0kL98wAGTAQ
TgUAqqxWOA+Peg6RvCqVL52NQ9y8+SMHVZ0P1CL+1EydeeY3/CxhgzY3Q+mdMeMEaNvEQRtlojfk
XvhLE0gRViLsZRGTs4sqaHHSHyuoy5EkW7P1BDWauDDzftTJ1UA1oG9KVc6vU6inAr32wlFO3ePU
ha6TQy2IDTqL5TS7fwzOjW9MMxtDVvP5AsTM3uw9Um/NRUr8/XhbvfbkHImXlHUIW/nixgI/jIzy
xfsRcFMSoz7mWNWTVqJ1D5CukEv/ojtyitP+3KTtb+2f4ixBI3+qg7lS9FQZ6ic4ujgPZQbEd9X+
vIW7PeyqUigOJLqmo+mlSAcS6Mg1Zj28a8tqEkywmfvRXjr8FgRHK2+zr2SHu4VzEUyufB+7RL7Z
DcU/ImKhzymuYaENBi4a/GImXGPpJUhlMKvJ4rjqe7VPK3QWs2eqhI5L4yIiQmTRVsQJuJTCpFOB
KwnKx6BpD4J1hMXtTrad6z4UTS6POj5W8sXIdxhp0Z5xc4dYeDGpRXxs7Vk7aPMPZC4XtDAgC0Kl
zsTp+yIL/k3Ao4SGo6WDHElTE35sLMUJBDQ+mM8V6YSPPton19ZgPJVAoZShtIvR1J+/FUZS4CYF
vdfoth1N61V7fLHxPaf5IvOwj71i+C2hvBLNJ0nj6WlV9vIt3DcKfXx5R9yW2xfL38qaZMnKFkV8
9+bTB/c+pBbEvnEUPt8pIOgtyKGu+tf4v1KbWFbQ5AJvSyHCdwMrtRJeLODyK26cLXP8ZvXpSDpc
TzNquAC/lWQUfW2K6E+lQPsHdwnws5OnRV+od5CZ+1muvNl5/c2/DTD2Zoh9TW1u2OjwoS3rwzNP
PT/0qbIU5z7NZLHVBgRh/C7/I96BnWiwXbpLeSfYU7R4ddHadyWpyxK1i+QhRJ69JfbMSwTAw1pg
0rd2ZPSX8Kp8t+JN6Jrn8+JT2TMglAoH49wq2eqkvgMOMKKWjdVZM507+KNvJhJdBICtHTps3v/A
gES0f5huttvCJgEB1bNNMkdjOR+FJQlu+1BXcu2hv0ao1/Cvi6DPDqPXGZL54kXmF232UxBKJHvg
9iv+FbG2HhXS3Ge7/cs0KpzosbdinRPJhLPBS0rWOubcgzB64CSJmsX9e+mk2Frw1uu47ZkoYWbc
FjsRqB5/4CTnkeMIRx3UqdKYb+LByRtHNwnNpSTKfpdUSyeZyUal8TwGokSOOLFKsjothVHNuAHb
5jIo48jKD44n4t5DcQfnRVAGyFFT7iMnsa0CNZ5FpTCXwoIuDdyR+YhD5DMC1P72VTN9VKASTQlD
y6Nx93Th8tp0QH0nDkeKxYGRRqrHMv8hrWUKH2Oo1hGHFAkTTqFOrDBV+/03j3DdRpl9IJKgc31Y
nh75lkz3YJU2w9fOAMsS3p9bmSIlfC/39lQlGwSAIcARGAWzjN+3KNMMxClz9weYdgvVzjhkZS2r
85i3Teg5HiptUbwKG5jVYQnq7mtDKZ5AgRmI/F+LYIc/MvGUMhDz53kzTUtUc5vq2OlVvTRJUXv5
sz0PzmyJOyZtJxtHxC7S+cC23r44vn6NP+sGni6VLl8g4852a/GUYTmd9u685hrK0YMxwKDm5qSS
FaB7I7QC8WJ2krzxgm4v624FAyT5gV5mavnO3NW2U3XW9aKYCflThO+e5cZ2OL7KOXVchmQ597YX
TQpVyNFm6C47Bph5h8x0hcKHy3k/KD7MSvRAFpzqO2NY5D58dCKdAn3k2QOFZfLkuDJQKvY9C6hr
sREm5/IEit4c/ljIGqgXnYJZHaXFnvdZjNVqIDFwRwwobbnKNhN+31HDIAxH5Qer/sZ6WrqXD9bZ
QzzqoQRxkBRMO36izzZAMxn+CxoKt6Qy43gojWKg9G3aFr/ulZtx0nYrAeqXm66k+LUh7R/gXxnt
jxa2dQTIZhF8UvrPtoQrmvVeqFqres8WaeyfzOf6/EgZzFcjWzNnSkQL33nnDNl1Zj98+v8zNFxo
WYTrcIFwv8wlDljWAsCRwnFvDrsFDN0WyGJH31zCPWPhPH7ikhRQmuXI4utaHx7hYjcwGPCtgXOR
EktPaFlVXYh3mve3K7VpgYxWluQqyY8mdpEg/6S1fFTP4CiQ5ejIpc3mRwSxm8LX1rQoNViB1i2B
0QVjd7tUrTkA96JtgPg05oIxPsn6L283iQHQAzb2k6T7xh9e1oJ0zKI1SxqyVxDmu5HX9I6eOZjV
m7kcU+U2h9L0bWZXnNNDA2rym6p8I6r8unurRaiyNESWPl0tqLxqc0sqjt+rHK5ymKCsxAgWhNZx
8XNnk5j1KszkY3Ts98AfrrrJrSMV4lGp/I9gOOtGx+gYU2YZP/uvyAJaDSE2XIy3FvasnKBd9Z8Z
F9d6Nb4j1HZYgWXJeQocCd9yY6e7yjnpvkN9+xv4pcV9KB3pm7c7RLUv6dIFyE3oH8xhe+MAk9Oa
uUCqU4uLrYhnlhGGbcYZ5FC22DhBHmdnEmimZ1mNE48h0Yv5QT5tUHkmj0pLIx8/6WNCO9S6zZCd
Tr+R1GwdH7OIjdVRz7seEV+MeSTexJ5HXs6TF7p4NX2H426V1YvPoSPfm3+MDLM3JFovK0D75Z++
IDKcrchnBE+LUXZ9uLEn76rvcWxR7aWr8KWGvYtchfrGsyrSgN+lu9q/je1H1qH2qDnbC005RVgw
mi9zWQz4dEV3a7ABH5+T/ea2v+LW394TIApS0xymNuxKhvbmy1RXjF0T5TaKywHbEbuy6+cs8iFS
WfP3wrhR2zETqJTX9Wj8oO5P+LKrJkHlbK0zKKZL3gnAaVWSmTA7DIwNEbdPKyOJEzbV48X7Sgsp
JhetnKXWN9uj3pw04+wSGRDxzBNepGVK56od0bzPTdBAvqGmtJYZaA9FrDDD24S4mX6P8bpj02x8
fV9VG1l6BL/RtfQBuGwgp3n18sq7qwWXr9shWxHGv4+/mLfe1RuO33yKSOJAKqNZS+Q+e2clleme
ObPLfDqeJaEK1iVc7MmnVCX/AT8kXb9SW3tuwtPhinE4DD/lB3bvmWOcSWrPnL5es5OG/4Oa27CB
JqFF6hbSpxTmYeWq2NIG7YVqnEvppxvMyTZd3792NmyHr/+LKkUeqpIkbXYw1r1vl4A3hC8XNkU5
kKnX2iQh2JBMqxTjqQ6kG5juzUaH0tHGwvjK6TkHiQwZNq218VnpJ129Vlnxbsw5yxxKALRQVzDA
rHMNZk42Y1wwhPOmRiApAFV/o5hr2afsYqzjcXl22fRjgRkiAOAGKXPkSbAV/16krRTjs7Q6RnbL
lYIxMz5vfas+UMiro1dx8OFsJowIt/3VpiSHJ27JnlvoVYuFE7B7TqrxmxwcbAbiOLfylU02xtPW
tezMpk8R1cDipNJtqZwvSNfYwBjKYwH1Xdr2dWX5OdexRwGNZPd9G4v6D/A0Qy7wldt0TFqTsVbl
3dwWV6/qTuzdvz1XihevTzAngmleMc37oD81Tn629IMAhFAm03atm/L2ibIEzCBrwF7fyejy7k0b
AiW2PfBayerFwJROWA2bY1mYZLG24bqL9XbQy9b/P10T0EnbBH9JgXf5mTk8dbx8GepjmA2AZnu5
oAmbnUAKOcPaxhA65tiHTHDnN24bsqmT5Y7tD484j9yaXZsH4UOLO/6EC8bFtlpWAGMdwxu7ZYKr
TkHzONhQUyw7qPGff84vQIzLSmThD1rGKBQkYEnfXwsclEz+kgnF/R9DDEVpGu1Qp4GIVpm7LjMA
eMG269d4nWjQrURXMkVNByH6nXeeGmhAQ2vuf7PsVpnnJGraD+CfB/L14PoqpNV1MqKT4YfwLGQW
G2kGrhG/X+kIn0TA3KJT5icfjcD1W9zCc1ELnorYwCvbGK7eFZsLsLls5esC9yvEEVOqgbSbDy4a
cPaXY/vlhJe6fpe2tc9GmtG1M48rij8BJ/T7KkrCws26u1jQWqK/EhAI73mqFgc1FgRfMGtRMohr
gWoJRnoVFtio2E9AQ/YzF8LDTE96smnOuBtnWv54t+qA9/fxH92APJSTrGelruc8R3rbwLo5t0ZL
nV6atobnqZguUfIFnUeWuFHqGUJZkBejAUR+xRIfJsz0g7LZK/y2NPtVKGvxrmUk2gjUPoahMoog
fcWq5L1fQ6bKXWxfNyqsYkc1YDPaAKGs7G4jwmwckbqsA+UMQxUl3NNfaNuX1D/eYp1W+OxL03wF
sOV2wtAHJ7IeSnTnpbsAeeap636/UHIKt0ioOAQt7gawTAbZF4iiWPcTZ8fxYnQNFFFqXbZY3gM6
+cwn34D5MR4T/ApuX6bFI020bI62SeAdmOPIMnhU7+MWJPxcy6QXmjC1MWU55WIeOtU1DVB39eDV
bwM32xOdyvk+3xmZOJO96EBLMR6XYbpsEpa+rA2CyLaBffUc937jALIzv14tUewg+6mUq3psbGR7
MJ5L9ktGjmkohZ3F8THNLzVccp6xSQEM/lDhe2+bo6MDiMJ2SCXCv7MUr3rvATQ4FXfhiews3Ufo
NnhVx8vmx9/FIBVBayC3DAisBD82QO2S83f7X3SdjW+jvKtJ63psy2A+/usxK+qHbaa3QwKKABAu
nUGLnpAPNZfTA/0GLsEkT+Dos6Nru/YSafUVJJAeQUeyb+J0p29qzh1TAj93M1cNGsM6pflpkgne
T3I5ui37aUJMHYJhwRKIQoEQlf83i7fEEyp1p45F2IT4RFqJN6n3YsBB+cfuzDyWmKn7wmnOlKGN
Kxl9QLyjj+MIRnzIZlgus0Pwiei+DVdz8wwY39J1dDT0YuHv7HWH8akgv2r+dt7s4tPgMk6oHy0Q
aPif1ukZYPK2sWHY+RuKYQcilovZLplv5cyyBbFwJnfCa4n42uH+IRqF7JQVdbCgZhrPHVKB/If9
6yqbYNArHSARjUDjpw22NLbmdikGbAW2RMz7S9QaECinfy+4MsqQJ09W0N83LOEEtpNjKFnVmVMD
0Q01tBgE/lhPIUwjI09fiiq+J7XPz/Z41zVU6LZo1INoZysxbt1wQ3lfjvVUUQ1MGUxIkD0Smqeu
U+RCRp/JHyEfvwznfJmgD09ojSvs932328gQYAJxBrWOQ+j/jfV16zgLgziP3nmlb9KZZR6trdi6
/+pBMVM2sU33y7S6FgMgVdAw7t5Q/kwUH2LxDfPLhynKkgEH8TdPU14oCuCqIRuAZ4GJYAcxgnie
HjUxXufiVvGFdzT/nyrJDYr96hFAmCmA/mousjZE6tp5yu3fbWp1+sriVw95mWQr8bfpdJO7lcaq
Ix4M0tC/Qtpd4eTaBlX1OWxhNhHJjo5XGfab4K/E33Gmp/28/OLOiflSLj63PKXDuDLACN+1WTWJ
09Mhm8pIzQAbDKJybMoI6FXxZmMtEndmH6lLwAVwhh7bICuSSPYseUhA+A785BykATeMfX/t4dO1
ydA4co1WR9gaHdHFsa0qMLvYhNGzSwqEY1887p6dhvCh5uycIqXdSIhdaxurD8CdE53LtwOkdY9m
t0s5tyWvtRfeX0jLr1NnLfWD1unySbDWTYWSnRTkjKo980Dj0xEVP7Fl/zrg6az7HoIYUjklO7de
PU8ziIB76XI/MirQhhbA3yGw0dt2XDNVeAjvBCts1qaGFW/QXlbJAlyy2A/gCPg7Laf95TIltD2x
Y1hF8hJX28rlwB2XdouplMpnIGyuRW/+wwLxseyENWTusiyhktJLoJG1E1tm0uLDLzZ5PM+8Fp2m
RTAO1rXfOK51IwJ3gGk488dT5jkP6lj5nvWErg3J720qQI3hsfNkTVTzMLkLxgnaZeJA+Xps8ZbN
nf1a6vYbat2CbomkcIiwwFbcTmIAIHv5tnYGpaXs0xceGuXA/7GbNjXaV99Iuaq0Jv6M3D65p5vW
5M5OFXETrY6Ny8s4YFI/ednRpx8SmURHX+ebXks3bzle0wDvzx4YaOwULvBNUneDbfa+D6fuJp6n
b+eaUX6agNzdpsEh7anuo6iWdwbY3epG7yymX4SXTXHwhVuLayGokXp5fAMPQ/d41g51Og+/9Frq
CPW64XekYku73FQq6RIkKPzvYZBTccesIkJZPjc8RDeAK5pWYdhTqt665FrbT9zZpFYppKO2Wyt2
r27q870MbHmQUhBcSmSf8VKqAbISj74AS7WlemZgetI4HDsc5mxgEMLCf1iCibF5eowqW/79KUZy
iBjQtqpLfrvZ4cld+gtqIyhW7ov3hpJDfDbYiCx9iyGY0ngiK+gf7Fw+mDjpqYmeGPJdLP54EwPy
5aTzMD3Zc0Z1Xg3wTByAJcZZqFZSN2nVcbXLY/OP9lijsdZeeaZUpXtv1fxKtiIMbCJVBI+Gitt2
5EFqunhMQH8Gs5nOpsgY+3sX6v1nET7r00AejHKI5dCzciI4iQRFrUJP+H03/T5b/SGBuvaMWUrh
NyAi+nd4u4fmzAh9K8xBWwNYM+m3KJnG+m+//9kK894GfMZHjAyrq2nfB8bbiCPm/J/QtUwDVbUt
Bn6dneaV/g1naWA5h9K81XDWdTwERc3MsaFXxQbFaTR3y7DKyp8+X5P3gquVH0IFxNOj+0kiZy4s
FbkvgE5z5QI/tD6KiYA7mdcfQ7e3Lqmi/WMsbP4xexXQNTvyMQH9UI2hZZyfYX4Fe6xKkCSsz4rD
GLlAxvkfrFoIL4PVI7+h4Xv+SbgWQxGj4GxRzKbuKd3cHrg6JlGncQ4E9VhsUw526avEgFJRK5UH
GzcJY7zLzUjdS1B/A2wWGMtAOr5ySayCvy6cLfkRMyEQ7b1UCnfXio15XgjMpQtiUz47+rBdpki2
GwTUCdjjQnFz3pOxxTl/reNVj6Rm7+ORPbu8zWsxnETTJwlorBg6d2Gha3ho9+OmeKZDNL9MrRHW
W1OoBCUwD7br8kgDdGkhEDJuZF+gmcFNxwu3T+1Fo9v0vwQO1axD5Dwc7kGlBPiT8tS09u30jcIw
s0GFJXydxg+/7mKBIefk2hOTerxfWCu05wPkjecQ2m5nASn33NVqqRhXAbja2Pi5G3wc+BU8v+q6
rzFo29txQbQEWXCe7XM0EHaqItZJMsI6yG5kPS38C2eAG4apBGGJjZ6moUrkfMxtCKFJasu+zsTS
xMuHjokc59zfHBQN5w2Q7tDPMEY2a+MEbiXiZCCcbuDofCeU6rjvftvQPaPwSb4qxjmFrhNeafuN
/qz/qLmpo98uUoee3ynM7/cTAqLHGMci6PoTVDUWvf2E3Gpi1LKiCLjVaDa+z9tsO3wLog0UmO2v
3xpKQ7B+60ug784+UyVAkH/Lr24KWAKULNGAhteH/JgNwCE1iHhH5lWfZQEPy8uXGoriIEYfURds
OMrrJScucqYchOpQ9C/pUptR4dwygooB741PXZVNsrejlagea3erD0uiwr9aLJsgck1rKM6T1du2
nHH10LVyA2Ain0zvSnOm8dQHyU8UYwcYdOHpKLDPD3u8DshymkNdXbnpRapTNuZOvhxo8g3uKjGD
QAa2gANAUPOsMTb25n02TbWgdg5tDVjoS+apEsVs2jyozG6m/VSoZ3DnSzZrRUfyDvcG2B80nUXn
0Q1sl8Ss+oUrnfyCOyx6fnlQuu5BD1a/bbComJUq+KOJmmsM0MM05sgmJ7Y8kQqcAgF2HE7aKuwo
ZVB/mOTEZ1cc0ZjKG+Orl0iXZnuTxtUsgda1oX80HKGUjtDEIkIKS/2ige+Fa2ROtYTWG7CfWJ7X
hr5vA6OpPhu0DrWLq7q6z9CYLGgG8bteKcFFjHeydZxYZLmXA1J2KMQqNoiBZsj/0TBHJI71A2zi
9pflpYVey/9O1rcm3lSl/hZ2vC9ztyyG+BfLjsBxovC4p3Mhsgngt4cYVonfc0ZEMzd6wrOZs0Eo
X2SQt1BHyRZRH5b1BHaRwKYjKMonu7EOLkAxfmoZUhDvfwebe9ulnjGBvx7SDK1hARBnU5a7ZUU2
0AVXZ6aPjLIU/8G8TDgN4vvdpeRBYIK27jIzvx1WngW5n+uwkkg7xChwNNTuUtU1RWBPCokUn77d
/5QH40mBf7ARj9sKjTgeGHjHPYUEmMpZkG0l3XoFxSI2KrGXU30Ic7icz2gsMaqBSCebcToA5Bo/
64MEjyqqLp2pBngT4hGjUTGjiHh3Sg238Haq4T0k3YZ6GNvghANcrZLkeKUgqDnbBZKZsxuaibMl
E1PAGcMArQeTxBifCJ3L+E21acMkvn+obl0YIs3d8BYZmtbYxpRBnCFSOMuf3bkmNA9b/xeUHnBc
S1hI70Us0wQfes3AT8Ew/IYZGu/QWIKU8pJ4vloK4JtNGEfWPLKMUs72nKfkLs+2jQ/ULgDXISQl
DQFZCh9ghL8wfr0dqTpfr2BLMTJ024MwAAXEvIvvy+0HmMittP+yr/fdrse2jeE66+1aWcS4EBKA
X0Eu6ZA0ux6lqaFzDPTKVXBN9bi1SqHU/fdnRQHV/qdeNzxPsDFxE0D1+1E/hyw0UDSzLNSiiTQr
QJs2DW+EnJMKfmla64xZuNGB8+U6bUPkYcfEk0CTCr8/yFSu8hZKoozGtWnjL6rOqCdxamBVGzdI
1JtGXUOYbGW2HIaSRLhNfoReCUDk7hd+pBjYi+b1bHo6yfC0uTc6Ys8JG0/77iINowi6pt+dKDvE
sZa5QOdhFSjA6ThaTy4mZFPMwcy2enEoZEbdq37GxC6jXeV/eCEkUq+CmZVaVp/Jz5MsXad63+2p
A3AxS4wrBaybsZzbIqzLkAsWJ26RnSwppofNyEL4qJtCoibd8mNLnu1yZzPD9QbyUrnIY4olAWKK
pKE8zZEPZR2sVCHeeO5m6HZJKIkU7YSbjQGmHUyky6VpfL7papicFZy+pXX9j0gdWOYLopRcgX45
S1vJiYZpJxUJPQWHef7RR0iblI3nLAWrNDOi3MkOoOZJ4WQYxQm5DX6H+H8qADH+UWyADncZNR6d
qFkKogBs1dP8kaxJ1I+j7eknHFJCsWJSKcYeTJlZShB2uwiw2oJgbUiOIxTiBd4wuMDbhx75ufZo
dpXCxYl8SYD1nZxC5Z7gJDoKbz5Vs5/AzFNz7P7q17awZM3WaMGF+xy4LEhIaUCtNWp5WCRpB6uU
/rJ/JN8SFaZ7/Q1t7gWmEz6ZASPJI+WbY/o5IRsrHjaHKz1NutB/vGvrMm+MCCWstXxFNW/NMv1b
5CMgEC1+5RBzFBS/jw6jamUzDV6+Pa0siPMWBi4c8NGP2Hh+sHq4lJKlgtyTx2nhrmH2foQdjV1/
2GLn0bCx0kJwT4632s/MQO8ZCC49vZ4V8Oe6V5k/AOVLR8XnQRyguotDAhFpnxZGpkUCjomZtNsl
24++BavocS5t+gugjEkSR57lYe7XpyGjtxbKkSEhIJhITcUtOZtbkEZ1Baw3SB3LabR97RZDNO/5
R37yIFYuUuXN1V1HcgtEZJNAYpBZknUrtV2khb2BalmTybv6otTVZww49yMPjt5QJFu6Yig4SmzE
Ec98MaCbwr9u0KaKo3rmC77wXKeL3yA93Hl9380nBPKEhsSikuxF3zCffi28yzdGEDxoeJYADJx5
E6zcP3Rq6oS3DPz7J8THtOyPXSSgs7gCiTi879Xstr8D1ru7wkd416LKMLReTgQVLApP3kohHK+b
7aE5gbIHemceVyam8X2viCf6USDL54DL6/yms9mGWio9RceascVnovtkVvduZFafJyZzU5UHof0K
/M3y4cBO6/LjfCVU+2mxW2X9WsUcVrRZx9LSuTN0hAKJCGTaE4Y+gjz7FvwYEUS2hbOUbZpBDQSR
j/NQxZrMR9HFWE0pA8WUgvHox6+SlbTKP0J0ksQwDPa55a3mwnGm4uCryhcBR+jHnJQ1p5czqzbB
WwphjEeKQfz5MC2X5dqScR5vNfn0qPi8KuoYMJfmmtT5e8O9P+ar1G/us4A0hK2bQPZXBiN2sOfw
nzozxjBAK0BeEPKmB6263X8tpCpbuXY/GtnlZO4iGtL1ccgNGZhW5vynY56jIWkAKMuW0+/eyx/z
Fwwf3P8BtytjC1+jL/VbzHbDY6kxa2OkhlDhgP6EwOF9hFgcjCUh0bwRfpZq4973RGI1koLzxLpQ
47EGemb7YpqlQfirUvAGxTol+YIEOOBeDQ9FImgn4oxXoh2mMAAyZ2S0sY9Dtqay40GFAJ47/Iiu
hx3OimsgxkhtSVV54zr+iCEMSzIiLmqzQIyvsGMeschCZJgpunoI4501EpHw1f8qDT3+EgJgEzZi
XUh0uuqGQYHqON9DHusri2frkqEnWtvxeyrx3TfSwazOjIvXvMQkekG2bcE52sdV8OCOF9M2II4q
rk0/ZmDq/TgTtC6vFumJ2GBg3U2HV1mtbIi59os2rJAOKRkkb85Fgm2X1ecKeEPGH6IFFOAYF3Im
a6+3XX3XIyGoko2CiC+azxe1XsteHPH0cYoUBq1eHO9TruIn3O8SrsXsL/fgfrnzNVXQWA2S8zYd
e1l+eoGGlo8tDGShVVnHkClf4e0HwvpQsvwW6U1WeQ0FkibAGQcmroTEdBDflMLatYCCPW+phHsT
iqy06/M71W5QMF+3N0f06Ws0+JLTxUmBxZvNtY7Pf8JfzTyoZcN2ZilfpjrQ74ixf1cXwXupY/cy
cGIcH1gF39UGpGruTC3+czzHM7DOio9A1MyUa7fXTvSbUc2tFAjaqr1j4hwLZ/dSb9AbByKZ4cAS
c5aTRe1WGaMuV5I+LtdturNWPM00oON4ZyBcYeeHO2dX4Nq4Fi7Qz5gd5TjiRenIXEw/UmkdnQH8
Gcn1WFccscZDo4P1W5IL25IiXCH/OAZtFZJpL+mGLkIvRzhdb9CwyQJYYY+y/VwbvoUiHFQ4vbtl
3/iJoLMMuMlmdcwPdtkeQGvxa0T4fDqxgblvLVjNdF23kPlY9UCeSZOeU5A6mbH2WTkyYudg6G1i
QfynVzwxk54F3Nebwk3DSa89muVQ19SilFkEEI2bL+nEUDU30UgV7vApdiWcVSQwbpvI4LHPbqP2
ocp8dKy5wzjBQx0yiIssXr1/EbFvlDQhnOYR7MZZ2qh5S34WuWVwrjur6FjPIy+O7kU/bv9ZuEOB
7OaU/WO2v6dRlCuEanPfc9FOfJpz0rEI8bpRelz/cc2nyPeJ5T25SF9iw7kzjqYZCJTK8be/Y1eu
JNCeOKe+Lv4/Rh322rcRFqfo78O6csEVeMhVo/KosyWg2vUzOdEpZAc6hJlMhFz/v5/hKSkbMCGX
c7IrsuRH2g1rR+OpNMDoupS6+4cHkAimO3iUVJajbfpTFN0d1H7vJI1fPrZeOsMGB+MvRYK1FnTx
tGRqWkC6x2UVMkVdvbbwfsr0EOGAk+RGdoA0LU69LnpRsm/SWxtGEg+1+eqNeiGil0oE9NB/QilO
n+MHU40y1nJyCR0aVVqC355l0i+NpqPYO1UU+LGayWIWFBVMVKQRNGTS3Bt1dY44EaZsepPfCgvy
GkJAFLaTNKnM4ZTUsjw3zWmjxSgpDpiYPfWVhFJ/EL1yh6JeGeMEazwhGweMa3EX4hZ6hK06MJps
W9fXjc5i/el8UIf0w7evoegpHpvJG1sB8myZonRSv0lZG7U1N7arOTCukBx6B/Kko1+0jf8i/mTG
I6W5laxQMdloiksryth6TlxA+hACX/HE49yRktyMeSKZSYHUcoZnpI/tQnjC7G+z4eO/NfQ+jm+7
AsAdL3v76ENxqH4Gp738VkS4NrAdNNEoiAjfN7oOqtMs0oJ7eFRcgry+p+n8agIAlANDz5vQCZVW
Tf/Yjh1n1idzJc1ZBJgtpt2HIEc1iqWZ9rxB1NAQkoEzXO7MUB/7rkrrilmmU4B7KTUNAJ1vgpxL
u6ELhRNfIk58M40PB++upDxmdO+0aMRuGaSdxBnX73cyz7l7qLJcE3bPaFEQby8+z1F0eoyKeib7
vMYnQtohs+ZWzzGKCMZKrcg2hUa38Tyyvzd051ytTm/gX5nzHillT2W0EYbj+0FLPt7h5ol3i+XR
pdojCy9HU7KYFktrVpWNtRM/5M0u+4Eyr9oOKbCVVpftV/OdIanLYr50TFt8dvoDmwBWec9bmexd
RTmojby0PfJ6/Q3LQReWjfQ3ptBtBVUKh/xG645re4oR3KlW5u9Rec8DSxXxOTy6JE0BbY89rIyk
Di9l8vIxunk5y2PMUQ2xBRzBm845zppD4iz/vmCTbgSIMuHdo7B2jw9CttNCBgu/FALG22gxzWYm
oIa4itJuCLPzGQpj8317nrc9Sq3YY7VIxCCMXPoU8/TvLbWMQ1ttS06P8i8ZbSd5t5JgD/vCFGls
aerUx0B7+iekkbudkUEmM8mqHCiA9bLC1ZJBGrNcRaMJPY4Z89fWchB/ndrcqBmk/+6877aIalyS
NarYOC7Ody+UviL/xNbVjfwFuNZuWtTCPa1OQzG56gcUni/X/0j0oA3cAH6is8aThdD7wfkm7oz5
kEdpHNm9sdBkSfZyxGlLQiH98kt0iXCRjJS5IqsILEEqOQ0GHzfq1yk/lO+CQ+xU/IuvZVcO07Gy
jblBVS8CbvzY79eXByE9d8eYozLRWGGPVlDHaZanfFrHftgbnFr+pdD+Ao+WSnX9Siu5NyCo0Kok
KNK0ZTgwZAdWXygElyLlWIEn6K/o2YPHzEVC9g33y+YWPfvnrpffURKsZ17MWkoKpHgbCAp4lSFT
zNmCfXVyarRzC46nYJ4F2KCp7L2eed7PK2MH9sFxLfheL9p/KMYP8rCBmCG2QXQFZRS5VdKSpdiY
kIa054pM1C2v8iK0q5HJYmkIMtEZssNENPIggrWtlBPDlnFVkWypxrfAO+cdxVXMMf5zUOlF22cG
788CCopfLsQPZVUQcpdihKGk0Ti1RQMuRThI8xsFtEdDVT/DpsN8IZT8X1MY9lrXn1wOtfdAHwg+
zAFcU+1sG24JLSaIbJEOpvPAUVa8EbVkl7Gi4/JauzZfSZ4uPBbTkmfv4tR/gDbn075kBlTv1t9j
JdXJRzWAm8gAtSdQ2MUsfHcZTnPaN/mYzDdnbkYArl4DQPfFbvEI9rouZ5DUuoMejO88kvy6Q3kf
wkdEZg4X0JQCd401c/ynzcX69GKDzLYJu79mEj4amo53nCu5G62eAFGUll+6Akcg13aVnWf34nBE
4WA/rp7c89jtf2FWOS8l1mzaoIOtTqtuoe2he9kdTzXQAAtCsomD8u/dsYfd94hMxf5ye+tGVq/u
9rT+A25g8WljBYflDLZ9PC+Qp44+UKDoX/TLGt9SGWTqD7EszSwWWOx4ktMxJvoogwPhj3q4Dyzt
xPVwc0Yjtf2msBi0WEDzjTQuL3mLzrEO3ifA3DBL+chZ/zpkqP/rYKAUJnc6g0jSCAhFBGatLx2v
1EfssdQ+nnqmlMZoT4qGkwFSMGRflB0ZEm4YEbsPgZ9j3clhb+Tkm1aliDgbSOnF72EYmPIbqY0i
6f+MvzNsZYWolK/Ncui7hFVDDTiu0Nm5jnRI7NoKACGhGhPj/uCz2D0uIiuLHTTP4q/46OZktytG
8CfSn1VU9DqS+gggAR/HuZD9pRd4UR72qQIxMzB7MOjW4A1mmABcwQQaPESc7pgURBbF5iOXMrjJ
xB45cdGoU9m4fg1qlE++7xit4A20E3UUMcEOKvoZ/GAYnQz+izf7qNIaDl0Exg9yBEk8ZHTHqDED
uzWQ6mVqCFxnhmgjCqWzgzR3Nqw430a4v/LXLEd4HtbaurOIrwOnbsVyz3RTldPEQ8MuO0rUgB4v
XtnNVIh7uuKP/0GSYAMOcqxzHXI84V2+I8y8aGQN7yTfQVlzAu2F9EpLlXuIsyowYpXZc6H1NHYA
veXd+uVl33a7mOVNkhjgl3dBfQAhtsMoAJpXTVSF8myA3eN5ZvnD8qkXIMiE5Rbvy/qXZy7BrTYP
EiwfYkXGPz7h71zRVhAAECBDYyw40SUb7Pwo1B69qTUgPWLgoWugUHDqvUJr18gLFJbmDQ3I6Ldf
E+Y/1gfQ4fY33EC3fwvf4Zu0pvjow7+fPOQ7ncCUfQmU3KgnR4O+hRzBZPQlhUtN0fKGHDSs7mUA
MN5SFBPra2rB8iI+k5P9Dg8+21E2JqewY8WEfpO4I8Wg3A0KzVKIXaRQD8saFEeKxTuam95Vutot
AkCYifz0uKaDWXzYQoVcNYFPvIaXgpEgfuUhe5zCfRXP0gDQy+OyU/ZUAv8pcVoH1sccrzxB4ExL
j/L1zGCv97CPTK1ksZ4CJAZlkzPpt4TAV1x3KEhZKHGxQryU/miX/FsLSNlDd+GOjHaYkwtuuBWK
LyPOQE+wn1x2TTkw1dGncMHyOQU5T8EHx3bwz8vyr5o6OP51PChkJ2EWhYe8x1Sbqrl04d+aIh0x
VHW1dpKAne70RVSJ2vfXVX3sGMOmukmrsyAAzF/t+NEdOQe+cMhUVqUUcYsxoiMsxUKBuBF38ZBl
AE5NmLxl9jg9NZKrty53XXcEwCTrjWoETcuSGm3ZUNqGoD+cnR6GWtL1s0zQGVioYLiGnBDYep6X
f4/M27sxU73q7PI7pPQg+lXY6nOFH+01oc+pyjhsmGGf+ZxQ8jFqPWr+pmJ/ZfDFoN995/ZY69aC
hZMtmOqQXmuUIsM4p01ZG+jDhll4dajeFt2hkhfroyYutPIyMjZyUutQfznUWqYBMTr85k9VZon5
X4PTS6qUbKR1znjf2Q8kcpl1t7IAGPZTULfk3PUf1N8uKxzatB5FVLHWUVxkh4l4XbzSpXuUWl0H
zwNHVbD5J0mzIHGH6geK2+qT2z4U3XAdV1n3KiueO8JI3bXW8JL2VoDNkPLyWcjG1UNXwQWe6pui
SbgEswRnPBRDkB59HLvj74wsqGdHT3YDvRVZVKquF9310RMX+/UcfQAWph6efXnr05fFX362QXz6
Bi74V/nwSKswIvYdbZQYh1M1RybEeFpIFaWYy8uEyypjkonuIW3sXC02qP1eqDABP28B3Fjh8XW5
tcmzU/RgYCn8u0x39tRlGH71nzCuZNGUA0wWrpMhU+PhdBC6BHPT633vVZih+NRV/4bH6rkj/fWA
NxoRECV4gT18agXbYpNlqIaOHzM/akTRjENS4SngYotH3CowjCSoQamorsX52nN+DsakD2IyPLZD
YU6GKSn3XwVai3u3kGcqRC7l6AcZfrv9ahXIKjSgTfUNP/8WaL3/TIONpmgq29PoHm7vKxqMENeE
7Nr2Q7b6wz6FmvMA5rQHh+Ddce265GXrm2V+IUaLkf1PF1ynDN18DuazHunE5kgObHCSDRvJgxwH
ezlLWDiIF3Hfroh6SLQhdeit+OEbKFI8p74P7KQD8O1j2sFZ9Rh0u9l/BTao+qJXp1R5ZzOH6rly
UNysgHSAO6h6mFh+pT5EWuAEyVoxS6qqucqlIk4PDgja0BE1bAyHUdrKeWLB3pRwY1sSv8FtbVgn
UcthRigs6k8wsKFkJ2kowBDI03hiamUm5fdnMPrT/5Zt23PCnMJUV6gMPiuMweJ1Qrh2UCQtc2yM
yAJLBvPi97rj5+tyQurYmJ2rJS6LTXkiuUNKmyw+HHB+LReFZgA+2QOArExM5wwQsTxyOuWdBEJd
iM7c9GvFJ5W0mMyYa1tR/ZZwcGMgkV/yxjY1WV96IYZLZoEx+NYlwT7TUbrP+Ymy0B3ch8OGAYy5
NFf/CKEJG+XkV5fTQ0TQOMgbDVv5ZC93DAZzA0SgFFeuOGNPUdTEMGlkSwBOPwTLsL0U2phe3Fvy
QDu3TeQsGJiiwaSMM0kbat61KsGkEAADN3r47csixi42ZV1pkg67rbNxme0ezDangjZ6CtjAGq0N
dLuC6oOAmbAkncqNqmPO5SmumbNE2F2G8wQ9gCwWDSCtFbWCACk7f+Sd0a6H75hNlAVJ+Xt1+pE1
pNPy4iw30OguHvoq/kisQnmIBF/tbjtGJtgCI/OHIDq1NXtjySPNcuG+oI5UZ1qRySBQHYH5RTOu
TacysyUBAVwZQYQ53LQoteTih0YlGAJCyJSvDmMcuP1x8bCN6fZG7YLlIAZNgTHzIAPJHZBNIbFd
RzR9ou8D4QQ8h3BwjfDhq+NXRiI6twZ0XitNzvAlnnIKkLqZpohG8vBzLd/D3q6ABC5ZPAZaPXud
E+N10w2nZHLB7hKcwjUqqvQXtQ7TnwFjZhkq3CdLzkQDm0Gp546JAUfytMOYtyi/wFS9G25Nx9/+
dJ8Df9BwDiHr0TucEqKOjEC6LJSrlhDz16Grk25sT0sPU2YrwYzGPyWY1AaHQbUTK17uaaQJM1Tv
BgyGc7ZGe3WBmLHZNDQjym0gGKZ0FacQA/A04jfRbLC0Ad5HoGVIoBwzEHN11pydSaoLzipv+pC3
LDosoVyUXvrf7ULJq1O4TO3j+/pbDFOMwhBLmjSUysODXLs/uM7cc2KENvJkCSbZhXb4CbC+N7km
9Q3t1jm5VDy4sYhn1iJrmwY8GJypguI9phTffNCDLQKIXroqRQoqT4NCK2cLmXzZDK2TZoFutqIX
ocuwcCRN5skTPUnIwVq7XDA2iyg7gVrWks5QrcoBBFZ+fcCoFboxchxN1GniECVDMGuoc8z8DQDL
WUxYklWpzN8cK5HQNu05OeVpeKXprrmZbrrJ4c0LFY/kVckl91Pc/Z2mPHsQlExjwwXB7HSzttKo
DETnuZNYAmY69ndffyUvYBuJYNBJKL63nu2Il2DA7ZJ6abuBLY2kTRFYVKulFXwkMYfdfg1gC5/U
j5m45xhVS/ePm0hDjXJC/CKVxqJNJcKByiQ/z98ByNvmufXCQ+kzJ6nFRngKAbfbf8T2fjHJYr6t
zj6XFgMt5rrMmc42WcXYskHohnvla6eIzGxfUwd7TK/1SispfgaiH60+synRruHIGOEkCRoir1Ct
LxvzBJpHX4AqR5rNvJjqIAo0fsfZE2pHym/ceK5MlFDgb0AshxfJWXNaJua3nUPPwOSIP43j6dO8
OReNve5Hgm0hSZj+YDI20Q1swpYrjetMxrseBvb11sKNenOJwR+7nl8Xsz71jax1s6ps6ltjvAzl
G2+Hmkr/2aw9qkPsOeoDdto3jFSIb34B99ce6zqhXfwdf7j9w4GEXy+Nfp9MUuAIGmQM49ee0GVo
hKW2Le0pQ2M2/4Z0pvRbqtsJ5UxIXTJzN0RQ9KUnoHMj9XFUa0nJO4OJhm1jBcsG2nu7w/38hqxK
g7DLUIhlB3hFQ745lwVLxI8lgQGngsBKcEn1QYP2JtFZHoentkLG4rN3y03YUs289U2JUjq4+RXQ
KK6P2QugGe+Tp6FUMXS09yKejoqjsO7IWh/NVas46bZYX/z7WQAc7VyVgpSeMy0IRu+jFkXQ8t3s
jKKHFZNaNIEVP+DqlzSTgPN0WMkWDr1O5v5sXSweEl6EmdUAbaxGn42Vyp6qQG6meATWGpMQ1//C
4yGUonSYpCGPdECJ/yeTMtDFyfQmdjBAvEJTFnH1GO4V8Tnsg2721N1sNCuTDjbnQI9Y35G65Cl2
eBeui0dAvZwjr4Xt+REgqHPKicOb54p/od6i48GMQk0PJPqmLeVnIQ1ecN/F9TCjLj2bWyErLyjQ
Gk/vVKkmLsdWeFOkxF5ZUtSTwlpfDywnMe4AiFHDtJiYGKBHzq18D/AvoCxd5U6HrgA2mc/ZSv06
1R0wDkaiGOR5hVgaIdlTkZ/bfU/KemsGnnNiPVyiYSaZGzwoAOcA088LWvSzQtOSml5zmc5jSIbJ
wHnYDu7SMyDLlnJeta2j+Il1ZRcU0Lhp8IieVlPOJeCDOc9WKeYZVYM6M8qrVla6gYtfu4rjWo7W
7ecD2AMeZL8oPUWwu7aAubZRB1Wcu+GPn3NjUcET/I3s0LFz7ZD69FduZD4g6gilyvT332n2xqT+
qWPgignXaUq/1NT3UGAdeqC3yPOg9xzV6anYo0u3iKil7SmcEBPUdi28ExAi3ZryZ1hAOQ8lr8Li
mn4RU+h93MrJrfCV/Jmzbye+6EdsouTVSqg+jehFftL4kmGoYGm8uAwup8e9lMd64UXUCts55yXp
nfUu91RA1sNpSo4K+d1+s09X7Geyzqv+j2iDhoiy8RBEOa3Hk25HdTDs0zhnsvtj6FbXBMmzkPz3
NhaidGdhc5GASWidHElk9GjMzfAd1wBvGSSoes6iCuSUx4aHVXJ8s1pHbNdt+22dBhF6KwmPOIcy
aQ2FA6mYqfR0ZcLif9LMa9NEqUIIDtzifxeuZA5heeeOJRwCjXRZMA5xbkvJUucMbI7BwPTEB/qK
OUhp0gbiC8tmjuKpKJGyHJWYkSKrXb3Fbsigl78rRBuDBfM9TWvb9lrOQPjDFM6EI48l6szCqxCf
ctD5oNSaWE5d49hvR/iBI7hdwCNvqWVqyf34rp62XalPz50DY2UZkT5row0KAorZuDP0Qjkv7faE
2YHZw2hxHzVzDmutnu8aQryYoSt+AZHZilFjhnSQf3QoabCJgxIaFowj+ifpShqMOynfbW3ShQXk
gkfwXgVf9SaJz7XCeyHDl1itS6TTzTD78qTLJEgEqT1NZ5Gcvc47rUovrNQQiCx541fbgP+L2ekB
xk2NWeVbAFVnY+A0FyXTfiG6ahd5bYHTDgyj4daV3t2GVXAnG1nvgwvk46fwyovoWgQfUO+N6lmk
yKW5BAZy9074S+N/EF8qeARY5+nGe9WJJkTP4HFM/BLlrO2gisgCv5U5hqs1hYJHrkSXbNHz8Ztj
EsweTVdGhX/THsHJMbGB4QuOghQa3OnsbilhpMHsORMlnG+tkP95tnHjqKjJZsmkZ1uv0KiosR6A
OhmTfbID2zF/goFgHSMxMUlwpVc2PVXswroSJv4XqOWngdJwKtPzXR6gTepIBhWBdPA30Vg11zjv
NGza/qLe1EAhzAsnnQZzag5I7tnh3nfCfwxVje0sDzTEvOUCvRkYZ6vo/ck/jkONSjMWXy5twXXj
dmdw0z/jtIRISvQM3favSe5BJd0lqZV8ITqAYQ9LFffzeuYST+2Y1je1kUHn1I9U0yuKuFurxSXv
w9xjlg0+5eS1S2ouHX5ZCSTw8Q7fPWW+cnK9Au9lomz/zdEdDjw8rtKox71uly2yRv8mw+FMpYMc
a8+5wxIays6QYCuBp990AOJed4O2kFTSYtaC2VstYHJZBx1Zrotg4PlX4hvt2jcgPRComb41cqS1
qmpUUkDuOHvAcMb942smk/uyyCnd2h+mYGFqo9LWQ1PTNkLumHAf5TSqpwXHl3ZGKajDF/4FUF18
QiT4rpUQfNuoBgLVTKGhBI/IALYKR1bMNMkryCcFdImkr+twc9r6OtVnX/1xKjFeEKvh5nK1fiK/
7Wji35LBxKvxe4i9qpjztjibQRrAaqxESAVBV1PwPCxyAAFaSUHs7D2puDrRwF49XDWBr/wG3UP1
jjLKmq9w2p+tPvzeDmc/++Hqrh7JUynw3iwALm+enZfWdZrxPdBBbY7ySBLJ6oCn0evdFos7h+Y0
lh54nt33QAxK61q0HXSU4praA0lKXG2/pYk3pxr2GC0zIN/KgC/FlD+G+Q+9NzBOe9A6CTnlOGHG
ONvjG++moKUHzR5EcV4LGi7kWkTHVJw3PoGh7Ssls9/F1BudCxk82maMy9cZ4DKLNNWiSP+R+fjs
DHaIXiVJ/grVgdrzlVfZxIfaG2s87ajkAUt7GZornxrnmXMGuiPdBcEhlFCbvxGC3011xu4Hjp6T
uPHYcrjJnJLsDbzJZxTrAVvhIXiI+O0E6napkbM2su4Q2FqN3rJtDPpPBMqSVtJ6XTPPQVB4zoVy
QVTpNZNrorf6C8ww0mOAiWQC9+Ah8OOAbSUyeYy7aeB8JWXjgqeQngTZJcq0VEK9GvgvkkVS2Hdv
lBdfUo8ftYd3DgNkpZK/XshpdOwZVwfNmf8k5RNHEJlRF5QfB7NtT/4Xp1HEuUM15m1d1zjQCx13
pQYyX5c4BG1/jYG7qwl9RT3WuwOvtypB433lAfsxjcTKeFzMEKTNP38cFdsD9FGZfd12wMng9ds2
A8MYBhU2OmGr6IvkkmRZOpZOidfvR40TsqzR4RmIpKAiQm89gHVHXVyhSCCwDQ/5kPee6e1IkRqj
yJwSnbPwxxnUB0m8VlIElKAZm2y9o38uZfHAEm5DpAi/KgC9teGNWJxBDOeulshtFItgXnvvdqca
4IoA2docgm30GWAg9rqBiKlEsHlpWN/TiM+U81FrvUZCViC3paA+hy5nXSuSWcC5eE/HMd7GyrTe
fxR4IEp2hVTqQlgieYT4ZaBixtBZf0h7UGvr9Vq55qCQMHaWu1tsvWCreymvYSARqcxiUYWIVYEa
FCN1CNr+Q4DJ0r/uPRC6QxT+Krewq1Dal6/83aFna/u4lvFpq3Irpxi1VhoLB4cFAr9swQjghM8b
JMvA2MTJI2L+5XDKN2uvtKk3+0/Vo6gbiUxcY+kfy49VCea40XRKDfD8aBlB7oYFR+khm8O2e9Ix
Upf9Chfmr2vBh2z5qnRbKUMWL9z2U1pTnULWXhesG+TX6AKOm2I4+i/uC9VOSmqvaCPN8EPlTswZ
/QFwSfDRFuBijH94a8a/M8UqxpgEQLnw+YDdfpmX9/KQZ52BTVRp5Ihsq3jAoTImCo/Gl5chLIrt
cr8DI+eqT+sWxqsK5y6QxZ3W2XHG+3LBi5eTqG4dDrY5iGdRz+1il/mlfxr1f+J36UYuBodyIfSe
QiQttbQSp448G/K2vNYNSh5T6nIXOMZXjkus4wlioungU2BkVPdDZXamqMbnsTnkztE4JQlXywM+
shiO+7FgoGSSU4zdXZKRPDl1uUUei+qpKXmfkI0zxS9T9aXbTzql9eGfoqmxtEnxNOBBSv6n6+C7
cbrjRI7UEamJTyyz8o+5/2F24UvjAKq/y5H3XLt5saJkHFBh1qjPfi8C+7qUdcDTf4vhsDxvJGN8
o/Kq2fJ1gZAygeqYDDmSNpYEB2Qds6bjYpcLe/f62wqg3CgyaK/fyahq7rQ7WvqbT5I9I1Cuu5FV
wPp5lI7BqJhQa2Pf5/32xukTv+Ni2eXKfpysgjP5E5XN0nxNiK/e218Y3A9o9ILA0S7D6cv7OSTg
Su5dzbYjBcNBGga6BgD3Bl3a5H1OBIkZfVX9hFz7X723PkPV2jDqUf6rY0aHJdjh80FfJbM2dE82
XXdD2HzweRxStDb8iwKbLQ76/8atMIFJqJXlF6Pvdg8ncZwiKxEOM13zcsfyPapYnRTBtXHpP5dZ
f52OFw7ZEopT2oSaX5mIisU8jpsuBr2CG3cfr1xSJh0vCIUPOy+njlM5kEqfLBsT8KNBhNlDyi3M
ZJuOp3EGCexsOKCFDRD/euk/IqX9IEQCy6NHAwn56jqzpoGDRpZ8+l+nZ6yfYw7rx/t7tnhSpEzg
9wuRQ5PTLnalukQzR6CjnGZR3tFDzPn54F5bCDls/fYkt2rprxSWzErJIiDzFIIASQxsv7vJcruZ
bFFwuJJwKjJzq0JHS8glHVv2SpmlNw0+ol5x8i/IdjIDr/LzRLYHTJNfCUMNBqUEmrCCGlp/psPn
7JzIGNSZNi73bk98VhsZK+vrsveCAxlN3xvv9+A4KMng8AWXGVAZkl+Vd25OxwghCmImR/kKnCcg
DQSITGfjYmQXTnfB5AEHIZdYuNtF00uroMvnJ5gmzNSQaYejKWS+9Nq1vpBzqd68zQY42TwVS4b4
AjI47B+MJlAo7qG3+JK1SBsaedQgukv22mMP8ATn7bPe1zznPQc38IQHXhGAkr5MrQ42N8mGBHh0
ipWsJtnHAWblOs6rUcUUWKCgI1ZtjfaZo5kjmWpRjH61uj+GmZZ1rePiNyr7WLA87vhOLxwFcQ1p
H0VAX/I67E2m8DVd+Ab+pe8Q1hliTgD7e9+DN6jeRqGSbIEE8UZbPCdTsOENLMCcjUeb5HSkrZnT
lrRqohF+j4VxqUFSvzeRKdYNuhcEeixdxzgUPhgkcCqR+7K4dxAWAaLp8NR+t3FHCaXPam5NPj9W
RO1JhERoOAxDeeAjKwMyltOUFMGmv/E9W10eERohDweNJvonohqnzRU7YXuFfrs4PCgcs1w7JriM
GK3nUSXrhpELlwi+n91Wg0LijLqi+NCL0X+zFquk8PCKK9W+s/MdTfOAYF4bOmGYvGhSiXpBMpsD
xXkBeRJkFvW71FiW3nAhOM033ST4cchALAjV2SVKlPCqyVjaxu6bfgUR0ek0RII+Pa13MP/oeZ2l
s8xHfYUEN3HnFAe5uUyPM5Sk3i0QygdGNm9E4oBcWzKtvgQ5Rv+NzFaIqwOLpGgGy4k9WeynbDPr
qdatqETX2izcZ4jqhqkpIlxTTK7Lnk+wpw8zL1COYZrqZ4uce248qfSCGil/VN4nOboHoWBxK5D8
zCIJ9OKBIuTLoG80FNl6072mLQWLKyznNi8mKroxykDW6QTVfnwHXrNeeSCntF04DP1f61LbF6Jt
m/ZdVGDzC6Ap1XcYqMPq3vu9mUFaDTOjp/RYfcFb7iDVFD9+cULJCht6fmVcL97mlEHyoiZ0QUD8
NNncwUMW8mWLwvpTE3nG/PygiDmNRqU8Fa5vwxxkv1J/6gt6j9xJxHzX3vBQ7Y0mumlgaWDuXh1/
IJOAZsyVtaOpoOu6PJUnZLbGVY/WNOzcpz8Y7dzi11gKrKzu6T/G4NxtinM0i/vSYcRRAr3qqV9k
wJgLaMwEs6vjSjKsUhM4+J0Oz9Tx2EcYdoiI1fM0TKIXHF/v+8ZcPn/5XSQT/+M83haQHVEqzFs2
wIHm3v6whFaPOjIFVMiA2HuL7IstyGPo6VlihtOCr+P1GLQQ8YVEreVQ8gNl+MBbMTU2lCdJ+WgG
7AYEn6pmoFQQinrKedBMrjV6ABLFTXFXmWzwjnIEPCyLsWHMhCQyitsUDbDlNn5HrOKN8HjNvGm1
AHxPICjLXnnIzn0jRIXUrOO777Ot8ChGHJHoU5ULBTgBALlXh7CCUpVguxXN8gJfXK5Ega/mG1GS
pClvlSQDcNBfWY5MXnJuu8LSR6Fd0UzH67scLIkUyeRg49OUY3rzvmKra3wsd8a+/7wqo1jdu3wP
HKfUfYpuR17HQxE465uCSy/uyCOpCrELFURjSXDGJx1JojO5j/3BpbicDUEc1NEG+tcW/KDwjnat
PnvvCN6TkMpX/wPOu0LoXuM2dTUTDCCG/RFWW1iMk0aDk+DisvFpckoGbKHhQnILaoAtB16iKJdw
EJTWf3Eg/a0hrSY38BbwHDHaIeh/He6jYacGFXtU8eLrzhmPzJBuLuEWGY64ijPNS9Ag4fwbzcuR
hjta50YBfq79js5DpCqQRsI7UxGD8BijeY0Z/Dk4z84Kw/iGcfO7J5hkt/Y2ImACeUGsYIRjQvN4
4uynmQkZVrLWuF/ibiKB6s+wBjHWzGc6mfjCuuWv2zwkRqoQgOABxTVCdebtH0uRxoM+WURndPLG
pDouHMgzp/VMzHHCWqBvRuLoPFAyoaR4Y7hEPTS+hlzZ81502NQDjqcX4bedLFKr4nLg6pCqS/2U
543qSgyuUWnKOZb1xX8w0Vrt9N5numEG0s1mzEXjf8piHxTobu36OlTtz9k7EiQscWzEglSNMOyP
rwKMp3D2Q5soVFVVrKg0usrbnhR83kb3+Im0a71d7vfuaUlPsDOZ5t2h+2ZkZT4cKcxfSGmbRI7U
UH9DSLpVz7AhElD10naGXJoUB0zZhPBrgKaJokRrTR6xn4gZ4/mMkG7nNy25mT2seMP6SspD4zaJ
0wD7mdAz1XW3uxJBpZFQs/YlvnFOgOw0FhT/o0d8tQAuTxZNdkvL5Wi2c0D5WLbI6a4Ls2+qGpBI
RVHFPp7Vlom3m/Vl7jTiSpp3fRhnrflHzdG092qsNa4HyskQMyuC3zUYIAOfl+WjmNe+796hlz51
FmGuD1fuGVevK8U4bld7Ez4aCxixSzlIR0lwiW6OskEaWQGZr7cEOY8F7t0y/UdDe4n9aAF+hCCl
e+UEZ5m+hOra+7Brx+e2sFyYJR27+Q5BZw7FVkTCFTkxcjn85P5uj05BF3QR4D2e0Fy228FtDV3F
wKtRMCg/9ijisN708xBd2u3I3X9MbXkD1indp9Ynwp+ciGZYc/WyDaiRR/xD68KNoPJYeohRiRaZ
Vly7XXJWpuzklWIWS2Gzh4tIZoY1zhs0146/XojQsfrlEfF1DF2PcsdBT2xE3X5hPOqA1cnRzzvu
jyrACL22t9GUpC3Wrr0YjM60NYkscyPTmoIibvRs80ObOZ0blOtpi+HDvBxuSlmtdLWEkpAR+Tjg
2Ft73s9/i+ONHlg2TB8FVZfpxewd+4qNh+Jti3hjQphwJBT8aEKbWGMN+0RE5HPTrmNxydoODQqs
MUtr0ovZTgN9ver5cFBedNlTvh5paEjIwVhjpKep9MQiY8EKJuZKVVxGA0QTG1Ba0C1+KFV+7xXQ
rCoq2kTjFkSCfgOS9U6086W5kG0dtXydGaL6t+DEmq2dkMfhkWkO21Lthz11iKFxqhw37oB2PO+I
P/qcuhOpnhvN+0edIP92DFHGkr/XwqVhn9rzVUC4CNWeFnE4p/rO6T3jlRg9i8/dqpSbFFmUF6/n
0eDv+doPdeNXNy1pwNqm06QY0fAbvQDjP7C1oNZ73GX2woR6QYdsL3RP8qn7oeItVu7N7EWvGgo0
tPYf46XNvHG9Q7tq+Uq6qVbcAgEygxdcaelDA2JoaWovUc0odz0EiY0TS3YT63XHt8bPyNA4HC0m
AbF9fo9paxawHCmq5crfdGAEl/DsCDmFGYeIQqVsNpVOPxuI2J9TImUd7rEd6R503k5YpJPgwStY
Ig0t4p4otX3XtrTWj1X1GaIY+IqfeKen9caJBlpjk0rouL9aLX+fAEa3/pjMG6Kt3W8uFaTpWshJ
LYJ+K1dddxU47byOJUZUtFhLqHTdr7YlyVkEAbNxh8uaOKbATaPkqQQZzLZou0t+cxGRtIt4lRRh
nmZBrEDJDfZ7HDPal+jZDmIHTenmXlTYzhj7Qkt2leTZMiimF9E6+bX1VeOgShYiDKtQVOXYsCb6
Nzbxrl3g12j/8G3qflsAO4cA0bG1/vS0QpXF9UJjMlOulRjNxKOQjsUVMNugnhQ8I9IuIqprbbTO
FrvNoVWdIvIeLcj5UZqXoPaR+aJTtr85DoWGbUtVHS59wTU65bCMEm3NEoRXpfA9u/mAZuHJvYVv
0UOWmar9FhYG/p+Kq3NwabmCWSB0It4jJfKmXZ9suWQIXZiLf0WMLCzJZansalIo2B7+rzjHxkbn
TBDmcA2QrTfLQ6r2NYQAd5HfYK9i7tRuPcNK+VCSmFk05vYdItXz2eMK42bQRnCYicIXMSN8UaqB
02o5qc8hO4G6uE3b9RJtcIPzYx04iIZt8qnrztWZnd7R9k1tdcq4rHhuE5qMFixjiy01Jk+U+75q
N+Zqd5gLpwVKyZHuVqdN2TzYqRTzGw7kDn/5t0kf77oOwBsCWazHrmnT/h+w6aKf4w83hWM4iM/5
coCMV0IzjhrR8GA7sYNlTGgy5IiX/6ZfkF0WgGghZeN+OZWdQ3r5KW1YVA6KyHCHVnhheEwBXb50
NT78VkJCtcVgauNmlBFi5EU0fk2zfQ99VOGwUlRGyXX6yVcIATcQqXmbnz8c5FRB+8Ppolp3rH32
tChSZSY+LKWnWJdiQlr1xX0337onQl83FuQfsS7X53FpYEQVH0bN1tw9ydkZghAbMdy6F9GreNYf
rr0IHmgtHkypZ32H46hBS9bb3ZMFnqfF+c3dA7wtRkyK8a+dB13R2H6eHU4HaMIw38OSMnjH7LMp
tmr+7EGErjTgm1JdHxJ6PLfw8b2ElsCtpdZF35zPZr6FPgMqZLvrVh6BVsLRy8frH8BKBfx2rlsC
+H4vCXzPwzBG3CcU/u8XJpybfMZ/V6iqWt7WzJ0+pF+Zn3dwZb0Fx8Blevvq8MU/zueVDH4UkbWy
9WdvT1y+1nt9PLCExk1dM+y0x64R9KJr25mfW/aeWLgV98WTN214QhZIeOsqOlPuWghZxROl5Z5G
udfFwpjDhSkaHP/9jNndfxJ/BKOhBicR43xpziJxNquaPyLV8A9RIsZ89FLMnQ+DZQ3HUILEf02z
gLOF25ErRhFUyrwt/1IiloWdtYB+gkMJ/+Mkk40zSvWYVfeh9370XrUjjUqFnuFrh9rmetw0XTwX
bWqT8whpDFjRMfWEq+xIVZC8dhs4LrTULqPwc+j0BptxgkUQeu5zKugDE87J3me0uBDg7tfkicXr
nVfZWTLGiheBygWEcJtfeVv84nTgOn5dlNk/2TTLe+h3o6WaItM4CyssA3g6R2AZQo5ahb+nh9Yt
NYLUeAUh9TbzGp2mzuYiMJ9XvLohpwMNzk6oZThMamFvrfqgMNqVJzKKu5p1r/JcEpauFk1TZubJ
10k71iU3vviVL7ybfoutZu3zFSpEci1+z4BjiRPa5DFauBZXRa6CXtyYAi9UafbJ9ibusee8ToWz
6GxgL5asoe5NIEecw3/ZxHhXtG1E2KFdf44uSxT0RFg6xy3J0NlwakQM/B7Ih3T37+h79aNtRSBp
YXx4HldaDqUJ9BsGeUfyMF5UDMlr2pBoF9DzXcfBtVKgC+rC1aw2aOb+X4Ej+Sl2Ns1fy9JpXWeh
47LKwWqAh1lGqgzMoRvEgEdHRkmS/N8WQ0JCO8ZS5fb8ExrfTBbk5oCwon+Zw0aAy94DOHp25Tee
qoahycxWb1UjfMjNsGJwFq9dp2EhY0tLFi0OeD4kulH2dQB+/VXxB6M9mhQ6DLmYFqN/AG3gc5Gy
Y2agSnjpMQwRdbdigK9KRarjngGlO5xl+7C5H0DG4fzev4sLWp7Pa/XE/oUF57y/hOThZH0SNblN
cVMOdboH0BtzkLjq0hEGCbFvhMpoPZuUVfBlm4Z2fDl8J8uZ9QHEBo+zpRE5lhxLA8hL6iHZDpQu
bb71tnXK5nAGg2LDtZr9oYMQTxG+Uiws57QUyrFPUtDabHng6kArP6a2rfOjxzvfj8ih+/Yachyy
YymKjqMIr9UYWBP30nhRj9u3FUit5LnHiAQc4P7a8s5ScFkqghGi0upF5RRJ/jwIpTlXlrVCHWh2
Wtir2oIZqh6BXT1kaaLiNsQ2Vw2UfHJTYT1ZzHMUTBKGNKnRgrR0CuFkJzwh4Y1vsxz09ybl/xjv
ee73LlnATB1CLTl22SmxXKafI5UVPM2nDBRRWyR43xz8azBfPlYAALkvi1VHYSkyWJwNY+J9KNps
pZ42qQlkjr5oUbFSK2zx+7lJck0GXexRldj4xjCXq2bC4hl2v2B7e7MAY7khuMmfihjvvtRLdaUk
yebhlWeuekE/1cTRPcqsoryrjdmwzfalNDk6XFjnP4JVvX8Tt1TkdCeufcbqLSss0CDZbV4P62Ez
jCoR4tfrGSlAIHFb+/M3dVFv1yLLgLoPIbeFpobhnVRXdtPCkwWrgEeD3nxe7j/zvDKI+qNpfkvo
W6zwuG3xjHUjR7fDD46FgXHmgbTOb9b1SLXk+awwA9wiUVXbSgdwUgnADopT5esgQTkb7yVOqwuM
6ekMaS9ph6LM8NwzOpEwNPY2HmK3ZUSBn6l5XD8pkX/pf1oY5gJFtxcMNiMG7/T9iqFzgfgnikyR
JNi1PGGVSRC40fbIZz/c7V0fub+r6xFGAEp+Y9Uam9OTwCC9MXBT55JXmIlIjcx5T7gMIKj+u7Sl
vBbZasH2pwAd36mhJtCz3styVwTMpoKRDmSx0DAX+dfbjKuPUQt4/UAduncvQVI6xaVpGUddeAko
H1nOZLaqgPgHERZRWAH3gHTlGyl/X2BItcqNvZGubbjlgSznnic4ziCrDIKAoBgZ2+gS/zyJpsfx
CPHBiATkUdaFRUsSSxGV7w3VEkNxfucmbJTrsLQZ+beZqDOHicVRjd8DiDUk9wsKiV/iGCNoLtqP
diDVDmnUsWxOPGErvq5X5OKsW/Zd9VczsOmDALsmiXEdKP9iiYxv4nig/ZJE81jV8KNyAv1/9Eek
lDmH3VTxUaJHJeJySzdbxLUvRjA+SuBZLlhWMx3xNju4Udw44BSixwilPqTEB9lkzkoR2/VSx27K
Zh++aown1P4lQSuWB3F5ONPI4YmEeFWFZT+9z7elua7C+HkeLWBnoNFd81cGtZI/bhnLPdlOdChh
gtu+sYbyBAz9ImrrI1wpaBhmMMuRijpZfoLjazKnvRl0rp88iY9gZbQnAJSKBEtjlh8Givd1XVjQ
G9SMYWiXd2A1bgHj+o7X5n8w4gGmUD3MjytqElz4btYYH+n0Y0S1Ol/6oe3PAcXOtmmwQj7mTEo4
ZbvkCHXNcRISOG0FjvHO99K/ZM6S77OclmFNlGu2tWcuBNIxCN1DVHNnQi9ROHhEA4xUunF82vyp
e/fSrzXQVrV5QEU3m2gFqSXeaqADj4xI3BmDTGVZjh/PnhGD1SKL84njo/VCkVAGq7L9bSm8xJ1a
Dnw24X6mvbcGopti1GBfXnHEr6FbM1KgSXLjr8MCx8ab8CJPwrQWJ2y4JElBf7Mzg0Vjx7LWoAxn
KnveAJAzoKb/vLjnVZbS4qAskBSxBc7siq3bvUyX/yvjZFia9dVz1LtwYj6jQU/u9c+a5yCz/X0N
+kQi3o9HsrA1udDg/v/sv3eJKN5W/gf9ca8aynrhvMWqIibX8pfj3LBxbEWfezqPOQWvMf1oO0ff
eTF4Ps2xzwXqQ2CC3Sfhoa1vKrmKipvjBzwxy0b2FJoXmd9NhX4ngx4AU7umV+OBToPydX4F688u
xNR86GSCECrEKSerqaHazGJhRWLWVqLD22t17IuCgxMUiIpcJuQ1XZUQWMzqyYwy0VoIQlYndpwy
HO02OXF4/KpHL9E7QG2EgtNJkYIbaFRJ0UHRBOw3MzdPvpJxA4Z0TsetcsPhJWHb7N+qnKvqArHt
nOrnc0UryE7Yzg16IPdE6T3D7k7zKhutQyup+uXwhAMNHnxEAOlr6/yhgBlV/+L7biQcb9hITiKY
9F5f6SkPqi4ZFxeZ2RInIJyovJUgWikgigeBWY6/jC3aGGyoAiziNvaoAP3StUm/1BE0r88NRDyb
zF5+AdATIc1nXkGgAcLVdCHd1Yh57SOBaX4eXrXbgsQBgMjUV8TTu3agQHZ5Gj9BnybfCnjS1ZBn
in9Ak15Gu3lepDxq+RZTkNeGIbON8u0pFF3Y2sNwKU/8kU1q4CvhSvfh38UiftX42wVRcdVhQSED
oUEYmC2ZJAEUXTleIdSqj/Eiukx4A09fMO41sniROOwQcI/Gb0L37bmHHxBvUozaEpHkQB35BUM8
xz3FDppl/nZ5CNzQkVxy18lt7VzZvz5OKzMflCIiKdUf3hIElW4hkk5Gx6Aghu+ntVPStGZuLKyM
R6ACaGYUtkq6tIrj3alUykBe8FahTvEp3aBHYTrfP0sJcMYuWPnf1gJGv7VuPx0RojW7g722B9gW
EfYwhuQxzGo3j0gJC1B+JimVKv86skNUhCZnxd/V2RlfUacCJh78V5rUPY/nlTTM8+RbizEwdyB9
4+ge/DDT4yQiO+cbr+d27PwVb6RzDOChRodF9dPcT1QdYdclA0qML0scDlFaKYKPLGL8FWqbdXF0
RhfqXLxMWfV8gVJi/WCfXw+2z1gPmRP+4hh3Eu9xbma96P8pDnDVVdJsOcuex5YSb1UebYx2X2U4
hFRFDNZVPmI4T6Dox1LvRaSf48foVp85Am5GN/bv1jlLi4nxy/lzR13/bxhjWiq4vrOgGFAFSuNG
freXyP4TPQtDsfBp4507ToCgfpLeaSVXPXha145GCDbrSAWD9nnwmqzyKz0FfrxMUi05vNs8hJtX
Cz0FpX0FRpqdH7lsspJUiaTVELTIA3sQTe4JyoEcvHKtvA5Gz5OmvEnZnI7uqEZsyXj81OXkylyh
MIRcPor30BpZeyWlKemih/kRp+RKs2OxQgkG9ULq4tnAk8hhRkKynJ4iVhSS4bJqRgvOcd1Iugfq
/JM+ygBN6R4C7mpljtOPslNbtq2TpVfnTrmtY9l3/ovhFe2kabUDQtKu6PNdy2LJ5GoNxik7ewiE
fsE2gBJ40F35haBg5WJtr91w9l1YamiQb2MFj8vQuuDD8QZqcrF56mk7GTZiPj7z+UTEpVL4pGG2
kMNEsL2lkDohdYEfBDVPAzqkbRFEYpGFS1ToINmrkPXIJXcRpDZJc2ElWCAG7WwPad2KIPy57sCV
UAYVrnmpeUW/sAcfwETGpy2nHkeAN3amX5nBQXLcS7bBznKv4aGgJmyQtQqjmTorOa7tMPXyKh5H
WL2YGOmYLaqQ90NnbS4K+9nCXTlR949NRuKfozdqMYkO33JVTG0sB6FzOpAL/ExFr+JjaUzaJTwt
O3gv6a8QhHCtvlIjjX9TIbPltIanhr0/BOa2EXVQv9/4oVS6Avjozgtf+JNCsM/5+xwwCMkbnQTj
ORG5TG1hx8VDxNGOlf6OzuS+RIF3CYERbMnaUJPRkcgGj2GPRBkF21oJ8jXom6uXlrGtLsNptK1s
17AdhAPqIc4vQzv0l7bH5ZaHPP7BfGyVvQlH2bdvunvwswvegK0i8AopXwuPagJTPsj3W7KfPDIv
Fau7UBY75LAhHoaIRJrC2OycOBogGCh8KFIc4lcmuXOU7lqI/P7HsWrioDfbPCGBU3VL35y4EiSy
iyTGQIEhWFfgVee3tiPuRcocUTygDaOL42vnlbxenqHaGRSpMV+lbuufrqUHHdmw3qfnJ82zOVWd
TgzqIIdn66BDjWm1916GXYLyeG4F7OvikWY8R5HTv40VQ3PzpNKhhrB73ovb7B80RWz2/AhRtZRs
bjoYdwE6z1WPT0mBaQgiC0iQ2cRwFLz4bw56deOOAUeriyT3HoPuho+nH7U6B5BqaHjiPwRnRdN+
Xfk128fGlygXAdquakeWC4knMtsZmvk4G8IL+8k8opv6dD7C8BEy4ACzSzq6JtDV7SO/j7PuUop9
ij06cONw4K3y2s4/urUGQkTQfavoskEWqfQ8oz5LGzJL97a8UL3qIqIiDSYnZ7LXJfEQDLUclis9
/FHqmTMJ3bLrIr9HmA0wkixkdv0DQcLRy3UqDoOMzUfpB3IU22n0kzSo3a52h/aCInRgl2vjtbcw
GPHL/4J5waairX2hBYplUDoYPFG0cOBMsN0bKFPxd3vm4asAfGQS7m3ox4u1DZbsxxhlTxQxKGdg
nZBP9DjVo2OUY3Chef+P1IqUq4HA9yzrrhGJLPmmEXKiXsje1Lk14BmL29C4nFEhs8t33F/C4CxL
FJHq6VsiJxO0bPRxlN4sPSW8qUxLunpI1R9uFQcXjRegLG+IcXqxE98fIKtn/05H8NQLmMim0Vza
KBFrDJLSBM1vCJjOPgOnfT4Qq9DTrqb7UxTCeCQsYEPeXkpQmFuBnCBYDvxMcP6DQTbjQJIea3KF
ou4I1+TBvE7yuFq2KaOJf5uXELBf3MO3fqTxnrHLMsCT+F9gsiYEDqH9HXsaZ0tComnXbMskVMRA
yHCCLyJH76OjwmRqbzQCUp/IiL90haj/61lL2pCQU7lPzW99r0sMr7O0yTe/w2DSMns2duja4HvM
WXVqbU5ItxOescqkaaC3FLFxNycrZpsdmv2pCh/ATM6YFMAtXSTkJqsNRJGXpB4yHmGy0oSJO5lL
Mbf99eGNONipHhsLy2LRf4E+UShj3MincDRcpHJATvvWVF5J2TjiyfSf5s0EIWfMguqNOjENLOfF
BAPrih9SQhAm+KRosFDAq5wTLZO+MGgxc9PDYL9HsRlKFHE5Z+/FnUgIMVrsP1EAN1AUn67OXjJ2
G6mmelrr5np/dZ5sLGRkWV0UbXWqAPfcd9e5lida+qQ2iF5Gy+X7KjDdiaFIx7NZ6ZCUh3i8N4B7
Oo9fcx5517HeX25V8ltTvTonUZeMQI5569Q+ETGuOzj2tvFas0bH4BWXCRc9byoVetPW6FX4oquS
R9el8G09KP+eiwnaaKcLVCrUzaHfKPE23+87d1a1W6KRDohOVUUDjawUK0J7qNHIdAyPBoSzVeGk
AtjSpNnrTVrwuwkzhw614J5HYmzb/hluQLuQrldpSCNKqyj8dl332wp7uqs+kv0SL68Nm5pJ1Tj/
xBvVCHIvcJR6UFviMRh/IRl7JGytb/epHduJR8gh/ZtCOylQoniwgzJK4CXttTdQr4JDda8OKieU
YP6UVZojGJQfmzySfVTRpV1cL60SkWCGGfdz7H/SnSApv3a2UZ5ATyej1q/NrgPtkrYSIBNm02Wo
wB8Y0NSA9tEd+G9XdPC3VGXDjs7f2xYDf8h70TvfW5IhEsygwqs0bOdoQM5tcEuYBq4yWbP/Usmb
+jPnEkCMpShDTDD0+yTD7s71A9bzXV+gVgqXou1EknUPQGyYR4IyZcX68Cd7R1eRBPoyRlF+UqOP
GrpgN3ljqwN2xsJ7xYAP+3XhoCtjmu28nG8UhLbKkdcMETem8WNx7E19RTRWXqxRg8OkBvOxmV17
DgOVExKxwRSGlcy3Io0rm7IZUZ/6VNviUlA1DhmN7Y2VX+bnjOFQVMr/7Dh7zYgHwiLS/3YzBiMn
8txDU1byRaPNK59wqal0yRJUWZaHUgBcnC5ZgPGj6H4lv1FspDgwQmfSPGQXe7W+O0qoSu6GESQo
YrkZ3pIqzX0OLIW2V1/oRI0aI8O5AC+RYTjiHLBjiK/jD6DDLnnISYZ26u1FghTXjuIJuQnDJRKY
ydl+yqojBboWwgbo2W0bQ7Z3KkFmfF0A8psmqCFi3U1VUBRhNo4qu1DkAV6Q4gAPIkBn3FUPhnDr
15aAYR9YW2yFtH4swMfokUfBEXoKh73l11XseaLxKvLgZC7Epqgw2WmuM98H6dDahm2IwBhZicnY
+HHFSHrb17dcBENbBK92MSD7kl6Ddv9moBpZdsLBgW02/q1iZgATvViWjZDZJDWpcIyRWQgvIkqe
K9SIgs1PDtw4i2gSxO7N5ZaBrZLE8k49vIX2C5e5mpKC2t1Ct2A6FqUtLRpMx7TueQzKh9Ajfqki
bixb5t9eHW62ELxDtFaGMkCHaVBXLe+z+Zle+XrgvJM/Z2JEs3HFrGtu+hY+f3z9528bexzLinsx
tdUMSkVydrEEn3hMkKNSN655QePDgyMpgAIr6cVqeOLYlsAwI8EMmHrFjMjrr/sG+9s3ViWMgCrS
gVKKWNeuqncJKmYXBAWde8vzaJzjWMZBlzX9l6K2HvRFB2Ln2ndFIohUk7g6vHlWlKyI1aXZL+cd
L8zFfE8uGoCCkTrKoN/P/j/9qr2PnP9iGltkZq+ORtDe7x4T94F08KIQHEwzCrYuVevQv61mhklx
WjTgaQSRcLyYCmND+EtyVkc7FbbshD/mfuvnfRihXxEn7WpEgFgC/LdHLhV0r3U59yanCM4yFV5l
6whmvlJTglbr/uC0rxTE7joAzdZbO+UzTz/WLdxM2h4fOTcv5WtY/j2CtLflSvD5Tt8oYzjsYDmq
87gaM4FELmpBISLWfSc/jTPwfbLhYHL/nuzVlwj2iTcPZBc1HMHr6I2E1t1DAuLWYCN6vKeWuTi1
mBJaiHSIrQ7FBlDtWwc5+5d+pFG1jmE/jkXQfVa/yNtUIAV1D6hfAb8iIFX8ynBKObP1p0ceEzv8
tIXyI5pKBdYPs3mp0eaTqIrAVPVXSTME6u1fRNc23KbsqHZyQGgzdkPMG4VT+P+xB19jkWulr8fq
SWKJyB0cTSRQmGXkVyZDHzplAvuTelwM+RSd8cziUycDsTZ9YvouQu75U2eS/Mi2xSllXQ5auWrB
sv3AX4t+HNHcQ2i/Kqbtu1Bqtr8vNHNFTIc0F2aLfUlaKQ3sgqacllHIbgTsGAS32e1gJI5DTNuj
2eiy3lXEuVejSEEKGB+noaUEvQIBeZbP4HHcUn3vtLHmum9SQUgXpviTQwLVztIgpil21lJpr9kt
eHDSXEuKruCzQhAhOIhjDojsuExhE5wUrqxIHBBht2fAKU1QZPffTgWWSzqPbU1v/sgcUun+z593
3goPV/WTo6W6u8IMskgTJZvNd8kZLDFDmuwbmwjjQFxspuLwjGhnWlFgvlc6QSSr3kjUKvN3FzCg
+4E3XZfL/QvF+4IQ8ZlDGed0Xg2EVBoJFY0MbS2i9vEOkgViYVYx5dDD1a5dn51XUgZyEKoxSfWw
wtR1nlpeIMVCJpGl0Z9W5h/0lHLs1PGDVbcsnB6Aos84bpapP3C3hsyaue1uxXbdSGWYVchUXOEk
B0c/dBGnW8KhrZ7lnSgFDyhb90qxmmDt94sV0k0aSpgVugbA0oe1YVfQFWqze2OBePIp8OiwHYF3
aoYsYX2FNWi1g3397P2Al/tHRHPKBD+eyAZ/S1aFuwWwVtC3hC2MpO8c6qNv8wgn16FZQgjWrVFC
VhDDB00bL9t+QeDfqwgjqrcBEvkEaZCKpa5JOi6O60teKnsQyrWln6tXRCcxUb6QkYaGastSyAvk
Po86kzzw2aVV/kfMqxWn8vq7OFj2TowVOcDiP02SXmh8CWQ2r74hbDcp4sQzd+BEh5OEr+oaPYFL
IlPAigTFfhvrVy1FR6pLv9jqSVo5/pyCE+W1PmQ8bzuBUQvJMLa/nYQXd3RaW6auXEFtglDwN2/Y
C/9ORqT+XPJCLbLZSIYuUr6183QUdqfAxgZaBotW+QffUmQfR6mMOAjtzhg5UY1p7W5rlH14MgPg
DHKCRVQ8JZp5uNxtRvECrVpruk5wgQzDpjrTkKuvw6IHNXYcMU7LWWSWCzirjqz8tUDi7GMm6AeW
2o9ksQ2Oa+VKF9puVOtnBSwENtWDl+QeUSwdDHc4mCaUJq6+rhhRMYI6mkLgi6tphemF4+dclv8S
QCPObBtE8etBIgAb2N/7IuMohZx4Ozaw0hNIEHhFgbiu4IK3JRV2/K7fDM3UaW4NrwXniK8dIuBu
FNQThkDbM1SNxWzwC22d2x6uI+zd4uIsYCaB4p+iDQW0+wnfXjJiZdIJ+camtsUGIVyXpJkkW8Qg
mD6JXbvdDcR3C+Zy750Jx+oFGsRigU91kbYUfrgXDnE0TKoyJSheLsr8rJp1svwCodCQGq2g/xpH
C+UfB7fjN+umkdWLeteQhC1/jB6cmKOMBHrkS7QJfWmQeJtu+ZKfrJGBNHxPGzwd81ku/CxH/EMJ
2IpbFMyXU2+cpmZsM0tArZp0A26r+DBtriMSsfUpqkgUP6oPFOS/zpFRiXfZANfhuWtzsYtRXXWY
eVlmF3zo6CLcwo1/abR9ougllhM2rJ8q49ordleQ/NjUp9j8fyLAqHCiVVX0vT6gY7QcIHuFvx4L
gPZzDfkl+tCeFBRTPJnQku+xXIS443o2Fop7838ziSV9hKYDbVvhLv5sfdBQ0+GoHBXI0w6By/dF
6erPdDJDE9+C0405efBehjIK4efC2R5sWf+Wc97j7ecKXWgTk4Qjnp9IcessFqBws1F+lMK7qi4L
2Ek5v2r4SPjoKPFE/siC4XBcIGX7r1rU26TX3FW0k9JImtpZ0ewEGwWP8hFQ4/ffC2ikYb3JnIMz
0KQmDjMaIAxzpaQgJDfXNYon1h5MxCERbJuZwMN5+TPW35Sd6FREWMGoYoanZ967IYLPyZXijyWi
v3gKZq5+mTPo9/kdX8iSjZQU20nxKgCvy62LNZbNzKdC4UtULsPjclFRTw8F0h9b836LjoVFJG02
qudwfWEgL1C7mmFsVbK1SO/9sMu0shNNT8CLSMpp77hwqY29ICZfdfkojO+kUUCcg9qYsMQkPJ9g
vTv2Srr8yf1nTMCrSxdzWabvbdyhojbOe76iyZkrKp3jNrqfd9vaF5mRQcbSvrFIEzIj4SrAtJ+O
iV/gU8i7ln8YKvonEedZsducNxGrgGyVkNjoROVkAl1iuML/oSv4nwm57MBz3S+ZjxkgPVuRxAbX
gz/NfONif+pmU3c2F7OOeFmMqRdzdqYcRoLoTLceENkcUJPoNj0jv3R7WzYubUuF2xpISwcyj2ZR
kF7kXtGR/HtQVe7bLDHn5HWsjx2amiaDYyMZr9dPmEMOrPJm8wIwGf9/qGRvxnk6g1lNlDL1gve6
UVb7pQkMbqWe3U68H/PFuoJ9Bkoh5LVrJEi6z1/ucer/gFG6eOnH/dbyHc8buYK6lHfiR+qDUu25
LlRiB3ZiPIKWgKIb3BNHxpaIWUtL6CmV2cdJz6FRXfpAI2qjlv+yNbsGf+ZeGj+3TjgWc63JOlSd
ZZfvNFuQ1jYJ9YDqubp6OaWf6H5Kh58Q7oBKdlnf5+BpxmZe7mnuLptYE5oU8qV56afq2pPLBzN3
Y6dIVomqsZ/I5GklAiVzK23lA0BOvDVycU3I/6FPUKr5JH8QuD0uLPD/e7BNI+D9RGbs9CxlZGcT
j8/f9VWteM32Pre93vEdok72B6hnELBG+ltimkASkkxMS/jQV46act9hQD3LYy2LgkzaTJbsPZSw
1qGLIqxttmnEDr1i9xFLiqRCzfdCR+MltnNQaM8Dzo0/m79BO/uF6ABnCRm3CaVCJQIBbmdwGv4j
Xo6nOIs4Grmdv2GVlpkZK7SAK5UOd/W58MvNyUlNChr4jjdVMJruXHSQyZEdf9rXOr2PNGfeNQXJ
gf/gMeFRn9j/BAEzXhqe/BuvY9DMSIdQroVkjppcsklElb8z5YJqbFoowS4dZhDorG2L0sBQbL0t
RV71LxXgzkStj07AaqMrUBMbMcEyUOG/WcFeJYxkuMwVbu2b7cr5JhLWfYqaVngFTBH2iCRewpIC
LQoU7cZ2XKVITVyJTfoJP1iLP9J/NyYKEVRv7GvH23el6TXB/hq28TFjn3Igp/+Roz33vTy6UI7a
ryFj4oSnvpyOM+THg0lpuMo2kLUHBc5af7ZUlMrCYK4ccRcb3QQE638t1w1s0jYBZLKIZOD15rDJ
DLy1cRthQpc2XdVxYwJM5A+e5GTVQNrvdCf6TW3w83jJZbvHKoVcQHV9ojY6tXbd3HK10Jiv0AuT
xECtkW+ME2XxiEQFjPBtvP5WUdJslp/ODJib6B0gAI/ynqua8pYVSPMijDuV0zld7/11IhjdwIZr
v+gt/ARufCw6s7dBJjELBHbKhuJOXDYXygubnR5sxyi2vbsP0b10NkgqjHM74s+txYqt5Xo4KREU
JlX9LlVZeBhwPvMUFojrmjY6Eo9uG1CsaBYhJdhvzxC/3iya8Ecv9CAy8RuZBNYjzACv2745vKL0
T3ErXcYTZqMQfzFve8HvD4jCheKWfNPbfurCXWegMjTydwOVgoI/TAQc523tmfXtf1V1yiGk57JD
9hCofvJQ4hccunufzLKYDQ+9Tke6eRurcKP0NhTFqeezbWXfWfLadQS8XwmnaJhXrZGDsJhjnp/g
zUheZkW8g0iUkT+YA9XQoBr2VKYSJTT8cIZzXoZmLqX1WoaTta1ovpAMcLLXDuroDw3wPf18mVcX
paEh5WRpAgfV1brubdAhm1QLheeH22wwlXczcHsOiiKhMT5jnif2dRXVjwz3C3ntCd9LQo9Bkx+F
Xl7Zy6SAjr/Ko2/UTsKaq1q7EjoVzzcubO+J0HxC+mfRRdzoWg6hBumTIA6MvVfjGg9BJrlOy3Rj
17XyvF11GiQ/+fFmExPLfD1/uoiB8WPR/GubHWmBhDKly/HIVtVg/XebhsyEhGcf7N796xBvKKI/
g6P7Q20NwteaQU+6REbKQUq5BMw2Gw44h03lH08DZPeltFBxrMgpBq+kR3r6cge52tTpuXSDzWc9
vrYGqkswvR+T6Xiw17q+ycaYM4KEc2S4oa9QSmFIIwWxRBv7WXQ+ZsvMfu1+cytOQ5upJYwNuwQG
UhhiufzwXgpg6n+HHCa8fiDxxHVRru8GdQr5NATSp9Ww3n/pgoQ+MPbwGSSTiL7BZaEuQsmzUrHR
U/OL4s4GdLmFqpJXrJkj/2NF1t8BD0Y7RxFYuJM0Z5hOOPuEUh9C2t0Y7uRGox6iyhgbWAr+RMBx
9IMdxFR2cFZgPa0MPb3bZlNmpiY/eKFgGQKFar5dUUInXSGJBAZHQ2OwsaQ2p4byuqQlm648WUnr
mOmMiJ2wKo2gNVkAgLdI0HEJKShef2LIfF14Ksk5RB4FZRTM2HNjd6SDhp+fxfDroSiTMj+bKiJD
XnK4Moc7w66ov45tew0BlefVseOokf+M1jkKxB5IH0bHIxWdYHA3SdTQbQDgFF27GN/LBJDbl/aY
xs51etUha4AogQSapzaJxOg8CMtvci+mLYFwxg3874rzgyROlitgOTQtu2HA7qz4UF3pRkUmr2yU
w0mC2UDLQ28MPtTtpqWrIM+Vt0gchqb1DX2iZGy7sPpnDrnfCiv4tFHfJWNj1HPjue68JVP+GpOW
DQjFzVnzHyI7f3UNwtAhwfvIkIo+WHTkj5eO3hCQzsZ+BeEEGo8B1aSZs9S43Y/+ZSYfTlaBGH5e
OZ4ys7O8CakZ3JOGIpKkv5UfwuC4RLAWIoFvVKNntCwy20kQcn51GOKwyVtHPCVjp7ZiHG7UEaYr
QV/TJgSzNN+cjKUefQ7H+Z8HfCSK+BOH5rNyh1YiVE6viqoldowx3wE+qLlfm3FfPrrG69OMTQRP
d/FzfI84BDtXEQQWsFiYStbcBzbKuDTUbhvoU+zwTTsRw5JfOcs6aq2eWry5y1ZIO3m7CMyOBzJK
+bllwyDqIlNBEXmcrbbqoMMEy+JPTbJZZsYgDt5BV4VZ7hPeETlTu2aApXwlxru7Kq0DFluIMnOS
Snx+13t9dF7hFI6P6OZS5ixBtZt1+jZWWJPoEfxl4U0PlAl3TfRcc3j1T4HL/NinTXPBwERiWtTL
iqBlvXHD1KyyfIkU1fPpqa0bQSqBlwus0TRLaF8XTdVGvBbaaep4VWtsydtoPrbYfS9NTM6jVdG0
vhs6KwmsXzf6xDq35Kp3qPe7Vn1kRGEXBiMqiRWNZn4dHgztnRifk6Y4Z46GUkaPK09hBDE8pMpS
E/bVozqUOKrbhP5rBm2IuNbkei4ZtL9dqLTR9+SWuM6fOF7Uw/A1M3F4CXgZ16NQdSIazLY5yrCr
hJTvMOgEFn5Yt3KP8Jrd98V/ivplGLZ3GzqiW0ffqkGMDrNoQj7S92hHIAXPZus+PPWS+12AB+Jy
xle3QcN1M255glxUW2t+htzvOx1Np+WeFpOlbiESny78Xq3QbfG6Od2ibyljGXTdy7Wn5zC0oA4o
lbUXr31QWCW4lf0WTSzit9yPSHwqEkJWTeWurhddi0WE/igLy1H8oh6jkzMYo6L1gXdYGqzk9GF6
I1u7fijOcwaXrPj0soDQmfkLE2BeepYEGAjgC48RYC9KsM0t0xfU/+aASWeH30Cc/EBr25wA3fe+
CglDHFvN5kr2+MBoiyqS9H1ySud+JCEKst4LadQ9Cuml7VAD37huJUBTr5D0MNiEhLEIRDrv+1Ub
KETSCfOLAi34mwzkg7nmJkoWcqDlHXqwlJ3sPsXoeSgic/a/sXhKshb5LPxyOxsze23t00kwc8FI
a9zOXp6Y5L6DOvUFYDxhe1ItZKqP5wfvCZ6q+pFXepCCLU+aSJGE+gUYu9YO98m8n+xLtmSuxUhd
IBRqfAouFSyUgZ4ofnpqzADdzdboA3xpw5OSNbimnH9g4cv7YxMJ0YYQDfVvkwXicW0MmEob1vdo
vlscLc8D847+JDtVWP2YmYOdVEbMbv1vY6UXfsMsVkzj8e/G3ML4MoypO2Wh0CbPgq44CwRRYfH5
GyxIsCQ8tNWkv2b4MR5pXfrIH8PcmOYr/Z2ELaarByZ4s1Xkhbbr5cHLtdvkxZa/MDilrmW6H9vg
YrVvsJGNf3gi2YrOyC23dEsro75nzT6qYvhw9cOTjQAr4vnQUtQRwXppuWAiWjTrgHm2gv0udWde
4k6WOF2LTgfUx2+dXKXfkRMm8Kam9SPGSBu95I1n3J/5PWNjtHi0ikPawbO7yZ651S7zux3dte7o
JnoIrBMBCFaCpiRFW5oFqpVIrK2NEkwn+5OgW5ET78UxcOhD8Lo+8Qbjb0ZagontoA+9rPcgVnpG
8wopKKOsC5eqxMopq8BwLpx8HvqEOu8tfVYtZSRyJN1rakjyPfZsvH1v5vhaALO+T+ol53DIjCSa
lzb7Tqn/ivt5xaTu9l+efyQW0++ZVs/nMvBS4xrEjNFC6+h9JBYtK8vit2XAcOeOd4t8KuDKWP02
Wc9Wx3egssuILlDiSS6tsPUBRig/yYLOLilXD0nNDaIOW5fPzXTymj1iTyNAUJLraij6T7f4xc3E
JUNW8ydEEr/I24gvJCYSUUVqpc/gxLyPYypEECAkPB4tacTRteWTF1P99o5heqQFpVnzEMU5aM6l
i6qgY4J2Mse77fwimud7mYykvWhU9+QOXMX2jUFjEvJZGAkRwwLIkoyRyCZaCXCwcPcNsoRpag/J
XdaphzARjGVCbGVZVW6ui5uwP0aCJelmddMYhid58wtQ1IYoB0pt45zZuSdCPPsufjPhw/G83rys
paNGX5o1alMLgckS620+OBFBPVvtQBmRycF1jkzdVFoByKKGbb43V8JWzPxWedUbqvV9HB7kgoU4
7BDtzKyweC7e8xeOz/hRgteJVhO5EFzN/z4gK8tEGTLI5sAgmRigdG3DcI8ayixt8I01/sMNudcl
g42Y9WJBS5bgajRBlLY+48jtxU8Z2UdGHtfNT6of6W60f7mNOpgQuZgGFKjdp6Er1fGVs2zCK3C+
x2ZWT61eCNAry7AA629hon31oPANElqjBqH/pLGVNXqqt2TBQwouV030xDITvdpHBGf0H6CSPIdx
dJy0MlYzFHO2FaXVRh5Uam1Hnfi4ySKfeRwe5ANb08cs6LR+idVFSaQsqyLUjjfVPXf3eVz2HdRT
jEuiU+E3IfvitmlVXxjQgQGOhKZXjT4wdofX9Np+s3NbH7S+wC0Rtwx+KOyA5ZVUumMed7MOWDYv
f2E6qckksZMNpdiDH5k2sD4l/qn5TrMa98jIsyQHPZTNfcvweilvrTfSuC05yqvMpaNcEWcE83t4
+ByeS0wD1VQAxYQWMxwogBpjKBhSHjN1um34SStt8RXUkh4v4YyD+FEWtJQciUG1KXX1UM05/RvM
FUk/ZW9oowL7zRrw4xATI2hdPK6fVRNjt/bEw6mWLxeECMsAU+Rl4NclzuJlALgZR4YJSqo9Dvz5
M+oogftorzvHxa4ICCTwepdziEcRrykDTCROhaEIW/YXlfl+bt2meDlL2cPWH63JmoEAaBnuVLGH
zXQK5fNephEVIiatoWP3eidLYZhQJZMWpdHPsAJbj6e8im+C1vGR31LTGopC5XxfQNNfa0uMu2+y
RUd5IYnJbqslE1VwMmzAOmDMvTOfKZR3Ll570P9fzhik2VfBSwDQng2C/MavBut82cqoFOIjF8uc
jyum16VOhEpcGV6AzHZCTspn/AoCsyr73xw3C9UlSZ+pYeE/gxMyOU3bmUNZIMIvja/qDCCDKh5u
yMEr+yarKSl+dUY12itEziVnHimPybtQmlq2xDFyc6U6KN37/DpY7V5tHFDQxmLm+RDYbhcFqyU5
/4oFsYbbF5Yv33WlRt+cbsAsQz+zlX+83eCzo/gUuB3jOhOKu/oVmiPS1x+Jn+ZPBBatZdL71Y0w
FSdQxruR9xi+FOYnmr+pNmQRorCzK4fYkWziGA6H7M7ew+Z+tTLfu5gKVnTXr5GZpPWdocukLjpy
O1o1fW8BrInRZV5qvsa4hHoC3AujLkH9BU1P+gcguNg8Uy2a2aDIGY8CK84Up39yss9lGezOEzl4
SlDqjw1JBs9Tx2ZmYXqUIpNoBvJZpAWn7ZCtGLZKCnxzp9esQ2Csxli22MMFEaet8T5EQhHOClNf
lpnOY3/ys+Rc3OecuaUYRTHJRq8AZ8UjwQqSw3KDCBmOqREQKZFTweJDrCJauXcRY8r3TvUoKaGy
3zInaoIBZmR7M1EGeaHFbzn87PAwjXNscGd1wcHHrs0WQc7lU03Nv3fvPty/71iYROE+dRPugcSy
oR0VND/EU6n7V5pn25HbU/HfFBZGg9aEEkA2BndZJJ7dIj7GuL55e5wudqZSvECtHN91vALfDVes
stgHNPmLLQAuAIMaz0VqbWa2fgJAhGTjkdFzkR2bHESpHvB0RFHZp5I0qkwxmIYb/dmmZC5hW4xf
ZHZPiFj0ayHk3XzPMLCe+e+dAcME07ulmv+e22A9Qw6NaYom+556WZZabU/MuhIwMv+0yfxq+/y4
k2bBlmq1Qhs6hlDcOel5+eD529hhdf6oTe+ObKxjdue8y4ahhs7IJ19zXp+MqYLeHNUfYJ4KeOpE
DKTQP86//0ukFnsRBOGWgDoWgExH6WQEYhiTNO1SGvyBCDT7xJ4EEG/1hhREIVb7kPx18bT7JWZr
v1qRouLkuTcFIfGnVZUI+KpGkT6Uq3Kqj0gsz+30Lk+Ii6D6LGvtSeW6vs6AUYwVtV4zJFBDo4iU
PNDEzLN7pzh0UQ6K93XYHaHLg3Lz4v57nWp3WiuA82sDCekf+i5Bab7n3bVxqCNK6gZWM2oASjsX
m5tr9EpmhJwhaFhnD0LKnYo4bYR1TWPpfj8jliaozL5L67vAUVz0vV2JRU8SN6TTzPVNW2/C6z11
cWzj7g03fZ2vMpsoJLoVHJCTiISdeDfFuI95PGh6BR9R3UhGVz4ZVusemLcab1kOXLadSKUQyTZP
tDez9ShdEs/vCsfFsOegH/JJpNi07LxNaMtSCJoG18kGshxSDl8G0nAZjnUSYmfnoAaA/sj57xus
LwsAdms+W0K4g8wild5FJDqWEOpwM931HWksUWZ6jUmte/erB6X3gw1Ci7TOgfg8oTxRm0tI3/rp
kYMwx/YbfLExtPYECd325OxoyyY8dcJOkI7Ev2fbK411HuEYcQVZLT8KIyrBIOv+ibrQ8ZxTOgHn
tSzCXR3Im/6iQa46Kev1+Bbkq42xEX7NGeSW27g9H4akXjCBoV7NqeE/bm6H//gisoJouDTmf2W4
j1kU34dc+XGgUN2uAXqWnh/SVuwVXDoOZ3fsclJGEjGBnDGT+LVYmYxYAFiqoEzVutofBc1AIT8z
weUd8lIWka+hQWBfrqWzkrPK+o45BbC2WwCEvX+wMgpchousfZVNXVOyV/df3vMTiqSqstdAoX1u
zfr7Ler71cNufeC9YFEU8e6YGa7FNwL/UUUltcL0kJgJ8YXuG0bRNCj5FlgaurrfE0HSeeonLe8K
k7dEFrqmjUEBd6afqw/L1Yo3u7/ED4qUelmIQ3bZFTFPomjbZrKGPJ56W8aVQ6esNpcb/GazfVMF
dIbDCapRK6FVqWDXHj/Ems97akJkhvcp9w3DK6rFXWlWTOTFCao1R+QMLyzJWI0uqCOvEwMd+b5Q
YHuwrSQh11d4amv+VNTfpeF+SLb3lO2t8kpEJ3BvQqFCBfZZqTth8sNxPBAOSMcs+UhVWC2dA9Oo
qnB9HZiyT2G7f6PhUepUNfQJcPBpD3ffEq/+eeLLSNTc6rcoJV2MB9rlJr1XKb6D+/gukoD39hvg
SUdgk7Ii0UXzhG/fx4jkCw30aWQGIlupsiQKpRYNOJz4gmN/HL5gh4pWq48tCcejLagYBJlC/vHV
6uQoZz53lr0Tt9AeVIRrXK9NZoQRBS8b4PYxs6iTfrkHZFK8gfu/rFfpjurv9dbOW+t0bct8U8Hq
jfuDzEZRzCugRJxCNKqYgA0TIEPmwQKvzXRy3tIrSoPoNDGHNr3PtS2//cgc9F1kPsiK4m8TwyVN
D+VOP7QI52PDa6U6c79bUOmTyHcw7jAA4nNoluNU5y7Qcuar/BEAQRxVZksTnfEipXZqxTbbMZZp
7NLMykojVtGR0fXIdUdhOAISk4EpYt8BWLphhgHCnPeliW9CGUXTi8ZzTfkP+mp0HyA2oqEa1QTS
MhlrtmFvxLNexqU2wyYml9J049jPjCTRbnnVXHflBmb7B+zwQiG+2Mw1Qj8v3UEgsZU/TO+4DchS
OB/IBvYci4dF55TZ6IZmmLo+ThLw7jFLJrjEdk5UdfintA2EZ85WgfcdS6jxu32M1gZXtnd8546x
+RBTj9kBDhIDxsSn8diHPqMkdf8HieAe8KW+ZU6f+Mp2ha7tye1Iq9ScUXjyEqlSfGCnxuy7bis8
xvaU03NbSgjkiJr043TPhFEonzS0anIAQbhimJfqRCeQRmyTmLPx5HNu6Sy+70r7VZfrihXtAXfs
ZZ9rFAH/Jx90boJOxDGWlYCxlZM6tsw0JUNuQB87DP8fc5tG5SHNE7CyGregVfsTkXzIz10bFHnS
/oaY7MxrWrhpYdNBdB+qNuWA9zsRascaCdpEYwqiVoNqRsERELyBF0rXJUSkrymoUNs77d3DTamx
7r1F5tv+0YoPUB9x/BXhUV5rsnUv/WD8MWR/nk7+DbGHMgp8e7AVxgl06Tb/nnKX3+zRS2GVhBbR
YAsaZK1b0zJkixfTsMmcz0c8BYTTdaYd8eLvesIRFqKQkIOoqxq1sUFJWMPLEMje8C/8NUzzbpA2
7iEZOnFokDtc/VxgNrlT51+VukObDuL3ov5Qxq4AV4VMf0YvmCE44OEQ1vV70kLX9K5jqzVx9fdo
P3cApUUs7GPBALhDeHfn66dxRmpmup701my3Rlsi3/QpVOCFBBp2K3rVh7ZPnBAgHEcgDFCIwvKD
ez0kDuehBfLDQlCPvzPefglTnlhQier6drqtG7C1Vgz/S31NpHuknZc+WicAlHUalU/brvClAYhv
jkLPCHeguxN4CdWkS6I1RATfysLAgXLoh0WCp/Mn2KhOkh9V1iBdlU9J65EdoATD2++EyGdyFgA4
rqVt87Hq4rUWVk1pLV/F99w/VKsdH8aiBjJU2kN36lLVFaVwpx8h/4qQXNzwUVvsCpCP4i/vqr7V
b4wEggP+NjcAba5+f/JOKindO2ddlFZP3M2W+hJ5gCM7YMM+bQjX5/CmBA+ilEwP8j9gn88u4hq3
sp2rTh5Mtgd0hJMOuHXbBQ1yaALAo5w6QartPky2osczxLAWDScPfSZEBa6iDENfsjckuuAxZ3cW
3v4Aoqzg+00Sgxy1/ShRp7Gc6STauzz03bXPa/Rn0+WeRHhxMZiDlQNx/PXMP84WvfyfaYzCgNVB
TFeHVkEfFALCNGS/izLYDiGcpOKn1eQOkCdUoNCDZ/B7OAhZ/m9KSYY+JqOl178lTLgn7sLNk31o
umHnpAjRIY8hDJK4scaVEn2P8ZEIqFBdlzvKSbkP3dzaQHOirKBKc0gUMrKUK4TixVAVfJKY3pEN
YzHsCSuPid0IARa6+4RrMbp+GEfU1lpneidgOaA7dmRxzHArCSxIqujxdI4HdyqcSigsbFOdp4z4
q5EOL5dup5EzABHpRTOLQyHt6kIf59Rsi6vIW2UYETXKDeMus2st2QOKTj1AgwUS7MSIR9iyND4N
PJTCt5J8p7GnR0sUawPPhTNSTEnjI9W8pzc6wy8xjXqauizczJeQDzXVXqPmEW855fSvNyLYy5Vj
x97gPpLLZ5TAedRpHT91rJlRnjXIg0ZYxrAcIEb86tkhmSSlI0V0CWtfpsiL4aimqKafaH9sxXx+
jVTVUZlO/cEmRWsIoK7keX8jQy9Wsp9Q5sKD2ytBTRbnFeJBGj3hFdqMkw48lXXQa6slEnvPKfgH
IsxCpaL3wb4fVopYer1t3jvMsZBvdGa/TVTrBWNh61llUYJTuWJvmukTDGHkpblrbIkSGN1jrxoI
Th7csMnxA1ssbl20ZlYDh774EiVBeEAEngfKwQ6qpRy2DLm1p3GGohVYdc7+bRe/0Sm4tx3dA5iN
KYuTZy5d5B0//f6RuKhceRjJ7cbo9MWrqnLDVb92XBoVv6jn+oFUWLeRXrhsGvaRGNmeEIAhNpFq
0C3bxi5QpdkwycXiPkn6xTjMdSDnUokvZYIcOLcuiAt+qijuJE+8uwEiT8cuy5b/AgzZZ0i69uIn
uzIORZiu7XiRUwfup2j806exCsDY9F3eufK3gXv0luTroHCm+JnmLN8evlnzeI3qLYx+muhTzxHb
/9qzZXi6pwDnmWB1CyJ8Xtl612cYYD8gYLILm/aumENpLRhqGBA2JqQEoAKTJL10wXxCyPvs6a2f
AoLe+A0XxLl1vBdl3zhqEG/zsdwy88TfsUm0GnbIt8ZMYGSMGLMcuULRgQZNjrmFCgKJmPwtrHi4
tZI7Rh/zGpBYsn89jcaUyi9SqfAQZ+/7jQSRYqADog8Y0yyz1pE1DU3uAXFO4pF5EKrw3LoBCrjo
HsUa9chHxfO0lFF8O7edf3k/awERHSQk060kC4jeP9XxbxivzvETNvbhR9f8bWiS3NM60Uq64IwG
04a/PlGfv9QWfMTb6VfpvuIUKTz5AdxWkdBK15BUsplRI+YfNtFWMCWw12ag1Wn7vonmrhpQEvcE
VI0AdbFhRZxE0aiIcq9M3x9HZaxR5WxFdjdV0dJzaf2AiFEwy2SpOmaPW9qN+UMLDm40w9q933I3
aMAH1afCHxUjRhP+OLpCEDePLvCBf+iVWioosYQ5TeelbeWCEUXWNnbOFMO2MYss50HNpG0wNTI0
Rvi6J5OQNDxWPDH6IRSgTBOChMB1m0jP85gOfE25vktSSGNS36947AgzqqzHLtl/m6vkNYiibCoB
5W+C314bc1/ACSGlLn6qpGq4bH4hJGnhgaE2++Qq2E2gES6T9oH6mdpKK1fLymMpnrjZnP12/2YT
IkZJoyXBrp1dRGmvSuo2P5rm43DYC6R+U3Fo7nTkQrARa6vAH3+HaFpb2MWsseF3p1JR7fJ1pu2A
gJr/H6iNoLNIp/Jyf7gZd+Hite6ZTmAR/Q/pdF68D5EJavhWmdHxB0KOi+Fmx/jL998g86Vo3FSC
RKPfYls5xz3m8geR1EvL1j/xGKuhkNc3dKtRXlbQIer5WXUlOmbZlgPnp2pN3EaakhrkPURx9Cam
VV0B2Et83MWGXBwXmMjTnFDkdekwb45N3N5szkyKJut3oZ1xfryKBpbFwfWyrvPno1OuTvffDoRk
QrpD7CsxgCe/rMy0FHL4IGVKVcS1ZXj2ruytkio0C6BZqPLB1nNY0N7I/hT4J7pmJSWVmkiNDixj
Roe3OKeb5JAUO1oRruFqErr620Y8XOvrX28QCf1qfPMu12F1qyO7uwei8lSK6/JUSRrAbyuQPNYV
3M2VgH+PzWqrG9/ygnTvHQy2EC7hepuIdU+i2tyjKRNeBCMk7bTSjrKAnGRtRjcHjzCdV5YomWWw
T6RcgL4wfpjf/1RyPYMjVhBhb58CLrMqJsMkBqMKTmzEIlH00EFIl5BEhIpHOCcTzZINS8Og3OT1
+zOfaTtg+UINRfUJMpGT2/oT5SnV5LHzj1NKtfYierIYGRBpoqS6fLJpiEQTvrWg+rPECz9I6xc/
BZkGI0Jm03Xy5JcdKx9SKLp+GFrbxX9xWPgP+ZqqAiQO+DXz1P/HAbqfn1fAR62dVncHkOfNqzfy
SOzxwWpe6eLY35ZyNwjt8+OOILyGkaiVQXQUBV4C+worKWPfBZIbX4UxZU66+Azjk0Nb+QJxqCBE
0f5b53kH4PB9b2enqpuBlCcV3u2aU+Iz0sB5VvvczpQ5I0E1bSbRVEL0JK1dwHl0Hlmb0oLdMNUn
eIAORLLLZ2g9sGIQ0JTI55Q+dGhSg43Gyyb159cDrAVejW2gp1nIa3XiQnNhaENJoqdZcamerMEB
/ElTQNYQO3cAsAM1qQ9Gt8fYNjbur+fysBSAmdqj8QxdFDh8ac8ySD0MxIAEAXPhBXJSzRdkz9AA
+YmpEekjbE6yE1c5Y8DlnDzrd97CYIORCyiBMrk6CyanScjIbRSnpIY3lrDuXwXcXYFc8+rg+qM4
Rpaao3SFvJ0urbMPjPWApQvCXvI9Umyf23iv+gtJ3dMkPLdOsVsrZDBhbnjKfyjvsCENkrzKTTKl
oUAwz4wPM1BXPqX1DO9eEawWtTXYBIkWg0+pByXNl1fujzOK3sknByD9Yu0lGefuf35xH16hP8Tx
4HPVOFo7WInPkbEH/PAfOIX40DXLaWr5utlIlplcfmjJFLLP+M+7bqyLOTiu97fUMYFdIUo3fMSb
1+O8eBnHQyNevGU1MfIICCu+3OHKJsBfa9+s2lXeV9SRerEpalp52vFwg5WHl1WtBCAY4dss9dUs
UPAanGMAfe/naImwQxvRZwoalO5uabL0lhan5G4zXOzCYKIQxqRSUqmDegXK1wf5p8HtI6lXYFjs
aD4EedMwSCrytV8KhdCiHByza7hP8V+27NZkrfakExTipQFL6Rfkp2pcIc/ohizPYBOzDpszvj+W
gbKJymm9E1AjS+i3zDsAq+4EJ1wiNdt21S6FxNEALzHKP8mxvam0R+VnOXlAKN0LCp4xJUGfmleG
oB4toUJWG06hLRH/DRqjUa6Y/d6VYMjoUKMmAaJ1yyA9YeFqmRoFKDD57USUEgU/bL0XyNZatOkF
zJTPK1wHYbskDCuQZtZmRwoy38lzwNdoAv927kI2WasuX0N6OEy7AmfIBKbmYppkmVfYQR5cWAen
PsC95Ja7cIpQBSnQ0uEg1i0HrgYgIIY8t0UEospmtn44AIorerbcFrX9r+iZPuWgm9EnKtyiCsL2
EiWQQCfx/248+DM0qpE1Zb7ZknCAm0ix3xQv1fQGJJTClzCCxR9OCCvYX232fngIhA3uVcfBTRER
WG75AaD8PADM7F2fKQ+S0EYGD/zWwkOV7YuTy0td2LH5mzdmVV1x1eZrI4XuSD5wge7x2SeX0LhH
tVvtlbiTvHvFLP+wEs8izZHSEX0Ue0j0vL8julQ4BaHlluhFRaoxnKbVF+TiEo6VDWG9oMik6eJ7
w/wBRVt0p5cGfoHUS87l81iuaNVck25vDtD6GTDVfLj0AFP/GWRnqqHPKv4IP9aiyxMptmgjLZHj
vSIwSM+pgMIJkBOUxt/t68rMPGtu7ZBWKObZhaGlwpvQy7o/kJJHIHyODfVToXiGVqaAIpEEfhon
xgQsNkf6iJZv44lNx5aSMM6jAoDfp5fchUVDKZQlfYzOm0knbRlwC/PWzUHIXawiHCgCiZkt2+OT
IqsGrlLsSeqqQyZwWgt/HpkxAzodabRHULuLTMtkdZDhOmk4VCi1tX9wPedM2cewZQntM8pjIIYQ
InOJ7GqvlGJ9r6BD5dg0cdY969wRzCiULJphOEyp6XC0cISQ/q6aXrqb2g2gJW7dGjqQnBGVbur1
DsqGgp7v6oypr1rmnD95ulLB/FmrGimeUsviY/SOXejqkPpn5+URJwMxKJGrm5wxcTD53ylB139u
+ePsHfw7OrU/G6+fkX4OME40buWB/WWihqhDWfkhuo9WWlYjoNsU4scFQyvwfClsZMtmb5w4o3Bb
kUQc46dkW3bSKy0wjzl7hfbmKOyqWoh3TXtYmWwndtIiRWMKF+CSBliNHwO9frwElLA0wf+Wagy9
mO6KSB11r6/lwpydDp8xURymfisqGTsxplt58VlDKhA8MrydV8HAVhkkB/vrUlnB07oh6O4s+th+
lQnBhJrRVMl1ejrolLS658RZO4DUchP0uqddnYY6H/rOIyFeeR8wWWXBguMCl7L2z/N2PapW7gNZ
zGvacDsXS/9xIDCglmY5qSxvqJ4rw07XYNEjQhtvAWPpRBOIefHbZ449nZY7otAr2TZh0WBLoROJ
BEOpqrm1QQLoJVuptssDjmXalpf8JO2r7qR30OaJxIPpW1RL1u48jY9dyM9BQ/zyrKx10ggWX8KF
tGD40j5ohg/vQS71TVAL9UHLD9356a81pXv0B8y1kCk4Phlya9CnOyPUsI4KivGcKg2Wdgpf+zfW
W/USAeS6CKZ26Hdc+UJpmBBfnA+bjm9dEGSUCXAkFHqDlEk4krSmHMOsJdZR+DAT1RdjtM7WihBQ
qcyM7if4OfRXBY0iU3eJecWfDPLmmZv5dQgVVCET/c6kxXfeu1AwgMaafpFYCLXVUbvvYJ39VWXK
2rxxIsxo5sZ/XpcLj+iq6gQ93cwUJw18/3XQALUCiEHcWAZnn+T/oKNm1yt/uAMaADAll7AYuG1k
joJ/Fj8bLxIY0hRMdsL2vhxbH961MqX96zuGreaxfCmusxGoe4CLzp1OrZvtaedU3vW3ERe+M4mp
s0yFOsshnMmFnWfwMmR+blR7qWWC0XSyisPWPsgbwLRvRtL9N4tjPzZsYQdtb5AHpp80o5EtyoE/
by22mzxovanmzMr1jthNBFMISA00kGk2v6HuzQN0VpGJuTxwKNgJ09d3/6JSipFssu0wnGa9v9Rs
Tx/CLPN/vqIM7/U4W3T1jz91Mf8WTk26t/dQeAlIGoEWFWtVfihy27Z9pwqANyur5G57syt2UaH0
wO2NDvw6NP6jECdYelrUBK1YUf032B4f+S2A+0yH2hHvxlBlrnZ19vRLoziq0MBEKET58t0Qqi4w
EtWQK1Fw0Pw53Q4JvUIq0fOHpYnQSUZRqAcNyvRJ7Tcnb/lqm+zNiP4slua8sOf2Y6tPg7HJfpZP
uAEP2hOxX03g25PGQ0IxrYEsHuMyVsNoHbVIHIWrI5o2KEqnYaxFMO8RqTO/hWCHGTXLASXeHbT/
8KzF9IZ2+xJE+6CctzWOGk2Pe0VNKYBg0Sf0GgiamWzr9D50icCqQd5ynkz7ArlM17Wb3s2cRtfV
IYZ/f9QQXI4Zwr5pZpQYi5KUM4ny1jj1S7z9fn8bM6dTOCAclDHowCY6zpOT28h2uM0ts7l+bm4v
R0bJjvivt9TLqC9QtnULP2S7TKpnffo+wT1k5ysvH2rgx0bcsnSumoqxDPfDYYoJCuFCxWJz4Vgw
z+Rry1LgdfzSil5c2k46VByuaHFxt6O2BtYzmkzAAOpwNGvjNvsofnESxBh0fS2AOeorkFF6+D+P
7YrLb900EHceHDCQ9fKH3DSa5TJ/4v8WEzMCywUkMl6yxtONK5ER51YcCuEzPUNsaagnpu4YqHC3
Pz8V1w2kwb8qDRnJ4juAP8rUx/DjeRkIsWuvdNXVPEfI3aQu6RjvaDexxCZVBpYhk2gtmqm18LLP
TvCQjlsDlSYO+iqBpFGztm3KEH0xLpJ4kgf3CXV5LXmg4N2PvMy25k9oyj96ONvLZp+L/IzTGIoO
paV3Buuc3+Wy5ZqD9MBrhnLPCuRl/o/djDjxoG50bTNLKJqeIN3DrLCRgFwib32Qc+6eBcKoSPKa
CemVq2Fzp/OSwxCZSy7jaqs1RBrdtEeeGaZaYiE+9yB5mrMRhwzUhfJxvft0g8ikwWGG9ndF/fzu
lBqdwMrYkJ5ra1xF8EnrbZdhQD5hh2loL72dMT9RNNLcb0YElf1ckPo0v1f41HAhY82aW2LelsC/
NnnjiX8HFXYQVcVaBX3h4m59ilC/oPRs48+EMj4i3jYOWsXrsuRU3N7JoO1wbkCyNtxUb/046BzM
S9q44HrpMEimuyAtW79ZYjCPhXzMakG8kMEeMXpEdaGtkapoNLEy5+dQziIe7D6Neo3jlS8HYnrG
qtgehsaMHQkJ0ZSfP9ubIMsNrWkz4JxcQ+GI7sz5KGoTO92P74fwB7Vu1209isv61ALn67GhEdy6
ysquwCi04gY/7RcAvKuNSc2Sm8FjWa27Ustql95bfFbogHelj15kCj2z1h+n9Ho+sFL2WydXxdaq
QT+LSh2k9SxriVrrSEKWNL9nXzCXMFcQrWn3jXc8+YNVqX6VhuZor65XwVL6dtzAdgVyZhBLWRrr
/e9uNp1WTlsNeFxNykJUG5wAN/B05pAIaF1aGSaTPP7qjXMz9OG0Nfav7xEsqA8Tfh06QeklnTb4
WHwn2Mkj3/+SAnldGY1ieKJ1i3v6sl7Br/eiIV3iQiZaINAQy2Vo4X5u27VCUxdT2r6Tj0HAmOuc
4S4HUHmldSJtzsn0dP101H2Ynq/Rvekp9dY3X3LOU6n+HNgLurTOod+aEphgAEFDEX2fZysRbSex
mxo/kHIW9QXCXNrN/6vDyKgo5609QRa1WVUxVFsxML8Ee04xGLF4GEFoUtRQ8F9IpZKy1I491bhk
HBPetFXtT2T8+BSPV5xtlC/ghOn6g8JpVsr/NDLPbjz14H1YQVZrf0Qt810+woO9EYQpv7KBQDew
heRlngXHuU2yur107+k2KvWnxoubm6wOsfVlmIVwmlsCQtUP06DMBsteZJ+W+JwfkL/rRLWhHZZw
bnd2LxqM2P9wEf7hn6cr3MiuUi38e85D7vKF1Am8cq66cOUWMw+xZWPKmuCTHVxtsz5yMLoF0SE1
27secDySUh0uZDOO1It7DrgptDmybAN5U3tRShXS7t5GoZS77lakxW4bl5V8xiY3rnjAdiaceMPR
Wepr9yWqUyFwASa4R9VRM1QgYFc6CmC+j+uUHBqBTr+szVLIiZVhcfBBVzjXRGsxkEOD/LEGfAnX
U7Q0bz0C/XdmMNzkaiwxi3H0ttvhS6JiezUd42pdYsxfrWz9Z88NnMUt67m2ZIgJCGuf0u9xxt3U
YPNu1g4WAcyo6UJMLL5zTYXNRX1pweCmmBzKWqGoqi1SQFbYhZhQ/jXNq2DX/Lsp4J1s1ktT/y67
kkcV6GsdqoDb5kF1dNRQL9XTT4/b6Ol1Nd2MjrYkRqHVils+GN6heHhM5qWlHfSLfaebe4inz0n8
Cq8ABswlSOmd0hoksAf8/WktpVPp6o+scHREZV/JFVnebO1YQsp6/m/Mi4C0LwLFoh0QISAZRKNk
xmCU080pcFbrmhM6SvQa0NTcxGKTDHJiWFN/nUvPzG0AR2g5U45baglhXxgqh9nmJ1XslE056U7C
niqtD6vrX2SUVA8EK2SL8wMr4ZGJMWDfFCPbjpIxBHjCVbrT6hnxvRbQdXB5Ctx5VH9bL8nlO8XN
4u3JFNZRJYgaNeyHcbXqIqvnH4k6NHjrmPgpHrKqc0/3OjxeojJY3hX2RCLELu++vW35V+KQyEdy
lmr/boQkOBa4bauOdKtEf8P0MBydGa9pO/9WuNTAsuZ/7tVVu+e2n0yC89WNW4G+dSqimps5O7Ha
HCdM2QE0V2wvYRZ+diRjvqETvdwVUC7Xv9QaZ1GFd4wWedip9O7ZQCb3iZqUMfb5kFUrSX2NM//Q
68XAC0dN1zQFg2dkYBnKF64opHl5VIwKeUVFo9wdeRXHs/FFuLVJr8Aa0pbii32dltsFus6/723K
UTZVZeJjNwtYfajeYRv0CE49/PuNktZDNMjcrEJ9/2s0/FU7KMoOcXX6cNzTWFkcgZ7FCNT4+2Ep
UvOqrwe5oHeHlwCJFfTo3FaKqizsYSLYx/m/g8bA8px0oJQw65etShaxCzvrErHPmXkU57PMf/7T
mTQc6W1Y4ieaLBR7flwanTi8xjPdkC5g8BMM2/YA60f8JVnpkNzNeWpxxvD7E8OcvxqdgikC8EFE
Ktmlgxwh51rk9iuWzZXPIjLhNczl+ITt4XKwEu/atIDAEQzXNhvKDc0x4iL0Q1qAjl38a97DR1rK
zYhDTgkPQsFmg7FJVrLPDterXNOQ8wc09KFJfAZPWfwU529i5WNb9FwH0XWq20AfCZAUm07pwFdl
KbSS4tpFqZtWcJE7enlVk3CIjCXG3SAClmXBCXvSgG2O2Qjm7SgGuyalifINUksVE7BlG5o5aMoz
E9q9Lv8sKoEw0cEaJpnc1egXCli/qRn3Wd3Cpim08dVDXTrggIScb7iahGxrto4Oz0W71urlmK5h
EeaS6ShGnju/NFYmsvUbWmnPetaawuh6zIf2/1Q/bhOdZvirxYKdAkZ7IgEOgEnSFsBPKJWsBdNs
ovXsIl0NVYLFoyXn0x0bjYcOoGOEt0OU4IMJUmvnLDaTOqtuSbjWbGU70Bh7eh9HLKvlhqR+uw4b
e1u9+zz89xZG70uXr6KSVA/reID3VeJA1LKjBu+tqlRbn1mRVq1s/FVx7Bv5wyI4NBPTLQ+5YFmM
flrfw5d6EAK/laHv+XSOIyWgebkuz3AoIJYOYwC2FNNWvURU7DdFdDFX2EhfjSr1YBYF4pPKef0r
SLNhNQqGxflvZwsRzoJcuBwLpe9X7R9JbSXKXetLVLx258UwfjWezxu64szwbkM8kwik5GWsXRMl
U9OfbGJGy85RaDmgB8zdp/yqKalrHH7LtPZHhH06FlMUezPPR8w9YppCzjURRt07lGV27XQxNlFh
Wk3NBSB4taQ0bjHSZWSSR5nS7prL/NhsQWUhGsDEKCsey+aDnC8oFfBNq09yVIX4PQuHXve9HN7G
KYbVGU1jLQfcqn2xGIOD6w25EBRi8FEnL8N3Cmo9QWRXl/mM7cyMZGmgbJxKm2kYcIRqSKZPu3XE
dPENxoZH/0/YQcRRl7TAxRzpqIVehsNBXj3SL0ClRHv33THt3FrLAgC45LF7XYDdZSWbOpORZ7r+
JVHqVGAREsE2UgPEE6Or9V+cwo6vjxJK+e9l9heRfYvNgPUcSW5iwMIkatU+P4zwXfGMRBX9MceN
wXObAsGSBXdpgB416jLKnzqCR+b3zsINn8qVpXqT85o8EP3vZqdxeDtoqXiq7afOqS7Ta+9v1vOx
L0Dr44P3UZB1kjLV/MaDCwmAMfFd6FSZW39CMH8nZ52EeYMiVohaiLVDK2LPMpSsBnlr66xwjVyu
iA2E7YoAu1tOPeoUwqg01xpJpa8huZD7TjiZ0LdzaERX3Q1qOHnnfzjC71amFPt0xfmI3OrLNKux
KVGmNq1qX9YK4OE16EUFLIW8rZ0c8LPsAgVutuTUdg76ijPjSzeFWjO7BwBW++tpyY3X9bXwfjLc
unIiD4h48xs2KpsdNQy3CXgLFcDvuzIgpm681mEXyh2/9yk5HyS2u3Lo4UxyomJyeiFaYsMqw0Oo
chuYZlVbv7JVKK8RKywEi++YI6BvQcurzotUo4OiNZ+wjjpNNNvUchFvBeRCWs1noDbzrMmc7PC/
a5V7zHhiOWeZWhvvnL/i3ZXgFZwNdneGUdkxjhXDCLXF7penf96zqy5VE9UBdYWcFQ9buYUZJF2Y
UGFyXFtgwvY813LbkftsRNc44AF5Rm2qgPK5wwKAqY8yDcFLmvrbD/tEA+sVhwXXjGVv0hARUbcV
Sp7evHpLSIq8hbA4snK9R+btz5qa5nIhhu6DeW404lw7tNsw5+Prt7JVFVcNSiqY21QNITM/xrHs
aF0yysk6aep6XJK7XJ5a1BnvOqyAobaa5KpJEq+Yt90udSadm7JvxP85WfGNedjMtXbEqT9zYzDf
5FkKtcC6137ButPBnYroSgYUFmza+n3WjShmq85DqshbTIWL4V+P8cORgwHE5CnBgG6hPSyMrAlN
cT7dwFgCT6VEOhNJb56tTlYegbWvS1S/VXtT/yWrOFLUkwFmoKWf/5pJQh82Ps0vIDrGFnhwwWoD
BGDruMLq9g0V8cC08QxfNjPP4qJDkohlLMv7FiMW6VIJN629iOZ1jcMSWnTTKvYCy1QFFC00Wnw5
zyJkvgjFsQcf+4OJgy51uUJhZFr8w2+ve/FsobUZb7JzpqgX47ikE5RPDRdQz4jFSC/DtEPAMYYe
S1xXNez7haf6dYzaropzUJ17gCvqX+Mnyjy/ObIYO9lybHirOwMKfLZcG97XiGiGueT1JRlKQ+ae
C5Am0BWXRaldEj4fOxtd6SnmQcWsxfy8jJGvK/zgKK5gcgDVvYUj0LGvkmnKCXyhKIokyEv+V919
KE+L4E1NlrBxOSW3jaQUi4xomfglvbl9Aos+St/qiJy00feQVDNktfhTJPXf0SQijNtkw4UerYGI
Yd5mUZbnV5oA7oXeIzbyjCMEb19hCDhQrEOyFy8rNx2/uOpRH0bBNQS2j3M5WgSXhpAe9n6ZnQoF
WXYylNi5HTFGImd7u2BuHlRfbtb9QIz3ETG0ougBA2Em10xoSMaoFxktzxbdvo1hJAB5yrWENRHC
Aj5y1L4yhmlGut2b+RSKkLTAz0xtciOf011CovThdYCvQC0nwHI5sZJ8Ownd3yhAnWQSYFfFtBRP
UePtixSpCxEa+/BDaROeEY3Gw3b85UHY+NkYtSMcMn/YK6HYmrK4L4cHDN0BcPa2d8+XSqPt/ZsC
OinQ/FBOmi8ncgtqwJis/SJSKfwE5laR+TlJGVxcshs/cxAUdaY3bWMDaKDYiN75RiRxJLZkqvqx
kMbJ26IzTS1+Ps/ui9h8quImDX5YuyCk1am3CviDx71sytjKF5zgRv6WmpuSl1Lu9yyM7QGoWBzB
8sp3wBpEvm26J1rTgNOBFp4yyZOE1zAbPMePVjDDJsKPmlSqxzLeeEtnDWkOW2QjRf7HhNLRPe4z
soBhpmExiJbhLjFnlEqEKusFPL0ilDYOrSydlLgoyqDHckIO9ouH9/PnAp4hMau1d+F8hFaXQpjL
4sC/wDaiw+6NLo1j3uKPuPu/WcFalL3B+rOlO6ccAIBgEAyYYOOZ8BPHpp7ADlTYAq3p1kGVys/D
V7EACq0H6tbhnrZTbeCyobSymDqCxaK7hUaBlt20pruRc/699eeibZpuV+iWX3Dl5EssHGEdSX+t
jx37mogrD0WMYrhqIWk2yAMPBBrzgbPccFT9feSjZwDOfmdKMc3eAf34i4roasqcpW7mAzFY+Ejo
Ah+i3AFbJ4EKFPZPu1xL9bmWJGAs/xTnbW2/D2/0M0hAG4xCEnwCEZB7j2SNZlXyKl3s06iSds6B
nlpWjEZ4BvqoKZ+oCt3ZEWHqttrYsYV02IAGegM7xuhRiggeZ4EZcFwp1LT5BmOQJ869wubbbUt+
+slTXRpDR0QQI7LgPDB7knRAp1Y9RO11OUNRVjWyNtaJMlZzb3liaMg1c6fmiU3wXhEc/r9l1tsR
wpmNeOcqhg9tf5QJROfSfeGbducoLpc2IbD/UeRZ6GV6IIGF5qHDLmj4TobtFtsaQAb/5xsoUnXo
kJm2zSmJb4m6l0i4FMkkmhFtW8ac6K1sUJyom9wiEFY8SS/c5Yyeb+EK2rF3hSyRNyxcsjf5IogG
LaDSweS0kdS12+mRpMGHbdHEyDEEocUZsjyws352YHR4seL8H8a9r9d2EaqDSBign0GItK2fIEgS
9yLuTLCErNUaDJRs64RO+8ZIB4uZj0BCKzNTfzgtiTdQGsSzv9OmmjgcoyYG5bb7pbT6mSnvYHet
gEStBiMSzvubv4rqnQfmun/ErLUu11PPVKn3VWlXVUKyeitKj9aqMZNW6U8YSo1NT0zdrYqiEWN3
eZRS3M2PHjVvzLfjrvkKUmJbSHdStv176XhjIIhYUJsWwzU+sBT4tpuq+5zhfcpmdFi/WxMaq+Ce
4VzMpOxCrggHHoI1qGTS7U7UCPevYzpu6hutLByHYV50a1xj6glSJhqS5x/BYHlvl1aJvgGt0fIw
R/y18CDBi18ooHIt0Q4GVVLQ/A74FHRuFjy+vyI7wwAJxJsFxWk99f5kLfqJeBWQKPxbGqkS9irN
ZrbE4HW/1YXJc0hPzekIjQNJ6A016recJ2bDMD7EI6mGgj61o+xONSTjh6JorvePA1CehvWBxDWy
T6fnkX0MX3D583eG9i+2kDaUaxILLaOUi/wer6NMsyMiPxQdTCXnlHwdWURlao5IZ7DzHGzILsZm
h9TmKcAL1HuAmDRPKh4cWM0d9uV4VOeqgegL+ZNvvPSUuonWh5sXYPJx1i4LExIiiodjPjHlrL+L
2oJiNDzPA+Qf6XMQ9TO6YdV/vd8/5dmcMVgSGTiszj8tFtS2n7x+DRveYBF/QdZB1HsrRf4LV+yo
p4lHtPZiGd6cFJGOs+14Jf6ogySeimLN6MXo/o4L03HXDywbFm80i23YqPGWHwxkKeJ8fd8tQV/J
H21b2/64ynZN+qlzmqweD9jmHsI+ohJSgpbnp4Ke0gqGrYBtyq7QbG+WTn2D9eoi3Bm9E7yojGJ4
cj+Wm6DIWWJHRNuwTBxaPGCQcG20g7j7Bh4V947qmUuceYaTkjjMsERlUliiFKMpop9Hv+vrRgcz
zvC+z2VfS1fm8fdeCua+4AljEJ0yRZrAfyjBDTrZUEQF4HIt+M2WVWxIJNYqpfwSp16i6Axjb5SU
y1D4Iv8KwEn6MU5Dd3s7t7pTE0NgJVyyGbzEkBBCVnbN6/HTXt2Hq7xyDvYxPG+8q3lh+Igb7BUJ
blDLKADOjwRYAcARc2P42RlIxvAixtgj6IZzdqkDX6tBo8C00KFKvwx9o9iw1cY2nDOCPCryRVCE
X899h0PmMOBVRrARcnGfRN7SCzvUX8Ilu1zXIVzkJxs4IQVpOPD1hGfvRN5cUXtsi5f0fQYee7Ww
i05XmdHVgsBEBptXTJAcGRp0G5wd6ta5/cLJmot26sV8dFxwSskGE6ajPXnuU6Jjj4lB4EA+ktP1
XcarhmH6X8jMkRkwrJEYfDZMLhtOUsftwVzw+dXiOCQP0fx3Bqow1KSPrb6F0MYg6ZLztFgOvsZk
CpnTvZdfGttsww1//ikVUmYnhn2pPGzb7N0NJshaC+5ptIELEpH0/+YDr/4rVj+Xkew3XTlh1xa0
91JuCsnjtvMXb6//YoJWnRfmyG7qIv+6MG8fQChsGJllQBakxfWrK7SkDW0Dutfr89rml2lJaEpV
jPJEtpRCGH2aXR/MqMM/sBbsWVWLITkjL15Z5Hi3MBBsWm4rNAHb2l6GXJJVrQmgucBVWF+MBUS7
O8TlU7LGSZwYEz8FlrRBZ7LJi2DE6liQ9W3gwofi14yXr7L4TpP3M8mZM3NK6rFY7OHS4nMD2381
9f8FkEfQG5X8EbO/wGraSEBwpXDiNgmzI3UrL9IMdG5L6QcKIvkzv400ylA8/JE8uTrewke4/6JD
rTld68ju/g9VVl411tyXR0FTOxvPP7qS1RbJmR5Bsrzp4d5kRy/jrBzm9ORPbHKinySZ5/W2BXqN
hhf1JLirh9JWBNJumvJZpO8Sv4IKMHTR93/W295MFsWD7KUVeK2Tav58UaZGbCwStmonYFDaUMkv
uKFvWS5nzQRFqpH/LYOnn7Fxyt66IxMsvpa+DeFT4e2BoqNH7THcUM1eEv9Lhg+1cp0LtukEADqm
n3dJH9bBeB+fXxF9S3+zfRQj9RXwmtlbxzlsT1vw9CacIoNkvB1sh2Dr8hERoROxRHNfH6msgvEq
uBf879HpmWrBRVn9b49GQw5L/fHTmGyjHVmBF/DIdHt0Mda0T2nbP4JeGZKfFwDMJZh/RkUo4lOO
zr0d4xqd9kPCgBGFhb8w6x8banMC811i37w0sySDWomSQ4NESVkJ9oRFLCicFSje0zPNlX7TxHv3
j0cxQGFEj3ufVx+l3TO13LT3dawW41wz4vVfmm4qf49OFkAWI0zo1dmdf16QW6wzUzF0228giwuP
fc4tnYeR5C9W3LAcJ0iz9mi7uA4j0/ZL+6DwIEUo5AjYgDbYwG/JCIQpJymmVFykp36sz8BVpfNA
lxFXy72rqKJABNbPlYMc3eMaTnBuY/F700rfHRT6J3p9ETWo8eyComUop6pKgPmjBU3XuOzXPCvQ
9A4yl+Zd65RGggfeEAheYRQ4h4bpUy5IMb++oPHhNZAJUco9V9mXZZbaPgZTaqRJkrel6/WAPWfb
B/e/D9ieUxxsTd6RZqBdad3//x806hrN0/XK5Zo3PbazUqWxjn4AXgBeherLUuGYHUsIjR/l+AA7
74btqI/Z2mvOadaxztfDbegqyNniiVDOayMWyBikmjIEMCBZoV60DBKdnb+s1636iTKOrKY6aEx+
D3JbbQ46hBQhRoWyESmeoW5f+i7ff6u+daFd/o5lJAfD0ld6s2QP8LF21oifpwEAl8b/F2lWbBV5
c2Pvlcc9HAEoCBoMObmCe3Rx3j7LQXVV2KHqbSVyfR1RWQB8E6FTo4GdoHmABo/A59cOP6epFDzc
MSm5aPfBAZeaHhYQxZtOX779ZtwTOZDFGmj/IbFikgxMQULqEZYRd2dGOqeRR9ksV1I0Cm4pEmqk
gj4RugXqC0DGK5icYSA6zNN8TplG3wS4mwFOXwurUUuMZ4bId06qorpaKBgNul1UdYEuBptMtNB6
Q5q5r2EUcapylKlHVpcP3BxJMKhY9TrXOUKLk1xg7RDYk1HDC9OTevRTDvSRMKyDb0z0jtq4h9gj
YcyLe125VDkjvNxGZ1ZKWWEsKYN3nYuud6jea+Xn+iMJE3qOhRaXgRClrSDLExiDvh7t5Nu4cfX8
KxDN4jVFfqsGmdzR372Jr1r1kb+54+YPmf0yNvGVjUxfF98u3H9fl4p7/5utiddlcQV7eAp+gYvI
luT32aDeTd6qxaUNG88le1vKDMTEFz1e8Tu7ytU+3XMJMUu0ACzczkeuoBGwq9C7EtGrpwQ9KHYf
+MtXqiRiUnTGSPDqsSpV9fpIi7W3+2el+1XBTMH7Pzd5oNbwKM7ca0GHPSntRmMhMgIQpqdtzeJu
45IQxidlAErcHpw+BKDEVwKnEtrnI99o7f/T0eZ5bfGHDpl4mmKwVPXdI9ntZUgfB9IWH7hFQRXP
3MvMDXs3Q4d8x8bb6cNzqGVOzKDRn2/aKt9v1VMWuJ11qeDrW3eadlG7OJ21oQSWMktJNIMTIi5r
lHWHv5Scp5lbypfuwsR/cC4pQM8QpIweBZyY1mu0rMpyTf01J1RS2SyKv34qzY0D8gBnqH5+MnqV
bUUNFS0+k9wZFQeygIvPGQ2oFPsy6/4qPFvM4JuAJOwD3VpP1QNE+KPVHcO3eqYS8O8JcIzET1MF
yJMfq8Bm3WQwTRvSBjtw+x52WpjXbHKiIbDVN6fQ2uTiy25hmJOV3Njte6e+l/cpSUOke3hIV4Yi
mcDAeSYBpTkrHmcdcrecPKg+xfOrloUUAFfMVb40cJrJ8sOWZDdUBC3oMGqGsNwfauhGaaI9rbWy
Aor5Tt04Xsw4ezAsUz2ZIMoAhaqjlNNu1+lpeqxeBiurpeotJeHQ46WMNF6/vRgQHukk/tADXT8x
DbUJnxyubRv2AFhBxzn2Clv83aO3r4W5dQ4zIrhTCAEUyj/VVDiJxkXmWSr6x/b+0fJF1LGTBHCC
GGuRZWaPfUL3MXwlj/lQa/T9050nkJihNv84qoEN6BrbLvbpaJT6f/opfYWGp8IyyATMFKzPT96P
i7V7hb1SmTFt0z0ah8pj4Y4/U/gCZZvUCvhU7PK82FWuUtilIWJXESetv3xouyMxnUdE1ACxd3Mv
tfaqI7KD0ZzRk8mkaGQmEFQHY7poqJBFQbr+wolSDGSIER8EufjbQ+5jS2pwPU6N+H3HL5mMPTz1
yx6JIlyBA04ZEQ7stNvd/CDv4xz+Iv9gofcfFEfon+swYqfs4VIPpNTH5m9BM7HDEENjzdmCFDto
5zp+QmzG/3/R04tm8uof1yYXQi2+c8jL7SksxpDWOWNnMgkUyhaH77Fy4H+7ZNwsACu2cxBctNoH
BhTdyI0bOG0NK96VyntKAtWlysSYStJOruDxkbyjFxWPhqWCtugBxD48a0Uqed0DmSh8C4G3OEae
4UuuSrEKOdr0qlyUPp9+hs0aK56Aal/XvtSc10kpSA/FKHF6Hq0WI7XcV+kVf57Nk5U1Bt7ebHCN
CDMaOcoUFLfQ3vE72N6FjVPIiZsMmsQ7ElbMERicJmgTjNH6XEB7Be27BdEQmZRlm+Xfk7EN1uTn
VSwLV7mKrboc/o6MUZDOZBXjwrNe3N9tbhThkeJP0PXPhaR26YKMAmTSSBlQLDyQyJHTlCSjNzMM
AIIE7WSddSebMDl+qg7Ir5vMSIhmVAbdlXFZV0ADQAGpWWwPQk1XL1txaBM1xA4vHBHDepD932Nl
+NuZ6JugL04iir2YtXhcTJmAl/1HVv4Io+qRaUqByD/jdKQlSGj+aty81eNjJD2/eaydBNHKsvhm
yXOiPIDMq647jkgFgX/x7GwnwuCZdAn4nf7JpVENCvIdBbnLyNMBWhOIAPUtLuG25ho1q4gkcRXt
ErzI/7W2mufUz+M0G3LekMMQ/OP37+Ck8ENeRX+by0vXgeSI6TQc6QaGLkW/NLD5ZjyTujZiMUh8
P4n717WXrd2npygnoJFT/izy+2ET6GuN4hjqR722GjyMs9YRooO70KXZH7JpOKvffNWB+jwU8LWR
AlUNJxKhWT2WrFNbvMoO7s8uB0PW+09/Xm9UexuXJfKpgPBtcFdHL74OhzZMUr0lG+qnCavp6gg/
FAoxhOcNFrfvSdcZSnuuv3W6NSB2a55Cz1K47618/wBay6yuR6leIWdaUT3VtblPR+Mq7Vdn6puT
LK9qhzs/HIjONUn6uJRt+1euYI/Vg6LABI45FKiNT60PXHFdYX9IByNK6AAK7/g6EapfvvXB4TNj
d/xYgnqlbWfa5lh2c5bfUnxX9ntxtMvZ2/y0aJtprH5j1NA889wYg/f/QQ3PAMfreuvXF1bPj2D4
9YDEngJluRvrtwi/drsvd0mnSGnUE4KtL2v6GyRh0HwiTkcdKo3G8jGwQgXSEpfbphG0T4AP3poV
VE1xRbYJ3cpq9u8B6OZ2KNQzBxoMbZue0RIZRYuZIHQ4v2b4QLOlFuKLaV1nu0rxLrXTUGoVOEtI
DKY47peOxC2nRlaR7P34i2t0O70Y6KFSEw3u9owySy1KMa/J3csQrVCJRELjd5rYf3c6fIBU3YDI
LFW0xLuX0fKfHA2eaLWs/bp/nxK2x8NpEjeeO/9N3YPE7YiQPU5X2rMwFqNHJOXphEnxbKj5mOu5
FRsreYArK/DwB8lGLerNb+DjZ5d542RcIIelJcshF8b1R+isPP5AO+rPFBNdc21Iskt31a1E0nFS
DiJYp6Z5slxIXYJbBsRwNOC2uBX+H4X9EUeYEi6PMyYl78O6scdYwUDBttSl4aYL2m1oY5vNfLaz
aTcpigP4zKItjECnEuNb2ZKe1mT/xbh0n1cfYj+JmWCjlvF1JQWefEr3zyXhwomMPxtoxe6+aWRt
VZSQn3kH6bHeTwBib0KQ1aYx2DbUE7zsVy9zwn0BiGT2dckArxOgpkKMwKE7QnX/fF14M92AT7qE
3V4sXJSQ++/W2Iyb8C4AWoOrKftlrHkobFR4NbrkFrNVLkapD1StRaHyvSG5ATQNXAO4Hyh2ufZp
PxYp8YtGJQrEKZhR2ZItiGahCuKW+pR4Oa7AukXUGZEDK0/+c7ZmVHVYWcsigt5eoxVlHNJ8S8Ue
0sLsYXOq6XBQdNT/4pCbHQmBahOfvOL4RTZ9s7OnHa+6Tip7JIl7d1v+MBaw/LLKLZa6/daujnT6
Q4fDGQyjL4cOBMcOAZOF49fQ05LA2CyLXnXTWYIHIjkaMkeMcluPetdecwRYwFoc0LIeg+b0A63h
F5O2EqoNR5p5RR49Zx+WlKA6QQF19bUbjh/clPUIp66GBS370g+g9DBxrvAvEYgcCiPH3nsSZmpC
cJOsLtjGgnfVrF4mecq5oZLaAWBYb2FLh1vHJ5OH+6RsK5zalHK9YNi7rQLQTDewE883ZpmItvMJ
KDL6m8bDsFjfgVDwvaUlV3E9rEtxhYYsLqVh6EFEtkTITGwY5cXR5FOxfD6/xSIh5ZW7ekWaBUPe
9oiYf8TCjVm6xZcL43Kl7+ocpVOpXj+vf3GIVlLVCKMTr6SLaz+X8N7v+xserE1sc6AzxF6Os90c
ohRW4mYrBD3FVMCaioM9Hw/nPjrBDVvAD/YkuqVzzkK7UFLttZEJorVeidEqlJiNpVC1aE50k8t/
BLehGaEXphwQeCqGfN9da8mafHMMMHFPBoeLXUuAKMyq+mG8JGT/1fQ7A4sSNIwd4P3MaYC4v38W
Tj/i9B+H9+E38xz+tvz3B1+gpADxiNGqItINWTzbzKTaAwZTAbTzTeFCG39rC3ueq70KOYi3Dndn
vAdwHzUAbfGAl/nl0e9bQv0L29O8wiEaLa/5gA+if6sNwOkN1MJmZuc9ikKYrzbWdaSlgVliTYjr
dfhb/+8J7RrwFcJRf/03jtb9pHQzML3Zmvd2eOVnrrOws00/v9AiiGJjuGLyplvJOqmiZ7jY2tE0
WqNSyqnpMgW9kYvpL8fcR5JfIItlmXeURfS1lwoQ5HNKAEdPbxOGBMTg7oBgHRPHQl0VB4RoOxtC
hlf0YV2D0pgrzVFoEOsEb9r8PmUBvIT2sVMViYzX/lK1rfo3YnSMpKHdCMQJxXR8iU2kqvqPYiyH
+1ewz9i0YSrCeKtREQRjmcnpF3ru1drqtGNwKJAt70kwwBUr0igNXX645OugCoH4TU/KoOcXgY3X
zVar4eE8pUlWQyQ3TpL12uSLiTbMLtMsVQLeh+SU73G26r2WEPyAA/Y5TDd5dyLYlSCHHKgifZi5
WmLaAbFKq0rYzvjZIAg9ifa3yEgplrJIbAfuzntBdp7Ds/LzNYyeJi3LeUtbGO1vtIr6vlLIAWBE
TR1yIoH4Fs5EVQbL90/Pg0bIVKZnOeDhCLFDnc1hy9AExhUhHAPmc2tCs+cwUIwS0SBCNW0aBmIy
5KB0UZhCuPELwgLWVvuZJIgBMXtiHyv73SWdmWYzr+9fnGwkS52Ve0J4ypSBa1SyYbI4Ltn+q3hd
e6djdhfoXulsnLnRAwaFzEFWfyOLkuiVew+Hy13wyGhQqqoRE60dQKt7NDG/U8ZePCrEz/kkwshz
xYyKlpM2Oi7qbO4Ks9+B5ZxTEmGjCYnXUSiDY/OH/0BerHZYJa/iWHL5GykC8BvEwA6TWSic2ged
hVLhFAmZNA6MwW21g0SD8YALl6JnV44AhCqMWbdfNs2/8/Rr+GUZ/5mXVrvArxcd9G3MJcccoxpC
CQE5WmrEmrdvtLfaXsBxl+HzP5EoLpNUcFBYp5MJqL4rT5KuKJY/ESlmFy99XAkuiIaVdn25oJdm
aF6ainqnL/egZAPwE1jtUgZSUEV7woPQbHRiqh6sRPHYxpSl3HXGCJqusj7cW8upxiMF5vQ7TOj/
yceHeV7IwMRtavD8VpJr/fWFUfbqK9UeOKFvc52b7/iiINUwvfbLTBjd4uXg3DP0uB/ZmWLDuhav
yHXt/aT6kthHDtJTSCOka76XO4HAnerOEflFqiIMdalDAqFT606IoQOkstolljuG7kLJtjA8qY29
XmlGAyGrVFO+bWE+L/7OOj6N/seRp3Vdg+y+LS4G58oNusEZHDJe1feKqvlufu3yZh9oUTnivPZR
5hCRODOFz2+apIIZybp+K6IaPbf+8WbVIMkZkd3sVYJ/ASlMp6PUXCggGg4y8lIkWr5Q9wqnSFmB
FP1+2saN1wz/gZB4qujj5z3auOlTzMQJJQ/XV/ErOd9jcT8RBqtVSz8dgK0iJanPxxWACyAnzMTt
awhD0awJv48RjJyOS8/Wb73rifR0HCkLgUeYJkdQf5iZKLh6LM835XuwlHCkmUwEjDhK7sAJpOeF
bviCIKRr1HLOJwDXBJ8l6wuAMEtDQ3lfefghVI4YqUWpV0PaJK1r0793xGPk2C1wk+mRe4hl4Td0
i78wu3b6wKq14+SKwDs3+cJvanr3968IYBLtWk8X+KBAyBq5k67+kN11/4aD+XMoFzlBmI/KWVWO
gvNJAE/NllVF0zoc6ZXpiIGCFQRl5jeuJKIMeY7LlnPKwzqzioOqkixZ9XMLZLkhVENDOaduLyJn
5ipA9DjbeCuj98vZnzbs6UyXkewqLjoZETC07tGn9BXFqIBxhTZswlt3N44CWhnQunbLnfyVCw9r
3WtiAYOiqEzxv9jQHz56BKP4L9Rdxq40aKRuGbCXB+lclHCjc0DEDg4NtUK8nyq6UF3gT4EWRWOa
1+5/LtruRTeCsTz+kFiHLthKGIm6Ygzdkjxf7XfVsBkUwLuTgOcvBdgKYCfaMF+tgxHwWUvndNkc
sTBa8Wtp4axhYJJpiyEMlofiB2zinQtszuHPc2nxqbBZHEFHeg1xUWLU1fUMkaAHX2vhAgL8gV+D
r7Q6hB+itslJGgsyHoj463HNVJzg7o+hbT4PpPRgGS73XyKm+vO9LsRuQbPiOUqt5qFAF+atnMvP
0zYYw56P3Fszwzbm3V8zZ7yz0EzlO0W8SYo57eBKpEjb9PSN+2x0d0PhUbFBJeBZYWDUOL5x/AnO
mFXRVJpg8iiYxJbAxwW93edj3LN6bIXKewxbk1ZU+ZYS5gyd92wxD+yMvW8BdBFuPUgh5NFDl7QF
SoZrqUbH5JDf2jdrzJDe4jMI/znP88bb5W7QdfuiCXSuaDoP3b0YsH7lBo9uxQ3m75IxcHB3wY7h
7h/VIqFMKP6t11SzJ4wQKVvuS0a1FStvpPaql27PnafvO8qt95k6VcuGCO/8AhiTAbPRXEXVY7lt
Q4ijzLoDujrS+DvMXcUVVnwgQC5oV4T8jIiBhrBeHWWo7jUtYRL/Mj1iG+QyPqWd+S1de+8yR6YA
XjYKk/cEHdM1kvjryftncN3tfCLCspEoYUyeM6Pp8CPGJYMffgY9dQmtUkkdbGv1e2wUSRoYBxKT
jiqbOj3U7Izlp/E2yuRjnmkeTdWpJhiNT17YEo6Aid7CJBHxf2+f1JW8lXQobbYLsjnn3bdbkgWp
psKnqPu92tNYR3SgfWtRY82ZjT0FVKKDTME5ViuXdTkBKiFJLEnAag8vy8pYblBXp+86+tyPQe+A
a/idIOx+13pkvTpmfLsXZ27l/Wn14dKQAeTfkJhXuC/02M4Odb6CKvOkjEXlzjxa1/4jcX/7hmjT
Ri/MOXFIBxwzoIQ/iggwIuZLVNHBBd/81PGLWOCfZnNzM3OiLlKd/ojrXQ7PCr4Qz+TE8GsERi99
0ZSGx0M9IJVxrGGEfzbEk806PZEe7Dyhkl3Piz+ssKI9NwJKiLGhYsYciFJlALVoMxCJcAI36JhE
dDk1Tf8WBA5igWrSccqCICxnPeLme/OoEd2gkHkevQqNyDrhhMZIfa5yZh0SUlAvhM63L3VD6RYV
uGbiiDsXAmriZnK755G7i+tBSFDZ3/gexco0gc3Sgp6NeZB3m82kIIvxM1HuzgESXxDYMWPghj4a
pxa0QDSX3Z2g+cC6mccLtOd+NyygpWNL2ZliT3i1g69OxGh3AXKi38KluX6tHTcvfIVVsGDsso+C
FYGYXi93qtguiJfNew3r8gvSxVFSUXeviDI75a2BS15xsrRXVFZxx719tPZ6BqTN4Wc8LWlN/avB
jclXPU01eag6XNxayM8sBJN0s6x9zj1/PR1nFO/I1vYYvG0Xj0pf5ogDZgGEqLNNawDE1MNbJW2M
f0p8UUUx3ia6+h8kjAGNoAs/Ab+r1KDPYl2gmDkQvigQUJAZsByl/vV2ZeHyA3Dw3d0RMAG0e9B6
/oSP2UclWyiHYQHng49fDHIJgnpnzA1KaeNMoCYpIXVVbpxPpqNTL1QUblzVUs9SNjWF7+Lgal4o
Q9+wl4YQR7iGS4EgWLgU49JLr6LGuOvnZBJe8kTbJYwSnLrDFCZfcJPsfDVTL/SsY4Q7LROiBD0t
whZAqwH4/YeXcNjGZbxWcxiwXq4AhL5G+tTwnYzaZCMNFC1ovlvNC7eZtz6uzukax7zrQfCWjb+y
2tBDYj26EnHmImPRIFKVVIlj59F9xDqAYQE5D4PiLE1SB8CKOSAhkSu42UKNm6Uq8Yxlo0a3uezd
DL/dUTAM5Iw6TOKi9UpXxKGO4tZnQc2ZpDSnniDJx0tDJhXejYp7EDaPHp+QxOrJSRJX49r+bOdb
aRtTmufaVgqz9AzgDxmHGSUZk7V+uJwV1Yu578mIVTBXFbqXP7Olez5gV7Q9PRw5qlMgbeeJLi17
k6vDyRTmt6Fzh+Jglan8fGKDmsC+WsWOP1Mr7KY3oqgXpPMLnwB7vO1AFc7Fu6GYicWHsn+xK8mS
8sjO8sgXq6lSSXStjIu+2OYuTfYVc8l9EfzA0skdmvyBiJalu5XwFfJm7R8CrGgegqeJB3hvYuW7
Qcg9/olVeG8aaCbzww4I4iUzFMoohZ3wXzzTiu4rbgJzJkYzN4dzIcYYcXSsR/xyiySbd0XGUdPZ
xJjXHQ2NKQ/zJbLxgEz3FbqT/OMMIBPSQNmCcVKjY6FX36ja2Qtwbpv2ZDFcvL6QIJjhfLdagZpt
pQVKlRj+7bnfLiugEzF7WK0jNMip3LtiMjI5NSoOL8KPoJajPLNB3hrtsnMKPYOhFoCvuagxyxxo
oOJerzeW6+xN0fT0KfHfLbiEywl6cUEuaFm7mcYvPujWyNjV7DebJURXWWkZV6Vosu6eI8vhNlAE
Xf0B2gb2PnlrqrxRrAc44kMyAUtYUPWXIo/6JsIZPSam5pzKrISA+xvHo6Yr29NkOYk5V92eV+et
6BMuFQ/jc/uEWZWFcKelVafGVlH7j08/z4qV88t1dGsrXE6NxOEfjYYUaAGO/BZltzPpz5cLUgV2
Y6nT1q62XJdFAdXsMQEhoDtuM3rnHKSwOVVqhuPkOpwa/1DPM0KRCounBs//TwA2jcLyksznTkBn
XuroVWp/NutjpcWvQ5yALNj1HFXQYakWFtoIkABdvWr1e+ovs4+JXaHRxW59RFn8qbIALTM69/B3
J6nqGBFpmfqp3SWrpxbRtoG4D1VE/kI7Xz81Mmj8ElbJq0JuhC9UvuVar3cDhmpnedi3HUZ0IkcX
4wR41QUgn2509D6AzyMQnL7IXlrEMANWF4nSunAgiJcYXDfHxNhYhfcsz4h6ZHTdnbZx7szr/NlL
HtD7oIPE/JAnBaebV4rq79WTJkOKPy2qF28ii/GyBty4doT6CLG4ySoWaA5lYuVrN8qbrywFpeGc
mem4bbZfZfe5+l03lz+Gl218LwINJ3+8q7iFa8aMhHhV2gm2n1++XLvLFF5qWUwnTJ+0mRBR4kNq
P9in3vkXwwsAATfvIR2v6Oh2FCHWAcT+wQqApS23Lhxf6mOoxyyY9MnFb9G80A+9Uau8rftbJbTD
D3hGrJmqpNCoNdv7ucqbWkkBOiZKnMxTqK3N2aDIoiisS02xi6F9tQZm1dNtTfWfwfQnFK7f6xYD
pIMwrW6Rv1DsqJidp7aUqqWYGviGBuDrxh7JAirDpYhktyp05aFBpQAChAhPi0GNlX+PgJANXyua
Y+rnabxYDv/uGmgyGm0Ycg9OwyOsdKfrON6j4SapnQM119e/qd4Fjo9qYcl5ilFfxxV0YXgeOpQS
uJ6s3J9nqbL1TYbaUZskm/z1WM+ijNh8ZUTDHM+aSRMLyYIdNvpkztAYJ9YZZ9AbyxohNL5IwRt8
YbvR81iEMXXqYvRt7QeIiCdhP94scBKowEDM+n8UIOHQ/TtaoGmBHSndk7QbbXdjfN+Fh/CuyU/w
aVyGmBRY+hF/+gURzbrtaxsJNa9e28T+zIzlv6rsQTFpOZdc45bg3NXQapIPIjiQQKexcd6+Iq/Q
4u8HzgiK784jFeJ1blYsyKqMDyILCsDIREhpYvEzl0KYp1ZfvVChCXCzmLa/MrRyl4aXWklFUEGM
+uBYYC0dyQLVskG2pTXJkB27mIPC5dRGumswIfANTy4j8kImAe5lqarZIK1RZiJeUmV1DuPJwcL/
sl7OjjqunkPwuJIwWcYCC+fRrYkTH1CG7PdTTGtq04K+Xy/ZgdO1LVI9dEpaTY1OnFkRH/y76PIK
2FNDJvW4D3KmGVnqqSt1I9sOi2LnOMKIegmupYXXXYBNR2xdpMk4Js0jn0TIRxOLPZGa+LOJT5nj
z7stgCT//9RfVHMoFVWInLE93cmi4hEhUkJtnKuSfljCNIX+yEfsDCb7APupVq58nskhM9ZMrK6+
aOvz8OXCOus7F9n6DuEmdlCkj4JF3eAJxIODjO6LUuKRydQTp0DEnJrg1PdvCWf4KBD9bJhgZ2/w
MCIgsRHgG3F6Xk3Bsayzb8nX2fZYVjNmK25Ygn4zArAKNJbXhYExYpMHH5dfQ6P1dlSAuEMZWsGJ
8lBGkrcxj2V4rGU5aV9TFhctFcTLm6rbdIZuPfrzE+QepCPTAaM/QajbeMDt8bQlKdBc3v5l+Qlg
JtNsooxvp9ieJcyaE6EUlvR0euwe2NL9+WJJFidu0zxjfDOGZMm+PHt1WiYcal/C+5pdq7l+lyG8
08Jr+uF0Ef4wmVLYgecQD7kpIZOA0h741Zy1dXTUFKwdxmGPKMCkdouM+A9xggZnkC7RpxTd5+kn
opYw329XtMlG+9rmM0rDa15Lq1udo3RDcuFSN7/9G0XO7hqFO4of5b2/HD5q2172KfFMbbkCdUqu
K4nlbms/6YFVonXadTBf6bSXotDq7T6GCFKqR+/aVyCadwp8g2SKvdJTxnXHwRSEbpB0lTAHwDzV
ys4adOniEHzThLyiTnzdglAYHOcjp2JKqLz//5sEZvXgyvaspPI7aAvSNVpDEu87OasaU4/Ut9G2
ludFsVqjHieUpqoIVdQQGKXu3ZZKbz2AOEKXzijJ2FjUTvxNWx26awoWui5COunl2x2Tl4/ET3Q1
aFXaeGHTtXLc4rqZelnSmNLC6PBhSTX9MQOTWuEO+GN5YeRNnY0GbqMoL1nSWPAXTUbZTZK6cmv/
XIEbKMm4BKJ7T6Xu57KJvTm4RBCjJjO1EFtQl5rvPsFfeSsRVhzZxus/vc6o1Nt+5auWWeA1BTj1
gM1ZxplQeuzB5A0zQMyijWTOpENCGDrBTHp6ZoGOiKXLh0bhGnmLHvVMsgMOa7zXc7/S1hMn7uzp
k8BipeMRRo62BDaVM3/3D85Y53kQsuIrbHsBOFMVvM3au2w6fuX7eGnVQkAWITv7mbA+eXM/mWsI
fLakZ1VD+igRj1kCBD19mxKWR5UxBswFMJ9s+thc+UAILJD4rUrJ14FYAQtsoqRfDpTycIAyoZ2e
U3j8RGCZYBVou/C3uTzSFjG9oySSztZ80A0kpB9z6yFkALbHzhDUrOTo0ACtLpz7QXyRx7+qJMat
r/RF846ipXmAayAGgISZxDVeDH3PMe1QFz5c5g+91jMCUS4xzj3nqci0dw3Gxb9Jxg4wnxp6g8eN
hz2/rLy5UaQu4pm2Xks/Lgzn9WbowcKQSk5TJ8xZVsvKDQ1wnmQBAgfuRTUOgqIn+dSpvnGMRJCi
/Uag03MIGEM5U3l+1UXmurZa8gmlRuVOpfCIzIPuuxtfhTj0QThJaoC3PMVCBG6CtMQLdz47DIXB
zCLzdopOVGL/PNPDRfvhOUFG+ausTrAtDgPVVqqMRhRl6JsAAoHM0WSi5GhXttZ+NVAHROn1nMKv
cOA7QXdJ6JNrWi1nj/Z/e531kHjYsZXTh2AoTMkahoVwFMrU0FmhGWJUhkrmFKuUiEDBqv49a7C8
vIJuoZWzjowtjYTVHa3OGLuE+503HiKiv0WCcOG7vunbynxQn2EqzO6frEsbAoIicai0Rd2OIHp+
wT+aN9ITiBGGsI+ptzVog9+spfHZ97J6nEM381CYRh4C1cBscm8ieXzOvRprTp+zokwa9ntZbQIY
1ZQFpc6xrZkXGWbPFX9BYtIcTPxs59ssClob29tIZX5QnUgGUo4nHK0mFJsZX12/aCr9p2Sk6ytI
DEq0wKEjoPaq1PI4p6EKZFfgIOkiB2PjhMIrwtlXET3nT2w+B7l3nv3w2hYJglyqqg7SLeiIwwkh
YDWxTJ7kQmHrVraWYjIXgAE3l9+PANIT8gqMNOjDDDJcCL9CuZadpIouZVYC/lEGpFdSMOK4XMk6
VdCy3AqT+/5xIPJwC+/oC8BT4dZ/ZAfK396546eNrFO+ZcQpjOYT80FAkdQl7RuVGiN7qLaICpbo
0iDj24XYgf5OnTINXBar9lsQnan9Fnlr72F1X8nRkW9IUlE6K9kJPUduaW9giD+It6cKdC3g1Qqu
BjiakgZuvxZEXx4cQabHgtj7VeiEF+EoTEGMFQaj/zlFSTuSlzbc+Quk+FxAmz83tVGatpQQ0ODW
8ga1sCpt5+XikubkjomdX9X8qJ0MVDe6CiI0JJJ7rSkr+KrxlBdS8KS6phN36Cp6/Aq+S1bgcSVR
CCJ3Xrnw/r+xrZ4hmyMVl9MGIeVmulHrxt5QiIrDV6OR9lnftOfHJeO5Q8xG3i/L8SuRw0xp0S6u
EdUl74M3ynAlBmXRSJzXiFwX4oj7OHFBWgq18ivDfr4fEUD1MQ7oLD7P4IZr37yPp1qXuiy3+wLD
xUtwWS/DUPk28iA2IufiNNZwfx8ZrGQizo73RTKwok1FVRi0qae4XXebrIZGukuHmEgQaBTGm/EB
9nlHkhijbIBQqykM/B6vPX17/jALHIxBaiz78p78LsZKJN5YJRK24z+VZEq6KblftWI9zMi/yTHv
MQdAxz2wFx7i9UW59Tp8pjm1zwr9uZ24SjDK0TGFIkQAbL5SfXbFDjoTT5esYP/3KqdrvJKYsd5h
RNWNxJeG8yXlw0f2IjnVyVzCuUWswpjT82RmU6KNJAVcSM/N0Q+zr4jxiXSwaNDaaoD22myF3MgY
PxMs6INhfeS7Nc1mN5w4Ov8aVopbR3e5POKeMGaDAkAEwBPeBoE2m/nTianEdKHM/4TzqZeOreIl
l9sPsnUVx79QI7jCPwGXZmQqDHlUp9HkrTEfE9a2wdeA37jQFxwvIGM14bH+Hq2YOWofJ9RdCW74
9i0yGui9l3XhprDSlytW3xn4GRiNIeM+HpOif5qilRBgArGVurR/mV9TK5FIAhzkHmIeCaZOLJof
PlPNa9kUt2ch+w9+k+dbSnzQHuGuJ5B66qqi+bj/VZcHZ5qwoclX5xxM01ffCtHPO8gyXE/QkRYb
Y8jRa1rS0kMKUPJOnHBwuJR7j+iCxgYRX0Eiyuvt5ccczx0tFK146zYudN/V7mkB4dDrUOSDoKXB
P40XEEJzbcRSukNj+PGccXpAfYpCxG+aUCuPc2/RrEGICwrvX7ow4DbFo9jtbLPVYd1zTB7UWJ6t
s1O9yUNtn6O8LstHS1dNghbQncE0iCIbqqZQFepkbhs/tmGAT+KA/LMWGYlsJ7CU6kHOMBE8xx4N
LHk9M66q0wSIXZubW+6N8yC06hAFn9GNw0MFau9qyCAAivTMyxsgZpbIrYjLxvNgLLlRi8raDdPu
S+RThRI2BrA5sWWQeiX/l03/kskYEPj9ehGWEjyDyr4N5V3ztKpYTjARqzNWeMpvjqkH9VogzyrV
AaiY9vGE+srFEmBsT0Kh3WL6sY0zB3Su3AJvW030pgaCp1+zTF8fCNjZrJj/ARdrK5iKC6B6Mhzd
+XnGKog4u9A/JuQJcKY9B4vU0NTCQh2Hxl159qaTeDPiZC7MYAzPbTqUEVOQkLCsM4GfXFJZhkPZ
x3DLTWiCG2tiV+T1Ts1hTNp824Muna3NkPU+Xr6bw8gJVKMRO3PYjfZgV7pd0sbZ7RauO5PHADyT
f09c824WezO+Si8wsTVg5ULwX5Iw2U3u6cl2ywPkC6TZ6o/R/3fvst4wMRFSkzgwOpFlujTDFgqk
Nq0uVzSHyEh8+DOUonO3ycfIs6cw0NTeo89g0FsQGvKW5D7iG9hwzt5ym1qf1WliT1Klu+e+7hxo
G1lIrw/Ii1eZK1L+v2tG2UagJu2e7VUGSchD8lHuhTHSsN7YwMN5OwxPPjecCk0GcVPKA4mIFgvm
HSrcYNDVdR38ZBdwdD7+U1/E9FT1g16D8Y12mBUjJECw022OAa1kznEjq7h4BhRoq7lyokXN8c95
xkgBX7tU9wNWbNWaUtUBAPUNfOChqOCdkz/dOVDjZIprUhZBxKmuOnZd08sW5nEinK2CpmV/XxMI
5gDdP6Iy7L9raC3JH12P8luHD25xfzZNzBDScz6Fc9YMbHUQDjoVHwXrV7yWoTT7jHdX61W1oZVU
met7wIrnT14ObjwhgkGlY7f4YzzUl5jKv7Ji1oSR0wEqb1LIf3XvsFfZMvtNjvN2LqCRoyyhiIYQ
6d/ghSK7gc/CXXLoEqwXH9O39Fss06mCwaOZnjXFfJfpa6S5CTAZyl2qi5ggzuSw2m1vbXRaR/0D
LrIVjb2Jt6l11sHw4k0Un9zeOxPPvehUHtB6brqkxGhPkEKaaoG1W3JP49vnk1Asc0mRaCo+4vVj
ceKSFxfFtteQcXlvi5CMtS70PPKyXPOgUlXNFOTMqzTXgAI2IqWOTOGnMaMksF1lZCqOtdqg6cGa
aTBZ2tJ3HDwQLHZ5p/dYqPr5VQVWcL1vIceVvwJ6uFungXphIphcnbWUDpGL41wb5kKafsajgwb4
w3rYoadwjHHfXc1jH64cxJKz5EX5lVyZ6y19VnBo60tjWC/Qn6nqpO4g4/jMo4v8j5+NhRhYJ762
hhZ7eLk5jThGLgZSbSFZgZhL2kdfjKcXQijdH5TBi7ZJtFu/mIN15Mjyq3I72tA+zzvr5ioOsLv2
Lb4Bmb0GbZBAg/S5Fqb3bDZj3NsWhnQ1EVZTBMPTFoC8svrEIbcCePlz9uNGNgENSJo1ho0ZnEO4
zX0iKUuaY8WU/I10U38h/0KfHSStNZBpGqjYs/aSqqQm4APFwKJtxLqd+hXi/sbtqrmXXRcwCNOA
1RrB8vkY1PePr6odFwG4BEGK87LezfjlL6xvY3aEPPCXfLH/kJxO6Q5AsBXz2gX0BVgUWyzPD2pb
fUogSsMeCVg9576i2Jc9Laq9/tUoBNltGB71kwXJAqAjXdIB7Vh5kiaxTblv/DHrZ/gAegYrQ6ER
AhJZYwW3B5wDqgXhExUAumtbQWEVyiVW5AQt9MuLp0NkKjyQA6SCxBKhUFYedELqxOmXog3h8sRE
VK7b4gGnWSzlJt472BGHznEPiE7iltQq2RWz7FhIezLlAUIZkzmjhbboThTWkrXcPe2MIKqluOV/
InLx5XXEi+S+PXtpeNKX/UPQJkBRUshwCHwKJhf7qonY4cFUWgLCyj5m63oV5ls9s3KmfVoVGkka
ZmVUXf7TnB4MK7rPlyt6Of5khB5GVHc2V1Ldti8wFjrftUdbKL8nsj0g8HAVSmGYuDWmX6hJxiVD
D/vasA2JNPidpbNU7W8uOeFW3u/EVcvUVjaRyw5s+Cpro7AVEjtw5Gkg/X901KnteP/qi65ylYJw
aFfLQcg2+Qf+iRwsgIwKiQObeVSKssFDMFLn4VetBJ6mog+8INv7NtbWcSBJRsF9dJ1Sgzz4/1eh
Ke31h9sYBijSzHv/FbjzCEyF0WP37Yqc6fE2opfbT8vGJ904Z3GAPQyH+w6QDRUFwXXU0gbgLWf+
PcpcPLr21jSLkFZWZswgKQKQwiuw8x/EFDhvPj/KXATPDJq0YwCqbGHj4Vcgt0BJEPo4XrDUy3PB
6Eh5Ep1Ig468/77pdgs2ksSQPaaV/8KahKM/dhaklqfuz7f19icS1woaqhofrCif1NSXoWgDbZoK
toH7GbO7S751Xim24pk0F+4UHRWykoXqrE3dq9PgQi64G4GZvzqUWkPjCRERrPY25m52xzr4H6r7
S9/+Rx0pIFn6LFUyjtRIbH/QVAIkqpuvAqmmRvzi3Jom6R8UCaNsv9zbsoGsvSLfPIl9sGQCijlq
BjmqYb1XSE2qX481NR9pd56frHzA87TTZBwemRBUIXJy2BtvYU/V5DI3C6nUcEabx+k38W7eOP1V
RXKd3Wdf9I4TeF1xaCcgoyvAxmRs6dcGOSR2RnKKy4Hu6d7Vej4J412vPjpQutxwo1iCi+rlTe0m
CIT2xBngaiAXtm/ofmlS4J5fxISFUnHCKgr1XQpMDIsRaBAOdqBuO+Jhjg6/k+J1oRCsJm/XzlxB
5T33QjHDAWNg+VUjFn3eLprnkIfQcqCSJuPfkutZyuSAw+k5ZpcvZpr5guHD3zXf7Yc7yoL1WkPG
16eLuhCt20cgfolCyMViIybJC0hZLZajZfy26yV2DxVtoMUDCrnKpuKr1sPxOjJnnqb3K1s7u0pc
SQCqDvsCsDtqfnSm1afwGESh6FX8cCHrTk3C0VmV/hainCyX5C2uo/idTwuw/baQKBMWee+PYj17
lCixMLW68wsgUZSq3ptOPrrEFsj6ro6MNJEA+7DFkhgzQMMBoRzNcK7yZsSai0KichKuYSFnBFFo
GCH1sq4gT+PMLI4h+Ry/dgOdd/UYRJWOA2qN4+4aomEEcnMAgBBy29ZHCK8980KrA5oqAeMmMfni
b9QFBJyfXB6+sxGPp1ixzuyXlvAeo0WmtvjUBKxSW2POq/KiBkgf6g71ORXdt/LhYkYni/T3fmfd
q/rmvsM/iI18s3AjewEXTtthMPSFEwyw2YVM/KreJpqn+X8D1/0S1USHFTQ2J6jxD2ox6fLreag2
FY00eIeYdeF8P796cmDD+gavbuxnE+oGjvAWS+v3a/4uA1qWJ/wwhgr5n5/4oxVO8tx7cuZpEaXo
e/IZJVWzv+Sylczc66Il78jTDJypAnOoTzh6X6fiC+aLLJv8DfB35dKwg18sKfGKy8en7RIiXLiT
pWwhqSElzDhC6JdvJiS2vlHEsdPpFF11OHcRs39xNLiz7DRo/JbLRgoQiLlAETEABBDPtwsbgFh5
1kcCpBiG5Xmah7gL1X937N0UkoBXfuzHKh75jyBIYo8dEVbZvgXNQvAYzn35rTmh1o41hiCK4zC/
g513TWsdM8uicYbX/lavZPqdiuwP30sS/TjAlBPuIqrpKMY8rvZQzBgahZKb06l3BBnNvidW9eOh
9PY97I8AZuQYQPtb+OUM3v1NKvNtrtiBIBuhA3kcJ55N/ni5ZmIqwL2mkUZa9bboWPs67rvQxWFW
99jGP7pnTRQtqqiYddGiTX+lXp5ae95snszvTuldZQovMyELmY5BtYIZzCpbtISMVyA2zmhIE4Aw
NudXqBWsMSqXID0JqCnahn9z+IeAjJqSmogjWzZHOEsN5BnHarwTBFnHRcbpfHYu5WrHpfJTqPaQ
6wRYcsSCjFM5VPExhMnt92dNXf9F0WI1RJd1PjeUqP8NzAIvWJXxZ5ZO6tBPbcLDpQm98opVxr98
YctLi+saDIGwI/bmogUWLtIj6Vnvc55f+9h8RLmCTqUm5VIMRcTqftjlKgi2KJdulNVyj1Ey7t2Q
fucgt7T5g8daTmP4x+osSWchYRlvimLrfTYEim3WekLHue87xihY5W+eSPH+NcM3Mi+5EaWG/6zf
B+dw5yiIUr7s2aFH74hx6dH4R+ikmhSSHy/b2BIz2RaQgzdu6106US0irI7vvk0OLi36dYSv167p
yRsnbi98m6n0F9YD7yR3srFpaH8JQffypDrfliweg0NuGETUgZWikkAgAfQglQQ+L5ShiuVPr6g3
jtkBpjLzN9ywsg5mNo24Pvl5nyGmZVL/PEVmKOovXVVJFMH2ifJfxNKq2yjAlOQBTzKjKW26VspU
UlBim6ANehNLMQCof3Nni2mflVAkEwK8Lqkqj7Bbldj182jx9XxV8QIL08pPtXcQsdGPxF105yBG
og4aoxjyNQLTg2MTA6mT0CmlOgcfPGpweLzBCnflTE6d5P0aBqaAbg6sb8WBHtclxKa4AztFmvsu
McpRmXdOGMpM5uH5jhFLVDMLArzSr8J/jkQkM7JgkQ/Z92yj74NrgYvKesFEvYFBpS1wpXSt6Shn
+c7mZJ6KE/w0lPnhEzljNuUs5Mysj/OVreF1xqWZrCcHA6aH6JszIiqW9ESybebWLqTjxj7ilz4s
kcUd8WJCkiffMP3I506sfNiEXDyS5nFORnzBDTKlyDR/Roxy7ZKK+6zUHxvC5PdK5QRyNJMQLQKu
pcjCXCunrBpxLZ9YR76r4Xb0Fyd3hr41pE4H/hAkqh/0L6pVp6TYo1RUSJSyvfjhb2slfa8UZTxX
oTPGcJzXqvWXTAsEpi6nyMAmAmEsde8Afb9w1uuQqiHTaGJIvHKaVKJB5EXdzk3mJV9EVOMfGx/J
BAccDq8h6BLILlSzIV6cgv6u4uNihTAXNm4LZRXD6Sh7jLML1rzLALQO76phEtYLEeYR2/YY8crr
bRTD678DqATEnxYCaEYpod9wVKKVlrSw4CJ1GmUg5B7I0yeOOzmo/+1XprGm3tGBLDwVdZyJzoM/
Tm8jICkrx5hmDQ1GgnNLf+cQLQQQ0dwQ5NVy5SfQRUEJ0tPGPnYzF8lKIBqb9vg7do8X74hoI2nI
m6r2hiKgm0F0hHXrtVaqOm4p+XzCgLz6mv3xHZ1oIbQvR8SlvEsGHyozNVkhd1JyVDx2MhJCdOlc
jakvSlJPa1Ym9EpnKImjKp/tLtSXOYqggZaV9P3UgqPf50U1BTPpODzYWJ1pv8FfqUoVm0aH5yyb
xm1xPAqYAA31V0Y8YVS5j+h9uAdF+lPwXuhtQMRo+Q6HBdQESlkYfhE/Wj2RV3bxBXi5nJC3FQ93
rynG9On040SsAmfO1GRFl03t9Shvnv5k8yUIkv9h5iabekFzyktDdkhjzTqDss2GiXLwfdQlomtp
Ktetw9ddzX4/gFJLtUupBjCAyKRj4nk1IiKTa0QDNUWjLjS1NrlFW19a6NSFNaxCRsttubyBd1Ce
MzxXOxgWNdcAFiGxnuhI77WLPwhoj15+5/JgC92vRbkwMaizZDXshH/MQ1UAAbn819V+XdGzl+KB
28H3LLHmjRg4uhMtxQuxW0zNtKD9e0RimmqDRmu/4z8HLfczGPPfu2LKfbtSaIMlJUaBWHnSEKf+
zJnEX5jpDiJPmxv7UnqJmEKDr87/BnNHeh7QDghzRBvRub4T1cir+Lw46b+/HHlXz7FMzoH/atsp
ezvC/BDxWS3PjsCKw3xYfjyG29UIlvvWoBKgtTeE+DIznRrS2VF17PHOUFYgYl8XyO/vGXGKXWk4
5mTGincIlEp5DiFih8O4PvuOJuF1pUE3jWEJhbYkTv1hO3TWNlRfssh7HnPg5e2Un+G9vbcaf7iu
/lyH1kn+odddH1OQhuMUXI7l+eBHjv+rzS6CbYFvSucpxQAAf29rTFpEmO/S2Xa1bOBgr1KtELhZ
55RhFpYrsOG07r6JmZKvTaMwKweuBVtBoJG5Xt0Wme2co4AYw7WlUTFaPEbV2WMyVDMW0fvgNei8
yz8IoKJZBi4937ksLsrF3ZsJ+D9Wpd/ewv7IqHkNqAnP1c+fCyEcV1fhnDjShfnljlyq6FzWlqfb
2QmjGPeu+0GQFl3feVkvH3ZWHcmII9qPMOnJ8KE6rnOeyl0OUGOiNwD+GKZQA1jvqcZgYagF/tip
6UMw7mW8uNl46OuadNqJu38UyKSe2IWTtTv0IF79rTQhiL16YtWp2h3uykA7gcJovwQA7FYrLpNR
x9eN8BeQ3MdgGKG/h2U4ZemOqBD4FKlR6NGa1PXc2yzJ9owwbpKa3Gay4mPnLSd21l2yhC89NubI
Ly6dVEwPoAiSm/2w6MDsgc4FSErIqTKv4f3VzkVRv20+KL9dZQsI1KVLWnxMI1gdrr6ximMWFAUf
metevhiV3CYwETNBnm1+NJKU+5N2J/wine8cW3B3UI9BqTGSvwycCTJFVdyIWs4z358Ah+TA8smX
yQgNAKFmLJHZBwIy4bok+9yX82JADetoxBXhFHPVQ3dugx+fF98RNZSa1IWDOpqq3uZfEXcRbgBf
rMgxpyIn95J6tpsHEEpjz6U9WuY6EoPl8K5dKgtfXRrMLqpdzHFmdjPpPCrhV2A445A7WmajsUyD
nyK02l5T18Tu7Lwl/GLbiALN2OQxmHhEL2xpQiNn23uYa4/sJjUeero748L00NPBveUT7dVeyi1w
F6XvrPFkwTnO+OqyZk4kkFECWYNmsvhbyXQqOW/obKc6bZxvNv+O5teApLiMzhEG/HAcbObBNUkd
D7VkFWFv5jDFGFwVZ3MhlfZOrhaeh7UXGliq+JUiFgLgDmrHhiHSaUc/YxIevC+wGpgLDpH8B8T6
NJCCVoG4Pa47YknoAM5QWsC3etw84Q4MJaasSqQGQW/1aMp8g6gQLHxU2dmCHElVyXdW+Xr6XmxL
UVRMGvZU7wKnBkj/6jSFi+C0BAbPGPJZcxNkX4Q9/tvmFHvxEqv/OnEDkutuKArI5M+wM48m4uFM
PKWXoxc1eJdXKjWKOvL3IckqV8muuVUpHsrWlkODAo66yz1iezkfLdRUbB7OS9rcSE3JlJRt+mLO
RRy3VuZxYGJ7XljvIx0yECuwzQDntsv4wqUjUs09pbGHm/4wB56RszSUQe8b0wwevmCl5HjtSMGL
MxfOObrjw6cXwulgUsT+U3uRIt3BO4/FitJL/dLNExdiS19DxTgu/R6/w/fkQF7jy0Zm3Hc4fjqR
sQSYPWUzPn/au9OvjUBDyLD8VKfcIubx7K4DdDs03zKg7wJeyNqvpll9WQFrB1R2zmma/BBomvuW
6zvjt962q1VWx6NUwWFWzm+Ojpou9VmUwMFL0LF07rjAe93sSqJDTWs/xpXiWUu7EA56GO27dviN
OddcvQUFJaiuKXHTroSJjqCqyDImed5Al56ux22AQE3CxYc0TgrefvMfE81xrxxHxFHRBJL9F14L
biXEhVui+Y4AfzKdkRp6YomxtpyCQ+l34icv11OJVwjvkoec863M+fMniBCiGc3M7vC1nZanwCL+
6loCz/VZphhaTSRhCc4KuDPgmtPuM8riQqH4NUQEa/0pW1gjFIr6rporVtwR5XX5jVk68pquXVPL
LGeMttgSomF0F4O/ioc4vhGK9xMBt2oyGUqZDOD8ZH8jK5Ng32e/FAa4BjdBOB3dRtdpIVrPaw+P
aPWvfWGPr5hUWwtCWY5POOT7wGYu1jIiXkdCjLeeD+VWNRIrl3jpkk+PvBNyYVjvyUhIUuQJ76S8
Y7ZGIoD/DeN8t7OPnG8fNeAsgkAJi0lHO8e1AUhSb0f5V6cpoEbz99/QG56MzhuMEXHTalCZHOnK
Ja4SDMqilHyGGNE6LC+i/QbL4zsmlbxS1F63YSFvQylahs2vz9+Akrjmc4r8gh7A5VHD7Pq2m0cX
+ADxCKiZbBHK2hQzz0X7ZyZBlW+izaPdoWZuPBfySqavF+WXeic25Exm6Me/nnk1r2N7zTAaR8h7
8q6lrIhbXdWI+ErWGKOTlzMoKqkl67wUcB1uSOAAaqacce3LyOImPa+pSD0Kp8jdubO4F45AH8mX
pygW5mYYWIJx5IjdRl8e76XiwJx1jMiWU0OmQlThNSUxV1NMn6A+fsHr8MA4NBohIQWK4Y89jO3K
l3jUxiJeOiCehUpTzdKlncIrbNIgbzG4AgLvmFQxz9ZBz1zgPw7+yeLNZXfJAUIUHvocBI8CD41j
j0oxtuGBLmtf9qivhKJoGe4Ug9BghzAdxVo35pZ0q7CY97Vibpn/4sUglSlGSIdxJPes08nsA7MH
stXanRpAjN4T+UCdtwDHIzIJhmK+37/iPcTJNu/0QZjdCEw2rCcuOstcmcD8ctl8DvrZ9CN8897W
Gh6Rnl11K6SgrqJy7YbUJI4KMIkayXCHt9R7jwnYG8H+ZemY/UB64n8Pd9N52DOi6AEo4Qfu6ApD
RYUnKxKIhkegMohM5hyNCmMPRoyNzpTww8i6R8BPwRO4vFLXPNDOBVOLtWnSgzXnFz1QHCWdKkMK
tjKfXhOiREbGdB537xxqoSQzCEmcbDATbXNWa8Ua+eSJV4F8nV2h1tYwS4qzhNAZQLgzIjXGLRSp
+JIX+1sKDfhcde+Puj90tlNh3BOFMZWzxGYbb/qyQaEHfyD6ppNFPrgHKcDOiqN80u62kjh7JcUI
w84navHqi10ngOVWWie9ip00dSkI/C7ktIF/L5n9s9xGxV3+vgXvdnUVGETF3TWn4zKcQ9SOfDhP
bVoZyMLQ4MDSlFMMaPSLYSFqn53hEgFz/QQNl4wV7lPDDKEQXibu+iYBfRO4FaecBpklbk6tacSN
j9Vx73DTuY3Nch8nhOMzAGqZwPwikcD4/ABSZOsKSrHBYT4aECy26R524YNyNsaM2sQeDJ1Ln/9u
JcCDq6rf4q+J7RjocefsluMIBoyhgZ6UmtoXvbKw0aDwhWNR3XTSvG8SnuBROuOMhRtR9/xpFdDQ
KBA+Ru04lJcnBALTkyvL45za4gYbhk/wlzD3EKFF/NDmGabKY5PwgV9U7WADI15qKOh89ZgWebpU
ip338dUUhn4A81rqTAdOKY25UxPQb/BnPlmqGOXQntSPWt9O8k/D60hKZdLzLePnN0avU+cbo4O6
nbrl2BPplEafFDAeYxNQBtbGIKFXHwja7WoZxXKY4RDaCE7+/r+RH12My69LUlSmrThj9lu6jeJ3
ZyhmMWpuYv0UxqNcGZ87pxy+zCtOmp4lWZC3Dv8My15/WBUSWVEjIVrC+BlunGEoN7RWZeY62ZwU
XpifWB6ZCE5FAsv+H4teN9kzm52aTdvik1MomlG6Qm+jL45JBdaNLemxP6+oaCMyZiV6V98iUnzf
D8PAnFHOOLTGCaNM5qGZpU1615m6A8TOg0qyrPPQ7GRqLrVnobLvIXiX7V3LWpOkak6Ti0Rr9cbf
2adeVUzw2s3NiI2lbl6s8R+Zq/y7qEzU9UAb+RKh5Rz03BslGKPq/ptW63FjvIUM0pFEjKVy6SFb
c93I+NPPTZeTATfi+DtqZPQyjAtqt/HqB+YxNy4sVwPtBAzimlBf6XFFgOtSMYr87Zaah1ynczvh
giwmqfYxONMhnfpjugWwlMD23k0cVbnTtPxnemrye+Lo3lI85YAm+5ihD8MdnOYgAWlu0TA0saXj
e6AWHLtUZXEdvv7v5Hr3JAH/dfRlDTfoug9mW6tm+ejIbqhEBgF4txY0UZZ6ZNtfLFftWVWNRX7m
f4SA5ELRUoVny5k7ewM9QzjGfo1VDOj+ztAwNC1QS/wSWfrZBWXIF2CrQj0W0KEe4ziWR/r4lifD
qt5h2OT0yO7mLnjvtGY725RvpFaegOrBRzQ1qNlEnDZsu1lF6tjiMd5vo7HBfa5ZvIsYBKnnEvDX
LfER91D/vu2Zrn/SMaQ1GBpx4Mk0lJBjON9ciGu7Q9HOr5HIxpDPeS+IeZOfWPVVFCp1YsyIHoje
Nqpe5OeirkQJY6s6gy6cT0C6fkodGO8ucIdrI3oNMUp1oyn3Cb0Nh/qXPg0lUFkiqN8KM0K9p3/6
2hEB4u/vW0hT6eM/Mi4+Bzxw5OaE9JpSFcF/LhoMYuXZYeygki41yeQ3ohq8uZxITRaZYar6dMDZ
NSg7ti/4ol+ch2RqWXezVK77dJfxJ03H7dlLSrvl2w+PuaPnnvBfeY2ijpqrT8rSgUPcOdv67mFG
phUND3quza98WOdQunRuh5XW3HsF6lwOZyEUJ3LPUmLxLeNSr2NBkvTN5aDGBbZGMMhjCp2WjFzI
bt3U+lMnETC+Tl8/yMij77gdzy1GZDMw+YGRy+lfui2BYhUuLV2QiY0FcFhobGdy9WIMRr0ZNYU7
Hq5YW2wpu5JRphcSuMnbNRYH0O2W/tQ0fbvrZ+JaO3GFLqhMfo/Ey32LurV5Q9+2K8F6YE/BvH8d
7SoUpVz862/JQMUYU/1YZoKs+WQQVzoKisbpKz0Phz6Q3H68r0yXMI67Unmgdwssmuhgd5PapiQr
umJt4BnxzPbr07/52iXKr0QjPK/ajJHql2+E4vXzl9cTaQBgCr8SH29B94yxOZVABC2Bw8yI9ilO
cAKqAfWyX/rwFqU5WpXzRvjHpomoSaDOS9ugRVtlUvSRdSFN9ILuN5bXws2Qqn/G66Ymrn/+hSyW
my+L3hyuSYj8CYmKBxLSSF9ZcTFsUDmR7fOVPcifH6q9VyzsGBhb55kySGzWgJbVEy7VtxHVCk55
9m+v+sl50UjVJtK7OlHHxlLhLJg2oIXg+CiS/1fk6Bw3gwZ4GAidEN2nGgmCr4rafeZqjHn6tbab
OLPNbzPT06rsD368sBl4ZpjOZxyZQ87ZAlwIr8VkJlB9F4zXTm+TJpUBsroQWb/meN68snZ4yKbD
cXpdRK+rrxJGsTCL9oZhi8Z3kht//5q2l7/mc2bGjwm3yPlw9GjIpJ30EHLNQoEG7wtIr8gG6xng
0Ipa3Hd8jpB72kltJnS5gtvlZ/J9vnTFvsaFs3+B9KFDwNdJC0wYEPujP/J6wwHoszCLt2EApx+i
xtrt/tsywPBLxQErZcA5kTThNTIlQNRb8eABdBZyiuFv57O/e51L2iYVJmB+PfFw586sh+o8OSDD
ONQ6OkudDEy//JYMk2663PLSrsSh0JjXqKZb+z5oylZ8heTpASE4eLIC23/sTyrlvOsi23fsHofE
lL8QyeUr4MHyYECXZUSTMGsLpqoEFHPfIM8sxklYRJfpUPVo9f7I/tQHZBWVhRRsjLzVxYKlNZDx
IjW4xMm6P0q9ctVYGroZNtNroechsHiKmNaHu/dSJCe+0wMplCmajMX8Wz7cHvycG/Vr+0WdO3/g
bNyEXcGI9qYuK7aDHcwYlep8hUni2EQxD2c5nkEQK4rvUXrb+CB8ygRPIXfUlK55CJodu+EQgWGU
1Fsz7CD/IzO1yo+Gumt/3sbl3xPkVns2bH5gJG9JsB9D9J8CDfqJ0fjusgRoSTLpJBP2aY6SPr6T
3WBJ1/MhzXOMQjwtuv1n6Fo9YD1t0+H4wxFGvZ8e7V4rr8cjgtF7vQLkfEcXGgGEaHrne91qt02Y
TmTZSaFTdWUxP7oEIBEf8MjwhDJYkDJtUe0DjtFFNKoAnrV1xVOyOKMq11Q98oSPrcMT2Q2GLv3v
jRRVFmsRZKzo8TJRrPNzpwrP0dkUh6cv8T+MNQM5T5Ij8+lBvmsR7tr9AmwrQVgpgsRqly3vnXiC
HHmYR3DzBcQvhdcL9ad0m9bqkqD5JBeiew6XyWRiA3fiOrwkDjqUR6sfopbHkpnJ+anfIY7OBwpt
i9VuOEMHQF2JNTQ0/qbnyKTg42jKaHMEgktBVhzIkLB4x6Wsr2YhkVl/TGAQaeUzDIFfLaMsrPSd
cGFzr3oL6NqDwHF/Dw22/nlXDLbvswHqLjbvJROXNyESh/KLrRsRhJgeeidz+YDrGIXqzkAU/iCK
PVVyOlwb6+pwC1Z4aVwQ8Ivg5FunhDiqwA6SCpFAVIjmh4fK0JiEV0tE7mLS2e250Do1rXJm+oem
zig/IdWtyPJT8nQaqy3xtoixjYEBws1CjxOdHTxfQT+cXKLeoq3Y5UTOTPcgD8H7bP9kAzpbR1Ow
fYZrM9AEs8k/0VdixB4BA+aVnx/eCVPNt/ySXe4Eu8PddjIAOmWrR9PoZO9dS4GpDU95TokuwfER
0w/etg9UJ97QBrjJUZUKm1/DEqAnCC0kSTl6tIVVTgkflT4HBnviWmnkby+pq11tu80crLlCfKMF
UnpOWE+oeIRt+cGaPOTd0AYNE9/TFELUiIthwMIkHFCVC5duOEu6SgK+Jd/jOeON0ltIDIwtOTeQ
sguUwQlcxy+9WrPKKsDpl/TudoC4+KhlgTP4RF07Ry6c0ikEoFq64m5LAYNWiYq/1BSlsM/bAZSi
EjmrZiwaqIARmrRq1iv2BBqzIt2a0FIDSt/qL+ZOfKfgKBBrevmXoKsZ+4RQUqdlHkUpa+wr0QYK
mW6wAQ/tj8BC/fWRhfbE2U8n+bPzl/Z/xG1Z4RM5oUPrtDy4qCQAlA/AbLZD9Ev1m0MFNTsxfcS4
MXlPeRPJ/3Wrx+O4icRo75mjilX6zYVpyW419wwzK9Ty5e1BlEn7v5J5tXyoSdQqn7BzJsE/Vdgw
xe+NY4yIQBlJCQZactllo3aOayoQ3q6KspMRivYggB1gkU3dxenl+hIzTqakQu0ySppcn710gU1G
w3L9N7qUL2a2zXxxNW4Tb3lYpGMVZH9mMqTT7SANi6AIfRdSp/od+MOAi0nJ4iCFQ7/4rEhD5c+c
CqQp+dtNcUE3VbYJ8H3iij0wH/Yo5dXoqxun20oWwzLxQ2d8Kbz7wzWG4awJ3AsrUzJikXAUy4cY
WuVL1OCEgrznIyXRKak4aRkQHvElWPWwu7jE8z53OsA3oQgepLTPsDmSdFyB9b9zmxliq/SSrOtA
hJhzTdtEuiH+ZhkTbQQQI/RrKQahmxbNg6Q5qTh//ihqzyYi3QJOa5GvV+Lt/0Pms6sFDyERPcU1
VuKlkzAqVhyeiU1tXVvTGe/1Z58jHD0jgUL7zo5O6oG3cqaByNRMDN934ssuyOdIdeh+TTk88QTY
eOOj1bEF2wfiK7n8nNr/Yimkdo4w/AzfxwEuQE66aknVnNo4zKns3PJSrso5PPeV9UBsX5/fjL3C
CI+4VAX8FHKwdH0yb4xrl0we8UnJn8X44CX4dEvzI+tkKnpJK6s4Kzp59MVsnLOxBe8BZiN262EI
UJnB7yjcv+O8ySEGZPIlaM83O+MTwu/oBFvbvsvrb+tLm4+gbFu7LQc4E5fsedz8pijokzlZFqD1
ctKJx4NRWn3NojNCuhiK4pg051lFXwSt9QLgmztrjAe82Q/4LTZv3L+VeJSZjnqDzAdMJIBmu35x
klDMRWzngZvVwQyE2EPu9NANdz3iT5YDuaXmccJhcmHhcex0R2PYp56J5b7p8WXfU7pEK1viCEeM
JYBO4KdFyJ5FnB2OSAUgDRxcATP/fqFqJHMQCU6QqAM9aotC6TNbtkjxC1492Vis/a0uMvp/fmvj
XufjE7eRuL4bHSiRcoa8BxsqADHWnAo5RjbHPoh0r2VU13xWRPvtxaNqsteZthz+/bIyqJ8WpWq2
T4ri7pnyCcQMzY+BSYN8gGiqhY+DYeeVlYQboqcYVAq2CieJdd+kBW4H4+NgrMDkixyF/96Z++xb
bOErH8iU4Cf077c80kR0AEdrENinazCN+yF3pj/UpexM6iqN987B9b9ZOkTof9xS/Jdihcf1Lzhs
QABLoDcq+lXCDIINfDlkayNHoAizU59v2PRtPftA91YvNb9Ccxb63dH7VmAAgbQbHjsa9SL0l0Rg
o4O7Bs4P6jQVtqBqIvCefrruWDwyZvu5kpvy2gyPJRSJ6BshIgmED5qud+mOFBvhlJn3l27eWTRg
XiwgFpHk2PDOrLhhLyHwMd25+TLm0OQw1LFOs8Gm9k9mFVJQ9WcWNBhxRTTMLmdsAQXjiVf7um0O
O+xuanPIZ8Lm5KO/ZQ7enrV7WTwFIB13UHNv+wFUZMx9lX+oXzmx3g6DGpO3YHN7+Iqqvh/ojuIa
I7LIjGuKCPR7bJfvOalD64HGW9LbFvfIkSzjgPcTw7R8vv7ovzFDhSmhAzwjZaoeQNeNX1v9NoU9
1fZS8CWcNAAwk3tbLFUYKbWraibRD/C8NpToUMFgGeRge+Mr/m4LPA4xyIYNRhTnBY9sbYdNolO9
KIChytXYng55VmwQVJIu5tvKJd3ifBuJtVQkBwhjJsRqqF4aYBxCxAM4WxURK9xEpeiulJ5UOtJ6
Vsarl+p7MgN022rWGAQq3SEVPn/kFX9Mp60EB28WyU5O7PjSA4ANY+BjpKVWd+MCSLMC3ZNd+pv7
c7J0IPjfU5Qb7sEgb9bghbgK3XLOAQmCDUT2l7yU8dQoOJ4T1h2vhrUHvSnjCH2VNLnOpbIuJ+oo
Ag6Nvhdak2x8frrVzGpeCd4OFPtAmZ33MLyRje1zFkyK57aCCTz07ztLo7Fq2l3/Wv4y4Myf2Hyd
rUIDkkFQM6tbig23VNYmheEnMRBvdSUtIQtfuF8ISb8a1aeZQNbb3NqnJjWyuQtEMxDiI+LtEvnd
vbm6+7Iy8brHXBP2nVea5ymStGc7zgdX+E3iTMWyVahfF57sWzc9ECbIr4SfoYKZ5ervVx2Kf3lr
yv8NidCDvxlEDoeSvH1Xjrn5S7JxqclZnipw0fwv/fz0pg3mDqJ+yKQLbbJv4Bhz+djUjl7A0wdR
oZ0dXsSljJH1+fHPdAst3Rqz39JPK66WnbHL7SzVQGKUkFqEKn8WiHJUldMtX3WxBmwZ31ilZrTX
osk20nZ5PDZhr4TtiahUi1m0XW8j2Lxh2BlrXxuyDSI6CyuqbtlavS+KzmIO54G0aK5M2fiCJMhh
506KXvv//PThObW+P8Jx+a/Ae3HZd8jUVZTTsPkbIklGwsb2wLcuBs0VKrTPEExeSw00KEMS2EWR
tLReQH5hmhC9bvgAe6w2JR94qOtWZU2NBjAaanj5Gu9yUX8pdW4wA7uV8gCcpp23o2ti+TjVXgLU
sSdH2xruFxsOmvW0miOjh7CVZxxH46En/UmCA7vYDC+eX4Ka3UHgo3H08ldRR11721NHbFOVaFC3
WbJpBwdxKoCx7sBvFySriYAy4oNuL3dnPKK2YeA3dyhnLnd0pPXlRtnvAmq5KNVQsQUXKdaVW6xR
udrAy+pSPY90wMZLE5TncnKCnxrM57KXKOgy+3jRP7LwBYIZfuF5aS0tHDkwf01uUiCrWK3OPBQf
bGTXM5tWq7OumWiTMKSPoZnbw001sYfpGeamxvLPS8LaaT4lVHTGAH4wR8xmhLf2ibKteLbfZT24
mpQkfQs29sCYloaj+7y4DsuVzNpa1XQpvEF06H9gEMBwgLqX4TjArSe3yD8CDNmwTgAutBshv1aP
8f0H2V3q2KSl03FXOB1EFFlrwD5WChNGYRL+mrKU7jGeFbaOKu9DvdrbnibXAPw+FCY5l4N1fotD
kV4yLgl8FvX6ZzxXoVcXeqx9nN12cdg3GkMDd+bxaUispWdJWyAfrV39IMBvCaiwD6q1W5imybrJ
F7GjlBkfh/k7SiorKf9qEyH20FRX/7f4jEb3wVCC0KNV8LYshU5ZZlJRalgxWW5TCCUf9ipgqG3h
n6mBLR/E4LWZd15W0WCaU0DGPtWsPeb3Pm3QhTL4Xq1LOxb0orc6Kc1LirgB5ncBfjTRxuvYfoSz
R+7VFIgUm0fRzJD700jg2xc3jp4CTpQSw0IiJk53lc3oiufihxTrUhWpZTCRCS01YUFFjIVwC0gz
uqXCqDs+fEZoLfV076nQxHuEmgSP25/6lQnJTKMrDvr8dFLeTrc8m+trnkQbyfvmVjwSfBDyu3BY
iN6t9DTRw83M3D/Cjs3Qd+frUPhLwnWh8NoB+e0bU4L8Tr0OzrGyjbKmK6ud9bWcNexFEWPywaKT
Mwadp8/0MX08XpzHKLSRQhwfjXaq6ZQhU+uz4CXoqVBB3e5xs8afi48D1rRUCWn9tma5uGpY4eDe
MGhMtnn3YYaiavnpeBnno/NbZ35Up5Amsxce3yTvzx39So573YiT9iudev+9vCn3/xLc6BUwpfaY
0E3OI+Ix2W85ZP6MR6vvF7OOJCzL3k+eIROS2Go/RiaAJUHaH/76oO9cZzZxSY84XLli/yDRSKFu
QQw1VJT9YNhxv7dddqhOxHgGylsb9CFCvW0wX5zq+IHQjBN87DbtgE3vLIIh8z3TM0d3iYgf1kD9
JG/6eOkpDjqdlDDqJNEUy2w8tg8r1bSdJKopsqFTpuBecRLng4pfhigLFStBdiqgVkQs4hM+kH54
jArWLkYb9F2gYUBUehGDlqwzpIDkOEAJlCOoZBG6pCnIr9TjFFLzxsPFVXMEaabs8BxBd0PNcDeh
1Xy50oVLMwJrHV0M5+30v7OGNx5Zu3kvzv+la0nNGr3DyEYxJvsITf/jgRd1ZnAAuD9mZNtwFiBW
3w9mXuNEvapfa1qcZZngfW0ji2vXrTmrj9e0k46twc4iXFiPhLQXg7pN/70IsrfBozDvqQM9R9dh
5sVgYSc+LQFbdjpkjFspAC9qw0fJjrK3iROoU/FjhZa8UMuHJSJU//9s+9V64Hz1KO5h7mfabMWt
Y90Rv9/3XYKU0H+m2+9cv6sWrRHmnhT6L7edcIHzFQXbeDW/WjgWBGuEXmzfORlerVxi7mHbfQVk
Ozis1Q6SDBsiZTuaLIgmPSAd0IfU6sR4AoD0FLuTzZA1jml4iCSnMnKOBf+MBk0OJpbJGCtsop/o
LpN0QYOafws5/Y7aMa2P98fYsW9tDBrjLPTTW1yjSuOAMG9PsEwplaohoAGI6qyctbgnHQ+8CWpa
CvXBf5qW/FY/SYMkhCSG9w3QC0KM3GfbqfK+NM+4YVvgcSkQh1iMdlK9OOO0ALa5dUkN2DWm2Bz2
WJFq8N48EBXNP0g9UrtZyXE7gJFfscilML59dg51Xh4JqlcmOSzIyVSTcGJ3os9lBx1G944pW3mH
kic0e1rUVNPQ//4KNrYnY3d7Z7f+bYNJy59Tbu1PWX+NgqSKp0UWQz3BNLkvm08R6g6YgRb1aUS1
PQJr/mn6wlFsXGJMVzj0iHvZnEsb1PShM9YgslO3JHfEA9IcNOMYhoy1yxoWLeuE2+eGe4ZEUCsr
Juu0Akx740DXs4JBNLXEXKOi0kC0Vbfu8kQuHA3nDIDJcf4OZvJsKsvVXTgGBwO3Em7KGxmA73m5
ubb3eBDJXWcsv6+var4iCLdqD8s8m4UXeKg1O97Kb579zukx1+xE+/nCcJmCN26r6q80tHxz2hnN
Yk8MXwMzIruQAahXQoRr4ZV6MdsXGZkkYWP8AgCqvPY7NHVWOfylBZXprmpovitNTxa3EGzr5ZOG
tOtXouZvzpNaiiDXj4iaXviCD7ujYO70QHLVMRVKbb/SQ4198C9f9YZ2ps1yKmIA+saDOitHZ3+1
VxYRMGPovhHqOItDx36JijXT2llD/r0IHNMTr8tS7VkCKMtDSgwzBYlCzFxcgq/nB36EanZjTANv
V71MVCU1NpHlMJQ6nkn0Vf2FpUGvzJXeh2SWjH+CShxuuT8CiZCl0Kr/xC6e9CjOeYaSTU7GEjTc
l4WDKw9nl9KtslIN8E8tbDjLR5na+0xXt/t0qhGxNqaeuCFb4AG9GMe2Gg6pI2s8oE7Q8nwQDfOn
PYBe/IIE6Q4SIP0zCTaAeiC4oCAKLD0GV3CBTdLx9pFiKJwrx9ptYgdUIsINgVFrgXffRonoZP/6
oZDxw4s78ek6fgzAanMs7BbkKqwN1mv2o7paucddA7ogqRd5TIlrR5KsECTuv2+BpmAy51eqCHtX
us2YHPr+UDzEKzVPPLuGVYEu2EBuVlZagia7hjGvMTTnn4+5XTibB1oth11epyvhii36Q1+caZmP
TRTnGw9qtRL3X1Kpf0c6vikayq9bPRlQEOvFpOH3d1czAR5al1y8BwKKXs9HRk4Y5GiuwT5xTknc
LUU4Wez8TVybiEHB9UK6V2j9BXJGe+PIGdsSsPRrsfgv3qJKaye6ItmOmDK+aRIOPTIWolJKWgP7
d/NVB134o3liyZ5TELV4CL5lvQHQcCRJuTs/hxg+W8B9sHNseXni9ZVWaDW8h9CfShFk5ZVetqPM
bAoqpdZIJ061lrU+R3TN5jJjLecZzwPmBViCCUgkijOF1bS9fu5wHQX/MDI8FTn/eH7bvZlOT7u3
o8vHEgpJ8Wzo+Z3LIPfuSRoLuTimqBBZEtXQiDt0OtK/DQ4/541JGfKj9lQbg29WBbpTNMbru5ru
+9xevSKKGt7TDeJwnNfpMlrz1pax+t4tmNN3WB7D7KrckN7i5mtck+3S7Xl5N4av3OzQjBblowI5
E3MvV1OdXVeLaLovzXnoBeCXzSMZ0dSbTGM2WMjMJnOPgRy6lHR1/adMNYKxqedq05eQRo9ed8PU
NEKZkjCNQzJjfk9jnCRuAWeY70/hlOy7jqNZfqhGAsCIjiaMFxpPOHv8q8/ExUogcrN5xnntfLwE
H5oDOkjo7Qz8D+7mGoiuD3w4sKUleiUCHpcfNdjHcOiLtjNxaDCTZMq4rJ0fItijpDO+yzWKcaSm
/9ju9KzcVIJZcId6/cMvz3SHo4bhKXm1/cfOcd4c5SGr0CrGWWnrEeXtMBAUEXvZmn6ps+OphM4Z
3BY2s2/hBL0OvWiAoBY0kBE8e9QMy3ERKDintCUWQfdC1oiulEg/72z+yMpYA7tF+9Cle41Gl3O/
koUfYI4l0PQhFYnabyxxIlmZI1bGNgtXaB8yx6EK5YTHVaZH2IulGSYAoxG03w3g4/wcmWcNs7Q4
OIDRLA26Qsub1LwTfHb409IollB9Rd32pVL1aD+3arLq7P7LcTa2Fka9qjVuZ9qCuZIDoBRPcDRJ
BMMC8wrA5xLMI1yTNdeOCcvduyPxxVEgDJ3CzWxKOqexTahwG8M9GtbS1M6tKSUXDdCeJD0gUifA
Uq48KsHbNuWvgHFonM/SiAgMUInQbs9HOecj4YcM+XdsvG0JlqZ7dOhYA3aFfPg+LxguqvavspYL
8S+4OQI1bZpmnftgWz8+FCyNv2ApGdxkbaHOxh2Cpy4xHX/8euhdP5dws1MXIURCHGziM5t9MwyB
1/HMhFwI3FDtK5f3wTd6N5JC7g3RWeVNVFoKBtN3G2V1A+6oV0cE3MUbB9xSfP3Qc+y1Snf8UBEV
3spIps9k85EoZvnBFzKa4x2hSdsS1lQZiMQxU7LDAidofdhc2BAfPEQ5JGMk2X1A7WO7ELsZTdPv
B4qV+aOgih94ImZHAdPbXClzJH0t2gYfEjkQ5jGA8asY9tN+oMwvlUmC5t1TUGQH+BoexWXMCzn2
JJVS0XL6l4Zq/con5sCqT63XiGd2QSFsg4oZZ2WXSxRZTYToFk6o9tqdBcIyqhyNX919zz+cjoPA
lDOveuvB8F8h88lpcQd+J4Xg5Qqx9iTGeWrqYIEZAK/ZTbZUpYwpnYOp1ybm1QJUY0wYvcXiIPnj
sXc2EmnkZ1d1oo7/AZGJGlpqimK2WZfeF4gurF64L6i41RIy2qboDg/NAN7btvXeI5z7dxIvW2ZX
8FDf0zX80EIkbA2X5D79cxMV5MB2yBZanf6u7IjZ8ocgxMIsxv2QidpznSMerLksXs0IGnfYR3x5
JjNvxtjupns0omE2YSO6XA6UEZRukgGeJ8Wjn4PnYiF0I0Ug7JzxfzJg2MP2mZzTHnugXvi77XyU
/fjutFjB1eyzzZrOFZbQB2/XyGjo7ChA+AYWfnhaRHorpfhQkkaHehbC5CfkKdmOt1ih4bwFnaWH
Nz7SN6rKmLZ/se94xaEFJBfETnkhQ21SCRolPktaQTs0mQABNu0hW73U6RQjDe1DDKHQIHuFMNfM
cxsYHzBKAICqLePdUBJ6BSEHKev9JnFPf19j6ECrunflza8GwgWc7by0MU/NDRQc3tHaLGaa3IIX
SHEaFpxp0OV1iGbN0Vv579s6yzwlvgrot/sCc8a8SmHBVT0MdELcOED7jC963EolHcCDyoict/2W
0Rpifk2nkwVN9kxJ1UI8Dt4V+DcAMwMCWCKDi21cqLPl5nAlSlvAepc5PcSopwvt31lnB+AS+hcf
ao/Jr0vi0KNjl/sofZUEHPK+sLUb/wkSmySgTfRZoegwindNIyjItE+/THlyp6Yb5ihCJskmoZRB
n+3kEB74rE+LjHmjX+aG0MLezIZx8RJXxovFa/dKRctGmO82WA895Ct+qdsMQOwIBCvPH6YXwOc5
/cgZ/PM610uNWO3Ggq6DNwJRELB2YEaaoEjxVdNZ1V+Pv/0zkE2WPbzumKh8+FQZ9dHnOzJY1s7R
PHAPXB1YQp8uOo51aIStavPOt/Z0qUbI6nCeKSQnExrhmlWKMBIPz7F/h0/8bpQBmVM3riLJG80H
Y+fcDHR4Rm5PhMBoUpa7YGL9dyPecBYozSVLGL+9p4ChAqC4GgP88Q9F1wfY1fnPLkA3FaM/o54j
qv9x/iWAK1CY0coH0nLN8AUa4ayM09T7BpBUECSAycHwMJs+SHJMQmHbIbJ97e2FvJ4t4eVgP+g+
I4JxuC/7cPxE4bXja0wdZ1/c3xt9t+PZ3eE1WTQn/liuT4epQVMGP9qPzOGON63AfblqVjmp4w02
lzYupg50NzCvs8QP8JVlKE+6yShqDK8VsUI2y5Il+V5vcHCmN4pUPxPGC0BrnX33kGuTAbHYbGkC
6WaNlSNYH6uSDBizKU5PG2V01cP9gVaXr9lpnLTveYfG/MoYMHN2+J2CuAS8eCIMZSgnrwEMtSVn
8P1lAEFq/tAuNQkdu/+CpQjck4AXUqRIFiq/+olDGXjXR4zfoXoWHBlFPY+FwpdfasOIx3rudHjb
uYz2cI+H+xCgEYD4nkTB8qPXk2EmoxCHDfOEJZhjdJF7r7RoEwW/AjwHCcmc+EoZKARIHBLP58sY
F33jz6fp5r4K7QVpqxP2RpAVzdM9fBXlhbOsnTzzmdoCiKRJH+IzptqBlwBWuoQW8OyuMAr+qDus
pYPHr5eJflDtpqczVYAgVH0lDuSGi74duQNsakEBMWDLXOf7oA5Q34TeYzkiEbPV1Lm/Pg2RqgPh
Fvcwg0/TL9sFjnG6a1JXPjCpIBzkeS5mVRyi5W6ZYX2EldyMy/ZIh6Lpwo8/IpD3Mhrc51dExGDj
H3ge5IGgw9j0Eox3URRwFagF8h+9ipZg6qeYTku9z6j2IJAsGZrelqFd9M1vVLzLPMaS7wIzRPFS
ocUZONAMdaeN+R6VDeNJvrr8kdRKTQFORZZWPR+3WjW9i15p5qHft60P2ujdWNmOtduX/pUK/Z59
8Xpe0t4WPmExlLUUJzHwVfs+rcMiWKaI2BAXc7Zolb7lnr7PLJ/8Qw1Y1zrVExgNOUtWBygjOSEn
Pe9yUubNlbM7RB4iUF9p9YaxoRNe2DGRAU3S5LvHFCaLbpRePfixbrgSqLI4XmXFgS5QIFxnofJ/
wUBgnC/dD3dLD+Qq/IDav6hiXqdUMvaw8rNztq3ag3XF4amZVtI7A0bFk6UbF2UNRkkMTHzAzW4+
cEAipmMhHucB0yMAhDOk3k7S8ukXJdp+qBhQQxWTQs+1EYaKaCIp/jVyGdPO5Bt2WCv5kcrVCcrK
1gYpxx/AhX0KXW2zltjhTRSqbybUkaSBew/u1Ye4yxlhQ+N2OhnkmiPZwvB+BM3mb8R0Zel/uTtW
g6ipqITg+/E6KOKLpg+pciygYisGBOYFtQ3gIO1m23ZlszUrey2tS9yR3nxZVegxJG2JIVl7h7NA
j6m/AQ1b7EzafbNjrNTAiGm3GCl8d+blMLFwqltq6I7HomOrLY42YdFnyThn3O93plmLcHsc6GZw
mHqYcOTFnft2TjhxNv/xyqZefk8f4LdIqvfaisZU8Z6HCAhcqWPANZ1yzKrdvr27+22ORe3Jd0xx
HrjXKP0RcPsq290PSjuX0OXuoZ9b6xvMd5Pd07egJAZ/1Kg1mmNRODAnHam8N9YqsNFCMwl31p8X
mkwnifNjS5uFzQJdUO9r8kQk40K+y7Y0wMZ0LeIK3XsuTFpK8aduKpRg81tCEPiOpLqmjODk6URb
UZMK9cWXAwpFggRARn5ikmuuBoY3aCsxOZDZb6jAWKcYNRVRZU8bF1Tbu8Me7++qNVXc1LJfhVWI
dmiKhjrFBQCBGz4nLP32fj81hNZ08nuzyxg00kTPULA+Xb2U1Uv6xCS7E8hthCLzIwUCTP/z+u9l
k3p1Ov5TQwvHAOK36C+2iPQ1kXZjx0ufPSqEZdDWw0UDzjNfNASOiHeAr33TgY0LXkbY9uKQJ1Oz
Uv7e6eGVhYGQupjXQDEes+zf+dDButcbOgynXkpxYByjS+NHmxHMClzZT2d9MWJFRWSRMETWW6Xt
6BzY4UUal91afN5QsYrA33W5tTnJ51rp5RzTJI9+4QEhSstHsX4EOr+MhaiIu3H3FAINXEotfUOs
3LVkqeyxS8w3O4w4x0ASsOXh4fMSA70DGJOOjNVrlonnqQ/TfhKrAwWiweCu3apoWwGWGt+hGiP8
ogK/qU30Im/A5/BNLpD+Jt+VJ5pqAqeSrY/JcLPMRPQHPyESa+4Is/15e92uyJVtCWDd6SSuL4i0
dWNiuXqkb8hp4av3rF9WoAIZ0UCeRp7kJ2GI3gxtF+kfLJ3BN74wTzILXmUFvDeIZBEjWQUYH4nO
3U/k0wnQwXOJ864KoVOzb6fVXncqIUFwdG6WvwmHqMBuG99K16NFnkoJXObLYU0fw4jbYZ+76NRO
2lJ6l1+y+qfmYFKmEWgXaIJXza81P6BvO8y/41VxvudeapEMhpvZ1VNd1PJSgltwLL6psy7x8oc+
xhN7ikhSh9JZIh/wjgOmdcnfPUSLYfq1atIEZ3XaFOEpOAn2/ztFZI5QlUrL18Aw7QNNGh+zm5TC
FXV2Vh5/vkaY4s62uM9OLMMkDyX41yNYI74HDNr04JZsnHzKwaRvlMKDoSnPPvFtm/mcNJ/4zJwN
vyQb+lrH7Dut7ShHa1amFxD43adoerbg366qT2Kgbi7ZQOveaQ5ZoTED7gn2PLbe2w4nKROGUj2l
RNiCl3VW7Ah3zwIP4X5EZFN+kQzSRO5DzYO7RLNrQRSdxovpEC2xglyH1oNM6IHSK4LkmU1Sk6UL
gOz4DPoxpnW4u2oIiFCRhhKC3t6lYHm90gl4CbJcwFKjVXR9JleI7Rv5zZ6Q7k/d3nW9BOJUuL1m
nRLcNq6IClrTbM4Y/lrusOTAeYUJUiF1LfxULVWrFM1wZfSS7Fv2DEJ0qHFwt44W3jpWrClIIITk
HEnjQOq6EwpX0tRySJwW5yO78Q+eVis/J07PGW97GMlQF92ppfFGeEJsthVKya5OJBNFNmtqVcht
/gwKxHX1ZOk0gqssi4+NAYvWJG2BkMsG0b6UoeXF/u5bnPVfjMKzgkqkzbx2x574INPEWJlE1vTj
VbRlKKPFhOKADg7bSTvMN+T3GcKbdgwj7d6zrL1Ne4Y2P3WoOF7+dd7Y2Svu+LifCVDI31YBI/jw
3QWWMfTjm6FayHPCL8xEolUF4/8XTTOZ4w/0KY8m6YkiHoF4mbGgLnnoausm5rKfkAbI3LLllUjr
KxD6KVlYhz9MSDCR1GZ0XJ6kDYMrqAK+E+YvAIrdDncOVCQmyJJ5Ah7u4GwNCakZ6lLDtFVOTPJQ
iRd2rl7ZQs2OqVAYODDhnQFmNlXebaJC71QZlI++2GKMiAMr49T0YfdUsSWFgd6hOMnvGlvzYela
b6iVyiR1ds/6oan9IFf9oo5m+ck4acLHA1/Bg8sm2EpDnAaxZz4fRJDI6XHkFKTsMLDiedP08zdF
pNpzWzztQEarlVpzH7ggBFUET6guXc7yxvCejxpJPAb8gqCUeELr45bfhSXplL/v1qJMhrld1DYD
STTwWF8FsS2aXeWHACVz3FLw/3f04vvxe23aa5CFNMInUIw81aMRQ3TTdL5s84g5xno6gsR2gql1
NoESmLMRg1M4KjdcqZCbMS1KVt0/c0J9/iTVizH12k2i69kNXuaeUJ+5niTqD0fERzrgJWRdjG/e
4A5gsvGOcQH3MQe4Z8YsQWw1zlzafdRoQCNjdzWI4mkj56Pm510qmzFOiC5ru8ihEKp7SuOpfnFn
kgsBd2uiyp57ol58ejaQ9BB8dyFmpOx/dobfrMpOvB0dD4q52PQtmzHzv5XTv1+4gcWgtUDC5RLT
cqcvAcSkLqChXiy4eMMSWzH+XBqbecy2Hs6YYWyZUcIuANEbH6Ng3d9oJIPD0zcKwSpOacif2qoF
redMlrTi3lvcMoj3wxrbSE0aVpCkQtXnbeUi3jyosg/1mHL0q53cFAQgnw2AQZqBlmzs8jioZmY/
jh1zQdBsMPtsx6IQBX6vYtwAEWpH2GqyHnVJ4Mh36h/OvuJTa7oCz2URF5j46F8yk+FGZvkhD/d5
rGqs2jUAUryZ1LuS6cQM1viU/sBCey1II0SFcb0b43q4xXP/kbFMs824ZS+A5Acva8k9yRSRMIqo
F2pyh0iLLvfWylGsMBNnhR26DjpxdSNXBRjVbp16voRU0dwQgjs4G95SmeYNar3JjzjdtY6NHKAo
dS1TFTC5E459lnIAUvxcxJO03X5xeMkhWZVb11f2JQbkArv5KO9blgdwEAdkgWpk4x0syRC9Rptc
w4rtyJ2ADuWEwz1zgNFqlATVM0A0Rhk2a21JOvKfVmsglBsFP2RUq1LnELoKomrFo3PsGWrktCiO
I+tgTvzf/n6N8G/sn2D78ev/w+J8G417CxzWOZGVYEsrki9hEUN1r+z8AyIgmuTq0qDUdaURNRuF
FiF31Gso2qD6MWhjhpJHMvUR3Y1iiQEVjBbADcGPCrSVIxUdQtzqr2BBJ7wwClj37nPxhkxERSLt
yqSCnei+5Yd0YQKPyo8JVyFmd3I7ruUkSPVIFGD3/L/QmkxhxiQ+W9Lya9pZNVU5eQ9ATiM5Zq3i
vdAP3eLcUOiW5fr+LAqSywwa4ccJK/PQlaB5DOCiTyFSOkD1aF23ZJHWJJdQtEkZspC6Wnhedi88
BY5ufFCqeWr3GykJAOWKSy/uMSqBgVm1fyuKDvoKiWuTUORvf/YxThNK/ExYFxN0QoEDvn+MhFP5
S220dgYidOrKaeAkoey/YNY68BQgX1+Q4qCevvhyatmmB7e6SSyyk2khJElxx7bZHlWVZMXBZBpw
v7H6c2/Ce+GhFNUrI70gugm/6j3Th7J48TfqecTIXpUkH2Gb4AC+TPmMbPKJqP5Is6Y1PJw1fRH2
NK5z5o2Ty1X1vU2G6hKhv/zU2Uj2IgSSOSIilhPxxGhYPxkhPKbOgZba8fViwlxe0Yk7UbwT9VFa
kleEPRew8Dyu+FYglCQRcDOqDROLC1hLdBXUOM/TH6tB3gCKVuYCpMZXi1E5RkN+FSrusP28U/cG
hMS/gOt06/zu+vTgilFjGAguOf0LCNSKyDfZbvB+kQaQkuyJnoLpRbSh2x7pUL2wMnepCYyvR1qj
Nqq/yE5VXZGyl1h+ft5adeyeBVj08b68VAuyYjDlZa2gqeh6kfQaM1h1tp8nHcTP8ixWIJqESs9M
8Bzj4Oy2fNEXHC0EVxK5dLzRoVvLPgegKww7mwoeGReVBJOZdT2DTIANsoNGi1i7i0kLVwxb9fGD
NijSrRItSxVq5dCZsgcne2UyyNjw2B2Bi3sEttPxI3vuVKSzbf/4JUjwNxrdx/zcmIq1OXTJCKrg
XR1APdd4E+Z+LmQukF3rUdCz2TIrKCTpW4AK1wucYbfGWKwp/rbnN8bCx1RKs9xBdy0Q1yOpL+aM
tLph9hrCjQZLuygohh/CNVc5yCe7PmHxNcCS/i4je08O5wClQpeMMJt9XOiqDKNLdcQsY24uWOIw
qFESK3yCIKFFXPcVbJir7fTYWS2RndlS2eprB1pLO5Pd9WZ1q9+uG/7mbqSeRwSQL6dJU+kiIaDI
6XJH0iV2zNlEnrNX97MUi8aMBAWF1p04PaaWgLoJedu9kdrbzakJi/II/ZRCjbkUVLJWqQljiFtN
Svc9mDs26ZXJ4TQ3oXC+QTjhZq+nHVPWENX7OJcAwPUhwtiecQbFCg5JvhW1dA/4Tl8faMCyA2aM
E4Xd0lkpNP2Sodh1m6NMtFdS+z2EnZXua7b3H5T7IgbmSNflHgPiX8f+RqIXwTex9ehf45VG+r2z
gF2q70ntqHboleYJHPL3r5NG0+3yIQEgz9XXXtOUNqxUiAWCfvajX5jH3NO9ixSgWo2gOXblK3Qu
yyx+e3CydT0uo1TkvyUSadcxPX29DYk6AmDVv5QAhc3N7KoMjK/RfjvnO/DJa6h/4Ce+jGn1I5p7
g5/qon2WiQyPwv7DofFAxwQlqBw/MNzprrtoZ3vbL4CYVdsRoo1O0EV6W3VyUjoXQUubpJum/e2C
ftwmmD7PShEmvv6vWcUUd0pcSk9+ksf6FyAwBDXgjn3OGyIjBk2LJ5v34fVz9nGJIxXje5iIJTBN
15AGY4aF1qpfXw+78qwT1RHSQDCCY52eDcX8LQ7WiKHy2XxN2748fHjpTgYaKN8k9tPRMWPN/USZ
/mgd4zf52wyHtulWoWSkDok6XiRp9A4zeQzUGYY/p50H+Ccu/X7t7zSw6x2H5G34LlC8QJ2xCHkX
4nuALMH44JJWG0ODZ0jXsE1ilP3ub9koZ7rj8kASSOhlFzKBgU6Y9ou1eWorYTsPTDx+Fu2RSfOl
/JZ5+4SbUnEQE75kE/6sPaOT3DeMMIqcB1gu0V85/tVGnn98n5CtYaLOLZqtGO59eNygdyewwk2F
mHjt3m4roeIu2D+AKxcGcbBnD/icoJwL9aIu5rFIx2Tcjfqf9ewRbIba18dM654FBUbyK+t/3EPm
m0aKZQlRuneQVoyuPmR01xbdOep/vFXhe3zmmYoCBr8ntUdsGdH/Qaw2AO6bblEYaC3yzdl1zhvY
hQQTRQyjZtXBEavHOaFouZhfIWXgCfWcZAtHSGQShO+V+wnPxZPDZKBiixYbJnBcVIlmiqIAQpwN
l5QVdIyDFylVfIvrfXVmnQ6IxG9tXyjmV39HoSWCix8v+tidyPRHLvDXUtZzGzK2WUx+rANtqhnK
HljIFCBKXXCkfq/SjUCx21LQXkCRqR1TRCvsePtUx4TN9+34Qm9rT69DVbO5ksBbhn3+QPG8QzEk
wsbMM/KkfNKGSIjyhpqqET3RYnMGxcQQQcnDjR1KclA1dVubhyygCBZqtPjJjYGgA9YFnAgN6I+w
bqYHBUlpLhs2/vZJF8RJQ5IRZPfBF1GvuYgnVCwPxQfkJzXbVzsBw6aixpNzTWAirv2Ey31YjNi3
QbssfLGDfneraEQH+gycNVZVJ5xJK4T+VcXbNjRKNK1hI6OWNoAvDguNyjgVh/Z5HP5cOFJNbgl1
M+QFw9lzEbhwugexGvnK6cCeO2QCVo0NeODXgweUkLz/ybOOXPgu4qmJ4dnIrWtJ4DTOd+xo1Fiz
MkwKHmmIrNbXm+77gJXVx8jnGboQse7kOr7Uc+DqhTLY/u2c4oKTUalEMrY2K6oQgsKsXMbFYP9i
IFJuFJy8SWs+6Ihy3dkHkm5WaoFPMPFQjAW8/55AIb5JScjamUHgSYlomTu7Ndbjw3Q9+7N/flQA
gQGySydLqsVWBRHJzkwFzApy8Agyq38r3HM5HbouC7QlDvX84x5av+Gq0csBKw4NQFjOreeC4kup
2iYg4SHr4MMY+6O+i/nrLDYpHQ0PDKxog7Eo7gYnq/dWaqoTPAPdQhM9ik3IgKRR05IsLdcD36md
0TmtEpPY5UZC+wVK+5WxxHYHnlhfZUFY/9fyA/hWfa+U0EYvs/vDcAGVoXObUcqYY9rFCwb5OKtH
WQdCWtKoiMT/QHJ1sjaoqwirQlvwXFQqbdevWaC94O0akPQqYxxJK+SktvL+GnLRBobq0GFvqAJi
Y8pbXGpEhpSqXXJtXyshOosh1epugQwtS2Z1AghtLPsazsgkWl5eTrMxQPE+hsbf7lLYWRcWAgmv
/zE64Fd/cLC3oBkH+k+mS0Lra/QiQ3gEm5OKD10QSZ3PHAEFWUWqGXouOZTjvne87tpNmLgHqilE
cpe7MNlt22qO+OExiI5ZUPNYupJXJNYxslBxA6YUu5GXgoEFciooiP0j08NewdOTZvvxetPh6psK
HbFaihfg8oEXO+xJ7WtNcMtFLpdaeki3j23rUJ1SZh0XOMB99aUpsDO36FTA/1D19SveMt7XePqG
idmMuWwd5+QmD1s1UnUsqsVAbFcb1cJRlbQ36WHaUIsvEKTA61vWp9PpXHQj0TFwqnQGUThn2dqc
jEg29aXnUB/LY7xxFSuTZ49uKd4or9D7cNoWAb+g/BRa2bLlpwBgFU+6doibQgXM69HBkrngcY0J
IZVTeLeM3i0OBcTgPueMojNVTbhkUrcgufcNy/pt+Z5NsNHDmUERpZX4ZON62pi8tKJoRDKCzPQ1
B+JorugTHURf8ji1qrT2Nc9iOIfds9L9TmVrHuaLrJQGSNMYyHTTytN7Atx7z3jEZLHJJ6cgXQLd
8Fi7kQv5WBfYtpgpmhvTdLKi4O1JAmocYhND0c202pSjRpdxzGZKYrbKQf+kXYYYpoeb+jH0yDIF
OkBIBZP3+GwnS2RWSkwyLl9/kgHnwoQkJTS8wba/ym2fUQcWmjDJAcR480ZMx/PYmLbXSodVZDwQ
yzXG1m636atrx2QmIX7x9SxbAq4WuoNjF3+e4/QrzxN2ew/79YVrpC+6uuLxP3qYZNxJD/a7GprU
wHGpuTDlZFMpE/8CNJ2dMrZeXojwZs+sRmbW8H0+caSSkRkvkcI2UcVvbZdpPheAe5hIAXQ8+Y4v
UuOIwRq1BbIwRoYzfHvtSVTTowXxhWOKiF1kZC3zuKSa/Tt7AWOSoYqo7E2vLQzKZZCSeDsOGCHL
mnaGSrQXrYffddTvYqL+Dn+5M1hISZTwStuXbdRgKXYcFnCtlGc2OMiw/DYeWsH+IqbFvKpN6ODJ
hk8qhouBxEJXY96IvsU7g59hBW2xD3KjbcEQxCgVyLLVyYLgYdin/hAlbKQEqKPhH8lJR6eCA8CV
ModsUb0D66o90e+B/Nm2RzJrZGMv6M4CMmVy/C6n0A30/7/mL4ZiT8rPxERIJczxLwABXWvpT4n1
+PnsUwgAtXeoCMQoIoeKqvHyY4ZOcATNSLsxEui/epytZYO5h+dbpOOyJ8bQ3ES7B4D/xe8h3ox+
3a9tbsFGsVdwOE1foLzNBV4PV0W8roh7MA4wBUTayYQpSOPI8Qjj/N1v4KhARMVzypoJuEhqb4Zk
J+u4vxmyqHfHGBVuF+7kfsM9Rg9BdCx0N1FnCO3q98vc1+vuMSFiUozhajjFOe4xxi+QscHcrtE0
yJS0PhwisQgad7LfbH8lswyVDTF/G20p4hKh5gm9JOfX6NImcRjvIfKVx4+f59zPhbSt6J4CfEWG
aw7RiQKCWg9oDMvRFIzpw+LPj+QHVlNxzqYhssUDEZKIGcOXjVYI2j5qulNsczJKJx6Ud7mO5gwJ
28+wFCH/DZoNAll/pqsomHWbqJ3dwv8+btNDq55tWCpnAJKWPph5fbg9yoQ4n23BcJhC/McNjeSa
FJnBVF7LhIMwY08d73w/mqmdinGDkFpe+t9gjFIWBqWpK4LoZpCTZd5g8xT1GGbc7dpgUBDtL/41
jjwbs1ysn2ckv8DR3MtijBYOSR2waTnetQ1/lk2dFpSoWINmGgJCYzFzEzLvGCgPsGjEVUwLpjXF
JxM31ZZHBPDJ6JKntDS3BfnBr8rTXxqskbzhBzXRmnhyfGKkLYnUtX0QVnxhxiHR+1/CzZtmoiIg
xqWRqNj4d+ht+6nM1x2/hiEK/mJsD+CwmgfxYu9+8EYbs5RvO18e48QdIwi71AqqqCzFC6AK6NyT
CaI+4pbYZMOxw9Y5mIkWgkbSgcuPTGzRkdL3G3fv9BMIETAVoljNu7yDycVz0A+8WVXlnzfhKCY/
rrqeRzZrL1eiq1XMiEvDGID7tX/KZIQRIlTpNUcpT3TpAqDU/a+wWySehkInG6KqCFje5sLMPd/E
hcNg9+ooe4h40TIDJTDlTC8QP4y7UxesmQJ/v0nEN3Lc2ee76MHDoSCyWmjXodcYoD+9xx5pHv7V
PmhokolpPoCSEHx+2FzAETpKHRCQYNZhqI3hmnUB56Oj6HxWwcOMBewPJluMd2hRM2Fgd8z2gFVb
gHrGA1NaINjC7Rh5WBOjHQfJBx2WJQNeOinmWKpb8witsQYQiI13ccQzfAQF3h1/uFctWKBlMUOG
Nvlxso5CQplag6PQZb183vLrWFAHLm/85ABPA846IAcssCEYUwvYLKjpD6MfzmT4DzPdYKypmkl9
7OP80w3+Bx75Lak4sIRBW0kFwzKJ+Dc8XNadBAARp36zbP6QriFYFvuCMkXUnqgyrlVr0DK863fk
4u7+32A3kZE/hGa0copiQOtzGd/5OkE7wROvKzaIPOUJQwKktSjPixrkmBejc9q2g+dh9++iGy68
JXwOXCLRC1tlJUtqmSepoRZKu8lAl3eXHZnatfbK6lniYv3e+lxv/0JZit+vf65eKP8VqE0ksiaE
TQxSGQckMwe9xYHdpJjVGc6AfQXsQMaMw3KcxSv3qFrGJvalaoLGr06kqkCGDCCskVKtQKKCazAu
WBR3EVdo9M0RYVK7bOFsnJ8Ycckx5+JsuLmn49GOePCYdjClUJXaS3WfTQgXTdB4t+1vD22SBOOi
kqKzwg0waE1coYc5+XL1SbY1cJtCPNIV3k0Z/Zrlt9tIV5MaCKC0/1D5qTMt9O39dkl8FWdcf78K
LuaxYZvLCYfiro75SiPNfrneGY0h4GlM9T+QoiGtKfNUazSUig2bNTrNhBM7eY4sgFozS9WPYGLn
zOy461nc4HfjZ5lqGybXNexMGoumXouB2kdfvx0QEBXNtZW83lg88EYTy81QpjudwMSQ7Y1ulC6q
bURkmfzSOn6HJ7s6lOateJAUEtB6GT4akYzsgBwNOAqtbxUXrmAhgfAOQIFXoHheVD3I0no89iC8
RIngVzM85XNtmHvT1lHqvTLYA6+qPhEHLcG09HyYy71RHNIXHN1ezp/bAoT4CfAztTs+4f2hfuJV
rQRAKpGhJI78n0epDb8OajMVYSvr4N4EnCBtIxUYvbHmrEdN4YJk5YIoqRUEWIlY1arSyDEb1WRt
1VOM6/nW12dlZOlxt8nfJgxAJ7/K91lEetuoiLcOBsYgbkTqjWzQ+SuoyI2dZezavMgGQTWvqY0f
rxvC1rVt/R+km+7DEDwHj17Vde3qdVE0tNxcAnH0blbnerMvEclKux6Bngp9T3wG2oZ2EwNZrNZb
4CvX+Oj/Sv/G9VkKUrVBwkvYlDb+YCknXCQ/RP6lBe5103vaInmMAw2Ai1BuhWPLCiUJVvPz5SZd
NPleJ6f/B1yh43eLuk29TzQH1HcoeCYXo3o9nj4hm0NsVFJXBfvFDYTpxfv2sPu47Xj++34Ap0l7
b41A31zsiR322+yR3C8Ci2g25mq/6AtxUM6l+edXt8dwSYjxHhvwuPyBWOgh/A7MfDfcjgZcM45E
kPJ8JVUUBPy8MXAD7SdSyOK6RGbsA7WlafpvJT4GRfFFp178eaTwzK4tzjI6DLCCfb+zt615op7g
G5g5zoErElfiYyPWyaD1qOyaVz45UGXPuDW9eBzlHy733onBiAlhKFBzsry8UOdf5pe5ZSIZGffb
ibZoTw2A0Xt2Ci7g1Pl1Tf/Hn3JIaGxQA/0i0EJk4SJo7ZKWnraZg4V7+A71ygPbSa8u3bzMP9D7
Q2msfBEwWuJuWPbwA/p9KapZhJO0W8hLbA036pB4hHtxaj5CUuVkgvphyIqtaOrJl3G2LhU4szmx
WOTUkXO6XyAuE1JA+mQk3KeRHZe5UNhqnHC2UXpEjvnxPaqemf5Rk0I783+xkPY27bexRJ6uwI7s
5huMXeLMngpYPhgYoDq4IDxuwn0u8+Z0OSQtWqD8z7YIP6Bb0AWj32tmq63R3JvrgmGrVyuBimYM
Aic+KlkITvah1qzaNZdiQCZNHG7bra++4N86GijARGm2MNsGqi2U53pVcCKRSIFYXCGtCJ5BefFV
aHSl3byejZN3lTIj6xaYsWZCpOULU22n9YSQ3SXt9LL4GX4sz4aQuwP8WJdO5/t7kTXu+lCe0TI6
J+Zv9G2TLLloJMNPuBUiFc8q0LnJ6QW9GQbdLH81A4AmGPUfex3INIkFAchChIiEYvqyvFjhS199
bwYZcZEjj/ioDQzX6Yuc+2RE2Z/0aX5dJuixaIz8f1nxE5A1pv01UU1Ud5Ol5bPdjHF3Co8HkL7n
f5swJzHm9aF6lH368MDAD6zLjc3GPuz2aSlJw9T9eGYv/XocSISwiBQqC+3R4hn0ezFcfuMQuOKp
UFmHkKO3DHGQHEGaYCSBVtan3799Y7a659XtQyXNw+/zYP/LoPJ6JL/QIrzsaFpdyvepfKr3JNhH
fi60s8tsE2Tq+7yWFPRu43lrOisPVLRpiiYibQb7wg8MUKsBxA/TqGroHtStLQKm7LWmb4KOKe6/
XnGtOVsbSS2Q1vGhgaJcpaKJOz9nNAZY74O9o5lTuw2BtHfKLidrjieOINW/6xnoCqIQag5qaK6a
0jwl144VSSLX/PIzmbY51p7H9UvW1wJJ6WNPaqb8bcyB2lU88ItzN4cBNwjIFcN1icSPnf44XMpk
kvoH/SKKKGU058FPELh8NnxBltMEzmdhWGaCdS8Q2KR3g+WETEWeYbOIx/AI/hOAOyxWdwZ4GQ6p
1CaQJuHPUCZn61lXPQYKTC8D4zo2RywgcHnYpNAwA0IAIHmTu3HTxvgW9r3A4uD5ZdbcczVXM7TJ
rObHChBps1PIDkkCityApeXZoPwoDKaXVWMTQVNeFSKPY+kqxw0Cjq4IED/vOmX2mlYewDHYKxvm
78v6vuywdAeeTpqQW9U0Zw+N1Db0U6TxzoSxoS2koLNOAb2clsDa5xaHvOLVyiLi9RRo0kZ9v5PH
6jepVLVSREvnIJ2kldcvWtX7wi8T3ISB0kDNOjXQKLE8ZmFlVD8ucpKgQuGaWcdhFc4ZWICfVemC
6G9ESChwJA8r4Hwbyu0h5y/HltCMPk5IOlCx6B+d9Qz6bC9xz25woElRMxi/GoJVTtWiMCTAvX16
2K7WvF3MszaoZvuopPUo48dkMgCQdd4juCwAnbHCQ8oiM20f8xnX9KYF/QB4UxQeXj1jpWpuypRx
WLX6dm4bSrCXFYBVyBUDSmYXEShuEziWBvGteBM1gIKOye2/tLklyEQ5NQnqRWteQdl40HRsGEMw
V9gswqNhPGyPeBc+Yo2sPe8FD0sBfN7R95iwOIlvP4jGCZgBkN7KENmZxpENlkQai9P+mrZMJZPw
Z5kDs3Em+eUaiyvQJqQKP1WsbNcEsuq5RQFXNrLGSOlwgl7TFW2w1FdTZtqrGFkkmDibdUIgbBg5
U1U8qRyo2LqmqV1rqG7JYtKLFZEV8wtXwQMhPxVy13UvaMTGfCrwC6pc2Umscgwp/mBHm6Wrz8mm
FbK5Zp2SEtziMO8sAIOf1Eo9EIIi0t68SmU82UO4qeuKGo1SNIzTh/qqVJL6qciA75hKzqNzerP2
aqmoC9spnejuM3G3cvWeQ2tkC/Ma3Akxd8wEVm46SeJ6gOI5/FJ5jgGyUn8Rp+mGbH9cJ4izQ4qa
YB9RS0Sf0g1c2Ht452Je7sBIqwH45DzE+ITwM/dzqCv+5bl2QLpHcX2HU1b+8Oz3TQ6Gq+mxGvXV
UsVkpQYEf7AXVIY8s9Bt2/7Xs7zO3l+MuZAk48LEwo7nMBFWTwy7G50ypwvGxNa+jzmNkbzjPr73
jtIvDPA4BdEWHK17+StE8Zm7stud+hm9Ts3K92UNzy0LJUe5UNTy9amYzOJx3FnBIB8PgctrUEPK
yyWVEnZfbCfMs9iBkxrSjeuoqG1q0u/SRvcI8f0P4ocT8s5csM+QMgw38InwjSaQ8Gg8z9Hkfz4x
xMrJaLpHtLzEk+rFUW+goiLqvY/qbMhTAq/VNztEeiMQZP9IchaQT1E+8RHJe5AvzKrbTYnu5n0t
zbddP1Si7hT/MbBWiXzHP22d+vmVa+WtPB7KnLDOZWzQWFRwoOigwmdbZ47VOOew0KhasyHWuUAP
dEproRExkpzeaA4U/kLjMrZkNRNnBgrxTXQompf4vfaL9mA2QurSDeIKHjYgfYo/LneBrMC/wShm
xnx4UzJ9mpWhSKV9gnEVjJAovrXDopXroJzeKr+0U2f204p4a+7IaF5Asssh7whWdGvu9bXow3NU
0EaX4UQVyX/dtIQSD34xniBqMfCYegTdAgYOhipNi4KvxSFmyskBSV94t+2u5PPblQsYq++liNc3
/Jdzck04b6Yd0L1xnBzPXEx90IsPGzCzJxyK/3Vtpr7GeJASRneJDR7yfp3bhTbp1bv1eHy24ko2
AGlXIb19sr3CqAnNMiYUHHpzJKU6tCYLiix9xk3zMom3MSD2b4dJILGn2L36oVpH3Petg9QNMOxw
27om1jBXUzKgK6El+3MeaXwKG6+/hpGNa/Hhf8WBvI8RrgpAVGx2PxAR/2/Nk8fMs8/jbpPiAzd4
ThbI0gpdaKZLYDQme6l1lucQTtP1lNN82swBGPT/3V40rI5+USGOK5hKUJFYHH2nXC2A8B4OhdkG
QXmncAkqd68k8MJRQTDA6CQ3ydI8r9sTfHZxkIwKTg3mhlw7G9as+KpeDowfCw1vtsUOFCpaQPEE
T0KB6UA7gQNY1PCB3dHsxo7XqN+afLtbQUK3nRCf1u3+6m4jDwtFcU8sAbjXGNFKi0pTVcbi6Nfr
753jugZKg1Trdm4YXYzh6189eVWglENUyLfeCrA+2d5tSQxo95k/1dduGa1H4NcRP4h6TvqU3zLC
FXpbar58SQlY4T9ogEuv1fo0aAmif+v0liArxBhqgcL2ZPa5AvDyAqXIixdf7NB95dOXmu307zOH
3e7JrjEf+Uy2ZEsNdF1nO2ksg7PpgNTCOjSWyN+O4PlgbuBMFluBLX5b9TUbiO008oFcOAFC6ZjQ
hAZ7Fzf8z+KG+1Bci1JoiMckDgf8JrE+SvHUfIp50Er01OB2FmkBSSnXRRJMIPcSOb2b/dSrnBfZ
OH/N+lTtmG0iNk3NsyD1dNP2lB86R3M3shiNW6PrZhSpMaAPxiWLlBaKl+6gpEIqd1nXxafaWjR0
UBo3SOXsUGpevUEkICdH4onnGLR0xfM+2PZkA4lgylW2oCRzjWu+T/VIfUJsu4A9ZFOXfvUvueYp
bCMamC1kvkm6v1gLxF9Za8pmkPnLJciOcKOwYhE1sumnN7kg77kHdMD6PwyzPUWJnUh9xvGKQ/IM
VPKj3wv6YJAjaX7Q6AMHq5zEQqYReDF90wejys5k0ry3sDlkKc73sQQnIBYSsnRmu6P4c4X0+1dk
bLCRJPo3s9sbMfeVv9kOBu1VwEuDmW9h9IjksVaGtDFfyU0GDOwuWSrBaMRcq2d6tufrMrbdZPLj
K+yzjkKKgTG9OcwhU2aMVO3gtdv7M3nI3lV506sEdr/KsMbjBKhLwoiFcVGcYwmLW8oE/KBmttT+
qIr8pt+ha9xHz0bPOG5CoMJ7yzkHDsue+1W38Fb06GE4azxo0HZZDljlbB0W/ZZG5exrQKMwgbXJ
hw+RuEXUX/7f3MEFViXPQeiYxQX22fxSE8QlOE5RoZNrieBXp4sxxGStLBMO9qi1MWiBrYDxgm05
bSo6k5TymlINQWdHa+KOIOeSWXzgh7bB6tjZQc1SbtfF3QMdcwNBG+DjXBFY2HwVG1eZG2m77QYi
hyYKLFGhXJ2OqBDbWP2wLh4BmEDEYQd7UIZOwZgIku/HCxreRF9ji4kEpq3DDw9GK1R1c8rGO0U+
VecQ7L8KtRq02wdPQ3vfWTHqJOgkD3Zu7JnqX+ovq05D5ldX0mZkRM6OLEGJykqwy5n8VftzuJGn
dyY4rKbZkF15HPlbrSsmRVbQ/MT1tX2heFderqlukMgq1UKjpgPZ1vTEyg6a0KqA4dXJozFTvCq5
aq3tQt5iYec9gqQOzCLVYOERS3/KzFqr/1f/ilMgtpHhptkmCJOw+AjcZljnAgh+POu6OszwIA4q
V/ftHKcPYY0TxHOFe/qRaKFNs52GBcsNQD1d3kqwzpe6WWz0xSsHzIY0Gp1U2VdGPRL6BTVPL9Se
K919v0hV8oVwm/bZR3NOoSWqJ6/DGyEPCkZnL/ALPH7+NvzcdJ9AzlogdBEgvSTiimox9uRI5fBO
WcahKWY++8aGYdxSDRLKT31GvZMtw5vGIQrWeCoSLIvZyLTyfQKNR/VGqY98Nf4B3occQYHUC/H7
h6VXYKwxkOkyKtPxFcpadbotwo/5NgYQmrcIsYwrvfvm8KQmzX2xSrFVxj9xqWvpMVxYd/bh47bN
9amEATVqxMoFXXaGZpJGdkU8XjPJ29I22JcCBJCkHS6djj+KAxxfMuwtcJdmnn2vEnKQ6XscBATx
5sHj/GzRAXrp3wVeaPe7EXqGFKyn1uWI7HAWphqQ1SWmNHszgbH3kyXxFSZ/4AlxV22BNra2oDip
iXMjAP0PkjFOecHEPYpZ6e6K4ieosWojhbKHbiNvMQ8hiqL2pMOTYZNElV7g047LNI7SGOvhQzQS
UbfveIgc1rRkHdp90FL/gEEZnQYYPK9g16ybdX6Lk8+xoIe4Il3acvOmzesGSabZY2QRh2D4Pn66
OJKxrsaFZlRG21ILbQ+gI3TXC9J2k/tYZzTT5HIjdBGvvQZXDlrlnnMjzugfdp0iJ8DDHR2CttjB
w6J1lRPviyiXtz8fI4/+aMkMIm3q2xPhJ/5DMzfcTzs5gE48dAFVKOy1R3QaCEiDy+BqnW5IH8sZ
N3sPisUHIetqupIH/SDN3pAGvZV/MkYmUGGFKAK8PewG04O6RQgDsZFj4GhEH1oYn7H/gruN4aow
J/WbnM/mHI8s06dSC1j2oPcIRP8mMiY6d7Orny/18jW5ytncC3k9F17CbFYZlYE78lweTrgEYhhi
VKikb3pDo7T4GXzAOAbpPtXd1pLOL4QV5FmL6CtNpRknQMlFVQcmfXXgYAUflaxmmagoxyNUb8sJ
YaOcJ4ye5A2EVY0l+Q1et+VAC2Ur/UvTGbGbwcJ+kmK7LFinya1AmLVJxfD/I+61j7L5JcptU4/S
SM9BZTS2sGqDqTlOeTUlE0ZXRcpx2JkRaFH288ZCKSg1xydObYhSFpX0pIbTovVHfuTPPJmzbjK8
cBschK+IefCFsxeyekDW0bSPFgJBo3UK/Pgkr8ndahnqcsEi/yM6DjvJRJlUqmvkenmN4t4h/XGE
z1QRhBfaJLXDCJAFil9s+E1gCzjVbqCRWa05GQJHWWQpdiIL0cYUdZDrxp0BzHCh9DBv2FNrzfhq
yQOXvDiI0gauzTsrPL4Silcnu/ZP8116MzFpMeEu67ohdaNNE+JgpeeUdD/60lGrZAUYaXNsjRsL
cOaDSOZLj4iyzZ4nMYy3400Uik5T+2GukAaM/qmMGFmY/zLxoIVscdqZe6tIwgaGYdNpv5CKwDMi
xEQyG+GQrzdDD1tPhRtjVyyaTxYwhVGcXQIau0CQFBoX+cyHRa/NvqFWqsQc/vgbHI4cEV7tVN+H
+erAsdRhPBsox+taEQ5m0sIA+MJmlLXt4u1nzSdxFmIpnj2jDv0mx44JUN7jYa0wpwwiH/JwrgGJ
8MCXjUOvvoFMKy61yh1Gsh5c2ZDIydDG9/P++AEXGXxage3/tXQ3zlzmctrAe0xebwNpK02JNYT7
J9ogE8u2DUUyikpG6rf0Ce3tns68yvfrhR+2mpskdg/t8AmgseBHRVtXbMbNGoyNszLBd2Yz9VAu
XvkmiEr92C5FMvZW5eJL4yDfLWOgQfyvL8Bg607GBk/OdS5oFTeZ7Sua+0O8Rwtxg1+UZPGMYB+z
OlQBPR40vquhUxTBHMDvOO1+JKuVYfdiw/CEVqZVAdhm1JcmB8g+kx12/0x+8qa29Bsu6eCDBr8n
uxKG/yCxi4t1Kcxu6yXcBOfiMXiVE+g2ASaVeq7Au9ExY/TX2y8vUsRzNL7eASpEaaODqHy0qcUn
JFt6BxZMBcNms49ndcjxjUVdeLvfZs97f+BX+iVbQnqfELA8HBWXc1yd+raTL5NHa7H02CDRKtxk
TMaDjJ8As+9xdVsKIDQTNg8Wgacf4sM+vpAU4xEQKqt/X3imzhtCWyH1l+jwNX+9gJHFdrKBPLo1
L006xYcoSKT9xBReojxC+9RpKlV7PKlrAdaF5FO+yRlfXKQpIvwodYrzPeqz42F2NQ5spXwCqGOb
VfFGrQi32xlmGCjXgwkRMn3bkqyfaE+CjEx9A6p8tKJ2p+G0yiav5vZmjNhcJfj+0hHOoVGT7wUG
vWQQjgVj97IqAi9Idi0Pb/6zARYOO0keiCRyjx4NYrOmCyHSGSGBKypgT6hihCb+1PIQs4gof9Q8
tHcFQIFOJrP6u2vNQjMsXlmXiI2I+IB+S0c6pZvjYJcRkM0nSSz7GocjM3Nq8h9CkEBtr/QftAWo
MPIVEHHSYQb/GVBZOuyoIh0e9F6bM6ISDOjBP/Uu9sf9quYscYTK3dB9AKqmQLGUBoMuK3FkXRoF
Ky6LQBAAWVuMj0RiZpOR1FXVMIpP4QAJX/YhxXwEY0mxcNN+rvfe5h8p8xg6zfjIh45AiOYRL2P8
pTXf4KHfYmBW+ct13YWhjhIN6+T9DA0+jkVSG+S7YFNszYiTFAcLX9w8YOJ6HxXeF7DqLdkIs4Mc
7PjlDcqIVZF2gWqloDGSLMQyTixUddxxJCth7rzOPPWpM4tuBqUQCuxgssFBpjJY+KYPvjXStxSG
MD/uzELrPPwLG7kHQYU+pC55ihu5GZnN/FBJOJgmOyH9mLz4Q+ekGCQjcmnNBEWxZP/6zPlSkuXV
rONzEv2uLv/bkkYnaib1mzAYhxk7eTH4QSRizm7iMtrCf9V9HU4+w6YOWHCqlXP1aT4M+MHPcjlQ
q/g+EgGgDaNf/HJTg+EewOtqP6eLg/Ifc7EzHi75L6vdjPOBUvKQIhL1WOO/orQEwl2UuZTxpGPn
70DFlJXjjz/JeVKw8/wkxkcLvnZNGLF40IcHBTEYJPYmKRZpSyUOZCRXyKRPp3KAiA2kjAMTAXyG
dIvW8mqV1pV58F4yqUnh8ZQcjtYlDuUkiSpNYvUVuGks8+ALNTqcJmYrfMMVcUkBtdCfOhaLJw64
iY1a4IGUn40uFs7dmj27ykoZi9rArRb/kYWGLRZ9pr0C33oJo6mqTWjUzLGx2MS4XwOHPMFeuN1z
jSGJb1Fcu6mM15sR56deFQ3ZDrJ0YzWcIK0aL/868SIlWm9eHQVYqmaYGXqX7uQVtFEgA8I8g3RS
RLeMy6IHSt4Pr/a0NWaZhQV7eBnV+hAgFSQS1hgFsHLcC+bI7nms6Q4YhjHyiD/s3+6d/qwsADzg
gdZf6PgTzotfHCl3uM62vba8mJNj4/4DjpND79NQnrVniKyYQqAwitlEMk7yE4y3qjuuHw8h+zbe
p1F+wBPQoEWbkRCYjg2BVe8/xgiA1ItepvVb+2Vw3AI0yB9LekPu4SxSboUjIMK2RAFaUvWzo0fQ
Y3YiKiz933o+gFQqCiWVnsl6eE5PUK/H8AyvT6Y/ozuY4zjvPAQJj4EpA7qdEpaZ3ZVDqRKWAJLL
2gAFxHHk+6KOgF9a/hNdWEJ279olH6/YWt/0J5yuaHKkxL7s/s5pENrgXYJdpKPbtNpOP73LpCoc
x4V2NrKYZ4K49BiVgT/LRNa6q5Cc8cp+NSV7JOn+znBY2hU+G2MkZ3FQfG+aoaAwZOKMJy/gW/yW
wKAez13AY7gRz5JfJ6EA7Xj9OnFBurjn5EuPyP+FGkEE62dVcHHzgly1h90AjUhkYHPAEuCy5sGw
pvZdVkzcDgclOpKOxHhYRPSqr/jAW5p+wmqj1UvYLIZcs61MbXZSUA0oItxGCQkTLPdy4B7pEsTp
6DZ+zkbxohJmtui+MpDF44xYRIOzTxKENFaqJSRBKvVKIxGZ8uNoc4FPg1CN5oG05+DuZU6IfYOv
kx1tO9J6lmWDqsJntYFTkIOLC1IdJ6ty1XYMuXHBV+Be+iRkQpa436lT6ObSoy+p+wR1F3RbvopK
xYBqkzWZuUyn6uYCiGrwl5UJlMoG1bKccwCzBDap3BzI5eYkuGW1QW9mvfqFuvzJAG73HA7z/Dlz
WEdwTwJ3sTkqtJUottOt99esMyNBlLyrD0cDqAmMMbdQmmicyDBhq9+BUutmns21p9SgKqQ9KhFq
Uoh7saPslwbYn/Qui4R6cnHc2/+YxzS3dVEHvHJ3B5JCXMSnpjklus4MVAhar55t2yYp1KFKiwiO
a2Afy6tnII0WpfQgsbxNAKVfnfAFXV+k/w7RnPoF8sKGzXi0yI/9ZMPwHfw4sjyhV8Lnc5P1Usp7
gNVqtJKg9+frw9qEs570uTQcG29PgUpuu+Je8vO2hgjxMGUlu1c/Z5oeLpl5zgR7EAbw8v/uplJ4
GYTAZlL78rTvk8CAIr8Swmq7cYZt2HBvkMbsTYay8hZyQIBZP5dnydxbHBBSOf++SLVifr2HBx5s
F/BVHfyKEhIZDqAxbD7IkPAzQa68mxZrw7zflwPaeZQv/mx9i/6wPfdwFTCaW5y4joDCiL06M1Py
3wis+wXaZp+nYEWBSj4SFEqLBlRmJSuA1LvIbUcb4VgUu1NTegjGmae+LNMaPNMvKhQTcVjFkLCP
M9HNOepWV10+InSzQpWCs/0uWzfAsE+AOL0XCIfUlQxq+++589a0wCLe9vpqxbemV3HAincvMPdE
FspmUXdpH+bncxsalwJg5dZzHX9B+cpWvFdVzfmsSATO0rLn02tIbEhhW0H9GRfkgo+idAJKut/z
xKWd629k0jSgmM0fNX6967YDVYPTQFqolMK0fRsVUlBIvdXYwYx6SeVYKkj/6GZeSoXvxNDxjkvH
VeMenrnkyR7LfPTtAAyqF4Em32ubti0Kgl0EiwrWERYs2HKsU3q85n80bSxk9jaFnFKcbyocuEiB
ZIPs+0YYV46W4VRTMTTBxJ++GxHN2mbIi+Su+zoW0zOOFbz9TWO0tY9bUkuRcPOOnS4hRNLfo9Qf
OsqN2jrqdFg8smwcE5rHfBWbGubV+iQdcqSLqjP5Do+WsP2auYztbv+6EmugYKwX5d3KGz/LKg8d
hpp5bGq/01VyzQlxTQ0ALifSZ52bUvU+JA/H73rYmWyII6Ib5RpMZQIIQeOT6zDgQcRQlcAFqkJ2
Gmag7R6Dml4sYwwjgncao9wElvOAZZBqTk7RtMVXHUJneUuScj9nK9gfpBbYNFRYuPtsQVwQH95R
oz6ZVyi17bm7HBldSlhBA+2UjxXNivO2wNdaxP7Hr69dYUpOvwI2QJ5wOshPb8Ybz59X+a1MabNi
j1KQuqLmHwm5++lEUV6R6tU2uNsAXsjAYm7y5zdD25v7Jk0IXLNu3aF7KMFuXx0/+dHU2UhKQZaE
FaqeqsA/Zm4JFxg6UGnUyBfOR4NU7T03a42LTxivoVQICP81w62dbtgIEbElSiU2MkJ854EZSYCB
IAQBZ96/l+QowXe1HujaMc7s201SWJDePOdWIjrRkPo7VlXBa1feemfl0bZ9sxOkOkIbMphc3XqB
h55fwVGgAfeBHSCKZzFDxwJmjN9lReru9AJ4hm37K5ZbUzKY1FaMxZghTZYFL9+nNaqWrnDgfvog
z7ZGSxCwa19U0bKf8Nzfk32bCESqTdHfpusxvt3k+JdGWNk1XOIt2uzzB7bMTJzroLwSxTVfMLYF
I6nBVyPsOQmuNqnpwOEDVnQ8c84y+vfL8HROQs5bccsXL+FsmEpTkmXQ1m7gEXJNQkcYAqi9DT1w
4aKdPbsAX5s50zOe3QoSNn6MuJRafypY/OYFREcya77qoyRSATczrzPMOGvDsiK5hvdpgMMNMePh
OgGqSh0ELA1OehjuQ3MkDy6GHcAqEnngO0K8GSPpypj1cKvoEVOclabsFKpbgyqg7VUyufThoL34
0iREPHhzG68wf2W+NABqiWg6rQWg0CGEjcVPsLyeiHKp4h5hoqbF5a+eg5f5YTsS1uiv6k1jQn2j
cjTpDxXyzu90bfQySVtEW8dmq5msQYybAgEZL9L+SYGBjlllp07xgquk8eODAw85tKo1mkjVJSCw
OefKoILDC8O6E+AjcLBDmUYLqCYJ5X1NrVNlgvpJgXfe3xhMNgM/Hzsh1YQmi2ThOYvBtn1ogfuU
L0xQWEWMKdi5gHemetdTHgrLNlufwzUZe1XbNjewegp+2lFLB9+tkHr9/jkODpTjPiDJeqj3Qw0J
YcotEztMw0t8qHSvOrqt2K4Su6vSUumul0PEeQeeV/Q0VsG6MbFNKzkXA2BaVr7NhPn2oJ+WnJuY
79pfDLt0oItp/cad1fKvd8ugS04yevPMjImGQYFU8f2g8NIQ3aa+LKZCeKieNrWmUf+JKaU5nPbD
6+PlhFiT6v4at1LFMExbNkSCsKbhoGEbSRGgu0n7T6hAbMNYW0lIw01kxCqKH4SoN5owitaVj1k1
kzwJqnB521myVhh/RLyKVLhPapRANOCkulPKyh1BEpTAmOKlIzZc3Sx33mOiyIbC0kz8gcjfcWus
gtDZlwaw53TBx8CxrRQkBYBeRt4gpr0W2fDSqDSqMffPuu9MWnlNUJGNp+RF2AjXALmLUfi0NYhE
umVhZ2JkkXKKtzlupMevrNyN8On2d21iNcjeQygg6mV+NhM6nYpOhOHJLQe3r6Ahen3xryWfS5Ti
MOPZ3XTBdkQ0H6MSfdF8Po1TL17DTXO3oopvpegLetbBAUsvlzmVTNJVRiWFLcF0IaANxLyJl9xh
vCI8gtiipSPuPhWvWoKW/W8EGJjm3w3NT8/xH9rNvx0E5g/bs8rMhLem8IxQCPMvWtUN1jRlsvTI
cZh90yZIxF5bwyLCuNqWC1M03cTXpnPqe7mWaH2rubmSaYHN5oPktACq52q8sBHbcuFq/ppuf/7q
X0LTzDbGQOg3PciuSlZvCrygf1W0H7dKPSqe+yQ+nK9f6dxZXCEg4d4Uq7gWt1j5lJCtBFlkjbp1
E9Oj3DY6+p01Oq9w5SFF6UB3ZPimxmgZaANML2TgPux7m+nRRC4O6nNBJvSBtMEYKbxe8hsfRC1C
jJ8JddSaZx/Pd1SuU/DxiUPN33/YzVF8pm5k71AXiIciurs1IxviWvolzWzi5O9rQwhmO07Jm64v
WiRt7jLFJ3wHWEa6K+tB10mmbsqnidEFLOnAnrEqpy82FQI6p8frPyyref/18gqZr3ziC453mNy9
xCAdfr15lV4sIJJp85/zeJWt9lNp/E1zlvVkV3D3Hwzt5k4T510RVVCH7U4+jpoim8rPP7BmoLwl
/Vpv6KmYGAuxMgeVR1AbfOf1uWjkEn6uBeYTh0jtXrZi9M61A+nn/5+SwuV2ADNPGtfXyVQyKgv6
MP0WbMBKwtGrcJSACaOQC9JhBuQCk9qfpWdnyfAC1lrIGIEOgan5tXJivtmZNat62MkLy/oiD9vg
naHKfdbh+sl28zPuHugKTkq83HygwE6QPjFd9544ULzP1i2LWXvW1tScSkN7skGmZussXkvdf0hq
S5JDhmiVMViSmuawqmRTHBBriTwYmECi8wbwun/7iPF9xZmCbfUkJDGLMRvGZmrSuduxwjiYfge2
y9diBaLvgL+pDme2i4AZptFyT9h0cbziUOKqVnH/okEUY8Vs3fDbzMi3N2ddlCDwxR5bK6KF4qwy
SwUqEwLjSRysmy3Lb2HGYTtotkCcQy/0M071CC5NyeJDs1steh82FNaVFumoiTVFRRssjzpEgY4a
4AHzjEpd4BQJxjjdV+SIWJuL6Ee120kcqbDECFtX1ZX5H0QAvvEaIE6zO6lELwvkMHzr2heFp3x6
e9RfIpypo1YhP4bqN5vLMmgIHsnR35XQNSuKl/XSUYgAT8rfdmZslvF5FUQzeyB9jwP9EBj19Mwv
3Riufrsp206b67oqTx1nVAJkxesq2xkQMO6mmzf6vBrEYRH/IDw8EtzHeFraQVKLt5Y1eArH93pZ
O+RcYVw0fVz0URHipalOtq2k9ESbpveK8d87vzpYYlGvTN5Qutpn/BJHNQcgMGNTyMYbhS1QaoPd
wYPlZCFlKXScfkcU/TjBPcJuxa+5zmP070k5V7I5QmticydiIC6E1htxiwEg6/Ji2MQa64KpIVMJ
rpZzxHP3X6azSibBXcawYex1GDaWaIUIeApjfGAX5GO9+YfJOucDzCLtiQPN8U2jNZBBXrcfI4LK
jkPVS5CaZpaDPn6Dl99enWc95Fnf8cFmE5TaqvTmNAZeJWsIJFws6QIy0fKwPZqs2ZTrVNJ41CpZ
SThnjpj35f52FVi2e7GKs7CnwmU46Haadwint1X5r036T/ZcsGp7ckTZrM4hO04Pyj0pVlnP+Xg0
WQWw606e3gNwV9q9Squ1+mNYAEoUumfzUD3Qe3m3JouGjJcZgGAXBu19ujVibs40AAEydsPZxsRu
Z9koErMLs9cgOqksPSV6aIlTO3cI0i8eFJpf6Rsn7YTvwFhk99XZfbXAUTTfhLZdvCy7yt7erysr
V5V44m84R5aDkCC4jeTSNit/5qJC2e556XMXKL3apLQsio1ppEnGH+Be4J5A3YV3UQ0ekvEL8JEr
uiPKdVSPnH74AxlEviIZL2vCO9w4cBo0mKgwilYHTQPEjT201ZiZaH9umoAVqItNMFQSlWCIN4Ke
sKkVjkp45oz6eEuz7rY8r45OqFoL/pfg04AT+aYsTDhh+BDjt8tbiPa+B7XEZaKqBzoFARrL6WIt
J+tj9RWdtAcOZeGbLG5/bMl+O9Myd6W7hVocX0ErsXDif520l4HBu3LWNvSZJN4PUG06aROROttR
hI/gpaE90q0b39QEZKEJQ4/HOKKdAdYPE3Nw53CxGG1AMO3IYqMMdgKJJUv3+E/g+2DDhCZiXI7W
bdzUFz2rOETSGb8JxyVkKIM7XAXlSRe/rOxSp4quQzaCVo4YEulQxVNg8YSMQU8PQiyA0oG2KFto
o0cr600gkG6MBcAH86IEMqa0ma5bvErlK8QFhMdgJUioSVp5eexHbH/LxkkSMYqhT8QG0Za/RuVp
TUgtJfP2zE8hRaDJFLMDLrCmefjHklO/blpdHh26//Pn2etIOjks14c9ET4CBwrhYLWZnCEyNV/l
a6O+m18DoejpUCChp0CQsY9PSdCSsPcr8FfXKEf1nEy+jT5qnNr+M3qQKebMeMtgRBiZyuW3YJci
eR+vHBxusrenazJ6iJNla/ufyWxQk7bN533hjIVWYW6oKN0ivrsd/14quDWbTru/re1JMFishl2k
gxKZl+YpBMJr+yNm9ayKh42AibRKwdvUsIhPCyx9dx+zuPgCSF6CbcVh0zXdW5OYUQG7toaaLkMj
PtEaJEzHuxck39kt8fNb4bQxVNjbfd7QZy9W+bdknymgDsyKkE3KXnvizsN6c8JyJeBWMev1JF7z
Fkk7+16oMaPLrrqZUXFSfANeSHp4rtlC//QqjyCKy/Hq+iyv19Ke5wOv/xzQhHM1+NlYHvLb4nXm
tyUJp7ivGA+aprfA9EiCx0nSt0K1m4FmwYQ+t/lTtOdG6w9s4yIjq+fUYgwuptODWGNkAPp67Nmd
S4j8QA7gH5Z0s1yNp7Jgg8xT1xZ4jq9mc5ZcMSwotGzV0z+Ha8k5M54YDCCsivnwfcdg2WMkE8m9
9TF9IA/MYGM5qKopkOu8bQ9kug+82CftiOhi5sCyP4FLXIm48p8FuYntd3MoZnK61P/Bc8WRtAF6
FAAhECflK/kg7h5sS204Ex3BtATpiuE9RbF76U9Y2syBAKx8xotmYOQuI70Yfr36ROCJO/mYDXci
2KdQldeAvXrGZZ7oghQIG2P79tkMfFAPR0F73nVrpnFbSnK5Bbx3ocmzFNjwVvr43W9CJjc2Yjq2
lkPBaG4hk0kAEX4z+k6XMCilQbjVu0tEhUHqypFIt8lBaifoVsr3z99t4EMDU0JSUKgdOKQrCdBn
zU8I2wL/0iKE6aIHIckpUanuDpNvq6yopkUFHhbSnQgRxuJPUbocczSPs9iOQmdtVXBtO42CFZy3
ETSqBwPBBA91ljixtQpj0mvUekWedXbXnGNVexZYXG3GMKgT0mbUsxcNMv9MP6vgtLG8HWuwmo/X
BqpbYrLIj7T347ebA+rJ9XbwlihshO239murDfmZKZLJXCXsOgCoD1XSaoUpxafpI1a3P4dV6fjj
3WtDRkB+z9RAZIc4V5Z4V/UaROs1kHPYX1rAqQwTJLnkCXht4/ZenwhtZIxY8stRJkpmqfXtbivT
RkeOLMOVwj1b9rXgdceHrGlwLN9JGPqO7jo6B62TZwHbPnJRTxkHipyN3sT0mqJstcm/hf4A94lZ
0/JEQOOACa9Kt+gBLyLYVaAGzK8k6QqJq1EfetzJMhL/0khZ33fjLOVqICkvIqFtzjhV2D2jAqro
zoNuxMXplfYc82kxGUwGhKtwc+dwknA3zCVhgBtDGdhPYNfM0ljNezmxRJgRhi8rbo9Q+r9W8msv
bIp+pneI/qQxfu3aEpG0hk2mVSWsJjzqMBvKJoIapaGDC/5ew8DjI048/oGoSWs01lZAM4ULTUpo
/YiY7JWJvst5h6xg8t1Bj1h+5Z7gWpeSjq1cbOTToUNp/p4xtkyYPWPbAjRWTFP4PcaupZ8cEUso
IgVX20ZE/nWbfmpryP8mNPqNVVs8ktMsKjUXbx4rmKRMYwgupsN+Mqdalfp3GkGp3EndpLzJOET6
2k+7tDKYg8fS+G8oc8wdpfjVE9sQiV02bJd+Wyuuw2blR7rRQoS1meTDJoQOpgX9dyqO6A2cN44k
RxeFTmHsTHYFCcdT2aloqfLQc4AG9dK7W4+nFtvDOHVjyqD1DjK26MAPhKWCLznFDbglmIpKxp8v
RIOeiLz5vKX35PxH2M7th3UQ3VFtg885uIMRC3BP+9OOTDI3tAKn9/qrQnksWJU/ejS1uC82j5KL
/tU+VTr/+j15q8xqKSrApU157Z3V02dnSvDUBnglmGify6co37yorYQZrchRVz5Dee3Upv35bgsg
UEojFkmaLs/Bfmz2XrnR18PXgnC0+khAJNaf1bXXQcgeTmca9YrYnpXRrqnx//4nbrZk3ER4Qxhx
8GW2/duZ1rT7+zOJlpJSsWyFbUBc0k+7m+vUaEYhC/xNuYwiHxzk+eBPVg3eMTXSCx2u0i+iI1Ly
7H0PIeKnxFaaJ5VRRaChjpAD3w5kaQtdeAt5QrhpDH2i8pzjsAseovD2Z1YALUbvmVYDgMCUCkYq
NwciJcGnHkf0dAYXcpn0ery+XfTKd0R8UMwQ6z/AMOBGaoIokgg7dI1Fw5Vx/vzz5clpShM4adGx
Rhx/W+hazwMxSvLjaQQf1FcAvI8qvelZHw9FeEETWk7ETr2ONj7xbD7XPFP0rrEm9z3y/xTESYkd
pALZUy0cTG59Wxb5B7BaagRw6FlqFuwFHPkPOBYOQsx+wG7hZkUao2oD3J+akMWNdYwYwhN6oqGx
sjvhajc0DePdFAz5fyVT9bv6DDUYMAfAjVbbevbGHB9N/P2kb7oLMmH9KMALuDLEPQCwRqaEOI16
IFJhft0rYGCFHzBfiHjHmSYNoOSHopaIU/2s/M6Ausxf/1JjGSWiBnxxtk+3r5Dz2u28E20CrbFj
8clFM5PnSwdOkLkAjq7idm2dJAbOqL1jctH9KFqW02dJqX3EkduqDUJtbVViVRJoXW4VOXm5ggmO
SAfiVZmacAdBQv0iWYSTC/6Ci4U8wZS3gpCv83I6Nq6wgmDtt1ojj7UlmlbbmjtFaLfFlLJNG/F0
8SjxqgQZmV0QJo7/hisTTXYs++ujHx+rakkSVchpEme1f/PRLHzzykeRoPqa7WHB0H2b2bD5mNqs
/kJr+5t3US5SGQERJO5OC7eD+GaOHyZtn1dBNAZDAqnrav+3j7xVrIha/wjDkKofG6SyyWB/NYmG
JOHxn8w46D2/M11cMNZMXLNBg/ZfeLl9v3/2ayz0RqrFWbxnnH5us55VZmPzVjRrzTf0tkiwJYk4
WQ7cAapq7xQo56m+OR+LNKffpBiHysivHgL5+XVKDVAUnQBCA0OJ6IWerIuGTBjh4VbRkGxN5k/S
avCG0Xb6SkI5k6r9fWEVUO3ob9r3pKPl3pu7502TQpMLmxdItQ6bazm8m3psbmMZ+UoXLEr45jYM
sOBcxF6J/C9lbrkOXjpgEURblIZJ01LYVkkXV/Uwq0mOe2EjLq7FVjyb0VjwGfu2Y8pA+51yQbI8
68djNpGOqS6mtpiQam+De+tx+lULepdwfkX4GqFjrCf9wd8KxFwq24FiwdvB4qvx9B2X355+4yYn
6YjK/M2XZwqlupeNKRDaoEPHeh7kKOimf29cXzY+1kyMurKxHmGrEGRHblL1eBt6Vg47VHKBSx2c
XJiThM2kDony5StgceTEGR3P81CzYSgKUjLePPZ5NeovpmaH8WgEdJFEx7+xaxVjXxQuZWJBwL71
uoLauIApLzejE7YmG1BKkmLwmNrWVdTvKnUQ4hKOeizGHNu2nCZ3yKfmyovZa8VN/BF+SK7Ex/AQ
09K2Yjz54UIKCjoL9vWFC4Ix0PzFKPmdfj/yKgXB42G/QIgvBqZcKUpKR8qVSdxm1ZcfUmSxAvzK
FJQszzHkGQUhJC5i2fmXDm6lRYWDx74xOCIaLejXFlkE6a9zYhJLfB/o5+bH/V9w1kBbavI/KGmr
hTOtUcRPEdzdQ3KiRR5k61ZXmoSdX5uiUWnw4shURc71dX6XZzGpgdVY8yYMFdpB+UpuTbX3QV3e
GI25je9d8c4pKCOJt/ljZ1WCaDt2tFbc84exfRk274bO2AzT8bxJ/tE79lTKOdCza3zh+VV7C+S2
LJNp3q8DEPmcFa6rv7fpx9MjAgl60hBUAvaApyjSWCKTSn9F+3FN1AGtJKQ6uQFIo8oKUkzH5GPW
BWa+m0bj2Y4K1YdhdPuNdMdJ7lnAODoIsOr5MsUk0BcB5xKJ8c3Ragx07o1kWYRonEs6CWlUXCnn
XldIqAivS0pqz+fZHY3Uu3XetJWKnD428ZWDbArrb219Yc4mNOZKaccRhE1CnlLM1YTc0esU0GVr
cicOkAaOytEySKzYfZY3nxuqvyMGy2/r3Je/BMQ9DGo0itPnT0PIZCPXgZHIRBzfnRvoYbbN73w5
zjl0mMfzecrd7m+ngsGJwkMI8B95PljmKgZdBnOVOF826zUH0ub6Vo+YLUQ+S4liuATA8lUugogT
3b8twtFywQ0mXFnpWF6VtpTx6r52TfzFO+TMT/wUcAw8KmQ7Fv+HEy4E3Z3BVotbJ7vES93cLkAO
X+EgWuwdWk6xQHj4M7OKI36w6zN7BZPQpfQ3mJdxTxMidiiNyJ+93j8lbzQaYMwzuxVseJQ4I0gw
ssTgT65PigXQEktlzRndqROKBL+zSYnSh5H3gGPSDpw0cfy7xzX25T0zsi6nU+IBr0i4WWqUiag8
hbyAv3lsufFvqrhQ0X3o6i4E42byC9VcC8VlVCuvqn1JTAxL+kvoF2kDbXoWunA6KyzE4WtNYDUT
6ATGFA2eS/KHBjMkSkL+aEMDd9qLK2SeycUJ3y4iO6wL/xP8iJYNPMoBZcvSAnyYxFKfSaeRgSIz
dP9xZXMWnk0Jkv8Qm63tfOV4KZHm2de7GJHcobEz6X3brztf0QJ1BFbhNqj6L2oRf6nZrlTe1DS9
uzSVP1GlvxZGDy1AOpjUghhiC/Qcaq5uK2XFKEHPiiSIyXznDQJ/8R5SoXw2Xp+7YD8je5oLcURT
P61xluA7R/lZYXiqTz9EKUVl+Xf4Z1c5DdwBtcEAlpAoDUJPAAKzccv9CeuvvqHZTdjN+5fZ3wYn
WH3xlQ0C8d1cQaTpWOb4f2YfC7RSQ7tbZuqMoT5NmAlgjhhiT6X+9VE/7zJ6GPcHyA37UiJAqhSJ
HlWfMSQYsQv7DtwuUySNYZqNubFCyrmAedPsKjwWKttyoJY9Ke9bEHRQInD4oQXFMk9dsTlgtW+w
Z1K4zhd3NjKN9q2ogkQvhg/JdwEo1SxGMJqJ4UUhRJelS6DKGEChK6duuCeq8/Agc0zIWcoU/eFF
2CPLm3fpNoyb1DwbMDQU4bOiVsrXBt3wgM89e47x25BFaynK7AGbUDC9OfpHUYbO/mduIHag3hvQ
DscB9Jc3Yr9nFvabSguHzfmKIEkwN6yDphaIJdQ12hEr6xJsk56UEi57hCju7iOZfa8zAOC1NypD
TWjF2f0uJKozqsM09YZ+xG8bA8EAh4DAHn7krtYa6+iFE5SkhHnCtszFInnthB+drOUHGHKVZaVn
A0bEUImAslUBIX8jz4uQYbJwoECTdkfh6bnLaR7mtTDt323kBv/NadmaSMKWlQq+FxOGyZkK3BEa
P9FX0YyquhvYCsvKozq4C66KkuGF3/7U9s2ARo+orTIw+qYRq9SN5KsjMK9wjFGpiHepuAt0jPNL
ixEUsPOx1GAXYBcY6D6LIYtN5QjluQloPT9DkUTpBysl0kkA6XKR4hVbju4JPENqZB95hKBSwO24
U83wUqnfYzvCXdjGteOEt0vaBFrZKT4Omex2KDrHrgvQN7U3Fm2Da29NJQLtqj6K3d3Uw88Q7a0H
bdpFrqfntIXF/bactLKOfZ+UK48zvHSEUdLOrfBgCo1/wVql7se3cUHVv6M6AIDMVEUe8OxvaZtI
AQwbjnjEww/9cVKGAbzgPgDkr+9I2MtSjNFt1nQxo+jot1HbyH+ztisA1ziKfRdjUGF/r4Og5bVf
9eAgQpJiRWNFM7wEHsOX6mD7o/SElLNlWaJd1Y+a9kPmUGOFbCThUoFr7XayWiQcILVy4lD3fN1f
bqWNQjD9nUIBXAZBc/Df59uT4rYE6cwW3332Zy0qEtdnMo7mTkpMHwwfQAaqe+Lx/R6YMSQ5LY53
RN4cctjI8i4AHJD0zNPBzqdU9tmAy6pfy7SJy6qqhKlgK6nkFCSfuJIX4eLQ4YCO4ar3sa+tIlXi
dTuv8T8B+dHMgD8Z+LvY6WNSagwNVGSn4UcVQpTaLZyuzotXmlHwu4ZSgm1Bsp9ZH6qjs9sW2Xzw
6PT0fxjgswKGj7pccKzkt7eQbIMY1o4KX4os+4FwaRbWXdKekJbdTqJkTh43ZoKTwF1yw2Yl5fMX
3Vs1Ur7GA0qkSjZfe4tabRTukt1suG9aJhd9h4TbR2SKLLtPnMqzBN63fIyzyz3xK2OaQEQxfvOq
p4zOSjd8JONhRI5VxMscKKM9jIPvP9SA0Y/+YW93oNinozCqAp/rNQ7HSTWE1bZ8ePjKJSUL75p+
BwA1liRXwysOzE/GXuYgexWepzJx7k1QP6950GFK2hY/aeq9W1etQXY7v1APN58I2J2MsaJgRN+8
z1zNzwvKoR49fpOmU8G03yybGFUc6mzIz9nUqy9Rq2E/tNQ9sLjkPsEE51W1yE/6qVZlEkEzajPn
NlMePnJcCqNSC5BqMypmnrhiuznxx2mu0ellBCGKBStDOAxnBb5MQzXfIVsz5NP7TajB0RjPM5Ff
+0eFNCWuyJp+grX7bRMn5YAAvi2ILPGO91f77JpMhyED3p/RsVKWYCkGEgsmXuMpCbC7Ve0WxrvD
fMHf2hl0HofJCTaEMoC/3UJ2p/0dXAzmvHTZ5JiDmNC1iRWedJU6Fdj4ox0Fc6wDModXNsFiJxKx
xYDCB4Ps13pPRVvZ4LcDf7r2/ToRl0DVxvDF0+gRMPLBH1brcgovfmF7lUSNp8NcapuqYtsRdR4s
MzuzzWpbfQdtE+T0UrjKo72spVZq00tKw/n0iMM50RkNfCVjJ3kFpAP9sjLXpQ37YMWRGBjn/6KD
naMjIetaSWmPsacSitxVYWpQhR6CeW0tHjOX4B7Cd8mS2XjKmLF0jIxVB/KMAC3p1DuodpoQ/R9v
sSYol0+0ue53NKnjHW4orZg28ThZPTl2T+ZlfF6mXhYeQDjwFRMJHwZFYUEl8OKvBh0Phq4OzngT
bGhNeguDef9rI5bCMUv7feXhdpubdtbrW0XRNjE2jrpignglxg9hWIVSpobziBdUpuvVF2NWUYts
xDg6fgMjJW6iXQpT2y+3QyvzRKhAhsrwTtBTxHcOS39g8tl/5NbX7yaKlb4NH9kCngg//7/ZC/wi
S7HCIWg0HPeZu5TxJGaGPPlbEl4ajdYdWQlMG220etc9sDxrZVOC/+W1vCnpvbnzF+s71n9f1hw2
EPduElprYDlAY1XJDdl8UNzmkSlt4J5D00GxkGH5/UvdJgCq7Q3PuSv4o6JNcmaMpkJ6qb3zmo6a
NkBvUq26bQluCbP9FRG3GE0dGslcu1F57EjqdrpiR9VwIMX5MzxL5etXmN495RHoip7zal1th0EM
s04evZ+KlTgyhP4cA75TA0RjsBLDkmIHeWywVJngcqIP5c82Y2ZZB/IuVTtnWynbuwyj05AYR1FU
bzxEkr6YQvFrxzRAiYzH60jKE2IMmmR+S5rG6sODxC9QG2y9lEmFSv9bh2wZ/IXCr3S+RDfQmcrU
hXxkROWwGgWHT44BaTozVpDW8fQt916fMMo3lk8Cc+0LcbMGbbVN2n6W6e8gm8V79uPnYxwjcaMw
nfiM01dinYn/C02ssBVGi8LBbRUnSE8ND4sZOQK0scGPv8cjxf3+lmGJIlom30uikI4IyuJIvobF
a2XekuRZC0Yd2nhxMeTD/+LF5HN9kxurKb2nYdqTPDEeVWUJAx35mfizxolbzHHImBOf/TB5BUHe
dLvADEHkptQ62Kre5t9isckzeqjP5wGNNTLvIg59nUfZL9dTpXQfIIDhkDnpAgxaPsSY2ZSeyHRK
cYj0N9YJCkfEd1N49ROkWOx0C7FijHIt5gSURxqOfuHqwsjvgynPuAkVyUKFt56LW9isVlc/amPc
X7zRJYkS3P9HQ5mhI1aoUIubSSrHvfQ0014YXIcTtRXnkQfOXOyi0SCsr0w9a+H2X1fbg1nagp9e
ZGD6d4XCgZV4N+Rh6ewfk411TO5u/ULOUBrau+wk2xda5u9qVKnsZD/O2mCI/Px2B4RVdKLzHsD/
8El9sUcoDDlsa8LZdcDUrTWYnX8LfD/SGNjsac1m5L7GsbFCMPy5hDvJSVpaxmWDIQTvmqRTLSjN
mmoMPrVFUCYa6WYVJbutJePOXfEUppT8tK1w9tRAgL/9SSDUtqMX322W10nZhWJF77Yv8fFqUchg
7KGxIYVAFk82oqkTLqqOgpBUNsbsA3O+K6PEZmO3QT5R7wp9hptnINiAqd1SEZxiDiB2T/PNFfOY
e+CE9zph/GxTYGDPANegYWhG1ZI5hoLMGjvrWPG6ZQAlVRn0rNytPGFwcUwfhU5y6RRx3U4jvOQl
qV1n6CT/hOveVMVASv8r3jg02BvY2KheFUNQO/OQ8lw0kxowGZBvN+EyUY9fboPcohSKR1PMb0qY
+ba1DjJJMd4hYB91x+rOiC8rrfBCfmGRRQ2v0C8An7QvnP+E3BzOV85nzG/1FkYOjkAVGzGVyo42
ENSkm76eXyvreviiE0aQMsPa8gszmvwYs5J1j+Hafz12fgIgt9jvnUVZ25fKRZMKNEQ7mqy3czNW
wZK9I0YWynChx0vEFKCIf2Jn4457u9dU0/PxZ/Cja003fLEJyDR7ob/8HP/auW+RFcxzN8vh0792
XE1RrWxymaBCOa3Pr3LBebHCT1h98AgpIMWELZ2ejWWp49XlbzCFY2Yl95zW99+qZlhzlqJdbXPR
RxB3F7R+MU1dyKsV+8smBFFQpjhg/kWla0UaUV356/lu5048F8I0FcI1YkcYz7YJ/1G0n1Km9y8d
AQAw8VwXTZv0kMH35h4YIDv3SLcga05d/u8BXx0om9ZUxMvNjn2qACPZd2f66Tj0IflgF1nPShMG
NrtUmAYIjQ2lgv2j8hdePAJkC1Wjt0In4kDr1QmbMQVpBptdxki4UHn+D+TYVj7xdY7LwJW3aJOe
mK0tdhBn02Y2nFUn9a/qih8slZA6Ox0HVOVP6FKYGCc3vB0r+WmUNvOywZL+ZvQUV1fh5UfXVLzM
PLnIvVIPDbmjjsWdbcHABH/9IRh4umQxRu3EYtZxXAVUitXloM6FXWvvsF+77WTpd/IjcgrXu+4T
DnJ+sbp6n7YLG8bJLmq2HXqGv7AZ1j6qVTWxt7lu7JoJZqj3o6jI364PenwaqNG16kza3KvpuJUM
zQloyIV2T/NjKl7MSH7BT0WStncGaJ+y+XcST8VP8D67dtAFO5ei0r68wks5Efn7W3I7MLQa3zSc
wiViC9TDLYQLwmIaj9B3LBnjv+xiSUdjeiZemCO0tNLfvnoXrWHOyNbjTHhS2xv/1O+ryGEP2Dk6
o+4Uqg6QE1wa/4H86e3h6egAo8CZVHc3+Vw5sYySCNEoVjKLc5nss8z91GCUdSwwVaYLqgkqdMPf
GlSgSgHol/qijvEvNcBs94CH05MZZzwP4pVZ/0zvj1BuYBBClX+KZXrhrV7Nk3ERWdXMJL9XRb1A
4bfdIthd8EL8/4K/7+5UUEnWYHfbTwmhmh2AfiN9TcqPTKEdx239A8JvPScayzxGFjTFI5RZmaNF
hAVlejC8YTIMKzU4XIQRS2OatZcnKZwBOH5nNE3LpJCaE9pYEVtKMdgTwOdHYckSmY4Nwk69ETQx
7D9W+4egOd3HIRI2iKBkgvaj33nZvykIljWkszqsDPLqasPKm8rK08GiwYu5sdW5oGvnzitEAsWC
xiis9gU/dBsdZoQ+N/5dP7CaqS6IzI5tHpOuwutX7AXyTyokl5y/IYw8mgGUuGXzwbVUJZ0NUlBn
g6vqGWXDDJIasqdCs7Ll0bEECN0mBge/lfsx2w+4Z/zcqqpocJaOLi8VDsuZpl/PH8hDpma5KeVp
0+yPNpM6oerdHpN1Is6OMK9ivt5k2ef69Rt+QIREfW1bbfjdfnEuxB3fJvvwctQRMLnk+hGRgmbH
Fae/naLJ7WzKoYJdiG+GkNOCDE4pr+tbIv7nCuR7MD6rYEN4YHfHYg4kRkzN+if5uTPnNqFXEkJ3
0XbmPq6eYyU7wb2G1JyHsxpY5aSsvggURTzcMEh8/DawV7ra/YNlPvVdoImITMIMZQ9a2Bn3KYmf
/Lw3XM2WSM/6aDY8JlnzpA6xpVb0XYJywQpThB9GXPm0MbJJp+lNjgREDrYIjArQUrfN/HIbLrDZ
ZxW7oYZxXrNgi1fdJ7to2IpUjlsRIW+tMGplfwwE8mgKA0d6PP+jduQugkjr6Kyxuw6IcXS/HZc4
coE5pJBErZLCxNAp3pJBlKn+KYqZ6p1R6xUAvRugZ2kUUzCQAdWWphHC60QKKtNGM/glD4gSq3np
pZdl3SAL58p4keAT0KmjsBUq58+z1OLdLl5wsbRegLHutrj3yvgPj2Wni7L/cFIUvcWt+E/NQWeU
gr0qHOgOYAVzjhjjSMRu+2m71YLeJIOJHaZJ1G5FXP2kV16PHAwXYqYwxmh4RxPswwN2GhcLrVAG
Ua3LPz+fKf9jFvsqgx3BXpR7b6pMOUqAGcx+/ET4WslbAGm3jOL5l2bxUPzWH9ikEmvJct19g6Ay
iIM96dLkGII1RxIh/MPrhQcWWiZmBLGzmQLV2avpKqePz+7tBVo2pOyPWzy/OZqVdfg04fHtRDja
RvhM5KzUUU963p4R/Lnk/pA3lQXDm/v9VGt2wftTHIA3hjiXapyPupL72HsJyzoBVn52hBSoDXPB
6N4MwsQezitIt6J/GF5SUT91rTJGoL5rH8lAkniHTuiLLDScj4neANlTBjFVrkE0xoeSEyFqi2Bn
az20CzhEu6DueWjIp0fcR10PSSVx80rOIfe1habgu+fwOEnyo5jDLhMyVm5VFXBIYgV9EFAw6Rlt
aVCcy4HBZZbzkPGrBI2IgAG4zOgSzDkikfDynmyFv1U92Khz69bGeWnh5lvMAbBOvUL5NINhGhbf
btgrPh2Zy9c7Lc+kbNtdO9aVabdggTaOUwyL7VUURZLcvLQAg8DucY+YHWJUo2vrRrQLlKqXlfcW
fWPDGshaeyJZRaNN5W3PDX2eaxjmr+6W/xThgVy+mEqI7DV6UlfBxQeEG4XtfTa45BdCZx9XZl2T
sZ7bQmBLPGcLYpZX+xmuhCEjvlsQeCnGREsF11Xl2T4o51dsi0x/sU845PhjTPI/5JdyMlBUaqdX
UOHnNwyI9mR7+VtNrf80VVVjkTJ9QGUTh6Oxx6SmZtNZu5KjY6/R51rtAfZ8qRv5V3i5oM8ms35M
U3p7dzBU0xZkI83lhVGPq3YY6hrfVZYmdXHOTKtUlMlJYXJfc2hXVHS3vTxGDHsTjnbMyj+1FVla
fEJ/Ldr71tqIqAv623Yc+2MxWt6kw+qjD+qWYRz4hno5HJWxYPQl4J+Ymq7fK5bsf8JUgkIOWugZ
JhbIjieWlO0ezGF+sd6nw3O/ZCWkKY2SAoRrETGJ+xT0lPsXZDgXnMn02wYY4FpLkKyD3sievE3k
N6vkFt1hWuzpjktIzby3GEqXzeo2JqgMMqi0tvDVhyRPT69obfyV5BkhUfPkoNk/uddLLRxA/nTK
5XEz+C+lxECJHmtosL152R4oGdkiJBavUm96CxEvDhh2RjHcs/jVntkN1T3XMTpfB5XlAj35rP1d
ZYQfqUtX3oXFjwREiEbndoScEmOKZK0saaehh0SKiGirZTgFovCmU2PicEHzSyeSiINW8suni9uH
EV1EM8PG91lvqxLtrBtb+O4ScJa6do8bdeUVAuOKDbBzSZ3IBzV5dZYw7MNGhaSZIFv+m7IlRM1l
8ud/yjSSnt2aQNtsitL1RTBl2qjwnER5rKdJVUs23xVGenHdvvHNTSliQbIyn15tLyUHRY3lOTgz
ruZZygxWUw4pTNHe7aHAoYB22KCrQNQ1BJCXXyqzDG4wmmnnXdJk31MtP0vUmt37z416Xy270ULz
k8WQtaUag4BCxZqWTkfQbHNzk8KCsbiCslMqq2uI3rebzdJlPStBSfUz7GVLzMpqNiJOhx6u+ffC
NRd8mtlF41fZCMzMBV6jk297HztLoXejDzfYKQduaKaJqm7X3Dj2nLspaVmsGerZ8KUsTueNmn2B
8Pa6ZdgDN7LE1OYy1oPxyoJyd2R/3UernO3wANcLgxPj+vpiILhBSUJNvxgOqNBi1UP824eUNiUd
EFqgyX+jxZZ1IWG2Nq76pbf/tP/t1dZgxmrjBd+wnY8Jw1L1uYj/9Eif2cIdeFrIRWT8AYpsM0Fj
fNQr70fBjr3eNA79i+Vgh4SEouRNFzPu+JnmOZoCWhNpsRSEY4d+mOKV2eB/fyQ5BuVsojEGd2NP
vw5Wp4BDw5rQ/5gljjNe4yDXEpLRZjpr6MwJbjGWA7YrBRDHKgM8pj4BsqJvXXIo8hddLDAJP2BN
TX8XS+g8fTXxnmTcQJ/LQUtB1eMWjvyGLqglwdhF1t//vckfz8bLouqL/ZvK86OyvRJRugIwA69B
auWZzN53f+ShIbFzRYhBtDEZ0//mNkgOKcxduN51WWBIlrtQyuOCnOTeHCwWeEEevOTO6qJVayqT
rPr40Kt9YSA7MUjGR62n3MNehSP9FOEEzdRmMcnmjVk0N6FgOewZjH+uhCvqaCODC4AaWCvosGIe
N1cVUR8/0RFhaFYoNGLjSi+0nVJ0CU9NFBLQoIO2trBEJpOAlcEdH6oT48s5KVtHbVI3phFA/C3k
KoUJvdR5Sj+F/2i8Xpmg/IbhP70OZg+wHRcQ2jyAU7Vc+UmYzRlnn8HsmCdREpNre/bKlncZ0God
UKaJCbHRHcn1M7Xz7ftgOchpn+X3/bpjtSSDCFy0C1C5oUifpJfGzrwNHd0POsdVRPZ1Aun437iF
f7hsRp+7O3z7V3wPAjoun/V0rciW7+zwk5qBJAC8FoLSqpUPOdcZ/3wqunbPIAOyFrjsGZFtV3Rv
rY4teNUrOVu1pf4JHV8G2lQX42fMtLLecRYeL4Y0koWBF27n+8DY98WvmiYE7xqSLzNU34SMgnLj
vne0vlCLk0T5EN1oRVsYk2xgPagljft9HiAkuzlPX8jhABIxazSCY0SemBNfU31AhHsI8nHkEcN+
+19hDbgBuYGlNzjOmkyr/W+SC61UWhKsoJt6AsnAs3M6nXiJcMKAXwL2SIKRQolhnfCq7E6dlAKV
Sq1hh6RjQSo1Q5GfiMq49uDsrSjk8Y996X4aahzppdzR1aIHNG2jZdhQi7e0Egt+zjaMLEtTcuLm
heBqiBGS+b2ieGykHagsImW9tJFP873WaG6lkVYraBIXRZMzlOEgbjy2/U80hkhd9kMOfEH+L3xa
E7BPv8AKBAnyIP1tkP+MNRNqoD13VNUD0KGQv7RflNvnvZNP4f0STMmJgfIcRBXWDVntEAroXBaY
VDpR/S5n7Vmj74x4/BvaahCEeqtvUeJhePW0TpViizJ6hXxkCzoQwgYK0D3qm3lhrP0w4QNxQCJ1
dh4HN3XCoAvKHQxqys3CtTQBIQV7gmDeFLVMkYlTsPNcpNMzm6RTryjq5AMd0HOJF6Va6l6x6uN6
M3ixsFszu9DjbzIsFtKrMwJRyMBKl696MwHF73HvGN18C368FOG+8tY++B+M3ybWyJHqBAVm54IX
V7+UWxN14Q/vp1hEh+VyHWBTrnvTOVqhGluAfi9CSxEE/Md5OkAqZ3MUePBk7eYOLG0t/KIq5O1D
p42MwjrxNCc2Iiflvp+0yIdh1AW7mxAvV5Nfy+hlI1TOlksYU0X+ViM58o7CT9fxWSYhyWONxFRv
UOINM75iAq+loKFs0/rSXPakXLES+LpUu3FFoQvWOduUgiLKeuixN3Vg+R5vgBBIDeItTAXTprgU
LqHAg1U3t4pFTwdx1Kh7Ovycc5XUf94kCkANzdF6AND864iOnnCQ6PJhKEDT5HcL2OW6QW87+uMg
r5nWNQQxLDvmOvmqGI8Pi/tpMKmVV4Xh/MrE3IxhySserBZ0sst4OScUOsj4C4OaztW9a1ukOGcx
IFA1YbDnX26o7lSEB/0sftOkYxAKZvDqpUNNPhDAi1T7YacHHj4l2HWAeLwfTy3AMy02ebhGGObJ
Sr97+3mxyDhgAfS2287PbaK4s1Qe7rw6HIgBgxzBR1QBZXtb4ZarXKNePlJlHe12/OfWDoys768u
mn2wse9rlFiCfyyRX36zQk3P27TAiWfKgk59sBlBKUmXa/tNg+ib4AJeRekEgU7/V2EzoZy1Idjp
nTjSH1qioAnKF2Xdo6E95hn/KZPoG9SKbBLnXmD4QF1WquKmlxtAFDDGIY78RzxxbPiC+VJkkHzn
7LHtZqmWxQUXGN1ul4DDmVR6K7rA3nTRtT2VrFidiUqFyP01NBK70g0nDm6s8y9CnQJIbtdOJvF3
d7L6vhC+TekUnkY3s9FPEr2hw+IhRgqazpe3N2cwBcuibFvPRlsaoa5F+BDH/wcDvVjsoBuvld77
hMQ/IyhcfZ8thKUpGj/wIHghQJEGpKEJSBfh7EKiuvfhlPqHB29dM/ATWlLwYtdtmzkUHeu1YilP
2ldGeMGAqGRvB9OVLIjN+HGkrekPjGh/HxJT2xYIKpwZM75q9VFEBNOkPATnyKfp65fqtJD6AbED
4rWgvfzkHc2zZqpweF81Nr6gNrxo0y7fQq4C9UOqfECrvfc4vqAoCJuRIdapeLXY0yEthlm+q4be
icDUbBxkoV+hhBeKvdaWss2ZmeOGYblPMx2mA9anpM0Z0CZV2xt06lOXmzH8dU9rIB1ducNombNY
yrxqkzEy3mJbPcQ0cejV2+3iP05S3agdDbMVIjG+6W55GBXHQEmiYw9W3isyevquas5Iniq4LDkG
WTSYsmjm0G26QTv7r0yyfon0Dj0plRiSy/BAoqTVdfljaK81F2rYEdCOdyxYCzB2UO2jJI/IoD5r
mBnuapBvGAkM9B/IiRnfIXZ5BlGXlzcZYr3czuNKugV2CQY+t58yFZ/BDDkQg8zK4IrtbPyGb7Vv
NomvXfGBvnNKsGdcnbe+yUIg5ESiZwXveJKjyzX5wUUSAiq0BGxDWIVG7LsEaUEq2rNsmynaFNUk
7ibyn19UVwG2remFhXYo+w0+T4gfo3ifEnq7g+agr1wc/SxYdqt5/Xq383t1XdsQTAXpmycyx7OQ
+0aTxisDLBsM472BFyPumV+P5GYgoaIArwps/LNWjfGptl39IyqMfTIXzKnpoivyNQUnfrM8aHab
j8fjMgNlcVZ/dtkRebGSkTovtlJ5Jzkgovs0YPKrpRdxEH7qVZoogdOr9EDiK1gqyYthQr7+9Ipt
Mv5ZDbjiUIQUtv5art8G6rNUlrNgwIxoi3GjInuyiDcpYXQMfIt1kXRmPJivNXiqyFXqb/p9HwYn
0+KHHgmwKFMU2G1hQliAnxwKlveSKd81SnQJulIxzRzmKrdloaCbzLPPv5ccXoB2UsCRx0lBaBfi
bWC5cnP3N7q6cEyWsoSFGRPr63unF1gz7QRpBJX9puYs6uc52FcNz12xKZkuxJyrl5X1m8jaWKN4
NxTSJHzzkTqzCqmgsjpocT7Qho0WO7/UOGehaYJ4B5SgWJ1NK2Aeijcb9FFG/jsLh6y+GmReFWqE
9UruvBGdcPCTxETw/CpfcgkvSaSJGDQgrS6fT6s05wPkHLCdLlYURbduHnb0xhs1vvkwiRBR4Ity
yFNSMFnKdltwCgxIOV0PK2ihu0VFMcpOvvuXq6I8mDTh7byy0ll6RcTt1u+/JTensh4n8nkEOOjW
Uaml7nrCuGRhumPVHM3Py3EY/dlsBfwX6euHqPNFsZyDKaSepsoLej9sR5XU34vVgzTNMZiueB+4
PCPWxc+6zS++d13N18hZBrME74G+OlbdFMPyaUhibCMx9yLo+QT0Liz51j/LbdecXN2qJBdvMPJC
9sfKg9jAhbiHpPZteTFt2nJiAoBIfk0AUacKNb3ciRnq7dqNZPmpwXksTwhGZuWJQ3revk8Hp9a8
wbUoMZxL3c4ayJp415ZERNNB7KIC/BnLy3YhYvC+4OCIDUyb5CO9KK3TXvY7nZqnBhxNec1TcyNF
p6Vb0+x/exa9mJq1O5ZP/u794h+NMCGcSN2hp1NBrWMhDNMn203329BK/eFz64payyxnFk2DdA5t
4ZeBAAgI577Dl0iLL9bF5mxBS3PpqcfO2Ov7T9FBtDthaJ1R8icoytBJQIGktVcaAS5dMOMQCrZG
HFKCcRvb32aShFil4d+pvErYF4xKnJf8+2H3t5WwCEq2WYY08UU9LatEQauD4ew0kuv5W/8pkCkL
KIVnJW79u7AB8fuQHvECyBvtD83CyY5GeakKYZTgAs9upZMaKirUsB6O4TzFgbWj4+HO26UHJGru
V5ZOF3r0EUD4Da4d1g/XHM+NQ+jPcjOcNy8N8f8FkDbaT+zmbTv0KawFy5sndp4q5d/ZZDTMNVJm
kD8+zfWszxyWpCwm2wnADVT2Ax+Ucr4mOdorvNnKcLbrV7Scb8k96qsmoNODBnWBglcR5C6b1aEo
/axTW6ISEDrNLUyU5/dAMzjyxU6uhe1BTJ+fmrnQpWsAGc5F6FlH5LF2apcQj47VOOl7YPdPkbIJ
G7FLSGZfRaozF+NqYyHtnch0230U2u0TQc+OQlhhCTUXdPxdQBHJ1yOfDjq2KRVWHLmKk57W7QHp
qrZzuEsLHz4yZp1XAXTV0r7Oyzdk1VkjpQCUAgOz+gs8BBgzdSTkPjrAS9YdAgMUDJES2NCai/P5
nhm9uOVygEM0rbeOdoj2u2dj7SUtyyYsTRt5OSOC7fwooH87WXFmVYRq2veup1oDkaXIv6EK3dny
nYploAYThE8VWIw9kiHANlEuMDdmLMkCyblsoOMvVEHyExkP5pQWFdehwX23IzfkIvHYIQH7Ia+U
3nwh6uZ8Wi5+xyX+v3INUSevAACW1SQNV4h6vXWcTWrvTQhlAeHdQjMlZ6BP6lTqRIfYwINjflCv
BlvAmyWrt1B7E22JWy/+uGHI2BJnxSzIvryYvzMe0k6ASMN3+4GNTMaR0KM0YEP1fQzwjZGVIrNk
f7wCxCnBLXR6oxkde3hxetYcUpCYQ4wRv5Sb8Hr2vDMhicUmcPzAI6BV9IFXHsuGxbn/ID47j0l0
9nLQE/MOCUCFA1aI6ofI8R6mxWmmtBnies9rLxx7qj9hglWb5xwBDgMhKjWaqlT8AlasSg7al8s5
Z6eIMhYT/NnfNmI3i7R1tGcEG5ddaeBPWfiXdhJFZatwQv/Kd9C1pSDjdQT1QP6T/oeIxf5tUiRb
p5PkotOIFOE42f+JzP15q3rp2kz6lPKdz5YDu+UpPp5Ik+Y1Ibde67gedHtzhyH28s3jnUD1Yhud
ab3Oxq3gG2ogMRGLXOwn5mwEMRQ61rT46/V0vD0GmIcSuZue07+Oj20JRQLkFcJcC6dpnPqy3Eb2
hxPwOMPB1Anw+HoRYA2AaHkfvBS8r52T8Ttd7XDNUgxexPMexB2eAdj+uGlkoiYlIgjZwzYVjdeh
FOrbYjJRPYbmKF8w+O/vb9bcW9vYSmR5xR/FM3tzHCSe3KyCPmB++mHEx/nxPVUdhz5LN+48IIz4
gWdsJEVXdyTNcYTMbxEce7W2VXw1nv3z7bLimVmM7I7uxb7lPzBLMWsR8XB3bV/KeFbCV6JHYhGF
rsp4bG8t1fYNu9Wjs1vuabfWxc7USRsNwnv5Cu1JN2T+/Er8qqkf+XrWN/7TBFcSNDdWvAB8KqbE
J/3OC1ypSAVeVMiDqxnLRvCJYOliYZE8L0vh4Cf5W/H/0HfGENoJhFuyyvyiEGywOFN11OJXgLU6
RfKoPAcL0Ap3qiJUvgaidpdp5x/2ZNYdRiMKed0riSJkfrx60SzzTwzfnOhFti6SzWZ840Jr9jl9
5Tr7+/odT9u1RW6G0/+CI6gJEbck9Ht1rr5ZiAVS7eIsQsFML+wPdGzGNZoAEG3CU6AJMXS7bRLO
2ro0PHIy9oKIkdHVgEUJ8OblJJyeYnPiN4uvH4m7Lfim4lmN4Vg8Ycxd4MgC6RlZpcHGRFmF0YFt
SWnjlVhl48sY7Q+rUKFpc/MgpvyIood2H30fnHm1ukQSTb271qe70oLnIHLCikNb3DmIKBY69rOE
FUHwF+qUPx70KY3ZcUgwPNyp+i88mAe47dI4gDRqiULey6lLSCjhXFFggikvTVuMyI2a1fdQ5HJC
K9YUHlGzTsidrREySW17pqSVkJjvKacYRw0E6/eJYIoz2avvWEKMvUVg+bydSvdGZqZQD35q106P
7T3iYUkEmQJcfqp57HUllB4csKGylhrmn6imu/e5ixIAMWUWo8QlGYWaXbcXv5hSw+Xu7NYdtk7/
0AnRGSlkR7pM3IWVAUGWE2KmU9H9sOm0FULAQ29/TiDt75YRtD2DOkqsqlkQYvIQ7ktCXNVPF0g9
BeoKejeYWiGbzVTaNTzTRzyFnaiocgV889tq6X6zZ5jRDYSnooK66w/cy63wGrbFOYY7wOINZQv3
kNp37K0z3tmJv/A79u09EvsnVAC52IgKoQKWUt9TsN0h7cjehxle1oY1hhEG0ZweRf3G7klMkW0L
zUaN0LBvTgx6MElZljctAanAoHoIgZ9g62S/RVzatrJ613bo269pfGMqoOYW92CVaiX1G5QN0KFt
y1Q493sWVq9j+3uFUXZw/FbkXWBHmWFxk6/rQD1MFSVAqGygJDd16CVIpfx8UPxyOBFse1r5ZD9G
9/kj0VLeAqBYDQDsFwOUv9280qn0qTbvL5z3Im9AtUMuTYsVP++kFGNXwIFw37MCoh9YbfLri+6g
nHelNHeV0OEaTnL3lHkwws+B2bFMR7oRXPogQcejhYwQDf7xrWq/E97LkVH5xFJBJSC0dEi1Le/r
GMnU2sQuiiid6BdY0iXYOI6Yr2l+da573irO6VZSUxY32zuOh8BfinxOaVA9sxyYRHry34Mia7LF
pc1eVJU1q5N3eZjLtPpOmhgLFiMyxLaCrIwelp/ALYlOJpTJb0lHPu+dcUBl+7VCJfJBiN5iqaXQ
G1k7NlUUfhncU1+uSvN9i6eXBnLtzPqe7LoMEU4QyDVuta6W1CrA6R9yYJNQp8ycPDmPQyiQxhr+
hsX+W2wrDjL9KzUH7hBb3w9Ja4a/TJSE974jh47zADNi3QK3pm4BYnOkhc/0ig4ZQVPByQRpECFF
fRJq103IdiuLVNCjX1hiF6b2BUJcQUEnh6+rKG68TOWXAiXaMgVyG+6rgVo/Oj/Bv2qWSES9DEQY
A820+dT16GY8tsus8Apae8NhrsPGvJWhOuxopYnFNrVHwK4gBPrEp7QSF6ygPLqs1AQY9vqlknVO
G+ZxMdiZ5nFMmFwIIYgO6yYQLj5FmO4mc3ZLS9rtTl57LeBYOZX/P5RQIoqvurRrwnRqOSpK2wdC
fKvUeQH3QxP4BwO35VzyTvEzgoCnHO4GmnLCi30BOWWU8XKJuAxM/MbrspnYFMPZKxp15kR44dY+
JwVnW2N2SFBMAcM7R5EQsGSzhH+mCmK3J/WqTU7QX1szGpAhM+e8XyAZcug+13uV11/HhkKGOdTI
P5ziqwnVEEUYmSOiuP2By22pMkukDuC4wTqCOHQc5xu73onHMLIs2vUdx+ttfKtWakCcrF/yU04R
+r/5zW2BB460OKnr4qOj8h+znc9bebaKl1NjobTLRhnOpdz853V77b0YCDFA6CWJbcPv+WzW1wHf
GIaYyI3UX+4qEGCmr1NIcRybuBNolmGmO3Ppt3wQU7KQ/miU1/uwwtAUdaNKw5E/6yLFGJlkq/Ja
KdomtmxQCVqFiD8WOIa/tAlw4vURfrSfYhr5yxlTKb7GsHPy2gYiHsREa1l6PnVF4xZmF9WSDMYQ
sHMgPNOC4lZbJ97a3wXIR5mqNPiGly2qVX6WOpiyRD3dnNMzFLlJvJfspJcXtVNmcOfa90UbhQhc
L0ZymzQxKGZLXY6dhp+IvvjkRx8Pawo5/TnRf6xAcz7fAd90lsUmrXyhl6u8VWB8kHczt6Z8v1vp
WpWMKTXGjDDaht+ikIo8I45pcPJX3Tr0rrNpzxF88hodg40ohe3yqPmYVMnqSKNHbplEdJONyOsm
8n5x3+69fBFACzDltOJlrkkLr/198xgb3Gs36QzsqRIVrms80+cJ55k6QRDH3y+lafGRB/6dQ9ZG
r/MEBSxfsw1nv1qEnUoqhJ4g9YYpXE84Yur0OJZmLn9Lb2UV4vWUl3nOdnXL3XGutO/4RJb5al6i
afDv2mFHpojt3rKAwkXgPMGd3PcsJQ6okAvK0ejGCDPvJur04oLXcdS2jUuQHOFpzDPVMurWazAH
D43Z0WSxoLI3IgW+HR43AG4xq8hiIFjW4zhaxtc+YpFMdaFamxYCoXerUc0bU6TpdeFM5rjN8OPU
D1w8Vmndk0AJLGHAFkYyF95U69J/f+QdYyyBBilDAienIkEW7oI+xJPAkRcs11NM8an4PM9i8kET
iHH9QTfziTlDLA+09fH5VGCU5z7Gmulj6AOdgPMU3ZiL5RTCNF5vB4bsxKK5wz/n3av62Gu215T6
XGmsXrB1DZizqDt1glaty2IKX6zcxZHSNmbHoLm0Dgy7XDh/jzcp94U2w/jLWQ8wNkwMtZjdMtxE
JlAK8QLaM5RNMzNMi5mbB+oCnw9GR/80DEYJZrGlndRSg1h1fI6ajs7sWstDTmA5L/B2oeCe8CTy
CCrYqDYxbFwz7AVlQcvEfOzs1S3TRkAGd/y0FJMTezZOLvgp5ExgU0YYnYlxI89nXwxYMHwZS66o
+C/B+cc8oqXVW8/WixMOqpw1cxt/f6QlEZjJoUQwRpBLFUy2NQDNav3Er6cSIfGD8OqhyZZ/lMQz
65jf8zpfhqgPOblOe5SXAsSaHH5Wv5uMSJio554nAPDOika9kLdixspCfco5Vc1UrkG8+ZdPA60B
8WuffmZNYhX7yuEA26gVEzFfjCArggPXO4GR22UjgUNSse8fD2SujiTpKUJCmYUR1AMuT10hvrIe
aT/Q3MB0E5jXXdaVXiRnvUtfczPuA3/mlCpYjrlW49dUMAcY8ulp0uFzYp9XIJtwCSizTEeAoYEG
5lTzvtAPiSMVkYw9NlnCvfiWQX16toIW+aa0E8z/CuyiJxp+Crb/AMEm7Y5jy7+BId9E3W5jGmHM
TniVLTTI3kHR8jJyiq+R06LWts5UPUrbToHlv43p2mSEuO+l6piH3fLSvA0Wf+Wyi7ax0h7MkDgq
o3KB2VzAGOTx/O5iO2oaGF5Y1WkFA8lBNvavabFI4rwjz6sgxQJOCdKtQcH2FHDGTrpPlzHPjA9p
XMa0dWLk1uUH01BjD/7qdQF7lKJBHli5ICJ/ffuQcUe79c57F1nJBxU887JPVY8xgFtyfjcnGo79
CoS0FwxHkYlocOj2Y+Mz44XQ0wqoEy84AAV1G85Mp0S0aAbrs8nLWi+Ns/xhaqb7LjfsXAQNx2xZ
yVBVii4d2FDIewqHFLVcXgTKB3VpCYjhlDT7hQs2TNBeW4ZrMBS3URg4OnsjexVxT3/qGsalKHlP
pmO2WjfVOfzn64Y5AbTN97v2RxCmxpbOcOnjnYK91S3VqlEw52lRiYytX8uBWgr7SoYltLu1axJ1
LFU7EdXBLza5i446hayBnp4bntUH+O7uG8lVXZa48h776IJQ+dVhmJdGJW/be7U+8Cpvl04hcDql
DLicm6RHkFJ7Yco5oI0g3tPwwXDA2cmAKBYxb7DtNqBpdJj3UqEYiV+GtyjdzZ8Hg6EbBHZXkbck
HORzEZAXeXiqzXy2iFDE0s3+vYEeCGML8klCVoK30sBwIgLRXm0QGtpePvEXEfFFSfjyTmoe8FMA
MFR93aWTrzA+q32GS9w2N8Wi8yDzXKCLZszKjlKHLaga4xGvBHbGqcmdIDr2r0waCDMjV5AfArWv
BojvKIwc9eNhUcJRX9HY3FXtv+L7BLxxYsb3r/wlpGQDWupCRPIgI4ggI3AvGC3WjaEq7HFRwkYf
jHTbY9fR4XFZBb8+YcMpB02RE1rxEL711gLT9xrumjf9gjwUGsml15SUR6ajhMqJCabcUR7JCN2I
f5rTa1bV1N6yqcdqbtCOePD5NRQvnQD+FABa/z8Gg+GQEMj+GhcVrYMbZ7kQFqu+50tyjGWLCFw3
ATnuVQ4WyfzgVYuZZyIxh01sP5i3DnC31txxABPLSdc4t17ikXS+JfaZoGKhEqiGwh2pPOVqK/Na
w/3KQb+629G7bC7sOdYwJAlCvCfliXTZwzo2YLZUjz0sZUCYYSI9f6GZXYPik0UMw7GrUDN6ckag
8SqbF+CmCofgzdNqCiAiq0Dsg2FLgjOPEOL23q0PA0b6ogDFLwooi2X3dsFKdXoVZqDCPTUlndib
mfbEt3sGKvVy7vE1v9HptuN16VxavJz6COu63G01kAg0Ocq+WjjxgJSdPZkS4ypo6776VTr+6FB8
IV6q2KUl5roO/6IsbedXE6he9F/5qleOUkonaX9fM1u789jpGSHBqS/RIljLYXa98OhNtlw5RoAI
IhPCtUPTas5roZpz0q4ywUSTi+dyMgph1hcJR33ySrayx/TuEkUWz3qqzFrcClJc7H4Ca5lnK6Ox
zr2tFVBeAe1nRNGvN+rQMBvtzng1ERhUMQ7fIA6gu6RWBRDZWgEZpuSZZEOiaEeqne158GO1ZVIV
/ojQJwrPSPtX39xHhHJ+fhfFS03M2OPxeLSFJLwza4N7mPnWdSplsxwVaCmNGQluBAS/hnzXpr4B
6xz0HL4jME1TX0Z+U7kxz9Yqw6nAiqQRmTlfg/oE6dm7qaVX+EXc25UGDk0/BaFt7VLu3YBuM0u6
8btk+EaQUDpyCPfDjqd1Hh+YfD+mP8pa/owQ+ISl9h5J5v5GXOMD9CLyVoiuUfYThRdOptirUTNi
Yomh+xUjU9IEtUNhHqr4WF6D/auaWl/d19tKebt0qtKiH8WXctfQJIxJzU7QXDhakWE/HgLKn9uB
zV+c3y9RJWmtQPRCCFGHCHk4DMiMiKmCN4FfFm7+qF0ibZy3iWbOKKSv0tqEo8gr6Uczglq1dl5/
L2BiNUL8gPhkkUxoIsi8bHO2urXVzg7F4CXS1n9rJv7Yc1xGQyv0U3NsnZoBJpFp1QjCQwXTSrqf
LNwwv0FWmqfZUc6RxuYEHtp4qVSwaOXjUQxY6jOyzZxg2/05ulHw7LUkyczpdq7kuN4JPxHwCLb2
6Yk5Ql5Q5agPwCX6jCyyDBccQvay3pW4RtySd5XDJcrRpSguT4Yxr9598ArikmSViYzFGxCMUwx3
NUG7lkAoAn+nJgvkT+N4k8rBePxhA8quPFQdggkmrGoWxzJYdLV9pwM4Wjn0fc3m2uzlOupAPEoz
VvAC1SkeHtSOqxNeUfVYeR/ACn/YHpAqmxr1dQ8h+4iLb4CzeyWtUoxTAZLpzNUIELQhvhy0kUFh
HCS0THz8DZXeD4ltU/R6J1JwWZm2jivlg7ug1tfuZvoKfOp3wXOYY5ktcSoJ/eAAEDXxeBqdJErB
tnelLTopQDFd9Tc7cDkiEw7XhuEImmXEQRxmVuCJ0Yt1q710Y/uozAY3WyW0Ws+eQ0AfmRyoPHkI
SCYwzmuH51weIlsYUpFhOg5tspvrgPjKSAP4qArnx2BZAq9FNN87Tga+S6mw/OiyHNqkXJLyv0HU
czjItf00NZA+ZnV6rkwGrxjt5RtjGSuHihgMctYLKApxse7v2zJdo6mo0xS4agZlZu3Q4zly0SXe
mbIA6JWFsyJ4GijrAzgDxr0l22sDgRisCEdtretJU4erckfi4E519eKScsFPZqi0c4xIzNP3YCrQ
4z11tbPIR18IRVmGDy8wcdjt5TSLPFju5O6D0tEhuip+FpfYsZJepXVtqpA2FtH2tSs4NPfTdrIg
fr73fzNcTjHHQ67GGrhTA5TBScW1Lsk/psvrP9ZOQvWjeGqCOTNWaFGQ6aBC3tEsFj+HIsNAyeJA
ysDHZ3iTV2XPzw+FOozyHiX5VaGP0JStRPp7BR4WXWP24HYPzSnAwnbbk1jJxb9830J5l1mLAWWB
/xGM5J9qVjZmCfiyHfT/btGU1WBTL/ZzNBd8Dmn9ypmUhZiv8TdMyCulLp183ulp28vfiY9NNfDq
VayN9qDUb09HDrvj79qwkwXozzkQ5m5jplxSUACmD52Xftn+Ci+5ECMl30+Yj54NCRp7sDnT/ZxE
scVzktsftbM23UmHNVKwxIASixzf+8yViVHP7jhs5hUEIyjGJTUC5E/YgIabS+u1L9QfTJaOHWJB
dom2ndRYgoFU45NZ04Q3lPhoG+VfXJGp3yMfEC1DH0Ug1r2UtXf93xkJbZ69ubItLTfF+gpSgvYE
X34eBCqxjZpXTPVaudywxV2eCfCGhi7lwf4d1s74V0FxnFwpnwZA0jhKGQ+GuGFG8wknMSimKBT5
aHQWD7U4Ea85DwwvX4Ue7A6aiTGC8EuIbbS/6nybAx417s41aaJxgAqknESTkrezFeSsfkQ7uZie
wXOfjjLck3JTa9h13jeM7oAuvJR7WHuzpORcIqIEYmEoAarvou+jFQ4PnPcNb7Ub45nuTUMn6eqD
gwq4tKfPEQzVLGFe2cjEyazlSkn0VB8vSDiwOK2gredkX2bEW4E53TWk9n1G4yq3+VnAkz84DmFL
BrZEy2931jduxUvNfR2BowzQgF+smPyE6HneR6wFR/p+CCul2pLvI160pnPLajx3m5euLpzUjac4
dlRWCvyqgF1s0m/cqXaOf7shjeh3RruqS8yrQzHVN6EmIrndEQ925UYzLZJz2sDcXuNAcUJ7U5OD
CiATE1B8wMO6liqba+Oy+tAYAUuil7JjsUaPWI5eyxYAbrPT9SFs8IqbQLL4mvZB+cJdx/kh9RPk
qSPd0wD3WusCbbhLa3ExM/fUgQGhhq4G358Pq/71SqtBB8ORpClUnnOsuSEgyADXnAbJkkLGfn08
wgbONPhTYyjB07H7wj4+ZYU1s3TAEkwJzWHylctL3PAG8YNozzdZjRzmkyrv9tZ55L4aVYLNITpN
D8bCpEQQqBpS6sXgdCA+Rgbmt2PZbGiA+1fYIVoEUExKkSmyxxyl3+tFR3c2Bf8tnUR8m8USK2KI
dxUfwALAd094DeWEAQrpDLLqcutn5L0p/cZkWZ9blGpAJxg42yXnordVGOHH5H2WuXIwS4i+eQw/
G+6IL3HwYR0E3JGBzw7gH6NyZDsF4P+wmxKxQQK7G9L+MJKKFTadsbdEuVMpX1gInn6x/EEMDZTl
UXe9d6ogNY1g7QQQK0kgE96lh6I8PVSbIZduVf2/MK0HTywVeEbvyZCgoZn48oz/n6X/4QdeBKEU
cJwcvgpeW/+GiKx31+IqJzw0oDDUB9KSk3kYf3ry1E0RX+XE7lu8qhje0ZUOEpjwNEjlki3ZHqtp
/oHV+HiltWX+bXtTpMcG1iwmxzEYFkDXU3GH9IbdZ4Nl0LQ9PAYZj+P5zumR3vYsh1YhpY0WQ0w1
p8MayLLE3UdaD1kWDxjclNuyv9aRKRzGVZxs0Zuf4JMLGiauRgHKmb1AZp6imqSLpxn/BD4daFOv
uGT3PHZDLK725B3uTr5GHwBX0rE63DBdDAqScM5S6PW14H5qFpJLys4OII20vQDHujMSi5thmFFA
uvByNab8/iXo8+nvPmdYh8RRiEkfYo2WI/3xU1CG6qwVVQygi+KvrwrLj6eX4JiJUn352w5As6Bh
h18iLBc8xKZty1W8z80f8mFTLzBEtm4/h+GYdDRmPxE4DhkGPH847tsIxAh0FiPlmwcOqBFVlInl
vyTtlq9uFMOqysSY742Pqnj4ddN9S+yaBeBk9Y2bsGBLomC2q6RDYuGnYeYdvca1o7HA1k6OuqWy
5eTAR/c48VVCV6+d8bhL0Ns5k8xWAvZedRDXlKNsQfBm51uczoWFzlhiU/Z6Z8gl1G6sag6EUfUU
oEN2hjqICnMvzw0RzXjwcDskedpUC70YcmzzfaiaJxBddlcwKoGLXTxmvlG0b+w1fTECtkqhavX4
/2OzRxnnhd7Uc/b7YJVeMUjfaHeSf+CnW7dIyOey1EYJ5zPBByNtPl+Rt7di+XwdVUZRS17qsBjC
4GhlPPmuHGm2Ijm6N57g2yuy8KUOy7yqnwtDDIOXOHkq9B16Q726Tjm84mTpAz7Bz27sMh1LV2kS
LSkFQ3nsb26cF2IWPuOUGpJulTG411xqPUKFX4VY/WasaV0Tzk37HRhkjNtRHEY3Bj/YIG+lF3de
d8y/VEgERQ9IYXm/stEpC8RsCFyBvM4/W2yhx0ysgSOFLMcBXL8ptrgvb2nu+h9SBSM3rGaVX3R4
o2/eZy31ol75quSlLVKgUywd29XYZzQdGJBLAKZ5e+UYQ8lziYoUfwTVh+HpyPaKp/pmS45KQjrQ
TQ6ylkRCdpnCkr3UpQtN+ZAydJ3KgSMSQPvIacH9KOdsB3bqWEuZQd305Mqd34CYkX9hLaMgBKO7
2x9Pv70Cr82OqsrORRZvexbCFof9YwLVCk/0ARXQOuRXQFciKNJKZxcSUUH82y/HDW4U4a9fJEg/
KZIkMeqe8Vk21fCHXj5a84BdX67UZXhOW+cZV342x8Pi7BoA4eM3R3qrv9PllSFqvL8k+Qx8T+tS
w8MLUUPeZKZ2qq2hPEfoz/78YsScjnkvYXY5Vd0aMvbP8QvshJDm4CvAqBv3GBKY+WVNG/tJf+8L
0upr6bRio71XQOHkuMf48kTqrBrR8xVtXJTNu91k3WqtwYl2hCPiFuBQLku2e1waYA6KlPioHHZp
cabjSPksuzp9BaEHEuRn17dW1r/prO1dFaW2vUV1ulpnxddBWIG1zgwX5/uP4DI7nt/UH2k6VIfO
jo0POZI+a2Xup1slKk829cXEWCes//srAOYIBK0yZnJSUYiD9s7psJsUswAFspAd+s1N0gLsCLC4
006v5smQfwB2yh8tgr8L79foJa5mFR5+Ep3agiaORc08VqJB0ftSyDYPedq4ij2voeR+vXHmLyas
Qw0rZwxdLuDKe4W3fj6qxJ4lCJt2jNpI8VV7U2KYdKtDcRvw6xBzAslrX/tbcawc8rAmNNdzyHEp
LLzioNaBqle1FmXuCl07D5oQ+Uzvl5W4Pzv/3ooEDKEJRKsoMnFLU8qtNs5XlZO0TMAGaLyrmfb2
/Lvw3NZFs8/iqi6r/E0c3uo5f0wW0dSIh1332IkoEzc1LiUkITPPmxyRC/kv+u+77KrzGXdl40Yi
1w528yMa2Y74uIF5vSDI1iPLHolu5QNJbhEzywAl5t1ElgFztjKwhKgFd5ToZ1XAE39BtVDeH0Lx
Iu4gOPfXSLExpkxFRK6akz+ZlMCqvUv5Xe62OAesYSSIVqeAXyRv/jZtxhUBPinH4pcSjN2t/A8G
Oyiha7iz6ynbj/M/WcnMSuvMXw2bfw77VuVPrIBkYn3EqkUoZUSh3m2NyFwcZ/Lu5VN2bUN0DQQS
taqAJJcysiWI6XnxIPEN7lwCQjChDSMSO5jwQfXdf2ZroBmE1STNBOVfPD9oZjRWCgOjqDXk7wLu
9u/wXIt4SpMjUaMY9UIfRZ9Fq+f8YPvXvc/NlZJGR3dQckyYjaOUUFFEWAvRQR1kI4Ks5UtlE8ji
iQKixtFgQticBdPrEWNdXwltUyAUzdqe/EBVAfgZVwGnZvQOf844v89AT+W4RPihl8rURzLBGzWT
qmYYrG+i2IgUXqOI4Wz4j5970UAlvXzGpEmABXlkE7Q9V1gkLGSjA0Q215Anmk/vzOoFyf4k91LL
f3kdHCmzrAem3f/FtvkhSFh25NedbZteNk9vPHv4XIsfLGjrAGU37+VQHn6lDG5M+f5Oynn8ZWsN
Ge5U33bM0NIMirQw9KARzucAc8cUlubMVVhIGQl8KkHJVjzqRIDKqr1OkKNoDb3xLxpF9tFmIwaK
Zc/Vxdapi9S5n2XJIf1W+MUr0hjwOPBMycataryvNcu1iOfglBdPkYJfqlNKQIRNKI2qJoReqGlU
dYxWmzhrjvR+Qr5a88C89J6DBkr9G8GXhLL1gGSWq2ALVYKFvWGrcQx7P0Xpwyigq2m8NehWHcTL
KtZfKBTJ917xn5+jnYYZ1pYg5+HiowGWoLstIANXkkwThsdzCysTUSVL+Yka30ySN3RwatpYU+mq
Sh/PyEVPHky9jQ0t3FsYtgtWbSCKeV9tHWguqyqRuNpZsASHcVlTbn6UAPshMDgBYunQ+JlTjc8j
ABVKessDfNqSTIUCYQMcfFrAGFApibkYlapzh4Zaxrmu8gTInJRcM2izBaxDoETn1X2Lg/iFqPfH
OXyzpT8xL17siAujMCYmbbyJR7bZ1hvenotUIb+QncrW2Z19oFiQ4m7FXw6lpxZOtFZJSNSUtSHT
hfweMHxytXMHSmxwaBgaOtBR7p8kAGvOUj4EjTLTREuaS0KqlF09h4kRxohqnRVqRLFF+zf73kMK
tg6xBcbjudMZBvsBwPBJ2Jld41hTA7EhyTgTp7BY/J5hZcDC4lWTEnEyvRb9MBc4xNCWk/7bFinf
+1NPj+OMJNRzhnwbfGcD41dpfoNC0cNlzA422ABB4dPUXGCw6D8sSEef/qItj87imOPgZ6dccfDB
kkGQMdsnLE09DBFXRK+xzUPtoiLDvIYE5lue1cKG/7vEuSRMzxdFQJJ0DxHnHjGZe5nhYhKkkKMI
8SnzlXLQpabESpfiBGH6vGDaToa5ATOtPJiIDN2dMG/7WRPQw2aTSX4N2nsE1C9sGrpEJ1iQ3Fvt
YU8pYPcldvYr+RCYU4M7RI2xqGVH0emdCInw6NOWlxGuaQCyvbBY7XHZAFz+gCDI8fcxeeNb/fyC
qSdde71MQpwUZJ1DjNoIzWWRiTNaRAH1Gl014z5vIKytCI0oeBiTTNoHYuiKGYrqV3BsV/LZmZV3
9FIocCPBm/c+CkwLQuoTf9Q+AbyIMfvoPTgOsUibo3tXiol3lV8+lwYd3xD+mrTzIZXuYqFcuUG/
oB5w5oD3FttwN81TU8XkOignp7cjQp1eeBN27MAk5KNDa9CvAEi4cmyH//5kyj8dOQbp5kNdy2i4
6hn15RGTSnU9/XUrdoTuZx9ZwWECm3rnpoVyF6ffBKkVEsdlqOVMyh/2ldRYirOyqC3YnZq0XxcH
GE3rhLi+JcaKiU0aW2Pq9IcjZnuwzOJ/3KEo095P/rxfWajIucJqyVN/nRGvYiD4tFkClrzJk5Vk
j2KEGo1HIlLkf4i2aEQrugsL31Nf9Q4sz2LdVPatvPaJes0xpfnJh7qa5su2zMMsM2gmBAfs2cFJ
RpdhHwTrfj9etQQpGHLcAknMvc5D0+fg8pG4tWVFWX7fyG0/3RoGxAnx/VZ7/OT+CYk9sWZbPLu+
L8FLGacSm6G0uIGTWKU+Dm+0IYbErXAmMJtmov7beTIAuAGZxwxl+gi4B0u9LIhtCXbU8W7Hb6du
z2upd8Nd/jnvp2LxCEbtp4FNoVW+fppFyvoUBtUT5vZr4gGxmjFdNWejy7UHTVtPMY32Ugxmgk/m
3o5YU9NHz4sm2N2aattMA34Qafbrob7RJrryvdyaRK0fjy+su0zsBn3bMcbYsH2ANC/AxngDeVje
XM01b1VpgHTWWWD62FNdrtZSpyjmCscCbO0wv6ZhWS11ttsGkxWRBIobXflKWArRF8hoVbc/J1Yq
ZiHkml8pRcOLUUVsAqGUbMRldOsKBD4cmRLv/Bc/x4ai20B1OQsZRRjh+rtYQKR/iAk71+hur7f7
ANWZokU7ovx47lacYav4jbKTOJaOc7Te6BtUiBW+sIct5K0QtqvCYyC4cA2lx5U9eVTGN0YU0bwp
Be0msWhRHX8WcvaucACCbtBRNOtveD1xMXwRdbHhScycpLtA5hKTymWKpUmDAuzVZ14g3IeECu5f
ls7eS77Jx19hv1lE09I+EPaVEOdHDypDEqTVHXPBDWEWlw16/1aKN2L8yz8bPqVpW2ZLrr49CjUH
W088fktmHoy3D/io+t/mnWu37xnl+kyH5Dq6o6/ydYxGTD0Jp0DiwxC17N3VekZ3J3OZ8yiW2zqN
mpJmuVBD+Mg9jnCaocuVPkVecx6adoshzpyMRE7YVE4bN7A57PWQ+zpawUTg75a6XBEGVNADZPND
g4S5Hvg9tcMiYtZJndE70SK7rRRLYlrvbUclxjFKvP6uj56rNShHY/tRp+RlENdVQhSD10+6nfh4
dgIQEG8XWMqABNXgtbIShGoI/CGfytonszDcC+8hu/ZkVeUhswMWVPatbS5qfphTqtRUxNUKO3Pt
i1rxmYVo4977UmiPs6+jth3wA9rVi0pu4eFyvy3wrh9PyPXTkBEtqhTlDqOAbqgIBgAkoFs8u6CN
pIuu/b5cixeeod6cXL5DhoohnVLpnjQQbvNSgRm/4d6xP2DLeoE9+ZcIRs50XXmkzurVXbde+FGP
j+86lZ8rFaVZAUjXnfVANKsMYOqQwrZPgrmyxzwqKSubD1Xeb7l1V1X1+38RaaFFhqsu+fXZCqeZ
e9jDddxvlVI1NJ/Eei7nrKhSk5QavE9wmRd2l6Nv5nqdFiJqew2WqZfix52TrlLPyR4ztdE8wiby
YmEPpfkZ3QG/gfwu+7vKGQzikMZJw/62BsuxnxU6aLtswLCk0siiVc7daZWRQw6X58rINDcn6psF
Q405mTK9qySFg6s1mk5EMssoZHirn9jwzkbawTJIDFDKYH0bOumfL1rdn0opdJabhJhbaQTQsf5K
GOyZupaWWn/loQSpQ0AXAO6phbs817QQas4oOIeHvXVgR+QsJKNumZPiza+Hkk4HlMOzDKNIc4UY
1Zu7vyifJ0l1SsLc9daJzbuLdbR2hKqBiisyhFSkUdBYQr4Qu3UWXuihktqON6GWOWgUsNoG+GEa
Io2UJBCNWpMeI5fzBZC3Q004TaLsjUteWWktwIp2xHeokMJjdYjqaO4WVKre5CgWGgG+0HeCTQix
/szhSKPtsMT4Hx8Xp2/vVgMnKfsteUwye678mC4ZtRxHlsv/sLZ6aHBoyH25TOK03m39/Ut93WvB
x2CJM3rnDt9rCtXt4/QDt4bFaVjzOS1Lti55oRGMk51WD6Psf9LMpv9DtXKARvKs4JcsHBbcj5kI
BlMCZto4C5tl4WvZfTRnLIid/SeJqnbfJVOWh+kBCcIMdTzU/iQHNS/RUVRRgW9i8abp5m2bQIKS
0K0G9Dz0OhyEZY4eE+lEli2Z30slrS7/oQ53qrws1x83rUzwJJdc3Jb9U4LSXiPtQe5JUK/EL69z
AIA8BdipCIhs/3AQNgdzbpOQE4d9+yNgO1A6WHmhlYtISiz3m8GWkC/yU3fYfZVAU62FyIqslvOO
maMy3PvDQbgGH/oLoVpTUMjGDN0XlDFNIfYZTFd90mobx/Zn4KnZWqvSkOASiHuILmq5IU33ITZO
0yixugZ4EHpNo4S1QGWX9pw+Ksv8BBBA9Ekp1e142mVcRdX1K7k5oJ5SVf338RipGg9x1LHBw9zB
ASyrFEgGNEFGGEhDtkhWwX9jRNybWQtxoPCPbA+ooN+4igm8T8T5l1q/OS2mUev/7fRv6bcRpVpL
5tkFs3+ZIyl2sG5r0orA4hUNTkv4TAE2w61FkxmRu4v5LzrFdQ1240RPTeotFLD4RiIYQWT0BEdR
pPnYnAV6tE//lhEzC6o4CthYhLGKQwkc/x/Mik2uHdAgCmnyXJ4A/2YIJTOD/2R+V2E2szzXbIHh
RozYBo5ILlA+JtwPF4+cwzPz5a2stZEPlHFpxU5z5Djs7zZweHBx4M0e/ZthJbPgwJYXIhhOuxzL
DlLFPqSDMrlSGREU8dJyphM6rBv730r4GoM5+xTxrd0PnIkYyvLyuT99il6CoIzOawSotLcq3KwP
ouxzl94axE2RQ+Lh4SA9I1OaPZ9i+tzf9AsmLJ4NmmipNwhBTsiznPZE499DLHz5zn/YRIx4t/gp
nFvoE0S4lCefBQRVwvn4bYWWKfvM2lS5y8XaEi5ClZi29ZV5Y7TZnkA/34tpD9LDeFC5erNyiVgy
0WkgLYJdSrfnJ/EFD75LFbWGHo0OgG4BrbZpBeb1+RukZUSSZH+rQz+UBsqCkJJHz09S3+wOMcUv
gwdB/1Ip8bkEawyA3CpBMG6dN8cmdBy2+OMsWtBggBJCG6veg+LUlznH1N0f0kAF5tPI+L9MQv4f
i7dG4xZvgtAMyBgVANgWPXN07YMxQcE2QNkanSAz+Usl4Ynaoti0DAYd8MeNohDHmsFTxU0gqjHe
ouXYsJQ4lf2p60aw9q9FzCeGq4wckOzMyaHrGzzWAaXuDgaMrXh9daIZ9+NsRSbknAU1rhoCAYJh
mVFJZ8ZglZ5SPqLtuzVRgLy1suMOWULDmq/H4noPvf7S+NuS0/lRhfaYBqMGAc9vzyia6SVypF9y
Z83M1r45bQY1yM5ouO3S2X9zkXqVLdrKHfN8038GWm3/fvYfuC44lvtW/7z1k2ppAQiJ6HIXtPXa
z3Wa6YWidJhiYPbwFEIrR20bpfmAPShzyJi1PTAouh6zQ/q9JgrAT7PsUFlogdwi0PN6Fyu3LuqQ
JWTfFPCFFu+V46ddFDZdfda4yxdrzyxon5NoFTThyDRmkT8fAOZG1T0uXww8wnX27an9Dc2PgLi4
pHUWZw1pYo1qPIaeWuTFPIZcpdEdLBe+G+VvnOplqREB8ne3jqtFnGAimm+RNxfDW637aAloKwqg
DDMs++z5ckfmRxIrzzUEz+iG2MUn56CXvuKRJLOo8V/QfqY9ILAUnFYFWMXH5l/7JvqGCXzLAY2w
23dDniZvT6YSH39BGI82/Ju9Lq66dyvIaWAkTAx3+QaT00etale3Ay+YxeVnA7eazLZIOwFMFr+O
9clGkVrV2ZRTWAGoGMPFx82xLm6o/NMfT6A3fL1Zwga5L/pKOY9DaT387BRGy3CVqcmSUVXnITWv
u3iFE7g4At1CQdCn1qZH9oNd1/wOqbVpDX68Gx8HML7L0zSGY3e2GM26CIdtwAVXo7IG64t9ZXmS
tYbm5T4GlYM37bIeXzgun39x+yPdgzfaJ4Kne8jntMz/U4qvnSd9+chx/UqfarNOvhlD3z1pwo5c
35KMRHOFW894MiiKRL6RayCoIf9dW8urTszWxlYPBEbw7RY91cUM3uxikRuompG6Yr+6cKXCMop4
OR7SY7e1Pgfgqg5iT5kQ+DJcnTNoKB4Zt2lCgq/N5W8HF6T5G5IKyOut/h4aQ6nHcPuAMlrFt7Mo
a5z78lqBTK0DgXyDCK/hhEsCErUbVeqI8xOCr+KQuH95l3SVWBdwRzTDRE9pTWRGMyJ9MS1EsJvM
wQkuFOP/b/lGHVIlZNfP2G8VTjn8BfGXPqqptm1WMud3xCnGS1ePvMdAHYMqMZiJEno+IghL3F3F
OpK8HyiCnzhyAbltrgjvyVc9rboOG1+/VyS6BIZrA2UzsqH3F9F4RT13AJJXra2QJhnlB58b+l3K
zPCU7PFKId6zYXSZYhwQfRPxqIAM22rwiq48UQ4gT/RCOw/NLroN1uaIVMotlsjekDOvGQf17u2l
eOFlMii2Jc9rZpbdNC9AAsoqaMujwpg0sFQ4jIZrHZGk/ZnqabzF9n1+YmeMCpOkhYQNZXACEBPr
mId6/u93SpSXbJ4bGY502Jk2eslpnVXuw1BIm+rN9eO2Cysol+5cNWj19ZAQ9G6MzYzewlVZ0PBO
GIeR3/AbfQFZpDnFndI+LSMQ56RKNcFC210fuKQtuzFZauGgDj+pQgb8UflZG1RHThapBNMzv5Y0
flIW/gl/qKgrgPrONGQM6QY8nV5aNulAtUo5OCvuEt9A/vPazUIvdHoKphvYSCQLJ/VwTzl48AP/
VqlyOypWjrq3xUtEHHvfvm6uv3u5P5eo9E4zoUkEvgVFVeBtVxilqoIB46a3F2EkGAwI4j1PZj3p
PstiqPxtSk+bbSkD+vBay7UDfvLXKQZT5Zk/tEqxP0srOD43AjIKpyYTSu6hgovHgAEzbFCHADuC
DRBM9DdMRqoEGixBWx2Qbyr4bMdVR/yEXQOgKLU7aH3GZKZ3GC/W+cvHNe2CLwtqdRsZK+Uuzyk0
EmMtbB/+K2+2NXKK02QIFlp7yeLVzHt9hH9pnPmZN1wygVDVS5j5z+p7TgqjzxsRfJ9cxs0aMI9i
9Ak7F+x2UoRl7SyGbeZAcfbR7n2cvRaG9dd0L02nWx+JIRhBPP4Enl5CPNY1fyyJHHLy1H0W7a+b
nxJ0xvoOBR6u+tok8kJkUMtJPgu+4ZR5VuxyQnU7g2iYRpIs6PqYeaWMT/YUYkucDklo2aQkzQVa
eX9LyWoS2RfEHHKdPwyn2G4inpPn8Io4RCmHgqEO0jD59O+/2SKQvVAVDdYTEAhSyjMCgULyQ4hw
wzhlRbNusl9o01xEen3HNm0b5FNFf0J7mIHY0j881pmYiJmYBqquLfmUjHPhFVB2Qbnfg+HWcm4n
eD8ORVzHl3Mysng+zGER6hOM0IGfHNW54R7+pQwwmAjbymm2WwcLpRMiNLRopCzMdd1d0nHC6i7d
KUJQ+T9pQqq2zYcC0MW1oD6wCTM4Fv+7VdOvV7Bh5u2RkOXhHwVafT27W2H3o7XZUUxZXVWUt7tj
dxJq8OhSFQ3DLsi+tS9LPZBs9pwX1inxK/PIQEE/X0c168/WuskLKwowGbBpiOIhmeIMrevHGkpj
FcPr6qw+CRlQVuRDic5tiYuJlKVLcTNSUFZi3SQl36r1mVTGPD/o9kwkAD+kOLfqIpUDLl0gaUcS
Y6qEA6TIqJ7828ILfmdym3jAH82UOl1au4tX/LELxNho3MtMXkIHmGZ8OmU8PYyhcT2KqcJWJ+S/
S7mQws9enPgCQ/BZU5lLbTvPse7IiQwgak1I8KqJxZJTlu4hHipcd+NZmbJS3EL/K++ePRrkRQt0
UpfMNvxmfGheH1WNoxJ1cIjj319HYaPo0Y4z3ohN8U44pP6SX5my8OONKxYORlF2eE/gR/a5eCKI
jaoDeh9+ErvJaS/E3PLZksF1s8kMYKtPtPLsLfODlBw3IyuBYPKoRtfnY4u+YQAlAJBbIQhkhjDb
OzNejTKzhxrUlmwdYpVknuUinRKY9F8qF8AT4sNw+51ccKjTNTK0aPkEdB/rot9t8mbfjUImDAkw
KWIwFLyANTQLTBE8dAM8e7cbCChxDYkmpn8XTecw7r+CTxUJoiQI0K6N93x815w7RBQ+e1NXa+Gn
xs5ftlYakg9dyRJcS+nlIUJ8xb8xoM6NQnDQbFEFdVBfQYEY0v+/eE2KaN0lQ7LL/wbWa6k2JPcI
WN4R1wUXe1hdh9LcFIgx1EDPYofWbgoNZAZ7/30DL2fDV/lDBFRIY7IGtqeWqCSEc5IeCvtBXo4S
KaqEilZUweBQCq50n3xa6pXe2WdTM++4Jap5x1zRvhSt6LrppX3B5ynQZV3I6brWcCaUirjMu0M0
0Po0wmeEdO2Ugv9CMR1Y6R7tlR/1V4+2EOrJW/9R7H8x4e9XuRnMVS5tTidhLwmOwI/7NYc0FebT
Gl5/egU7gKWiUuomSS4/1l2JwD7WzbDxGvxV8EFJAnGY6z9DfgzC2qHvXEsckjhb/MNXn8FQ83zK
CevG4atOodAATS2fh/J6dyNvejL5PiWFD2cAg35l0Afrn/eLumU1nU55zIYBRKqrJhkH0VrgG1ju
Er8IS4yd+PoqPOS3ZmMJLk3yXY9vZ1gAH84Gjq+zQmgbfqTXqVDigR09cm7RcNosXgC8KdulumR3
HnKG32G0SJGVUvDmhpx6uPwzxNysRfuwH2RrzZ4x6+p0xv916/WED9YBpBmEndHCYeJ7AWxPnsHT
YDe371YzYFxaEyKG63KBnpXmCQaamVukbF0NQ68GnWVKmvW2R6AaEsAgQPMVQVnMES75NwLepgFQ
D96dfD8IdSezb0T0UguRWydf5LHrmNTG8hSHPmiQCz2R0FfD1s/hrbwb/HBy/Js6qoRofssaUr0R
wpjsMUZ9TXXvJxIld/9mhIxNxAUc6nh1j9RKoxMlFgUZoxyEZeczh+FC+aAQUdI98+Cw4BdY1V+X
j0mQj3QksrXUZaEQ13/611xZyoTunmxunV13nrvL6dN6NGqIRackY8mZVQdxQDJ9nJxXcsdjkNSt
cjwkQNwK/zqL0egXRppscf1PsUasjAH4Zqouq2bU8yHOPIk2zoCwEHl68KJXrL/d0AmXM8iK5xCg
6sK3ZKhZx9YUoWmgnA1Ak2XWY+9Ow9oQJ6dKpmA/9F/lzuLxKW98e871HPqrSE51BW2Ilyj0kk7m
nVMQBwewwSNxQsRX2Y50/IqqO2G0fqMO+PFaH+00QJCJk/FGpTQE3le06U2Cqb15+hN8T0fbsfz/
r85wwIeVTUrWjmYcQgG9in1RD13jGde3U9/sYflEp7CIecu/Gyj08b2XjOXOFpEMYkU0XIlJieLp
hta9Oi0IGK5rJajjeOjv8H8JKIEZw999K/zo+Rvs9+HbdMA4lE8NXqX/x2gqNy4m4sJHPtSPTY0H
3Cc8oB2XSZrxRkcbBXUUo0DFkxyeDs1Rbd6lRaWD25VbGTiX8aejLFhw1jmrMoFruR9szTJj4GlE
06oIbn330YbO1cugBUTVuk+4yCHXJJn9M94TZsK+k4mqRffmWEheT8Ls6YN6kcuuJG1jKfmCDaeB
gcgwSc4Iof8WimEgANlB2h4hjGVD9KsQ4nNThcBDDEehPKy4CRRqa1AhjTweuiZJp4q+8/x30rxK
GBGIwrDDOVCg7W8oUiTv/7ZrWJjEYWvqTXsZIv5hZvYalP5VT0FX2fdDJT3T12CnhoiP+2Sx8YMI
TgtvINXWM26h1RKGViJrqfutwQ9PqCbfkMqitcdxeMvUugdz6ivt89wg4wH8vDcpx9wwZ2n+475E
fqJsGEdbJQl0secU1E7z7w0AkOuCBMVxmagijb4eoZicVtsOJLFd0qpIZhFJASnND9p40IqWaf+r
5fvQOMt96OON80uDXUL2I4bDDhA2zMHRtrkv5w3Q+SF82Qt1Flp8dQrzNYJsrH6PzXJcNfX9cAr9
P9lkLfqOz8xApXGV1mxqz57G5Y01pIu+DgReeD9WFjZHBBmhsAQofrAKufycuvfd3eSARXCZTwSZ
JJ4o1nCVUrFY3J40zBQ6P9ATYByIibfwLCfpZaCV4eP+yTMI90tQh7KwjmPN+iNWxIftSgqkcwmM
2nzxdKoXppumS95eFhBNFMjM8/wnq9VMhR97HTHhn9n+PRDfDyvHN0VbF8rfP8ceelIwh4X+gt1/
Up0MREUPIbt12ZtWDSz3QVvkr6+b8XvOh+4NgSeuUFz4Rjw0rAG2O1fkDydaBGjpdUbZoL3f5/Nc
wP5blS4t2DmtNg5qiK4+pKeqdpy+MTMEJLbYOmx6FqwxhdXH9wLD/lrr71R4Vd3NmbMaR1Ifod9q
/2/+2MpEQE0XTKM75Evposlc/h23kPmK3vWwVYjYclvkbrLu8F+Uhlw2NUBVphZYQJm+kDpUW9XP
mV4qNn+csPUoUHuvNOE3/M2Zcn6IUUvkMyeRADqOl/aMkuPOMKS0rh2At5aJ9L9YRp6a6FeFDRkI
5hodbGWciKtKDH7LxKxQEQinit0KTSEOFknoPMqvS9R9JJelfeeOfO3QTvYTTscj0JZGercBC5v/
06y3wV58WWKzuZQ4q3Va/hod6aLvu71c/VrhasHVmtM+3wWkPMMRI7Ty0uHZMgvko4G9nymt13FG
Lews+PzUofq2EhMAk4EfXXqLIERBjL0IELwyS+tqoiPTv47tCRcgb+SGoBrt8rX5bl6Hh+aBfgn6
fIgbqpIQibediTbXMBF5SStGqAc0jzO/4i5mQxUOKtBF7ra9yJ7I4ULu6X0QoLA09rvMfQ8z/01x
yq249b+XRKQlgwkXYiO8H+kzA4D9EQ1kScK/J1Wti9AFuAo5Y7gBVDcbFrMNeiOv7/kTHBtfLCEM
QOMB6nSdsl/bf+gMtYYzRRp+QJ9QJ682oFi5SruK2zauiYuZdBYc6CwbnB/MuXfFzcv+Zpsyb21f
CWwTr25pfkPvjVG2VSdQZiURtjMzUTyNr3Hz1I3jHnp9kwyZtRs1vkGpOnOvPdM3oeQe8BbK8Epe
XEeA5+3Jc9yIuUYv5dq2GQAGl/uiIZN8gqNhNUVWI6hmbeTwA7Z+73ps3Sgk1Mk4YMwB/I9hFJ4B
2ym+nNzOiT+PmNO/yj7Xr8GLrq2qqraeC4Y58njnlA/Yp2+YgKQgUOLIAggN9na1IQBBGP8IMaZQ
wbpIowgocVgV03/ZfWHKopCDMFJn4OTkTEhE26PEN4q8+B4nNm9fhc8QE/yHvxO7AlMpZIA2ix1d
jseQnUT/mGk3O6if78pt0W2KbMw12iWuX4N+drz8pPjA1yGx1cxDJO22fAHk0nXStJIiesymJQAi
78HdmJSnTXiIxmLV+AuE02u3TYHFW36Z/ZYD8gbkjyBFvjwhu1XEvnPx1SOeDdAHGH7d15gAk0np
xgZfwjg7KqY2xSM2UmJbhIM2d2jXqieyUtJb2aGtNXA6QSklbSGpq76Lvet6WmvUGErVs12ZOtPz
hzmKYLKC5FMmMmh9I/Fk8JWav0ECr0QyFK824N4yRCIvlvRuIbINkWO6NEAHfyS+kkPfEpt09qp9
lkTGH6qcxdV87EM4SuOE1q8/fV3zMXuAnyGmzBZE9hdO4J0805Vq176Q0DlxSmUWJa63zeQNPZnL
DahsdZvfzf2NIGo40DMZcr7S8S/mdzbunH6xWAgcAafp7RJ6llWliAGXMdt+wE5iompMXHROhFYF
yEYxr11xZ1jW5aIbAsrbaVN2VUwKF1GHCG9Ln70rIrTlz+eedKLpsQ5vz9JPC+iwhtqLo870kLvJ
DvpvSOy0W1Wy2b/BTtdMC6Krr3B5VCsMRtkivZVJ3S9Abp5rBZ1J20CbZ28lUCkaFLRvEiUw38pC
uGiNP+RO45rIO2w6deLn6w2OeORK1mkgQ/SzwIFCpHvvxfjAVFV+WagrrebKs/bF12KI7IGM/o/m
Kdsq3kBKDXJP8yJR/pFGMK9nyODeWHnX22RLoz+Jjn5z8fwtCqIQPoEYqPaOJGXNsQmnJLKCKrio
wyW6t6fQCCZT8Ex90nwPnWHA1ZbWG+B3VJaG6ItwbnKP0rskCLVvV6g8eWJuUiijUDjB4fzhcNZa
vgzOE0M4izOQCfh3LLmlOp2r+/5KxU0VgAAcMhqcVhdwvnFhgi7zhjkXYG6+nLaQHEAEqH9viH+k
axgs8+M+5dHEjmxGN7IRCtub88JEUKdsudQUhIonO5+QpP/RZD2+ws3vzHvpvFsYjhje9De6j6qJ
tZnU0I+jS79j7Gbi3Ih2G9VQtH09Ona1TOU3Knu/hvYn7CwCrhLifI9PREW/QIfDW8ExE3uM238G
QKjeKZ67P4wl5zjMMiUBPnalXIFMoLMJ7nU2ago6kaS+C8jLWaE2Vgz9OKUrYLL6rXsm070J8O4m
sKc/GYyw28/GumhvSR0pcbuz5o6TprYKsUfXi+DJHFUHQajzwRMYfVoJFDS3xALCLwiXus928oQJ
tOeC6BAuLFfCW2W3ZSURZY4yxBHcsAYBScX9QkrVqyri8CtsMo8SDU508R7Dx979Mno8K3Cns3SY
DICCDBxMMW//Yq8jrTd6NF8oSVnDy7lzB9WBXJuY5/lE93p2X7irJS0IpFQ3UtoySinUSSZp1ZOm
GsER7OvERq1mOm0USLBiDw3b2XkcMTsbtxAw983tTuAEAp372iQHTTkBODqLy3iI7sw2u7Rkq5mD
nNEfZau7O58qpwXVFE8NOcGjvyuuKm61roBtoBAbeTz2TTvnmS99Cdrqg0EwM83pVNzR+rzizshC
GZbyiunTW43NoDlIK4j2HLluxAY8llYTjs+quD8s2106MEe61uSqk6P9AUKlcvBBFdt9KoDusx5/
wybowQ3HUi0AFZvZffwzepurV4+2uWlcKY6vbapFVDz/XM4HwGfDqSNLrKFlpru39BQF+B5m6L/4
o6WiCSPFlhHrXYpFAuRp1ApR9mo2905FHsrKlW2Kfh5IHB60IU4la0C6Y1KoUJVQni5KY/gBolFu
4/F2XnVWZBHbcmZtjRKXce7KqQZ1c+OO4bhPMjau6/ayAsJUDGb2rskYVHgSP4dMJpOshkvY/C/f
5i7laVfWGoURQgMtQrZ0JtNRrn25dS49TkVfqpQ9djMndnmxYn7kC6x1skPhD88zphPgvOyr9mLk
Qt/9JvHrgRyYgPuYrdLijHbTj8w/obRTir4grOtrmmarBO45vLjOnYy727+M2fwBomIc+iLc6AOc
d+XwGw+dhrzT2xsqP1EE6LCYCci1YYOGuPVReChLG/1++MvwHHr+d3fAO0TkFceJreC8hDroWOb+
62seQu9+vqlNtgmFWoaN9AfCFFJscrFZtWhoo/ZeyOybQlOXSahCr84en5IHcTWbWaLQiAn/AvRI
sesFmFJY44R91F1q1ZP3mZ+Q1TdMslBfgX9i+Iu5ZXBAUEH0PZWKL8CLAym0zgMIo1PwCcxzjfsP
J44JOLweDTh+irfDaEl5c2qJ+jHDhxmj1n9cCYGYchDBpeQy4gDQKvJsoBK5PAqgMQYDHL7Jk5rU
UxImULkkEhyk4t3YrOvGTdQsBKsbMZAJ1nApAPus+NXWwMgesUWKv51UHwlk2feIMqnX820vj9tp
qeC7iGidHQJvs7NVJebD6EXfFErMdMNVe7dCeBY2BwHOzetJdV/HRliZ/UExpnsATV6VafWJoejs
XHKEuJj/G0nI/cr29ZBzkRCfg/2CH5xwRDPz+FBXg0reqdNarJkoqlQ3iDbgkLkQLvYV97LtOMG9
D5kOrl/hZncE5WXmluVcmGcMt9VB79feCh8of2axyGa+iLHxIlh/YSetr8wr2v0HzAVPUup5pyOB
96ncKV+UkmiHNnv9pmOB99N0zTvUNOGojDQT+fslscIKh0V3ZTtiKMMHJwMfVpTQ6+G7mJNfalC4
UMZ0qhLho3rC8VllJ/hBvov26sQzGq+lR0EcjUmWXzbZVEDgGwkcGLQ2m6CnsvOLodUmK/Vd0TPq
IA+X9SNeHaz3rMdaUUHfQdbI6t2xtIkvTINPtDLuL20ulPGPOTZEmMmUdC/ew0jJyvGfj8LPKRAe
65CZPW7ynR1bQT8iVx3eej+PyOKaB7n5MIKpNL/XsayeO1XD37Mrk802g0O+KtLPOkSTpuFOMpNh
mRevfhKpXv2mdKiziW/1fmZ0ujiRMh3YZfTUqHf6T/SUgzfZ1/V3o+ASeBdoCEvwgGyRxrWq3W+d
Qx6e2q4AVK32ImrcgmDGA6QXYrhrTm7lC8A5Tutp4BA4JyODzLnxnr/BDjAgUY2RL1snOYC2KU7T
ZVli/q4kMhjOWrMJvBfUSDjeF6z1C2+ex+zRiMbC0Dz26IIT5bf2uMupt0wGNPo11n0wmoo4iaFH
UPLhZwRsNX3bpC6DwVwFcS60DkTSVvsyqi8sn1KMAdImInrZqfO1p+tmWioJlL4RSZPzMhOyrYky
eK4Xc98Jv0m8iKMhX/ncjdiDus5ESIHXBLPBQLurcj49I0RquSkkpkQdoo9RNGgOWNihLIe0wKx9
K3jykNdfITM0yFaiFeS8ODMIFlBj2IAmUDzKAwovXCvxbOLuuy7y4RL4kCQwTWndZhnNyeoVM0ya
p9k0pJsVxjzN5tSkqSMulm3fFN2mEEVzpuuhSjPVJ2pwoK21xuNxK/vljM6BCRZfCU7clImO2is7
XHbzn4nz8XAZ0RcGjOgINIww/jC2U4fvrUOm4Od7UYsWCIEcM5Ji1NhIwgH6mxp1BeZp+Q8ZhY5d
kVbiD0eKIB8TwqVxH9uxy+DAOcc/264AWUf8SSuJqlr+nWwEMuYQGrzArAcsLOWYdrs+l0AcnMTi
Oq2PDyo7m6JUX7Rgh8LGyAzu5ndYzM4rwV/mcqYUA3PVFoM218JwLH2ij9NrJF0QEuD9z3o2NS3r
fPlQP/OrihT69Ct4L6AZAnrgGqLOXaW4/XHxwRZoOUBvmB8DC+rUuKs1FhC83LmBgmZMfJGkY/5r
CE6nf8TfyBIHz4O0Zn58kAkXuPJpz/yLrxTgk2nlT5wv9rCmZ+UNnuPA5xQA4DvJcJxYUPF3M90O
oE0TlZVw8GLqugMWbMAu0Jyblu512bVdg4U03pteBEK68Fyg1JLO6+1VawtS8kO+/Z1BPzskllKk
SnUwU1ME2zLu2e0urE4/AE0TTeiwZ62ytZ6fmuVJpbDZlEmsr/q8JwLugKync6Sd4isjxQ8puNjm
LYyKfk+JXnONzuAxolyilSmLtW7m/cqQWFrQ4f6nmSc33UTximD+mnxYlDuCmg1aGWA6eHK3jK+o
FMuMof0GhQxyCiO5TyvZHRRzD3WmIOggn+DWCvM2SN/pe624ovTysksBjBR0hx9rmeSXG7n0ites
qU7iuQs0CG4SXwAjQzmCtXZpNyTvH9REsMoMo5KXw6KRER5YwgXr2QGkkUKniwnkBILlAFYlZgh5
5jKs1cBjv8bZJs0ZhA9Wfv5XFcy2N85XC3X668/oJSqO+Vvfylym7AnANv3Xkv8hXAIs0Y3SZl1B
SgD9sMYbdelpvtS5/PU3kQ70xijdGnd5mYCu5cjKjL9pC2KrJysxUrDNNhllzX2GqOMTUIZDUKQ0
Rnk4Xh+gwSjry3MRx6eEoPXr9dP1N+z4+K5mgv/22sCGgBm7YXjXmazsHgW2fephzK+h6L1+e/nB
htMsLd73YctEkG0OHAFsgYC+xGal1qCyhk2QZQJDxo4wGcKaIFxFka031yjH2EWbV4nkb2er4DjI
VgtmD3E8CAX8/6zr5E2A/jiuHIt5z/xkdC6GVty2L311VjD2zsqRakphtRPke7rAQt7AaKVNEO5L
E2HD0vyKI4gjzMiCq8izMMnXengD11/5O3oMWBMI1OYQLxbxYn9YzfnI7T+mtM7Tn2JJxVBMLEyk
TByofYnkoseoRl2tF3vSxlphzQE6o4pYJ9Uiwy4CrkJbPkzgTEzjhf1GRCHdtn6gMmo6jjDZo+w7
4+dQp3tTDuk/Uavd6Ox09LGIz8wHIczlx5z/Tu98BOLEddo1TxGC8ihs5enheS5NvwziiJc4av8r
gKPnMW4KZkXdqS31Td94kji7EwoR50SA/20mWncbP96k/7dm8k4ceK0Fk3SxTEbw/holQessPyX+
SAWxCBCLLDa2GepHkF5fE2SrUL4Q47EG/dtWVwB4jZWmc07ItT2mW+/K+Sc3+5dDgJMJyAsgKMJ6
cHQCDHmDK+JRe2lDQz/6HdkmmqTHopXCgPYQZzMKLS9mo//n34e4vLd7obGQ6ZQQngwJQGfC2E8z
9N8IaC8N7kQx6D7AuJCHdSwoBAyNmXPMflQEb+7mpkOUkTWDJZXguJgYUkUYKHWOhpBP9iJJ8JPd
zx8ui4ogjfyXJAPrg6me3Oxym3xtKDNrtyEdom102+Yn3DwLvPOWuWuKgqiH0Ps3afRFg/ip50SL
kCYn0eZN7YCSW2eNSi9MJju0vs9cWtj01G0DYr1zIARA56Mb9uWXtlxS9VwWe00x2NTzaOKh22z5
XGCHoEmpaBLXzIHMjMJK/sHMQje9UGPweagOEgyiOJBjD1++RUMMCSB2lkJje6L3eQ9SqKqH08Rm
JBPWx/aa1QNwI1ou05CIGQORJJ/fSwFtBUoLoEwVcwr+kZKB803LyxH0A1C/5aj2b1t6m9no1YuS
1VCPtnvbIlk57zqkDN/kG26MBIPvc9vmRA3LHChlqzG/gHf6176YtPdptBmCE6E3aWxRpCvedHrt
T/EGHPNrVOmt/T7EeKYWkCwhla5q2/DlzEXTBvkH0T/NmSvCQR+6i/op0571YHPPAhscW8aTEQXw
rhAFMv4OXnMLkSYXpPUSP6ujBz+/prObDiqbL5WEmjWpBc+Mv7wC8nmhPEI91QU1nm/j4N7w5UlO
t3twY6yQx1Jw5QkH+QO0CZMLz0WezMG/BHWczZA57Gz1GX1XHrQkFReRSqfEGfNz6t4azgr1JBCJ
Hk5ypl8+z+3J4XOnHM1hEcAx72Mtd7w5EZwoxQ7DdVbsjqtrCnLCnAkm3bfneP+uuLv5oFLSXVBo
oIRiO7hydlU9X0Q6UJ0eWJE/4/YxjyFuoFr+wUPxxDBc+W8LNdbEw2h1gfvQrXbxWAVlRUoNKeKF
lRXaHrGM8bqTsmt4E8S8dZCY/tlaSGVjvP+IUUrTnBVGNwi59kMVk8I0WSx792l7bWeH8VAa4J5I
MN3WY/p4zNhaigbgh48dNq9k39vmKmqVHnji8WAdMJRdmr8yvA+kQPipEsPgP/Iny8VU6UmsAOOI
kpBMbhne8DRJYp/ZvdvWP7lyC3RiQbknFLwzvsoqbKNddKsfMgHQXdSSxSuVPnQzVFuEOoz/dVmW
QBCITq0urJIs0CKUREvuv11qzUjgZsll/ykIbJdlcjOwYlrTkW98S5Y/zsGHBFZ9/rqkflXflO87
omwUqJsV96/3pc0N/r2orbm39xTH9/L3sLNdQ8Qzg8PfElQhARwCJH8YHJoD7ZNn/vcn3k22Ymdz
9Y6Z3sG1powPgr6/HypMizmddqEYZyXiPKdE12QunEhKTHlVXvUMGaSvRTxkX9OF/TGlzc37qL7S
OcW5W2aN56EGqFsLcOKUnqvyP6FaGYJ4XVpw+lDTcC7JwSV+pGCRNMhZqtsX1AfzOMQs2hIgcN5E
jd/BNPipwxBjPJ428aqaZKX/bn9u4dvOZnWLU5+5U68U/rgmMyNNdvZrhmo6WAcICGobODd6LSRp
k0QIltYb6Wcin5grxavLgCjpN6tnffiGwZPrZZ2WaVRIR6iIxGwBTSf2bDZq/EKXNlef04tawnWW
0mWhpWBwopo8csWzPWSoBBuLlntkx5TcNMSNMP3cMaFYQNQ3S/0E7Yq2a/IPzpUQNs88Nx9yh/QS
/NVOKN3XmWPZi3xFjuc+t+VpJRYPAQSwxRNtgpCWYsGDPzUPdqrB/Kr4JhIwVQ12ZMDDf8Yp2MTj
8mOyqZvsMyGLAoU+V2VuiKicX0w/dEpGFdgcm7DDyD2M3kr/DjMR96xEECqIhmdKzJGytxfO4kXj
YMh7lvmFF+A9CR0FnmfWXd4FDU+eBrCM7wxHpII3lDiwMj5+pmcO895m+E9pQwPuK41shunuTG3x
pG+eGVVtvzZRbkEDMQKYLqOpJIGpbP5zncP/GxIQSKhXQJ2JXcxLsNFj8Xlsfku4xM4CINIC8r4V
t/0XywFtglM8lLHeK46I9I0ytUGT3OaxRVsSpkjJnJDTHMf7FtymUqo6RIeQwrSWynvG5/w2XcNq
ERvPl+2hZHFNSbGqoBnvAFKaUzw8O6K1x3u1y4/3HdEM5hgfHP1D9USiATiNpvdujJ+YUQeLVyRg
Wlnb+62eSpzXkn0YT9O3V3xYBCWWewVVQEtLGAG5Z9xa9LdhdyhKFCGFtCWMNAHfFdXtkkfVdboH
I67uhW4IDC/hvoqUkjYqw+BX1k4bTMYLDyFuumoHfN0bUFoylWYgP+qQOFiQ/vwXRZXNipu+PtnS
DDVl+Vtrx8RXIceyjfVyA+c+VMOxgHPNX0VOMfPsNqBwSUMxeibY1+/clJJIqcmfA+2JMiaXh0ri
UtybHKf2nfOrqWYbQjFPhYtWPNOa/vp4ayNjU5aF3A8vvDBSRq8yLlirm5QTzkB+QwUogsqouTrt
0E+PxFgz/1P/4T9zoxQDf5OjvoPfhqC6hDmdSlSpTpzPuyroLgCIcdkk8U8vIdL8WmrlWHbErhWD
BZeKpvZDeEw5x9IPJin0Ci9wzCt6D0FFQCgy1Hdi2C3yZGv4F65am5tltEX+EMwnH/3W+VXTwnIV
P1UKjTAnvWnUXiKu7g28U5+Tv6n6AF2cdm93uNZ51PngoSR9+7+UsXdY2YTbBecKsuiUXaYESdVs
90YYZbcUsw88a34eB0L/DUrqz79cXTEosTs6R2/qWjA6wISbweTq6OiI1yt5S1PcNfhRUKXJa0+p
WZgZiujbKU6P9atbXwqyZb1vHVIpFnaY79mVbnOMGIeM/hFPamNWYRTCTVur44nxA71To6YhdwqF
KEUpaR05iFue1LNFpd/6nGzI9v1pt6f+0dlvZJ+sHi9zEQXQhHNGDaUnnd4sVilntzxzfyqIO3sh
/zqDNj81CVRv1TLHgBVCl8djhJ5qJrqoEolKweU4HSqUnqyFwatgRFfpa3zKB4zYojVbrUdUuJq+
Z5kJr/ooi+PDKtpCtmAZvRv1LNkVtOygAS4SnzUeQJeOrNm9DIarMlfoy9+XInEawA2SkKrk4aKu
KccQtuaaezX1twappSX3nzH4tKCcxA0iat2sjxzhiCs0fAHHmWtIlTUt7mACu5hnWku/jmEb1rBk
dErfmpqtvv88RZ1P8E1pOB5vOzGR/2gE9aNwd7ZS9y3Iv8JAqMi0KqvzYA0XSoIWCgeg37e2tFRM
UD3+5VQtnX/PDEeoC7Bw+WZgz0lLHssAwn6wu6yXcz3X5n/w+YMoaffWa/EBpKNbrvO9Z7LhT2FV
+qR4t1VDi1SFcpdD0tZ3+qpa7uHi70EO3CpvkrOJga68eOzzdDlY1YdHp9xyWxkl21GmOsDjVnVV
RKsKNWa/xe+tkKTkiU14usZb3AT8Z5MY8UdZOexHozX1tJyKtNmJhi9X7UAlUSTmNxE2PcCFBVN1
4P1MuM/hvT3i7f1S8FVeRo/rJBky7nKiqj7uQoIoP9On+gYaPgYgeP331lBA814rZbfeC2vSbfGz
oxgG5ZV9bUkXI1l+ONWFXlzSiXV1svH4zQ5MeDfcEpO+WIkAkuZDqRv1F1rDsV7HkFHzaN/tfLMI
3k/F2la+otB6tw3Lx7lBgSVRsBjBLo74OXtqGHYHy1kdPDdoverXeTY0gVr0nGe3homagKhhOppn
3Ez6tcTHJCIPUCOfO1n/FwP4XgRIIUql/SloLp+nDRzpXNTovEfi7KDyk7o7MhWSCo7hQ8wIWCTc
gaoDPlOO7OQj5lyNNghkcvFqAnKblgiUmRluuIX0rmAxUKNt4LJ9bRl7Zkfi/+B7CMPX7xAW5fFC
JK/3It88ISjp+4Tx7HqSQj31RcgbTR57sA7jo0FAu9TJMicDmpq/zb6AC0tBE/iht6iZjG0qGpMN
/93RN5Cq0hDRddVL6tmCZDZldC5VLkZAAFKbuUegrv60NICJW5qPV//ArRgawkBou0mpc8zKMzto
Lixsl3RC41fjrotTUosntI+rd2oO8hU7x8uqY7gOV54UGIGTBnTM5U/hj+AJNORV3S3r2bAlLdTI
/ulksMFPoRfuIVWFAm6HkMMCKdUR9rskcg6gEguaqiPv87b9QedQWdB2m/B3BL3rdXpneZQBG0iw
Xx6cG81QKYZSncgY7uwtNkMhF2JEE4KR6If35Mt3bZ0F7UJzLyegNq4a1Wsr365gZN6V5mLP2mBB
jRHEsSI+Cent6zK8EhmDfXp4d+We7edkXctVJ/jvwo8s7yyajfuF1ZbEPJgXMYd0f31H9IC3ig6G
KduvqmBRGJrHkaKU++kZY6434x8/yEpGeUpeB2jtGQ+I/uKO8VywJuX2TXsked+12bbWJyiRe0Ip
aT5smVcvUfNHcbURpbBTOXVEBp8HT7xjhjh8uqtvrLaofrL8IyMxwxDVITm0So3cUnEBm2xRsh32
QrLkQThY45kEdtU2KJ8OVX4UGGxEYQDjUzUATSMbkKJBfo3Nk4xCBF1NaK4woe27Aj1O/+mAPrHa
c1QoFuHNq5G6PpJtKuFWNT6ba14njUms1hOezUwSacQgbU42aa04CsPgMTkOi7smk7Y0RoxkQubU
4IxL3BzFZ+OZDZnrI7PGqkyHci5aOGj8QF81dHDNdMD+S+qpRkkqP23Yxc/B1LGSGOLFsjamHFu/
0xaS96RWwt7dQ3Dsp5bwwBe80gp5qqOUqZ+L6dR51KXTpPk5NccifZ7mnkn/Hn+Ur23lgGPRn7+U
aeQZcsX/MUcNIzT4qkERYvV5zmHEayyiLQVGOCN4w/DU+0RktDXc9rvKKd3EvIGCQekhMfaCtaok
V9EvtWbNYDVT4ovZNn85XEAzQ96vtlcC74elO97BmyJ546Q2cnxNmxyLY16veNbwhN7w1Tba0Gey
SVrGsrgn9Ceqfs2yEroLY4LafGuygMC82or1KKK8Pw8alUSEoA/A1LyKvCz9GtwGGl8BNhp6Vydm
lRIR3y/+l2LdbDdI7CWqoLg4+Kk4FTh4nfV7lnOd3D+xOn11kuQTwMoxJW3U2di9wymQJmWAEqLb
T+3HX/Ff0z+dI/pAMOJ1VxJR2LEG6YpKWoSEj6Tn5Tm7L6i+qlGw5FlLApYofZZ6DgHmBTCgoe8C
6Fay5MizqnsMFIQVyKwITdZZkerDZj/mtwYs/o+tgWBUFRgkmzzqBYIT2aew4LiUVgYWt8IKwmiz
RCCRV0nMAz6radghBhgYVvTn0wOcEc6XYsuWXLcQsOeeeYsDUfMwJoZH4KdFXR8HU806SQx//ww1
LgN+IYNkIgtGstt+Uzr0BSQkRQPRiNF8W/lw5bzHTPMsdkWFv951EmokJabE6laERxmLtjGSkHv6
INaB5Fx1MjYGt4gCUqdtcRMmZIwPCh+v3n1g0UpgZTA674fYgPRf7RnnWCH1808wEhsmY+5Jt4+0
PI3DvJHXrZ3vSQTIYLgzIPuPSeEodfd1+ELfiifyMwM6adpM1UB0b3igWjZ4b986xCFRXrFpzzmP
fEF/L+rBIR+bY+GfyUlyKF1WO54ziLPU92TtjtObNBXq47SoWk5/6lVfmgGk5jCI/yAQtWtvT27a
wEefrrK4KYHNXgJred5KC+4LWKQqSUESoClN/8onu2iajl+bCuPn5XRXxUv0nlH8WSY+SZLBHzRK
t7vq7D7AmBZ8Lk/c/BJAIzvozZdOVytmOlV0ElFhoL9XH2egCpMzbGOEJh/Mu3OpEv4YNrkm43wm
/z2qDy/0379Y5DOaASxvfKiDxPL4lOXpUUZb5vs6Mqnmbp3rTXXqBpEyB7hKsXqiwM4RXhjvA9kr
8uAbo2/oPlHJ5XLmmq9XX7oRpPKICI+Cek14E0e0iUC6hfqyAAVRPEWwglg/Klb+YyOjD4eQvS00
KiPSD+XM18p8UsSsGmjgqzbWs0F+frup9mHnIS/BrRj10fyGnCwYL2VESlgfgdQKP/23F9Q5r/YZ
xa2okQ5wlzGylaS7DXWZ+6RpRzRqOaXJPqw0s7OF2iccffePbUwO7PNruYcd5zqof0AXVG1PC0Yk
mtsiMXY8EXZduOVgtg3sApjNtg2V3MY+onK2Z5asuOjZJ0J60aolVhDSxc7zaLEje6xW5WYOxNo4
UbGbke9O5JPrZHFEHoRyx6UPoMyF3devKl/YoSG8Iy9T3aZOBPa8AiYmqvSazh1XBNyci/+W7EXO
E2LkAyk4qk8/Fymv9YbOVHJdMtrQh4hXHf0mWGNHNWF43/utMr5VLUIhF8vlodMritH/dm4sebgM
7/M0W5UfOCZMFdKSPWpd5mP5zp+VGRh4CfYXDBKkPV7/MgwI/UeJH0GzpO5pXLS0xytyS+HaZQSb
BH9PuwYfJOj9L6R3/bfyll5YsbD9atmHQqCw3WUoUyPaF/aC52LNNHD7H1sXOKOE4ttTke2unNiS
4Su1AdUYeTlG01+U08Rdddlb8fXYe7hUTZRZ0taE83EYSmXAS2UsPNNusqiiZRLSODNAIsHzPTnB
SbIyVPfvsULvm00fA/J+/slt9NwjAlQ6SekNT1nYPBrxP0ZelobkLvnaJwgsZ/xyoMOsVTMbLqtk
D+vT49UF4wdqiumU9uc2mQqbK1NX1i3cJOTpEdXit9yxAR1MJZU4c+3OFUSqSQAfBZtAm2s9bYle
rerRe90FQI0Gn3NgIERIOwzDoYois6sn2Af/KwAIWiyD779OabrWer/ne9SUtIgPnyzJJFOvxQsC
v23CgtmWJaz8IHuBPlDqVS1RceNxKgOyxzzjW0BgWLJYuzA1eSdBgzcG+LCd9mC7WNIJYhc0oipK
4I8G9y0polM0YC4iD8Hg5ZHV+5Zd6hknv3rmY6tZTg1JXVgInXm9W+a53NTHxELZNgOi64iuazMc
Obyy8R/4X+0wbzXPjcrnuIsJjD0E4x/N+vBNfx6xhkL3op9pvLmn0N36a280xpj4xonH6OnRgZl1
z2r1TxiLh+FfQ9mm3YSELu3hFl8oxfIuFhGwFFBMdudgW5b0DGDRtPf11oWtajiTWWSE7LCY3OQ4
RuaA+u7ouTdNB/6Aw66eJuCyDEDno8S4mqvGHJdXWxmAaX/sJNIxYieV9Rb65Wu93XRChh4nT3Z8
Cny9EV1QNtKQwAAXMyvNDPC8nkwKPU9W0lGmnopHUuAht8d4LNKIwr/6rOX8uWH6Kcdjm4IUSjTY
2th8YcvXZ3uFj6OTbPywqpVtYAlM6lFIqLRXTYVDvBTUHcFgR5lpPOT/b/AKLqI4vAyu1BEwXgMI
Ib50YR+WIGdhUTew5hV1wlyJ/ugpQu9BTw6tVe/5UdpXuZYFzmkoHTlBt0vMRn23fvoceKEv27Sl
krGFto1BF2zCnSi3Hp/jeMfPGm2RUOrVCnXzQRelMYADN6lxPMryRVdb0Gfr7z3ZIbsLYHSbk7WE
Pju1wvrTAAE+R1YCv/n8NglwV6SbPD6Dd0Ay1xA8rYFzvJzwBWuDcbc86ptwM6zUXfUNoL7O6rKX
RH2QlUpQWWRhMgwVgDvaajzLlnLlXP3l020kgBjwn2Yw/nYtfRzgIa/TPbx4YTtSC1uvtCpijtt2
3zVUykMOqlQh9B7eExe91WprNJ+yOu1hpYv6P93hUcqTkJOkM8ASgOBMvmNjYwEKhBRJdZcny1OB
RQr21JZCcQ4Ld4S9slAUmR5LVkcfDVPInbYrl2ohkSBoWx/0a3rJvKakzpWtXP5IxghjT9pCo4a5
oeIB14c2ypW4y7NZREuyCvP6SgMNgS50jsnhD8fKtqetXkmZSzSclL2B6RXPtxxcv+cpaLXTEz47
O9S1wZElIJIzBCkGqaO0uJptka8x5mbQW0YPAsDqOSztrj0He1wAfbjFaQdMNl2ydpu+b/eK2660
BEVpg7/c0lqaobAWxYpvpZepxD3gkEPnVMW2No27ILqShtkhykHopyIP1iF79cgRvowwR2a8DhEV
XKWDp63MihNL8A+j37ydDon/LDdK6MmAAwANj03xxTx+5OinmrneiXrKVVvXubsZQAqZjx+QvUvW
3yUuY7hr8FCRc91ia/E66ewA9Xv7JT1gvZqM2cJN0t52KHRW5capGIq1YotMGF+xbpRrwKxRxkOU
cau61cMc+OcxM6whEWHeJzf2ZJk5NVJyqM5kB6yA5tSrIvfQ48vS4FlBqekfxb5CJXienIAjr/MM
XqzH9d+4XNtaPbA2NrseSjpv4sfGQb/YPk6g4TXxk1Zv9VC5moyiZIzYAJpsN1ztv1pdiJ0hNb7Q
M0qushDT0arQ/eg78bw8Pg0Yed3I1JPxY7KX56pH+zXb5KsAyZ8x+xJQvtPoGCLrnnPg2ZW9sqax
omlzcwXQ9+zisjt0uixHtshweHlgaf6uJZFCyIyVa/fUWMGir6QM1Ijrwe6TmC0ie7O/295/om8o
UUYDnpo6woNKyNLp8U0PaKM66G0/wdhNSk2GncLydzXBi9fycHabxBZrJofcFbrHL0UJlNckNYQq
U8lgry1/6f5SbGGPqZwGm+o+YfIJmZgjVPYvSEmE+L0pye0S+XybYIUQP1HEddof8pakcnX/VlqE
UM+BAfqXXC+ME+raKS4hSduGM6HJ8vSjfksh7TLuYhv2fOMnvrBzo3OvcsSUQxB4rx6osGwYEnt+
JK9I0cxGsODjZl5GPGW9YZBzpmlLztrkiT3XuSjepV7afyCrBPy1NPytJhntZ0cHJVuvFdvezvZg
3JfXIEpeM2lxbUYp/aXgE+QxG/dVd8mi/ZkjvdJcVY0vmt28IuqeuJGNSvW/J9P5bVgXotR2Vgl4
wwpdOkDy77YOU5LddiiF0pNKjj9PWNagn9hL7ftv1jwg1185QGf+iM8fo/kmJc2jdNt4ML33Lnct
EgE2SkwQvqY+dN2qxjqylXBSH6YYJUZMTidv+pJKU1G5YF06JWcpWS0ypDzRHlYw51hVrtXwrmU9
H/Dxzbz1ebkyQv66z1zVWkxS1D1fyFU9Nd8rAf/guRbjlDCemTYFlinCcYmh2XqzO03x+B3MdDFw
Lc+BA9WzmAeVPVlDHBufoVX+N6dn1tUk4UP4YtRmbnXbJpi2bE4mZ3iViUMpasWmEezspE11c4i1
qoZu2TzgGci27RJx/qEOONG4tBgy3e3A0TDscJpYbIgpX21Khg1jFThEsv0rj4zWGHI3V+M/GYD5
z624LlnJNCXSq1kWbqOdsshcsO5dBvbJD6j3Kxo/zZ1SeZHHqgWMdwlxsna0LCIZAEJCTT3fqXqq
Yo0D4ZXdj7/+LtFFQj197qWCuR/9ULo8AVcWokJQrNocXohwv62jF3DM8R4hGcx/oWIKAarVSsYC
Sx6PaqovC2UwgaAnxaGvWgBOm1CPLHiELHV4rx8lEtUEYawkPA/FW+uWOPP9ucZqT1fcuNucISAh
xVPOg0E9NXHvkDdkG6IvpzaGrHCtFXlDkuak3lqba9/pOWEVjEjz2jrTkAwBDKIOlhhHChKJCeKD
8QP6YBubTKn1UCrKKX1sHg0/vOOgfP1szB3EEkUqYcbxKHj6cW5Ui+t+V5udKIPpgNTmD3NloXho
b64ME9qA6siJfFSh19lgwDtWh3z1jp3Zwyred29Pd+saVaFZVcDEvtNgf6eZKMPuKWeZ3GO6aFB3
pim6u/RS73U9/Sk0WCd17ma1Gz9v2ybOnA1YpVG7h4HUyKFr+z08O+hNekSr3WLoqFuxGcCkGHx4
kk6BiuqHj5as5vsaPO9CIbrSUFQzsg+nC6eK6Nf0hGPOtlRHctiyxGnIacrfyp+f5lFZEejSCSJS
58Ty4JUNKZ/ECDF4VryunCAKE8FumBEoEH/tCdZF3Qaf71XZwqETLZI+u8O24QzNqpBf8deKISiX
EcT7nkKBDTBV589CWg3yoczfSp7EtQyjSz2bDbK+2qDGAwtOFrpOBX7lDalzVZrgxy5T4CMNkQdZ
7kkiERQ7D5k+OpEHmC7dPCP7Mq1fWuXaPBItHdhOSsmZMRb3n5hQiNJZKfo2daPWbghG82oqwaSg
SteqBsnsvPwKdkR/PZpmzkDQNddcEWkgRWglNXP2JDatKnd9TNrGOEI53QO2iYNdL1MPSDlzj+mb
yKUNZzoMegvEbVxRXIJqpL89wVjfEjsYb8eHxriRj0Cev/oNqdTlUOJUBL38GaVxqirmF3tkKzdE
kOxYtq5K9Qc+mgMsLnJnz/0AgUw0ecyWZwnBNSq3cZFxObtAWONckF4gyWFSV2UN0mI0hcif0TSo
V6G5fYkCrOrylAI22M2h+ecxvEObnTqN/UdCzzb7HkjiPDCRTd/5Idr1/G7hILMBhyU0buH4m2yE
U99BRYvIIVcnYQso9HIYhEcE7haTR+8wjt3LBPN5R2Rk3yXzxXOZVzRFHQMtIeuAyutCSazKK+Uy
kR/jcjN1ht+QpsCG4K5xcJx1SARpKjQdNYVM32Saxfb5LmxPBEKzJjghbyDvh1Y4yXwNdcK4OdGD
BjXJ//fKDoSEuCtIrqLt4vwXWUJsTPsbUmC9E8eC4jghxqC1RTvgNfx93dQ9tH/aBWdSxjBQqzJv
BAVZdjcXk/kfn4VcWlTZw9HYKCjcx+cCfjPNdPnfdp4Wpkd+bNNVdyrmAJwsK73TJHiXwpHQp9mY
ZAI/8MuFLsThZ3K6KMBloPtzN7W+3mIaHZzmKyMGwTcfrX6ZFzM8CkHBVIGZt6maNAy9G17kfIdF
ym/u9J2MEj73pWe26xWT1Edz8Sg7XXfEm9HYHOFk1+6scVGK0LqBV5ngy8q1GEfH4OqVbI+FgfMz
KY3zPZuxIIxvrib61JIIOfEoyRoye2STpltLWIbyOrOXsiIAqA1c2YIgie/xBA5F/BofDJq11M2z
VV8hSxNlLipkvHjkjkPcJdjEE3uBj+/dYdfgvYaLOgqDIofrSJSKw4xEM5q+uXB1bD4+TQhlDIsF
EA6z81XQ6B6sV5VE1rtJNsrXp5Dd1U4tKYvErzXjRv9zySyw/EkIgsJcWCTFOd1V81hsCYugZvKM
Jpxuy2AOEyznVSP0OFGfYBckbbwnTdyGSw6h8aUgC8iKi5jeYJLULKw8oQID1zOq11UmYQtJvp88
ie/itJiNXZGwA60RSe02pwaen4IBZFsty3Ld1jiiap/yBYf3FAN5aVLzJMyrLpjuui05NAStweVG
mf4J3usFIavR4luIy0F6O+KnhGk5fmfwyHv5AbvdqjFnhRxkq3Ze9JYquW/q9fh+1vJMVLuM+FK9
1G+NnQkbNrZECYrqSu4pxV/vL0XqVh6h2EaiyJepB+iyygQO01Tll8B1IamyeLXzX9lYquxTXHt6
P1wdgeAQqphWCu/e/whSTxDE0YN/7sqgPlzwtXO6oNBSIPKkGrZ6vFuvE7lu8mixpp72gtKCk1Ai
5fFr8A13xWMDj0OiNgE4ycb+xXzIEjebTAG1tLzBuYYIA3exGC7x7PbvDYYwPlxNpzrjAhijOxSG
2Oq0tH4uxmlRBjh33pnnSwhlXJQF1qLHlAkhlT5qcQlOHLqZ+METx1WrBxRVjcOJGIcWes7XQncU
wvAEPU7gk9pvzof6f5A8ZdlAyeKgL/krTxUI1vu92/DdfUeFRVZVi66dpHD2tPBoblwBKnqp8m4c
6foiCDf0BfgoELW37VDTLWfsC9U0h73sovXTIsPLLlNuN/oB3XCEKtS/gtfRyLothzMNgs70+P4F
zS/1dIaMeeIKE4DcUwKieyd4asLNX9Hd+JY6d2FKfbLvOLoaecrnVTXydX2pcB5+7g5hGXWF5ePG
zfllsjJzsMSAdXWLLs+1AM5eLZB+RDAFaY1ktPWBM16w+hA4+fQmzoqXjzIeLs/b6MjdO9/BM6hP
kvlJ6tV7VfCCFke/w0ItIvFvL7cz1RdeEXdmDCkn+ifqsk4qeNoKS2M4ajNWjVKJU5ZkgGeswpKP
oeOTSEP/AlhUMrBskoFOxGD/jzGL8B8/CbOLWpAoMboMS1YWHEbybU7RRRxIQR8cmAjPmOT76Vm+
ZODV4O5gheczMasYU2+r2ecisu+YBWrF795TC4JSeOoHO7C2clxk2tsNzclblw2bRbbfnDpgTiWy
mj8RvJE5XtzAPSRz0P1Fv8vJn1fO4SnVfO8dSY3iN2pwiLDZS3WGJ4Bpa4W4SlzlJLlWOMc9sYVz
QGZaqMi5TmYP6ysMKEvBxrajfT7z0RoRf/vHE6shTpMBrbr8Ddb0Cmn+Zj94McwNENmRb7sD6KGe
SJUfjf1xRCnNn6V67JA7gTEYmSoZMZ+RE6o1HktMVWRMtGhVY4NtLALQLjOwL0DFEJb4805PH/Fg
aLlfE0NClhP3Dkk0ThEMvEWiEt/EmpF3UsYlBaC2EIwEkXc4AXpxhxMTlMMjwAmR8C0BUhVRf0Od
2ijPOvLTCvZyZWuMu+4hQJoQJ5FiHVUq5+0vJj6nCfbd8LFFhHEqLHs9jPToamjoPIBj59CKO9a8
HkIg2A2ZgDKoG4OL7Lu/Z15gA0f+BT7oaO76cRQsGHkgEgLBBqC1n3P5CjYbCSe1pyxhOLaLuJnI
VoPZ1PuVNU0Osve3nNqVUCxfoPENsx9u8GFFHBe0opXxbn4VxTHhQW1YXJ9/S+jhhst+qK5faOk3
LRTJR9VSzoS+djmRzVqua5C6zuGIzJk3fSEA/qDVvX50dsDFig/FMxbd71SeSDWHVsSkyOrSF6E0
QBHk+RL6XS2UuEST9t0UtxEv7KCv2UK1cHxpuGOYjfdAot3c1dL+CHggnbux8FfOMlG29P8dAw+6
EqKLOnrjyYXtapj15lAM/WWdhIJwKge9voaddu/D8A8isL/csekZgQCldpvkPx72T6klqRqvEZvv
1KGPvFnwsDSCEak0HuBfinSuitJ77zmD18kf6EFI46pREv81YQgC8uzdLdXxRsn9ec1Ml32/jXDe
TrdLu9d+7G0QzB1WJh8jmThWpZxH5bXHp5hg02x7elcTvqmjFYUffRRQwUgT6fB5+bviVmpXV1q6
clv7T8Hx/zm4MH4EzYx9v90ZIAoIGMZUQeFWzzoEdS09G6IOPAc9qrtjt3yhC2rYAIv5nafZRPJu
ThrCrNrTsY8keP1h8vkp7laKytaZRPtZrKA1GM1/3vtrQK60wSWMDizmC2xcrkJCWyJ+WvK37fqD
XITWj/H/OKCtOOdmZ8jOebrfuCcHwLc+ij8ISDxK5bWWlCtuYEE/4bk9fegbVXD353mISS/zj3cP
E6AJf8v1FztT8kOdPn1CSFRVzYGHhj0UFKHyYrN5NML1GDEN5RnPsnYpf2SjchgQOpwo1g+KQbKL
aZJqn2LUtptjOpNYqkZ4X7s4cTLCjQ2YpHhr7AEfUIs/44J4AAowdUVf5fs21w+HPD2k9HEcZWUJ
3xLCYetEOkTd5ThKtm788ym3t+fpeqnWpMzAgCNfUZZEx2C3TUhQJUli9QaSWaqvksOOK/1Uet7m
uPAjo4m5nm+KHH6EXk9QZN/LzZbFEXvFA0m+3DP3xOcYDkghunzfXlwkhk76XhUqup9+AmflslYb
766J7u9ylfUGDb+xoChuWkzs8VERCFMlpr2Yud1Ezql7VcMfT01+/cT7m7vGYdhFhPVy+UuyKvnV
RvHwDcOvnzltAiiGaC1yO0qz8+7jNXeq712EQHIL+A6lUP+HtGDdXtTLWD665Cxzb3XnbP55IlQq
n8blmXl+Nn7SM6077CRpdP+SdlbhVQwvHCTlgAT06BDH/Hp7NHK9txPQVhloj8cQuT/DCRzz7Niu
u8ygFJP/ugdrR3l2KkXP0IO3LJcRRMnzBfK0/XgJmSBQugrxK5IVtNOQ4+1flvisVzemgn4Ad9wX
+bVhrXDATEki8h1U98xbP4PhDz5y4BcyrB6QIE8yhPJre1oz3yRGnZ5XxBHdGm8uy2C+Ag0HLsKN
IAFcz4fFqyxqJWEbRPAlUNdN1zFmFHhLr+iBkXRp/NpriC0OKNFhsL/tsiOgGbyxsVwkFvLpdj8o
ZgpTuoWZ8urxz8hue12UllsEt0fbjA07YrPPjw73+MBRtqcnwGOwIaYWdgHXNeuzHEEySEAgHTPP
5/FkU9JKhRF0HKnIHDW9d5iG8AkTk0hUkUEigDBIgJzIXtI3sypcnam8r6ARKy0o6L54JknVybFV
7VQRiV/Fg8y5TKe4Muaj+O6IMLG0qm/t74cFiT+zJFORF+75E7V44OfDyVbT6ahoFMCo5emoy5mT
Z+3CaigYjuCzhOTVqP6Ls9N1ri/EXJeUqA/l90xcngzZa6jyy8wlzZOpvpAoUttSlrC+kAIRc+TB
s5BbhVTueZMtgKZ8dKUulnV0kTKQzmk6RHUK8qscfP1w3NNSEyXVlLFs7mkLTEj0U8r0k74s1L4r
6D44ucvV64jDbEcJ4Jl/GzdPORGW0hDpN0iXjyXWnBmf3KpC5R3hUWynw9qJ6KvkdnlK2K0uC2xv
8pN3yxtSLd9vX1b4uLKa1ruelXZWHxnicCDpNWH4gXZzEKsmq+4RDkGkVZepqMm+Vnd58NcvS3Gz
+u4IeLHtl7UKvwdUy6VRohV7KWuDi8A2C7zQprNbf+FwSobQsSLgUjrA855B9q8rr/38saJdahKV
wUVgxFVUAsLOUIpqe+M2C/WDNm0D7gIMOI5vI9/zfU4P8YDS6EH+KCZm52JTU6jL9VZWcSDtWk9T
cQtc7ldpczEiQMKfMeeNfSv9l9fAL1XjOh4ZYf4MJvpdv9/RMQRP+Ek8BErrOqJNYPcyFo3RUi6l
Q8XDgFk3HrEpjg90/UemJ5IZxxEVIycO6GOXI6BiLlP4L7YmNOjh5S9Od1cgoYPrdlSbPqvnA7Qp
g75oa07uelpF6YxHaPWL5Ge/cxs9iOc3hpnk4kZ2mHfKzrtuREnPFDQ7h3HHXZzRUEnCl9UY734t
2kBhqV1yEBQ1RDRhQPJmTLchRIN/AZG1PpclYA1hvznYfw5bqzrYwRFenmkGywtgNuJiFLQy2jD8
KWW+gm6otP52NAhedGScAVTVuYgfuaZigMXcG+xJzOj+KKVO4wKZA4VxfsG92G24gz3Uo4dvdORq
/+Y88EQTKeStDwa9MgUxWoJuh6Fj8f93HP0MfxBONgKCH331vtD+jk8V0cshIgfFcSqmLX4HyQkP
UNQwq1J3ERsf9KFTDmJhpeoJaTI3lNeCu7/IXUWnnvgcG7fGXmdcpd8WctyCHLynlt58z1n+6kPw
LEElRzt9J+YXQ0qxdnxQeEgruz1LnaoVB+dR/GP6Z2Wuk/xra+qPz86pMD5m1wvhs6bUZdJTAsM9
EALyGZRGqoA8g4cJoqN9QCSJM2lFQm9jyGNPa1+5oQ6MCzQ1XzV9N3ru2wT3juSvfu8e4znCgzIR
Th/QjOr//yArKE5wYCXwkWZiJEZfWq0IXwPXe/fhWPHS9MNuNAjM6wkWd0OXTWUCE4J+Sv9znnS1
5yJA7YnuAHmrhE7i9N3X355CCtthO7wG7dmnkOJ9ecDfFE6PFYeKPVp1uZiQX2pyWzGuxsheO82w
8tfMAWRICCFZ5pzXmcZQ8UntB2RxkzHP+uDHjyHJSR0qaxPxEtcb81KAg89XSSazmmusTAhOdpCZ
w/Vn9ZXsD9KlQHb6l+vnPbKyEqJkRUYzc9kaSgF2fEgmQkI/sjODHXHi9Up+S5NreRBrL5v8GByx
qtchhGJB7NPEVJJBcGXugbes49zsdvE9mLxsXWRhWrbbUuU1DwHExOeyCgmndWe8lf5crnbkwNRN
1i/zRm3cIRmPxb4e41iR6baBLVz7Jfilna1/fP5f/mSD3iNh6uJ9Kw3a/JQk1wbaeUyAz3/SUs2/
F27khj5obUma+JIotJ2vqiM80+P9ea4fRVf6yQUZz/aiNNNqde8unfGzpxbUx5mO0kx0CXkodt3p
vD/i4y1oEunsjVkeQHcwrnb/3P7TtEgMUpgaopsIxZGSMXRgreCgYfq2LTYX1UIpn5zV5sbveuOM
9yME7hkT4F8Dp1kt7uCLdzQWT9hkccrj7aP/+pJXxe6J0T63+5xLMTU1FRU0tUW/vA9f3wNgQRZB
/FqeGP68sJWQSYmHapM32Bt8tAxcg2yxYWRjuVacdRSnsQbVTwIKqBBGwELBABMdlz2PXb3w28e0
AEr7oaIwEgwa+lJf++ooWFHJcoO1yvwMPotN4zUc4OnfRMS0xmXHPjbidDmUApusAY8vETDITe5C
/ZNvc9NTZMqD7hjZv+s/DRnQNBI840sbW8838wZcfjjydMZ+QOaJG0hFw6eR2IoC13g59x45mwLH
Vg2i4aqeXaXwxoWmjTGV/AdtUvcGoyNJZ4aq+z5J2FXAniB8y/hoEnr9EVZk9vj096E4YSEOZCIV
HM7BmuKIZ/P9dgIZ39NhBNu1E11Uc+5XgE8uFStFzX1MyRJSHhW/flMkYYG9KvNY/qX9yMAYgK1R
niaaHxqUKur1jvzO1vzhdCFCZQSKP7MIbSM9f0NLTKnbWdWTtRJN6glaBo4XcEj9nl9/UNnn3S4W
7RRnC5IccrjGBa9PuhLgzES+BhZI8EQ4JUw3Lvlclu2758J4p/fqZ8zG9tMZd/D3vuUTf3iP9/wf
Rm2xvDHSwAo/prOKTXqxp0bogGBAeslaiVwk6nEKLO1BJksvbJz95WbgU/ZcQDQnzZ+B2RFaBxHR
QFBTcby+sn7X/TnYcn+0JvWn5rERngbg2ftXDtSPXh1izOQvUxn/ozuMOAONXD4PuK9K68kw7Mnt
np+49erfA4s1lH4c/vU2r+aO56zl+OQT8shR3fRC3VPp5Un4AcSFrv3t1cHKyjPSl5BJ0bb+9vB1
qKH4jLjCkCAQYJZcUEL4CAx/6EtsyKeh1gpO2hMwW6ppbfQ2+Um6dyI1mbAC991XyvoeXZMVwfeL
qi4O7IoySJB+ugmfkhbCIcqNwSwvV5AUmPhbv8dahMtPjvTDRNXoFl/CuFAlM3yrV23WqkKGE7Ji
DHNnOur07tjNR3KNc450SG2dTmGVbmIobmnNC2jRFwgire8Uv+MYGQpnSKzHbt99nE5ARNYyPAXR
QsvOynoH17FuYIks3Ca6m6duedgaMYzChRFuILTAuLPCya43dYGDf7GipzBYPuGaB3X8/rcaI8FS
hV3vEeiLDd57IXRdOGjTX8FZ6VLluzbHLEWhcezn/J8Q8pHh+dVTkN3KymCnCu0WWC59OpghcP7V
UjYXw046yGpNoTD156IieebgenvSJonFVU3WlVwhgzYvuzSiFOs5laK6uGZKSVyw5S3vyxj9vB87
D8z6/WwMGiRu2q6MDv810y0Y7AvV8OXIiWtegGdkHpqIginyNLmC5q9q2z199FK1A4aDdBbjv6jd
vwnbLL3UIZHOpRXFSVPlBLU99q231oy4JaomCMlXDBriVov6TmYhnUxFXTl9oUlB7QDptZ+QlYHJ
Z0upju9dHoXD4+6itgZt9MEbwQ4QN4iMXyeKqH4SX8kj2fxHRhxUYZQaG3yiJH9OQrM7+H8Dhjzx
Gy0FIKmXAtYjrUUD9u/NZcxUdzkdwL+oSchJQnY/JYseE+yEXkKn8nbnn2YtDDtHKfyval3d6LuO
hvkn0xdil13hDQ2JZ+sfQGuiUhIQrly3LePA4nOlIB5VArD594Ll4JHJn9MRkkSj3XrOHle1TNCU
FkOkPm/l08Ziaa+b5x+Pb2Dho7mYDf+dywNCeC/o8Yg9fgW8qDD4a1B0ZTdjSCkL7xnqF2CWMX2d
8eNGwSCul3ymICmgV/pMPGHuS3juIzby/CeqJsMFZ9vFrxh0gpJu9oXi9NFf5nE7SLEonAkdmmsE
6zAb6raFBVnA49s4kDgfkYUTOr21l1XRJ95PeotmAIAVJdnU9E21QkFUW0WD9FY7j65uddVH4nu9
XgNbxNvlE50uthPWIyBJNTxcss1yY0KCgtIAkZ3VmS0jwIrzP9ETuLa5tzCLc+E1HY3yJGVA1r1U
zO6Ktc00STmIOajajK/VwnTMUnEkEFSQFwkSyKbF/uDNKdzaMqsXfENrhDbJfY5So/pz2JURnktF
HiOZzHhTL7q94eHj3lNbI+On8bRo8CtCUOqlyiLxhFZD8r5tJQm+TotfS0bexY/5gs9sKAJuKOKd
hbRiwNm+ZNdkrvvWJwnZChfhovwu/OqjVazdOcygHeJUJx/tzc1Jzgu3oNIN/DiMCuRZkE6BAzme
MyZpDENRFv8JndMrQJ4+DCCzzTBKv+Wr5MUUIDmMZXd/0P7skOOOLSmqKUOvAvXCywIq8Fgx8u6k
wQIWyCdiEOasB576psnFsaK0AgnTf1y72WwOlCY28PlaBRE20ta7FpSCWPFgEcZIRc3Ap1LredpU
yUG3iTiiDFz0ZaZa4HG5kToLRXAoywovBoBq8LIXO/7t5WakbKNr04+9BgBwpOq6xmb6IkLhZGzg
MNTySfmXtbfB1FoW3KfyMlZ2UKTJhE7XY2oetL1tYm1O4aAGyKDS+m8QjZI+m4ZHTyIZSsErjOP+
ncnpfRyvwPoPWG412eKNxUtRNH2rj42hdocor384xPjOniez4rsFr7GzrQQQxBsREEBo4KoDGAX2
wWWP0GsZtXzEPLxhvJOdlRhnXYBYB8Qn6etzYMWM/tolUMOKVqiPhvjW5WGZYE6tWJxn5F9MoVDw
62+isWSp2djofv8hkrOIr3U/IuWStO7D9pSK2ZWF3mYDm3vgpc5SS1gBnEYkp80nTAJF6S4AV0px
l2vrUo3bCm495t3nqleKx81YSDwJo1zlmjr5CVo9pYVN+nQeSsOLwOclnpwqtEwCIba60zrhi2Wl
8Dva59k1JMIYT/IJxoDfIrwRfvvPaUXxzmiD1Kqn+QTkPX25WqkHLC8vwf6fcomUAox5oOHLQb76
iR2WCIUqyJSfLM+fKlEzdEVHssdluZ+S1IUqNSQPTvXJjdI/i9YbXRceA1QFFX+Y3FpKqf560j+C
pT1+camNIMpL6Az3hYgh3fJ5vEJYAUbgGFbEEA02h3q//UWp9+ZPGIV+XlVMXXFEiG7HXdcNtf+s
cxfIyWVIwg7EqDqJnIyLa36vupnfqKuvx92xUoB4Wax7vIj/LwdHJP5TTG6OQCxkePnRC8JoJ5q4
CC0RVhGmLe3NQFqtDT8r2pbfyNkhJjFft3ezOC/BkVGOaAgH8W1ltt3DXh0k/fZM1WIcQNBL08jO
lIc4H2FIfpbpfG1Dui9x+oZdTNn3NDd5rtjvZvjsqa8mzS9nyCGZA5/V8q8Cyq7+xJKRiEZIjHUJ
UfAmzTkErnEklXqKhij8MiiZbfZ66cf/ewF/5MlIOw26AqFtt4EG0TGDahyY06OVeQOYOfIm/KFt
sTP8hqT9LSGazdYUya8oWb5JfdC/TsMB7tj+hD4jg36ktTkAGgXhprbqoPTtWqVSDdOlLJDMiHO/
2AkzsTJrXB6dOdNcMH6MiFi010Ec3aRW/BiLZZuHh+sTUzW2anqmjaL0vV+emZM0h3DhE1I/WAR9
aMuVz5TobCPFrnCfI6vp5hnRxMdEjv96qRVRhXa9evibDQgDq+L6nrfDuHWLeNIJgTn6v2eVptV3
R7uKvj5TnFU0de4+H3MD0bKcC0jVFjh/ikUH9QNewHUqRBDr4KzlgmsyGYK95ca2/U3re/Cn9mzV
3idyHsnMfhWAgqiLcGbc6MFWD5fmbkMUJFOiOLIhzDpRSuhaj9oz93WbeBaThQN44gRy0LSLlL6B
H7JZ+jay7RJXhJaooOWf9ix375KPAFMKOdoxzlmlbJ/4HNn2CWsuprgmGCfH7bXevZirA7z46Wpe
79dxajYVK7FO4Dnxg/PVm1w4rbkgdaSyFOVIB/Iq+S6zkoOOi2nv7fp1879dAKVQvffI3ZA0hO1q
hXOLm4To/F3DCkAYMPwtWn9mIZ1xJ08AiaMg2kG+5o6liGBQ33cEwmqc2wXZ1t464QW6VbNGOC8l
MDglN1SnILAM74+3Dc7XlZyQOCFE0znSHBf1M55KawIHWPPWvjOdJK6OM9j83kgEQQjkFMpuZ/yX
jbFGPJc0hp7R+L5bpUFTK+gYXmOABtq1wMn8W31ipc4jRN4FEsvDGJJ71/xfTVARlEWFAjcu+jCX
C+Uvz+xViYv+1Qyvd7OLSdUlneR3mvl7g5Gv8p7dJtu9yTxtZxj7jYf4nDVGv4B03wpmLUvx0xQu
yp06xZUDoZ1rrJ34GFrlT7DpM4ZUJYIgw9RnUvEsfpmhmV7yRWaUekhDxDjdYn6M58kXhRvtuVf0
yxRLWvTy05c3k7l+Fkl47hFmzf5IiNx8dGZhBDez5/uP8v9np4DNmuaJaGywW2P3vo7vSm3WWkR+
06mX0yiJWIbW9xgmD+Wqw5u6hBycBn70YYJOnIu+qf0NZMDXcYtFZvW7xskb4o60CBRoEMsMZMFl
xHyz3G9553JhZCnsF/qsHAwQvGehaIibxljmP7hBV/E1cdA1rThFVT1RduIPXYKVlqTIwMPt0Nje
cbtCsSndU3PFs6deyIC4YxtcgJNWq2YojKaBddJZTA4k7cfVhsYZhtQ229zADfDoy0ivYk/srNDU
CumjeAfK6rPw/MhqItCHBNF4iWga0lB97xWyJKvF78BxAOXO54i97csg6dgEA3EoHo06pzkTf1Jk
pVi/fmKNQcpBXXg5FyARZz2nlKOQfgCBXf/YeMKKmD9T8lY/Kv/ad+UdfP3r172qnV5jMLuHvMio
lk4q7LTultNxBsnKgel161jfnFrXfaf0fNLml0BfMjjdk55DNFlHKZDppYcZo0w6aKege45YOZmg
O8BxHIix2WB0JNC37kcjBtb/NMtH/pNKQVng1vV7mCX1Bc7hbp1wUXxOHUknerzmrebdDpQYqXQ9
lB0k3UJ/i07ov9DsfPlJ+Q8zWko7Clo2rSd69XYInqrEIeJf4zMLK0GAzo4GAs4MlNikuM79IdO3
rknqElPmBpQQ+pnuRicFAqTY73HgP225ZboWJkcRm1BabKjE1IYyG/DJma7Q8C/LIlhtWcUQw9sw
X2kVBlRDSlZiNLgXIXl81axFp2tn+Y9/HQ9TPgRm2HLyzm1Qo3NGqlcgS9AtyJdth27J/iP0OrNL
jeC4ywECShYFyiLKEJCSnIBAklfMPoNgXIjYX+jBtYYlUtYwETHY1AcENrZROH4xCVd0FA2Bo71o
mCly00b6nMf3jmvwloskJ1YwKLjfOX8RgcYXIuNdti/bzE81781mLsYI50xiiSMBzcARI2DUsoKy
VBi7EuL+GLwuLlzl3YJszd6MkKaJW11IfUFDb/d3oxvAUD/GV/kixbPB12yaTX8kHx+/g1pR6NEk
bZ7iZrwdCyGHn6KYnqkNHOKUJze2BCQB3rZYm2nM2VGdJW0rSBSuE8SSCyN+pFJHMMK7OS+7mzVE
kYE8XWPENaBCr3UvR1kSQz94wSHn93W6B4X2SNS/8EhkqFp49Uxq9EZ2vO7/GCsdTKXYAyUVW/y7
yqs7HaIsriwuqK9eku06ROuWixxxcWbVeVBD3pcBuNTT5eF8gGRQPKfWRTtT2Ygk6dsdSNN8UROD
j9tzkxFZeV4NrCz5wwD7pI9eaKDbMkUF9VCWqZfsrYgJDp/vY5Vfjo+S+BBix1co4wC70AoXudcE
joTC0QUt4wzgWij+werVctbasmqeJN2mwe7RlFsKn1OGO6RSC/CVvoHdqdtvO5UHYevDbG4fG2QR
VJfd9N7LdV8Ezq3ZFQ1pZuKgYsu9e+Hjeyh8COYHCMdXKJmvdo+GJCk20H5pOa/Nud2eNXwEUbOP
n3N5cD2mx0xArXg3xvs+DTX9jrhV+vr6nuNZ4Kl8ymDP8cjb5eVUUHC9wiMkkjvCuD7fF8RefWlU
KKPAld1/qG53zMIbz9uZvA6FcwO7PxGNjxjHTFV3gaO7sD6J6mqiZVVsPByqUq7FVNfnLeiYqkHI
QDmD4vkbvWrvsTMp5tM8uyAHIVycJHZYUC1RgcJCkUWvICPMrWnCkoApPX+7frt8s3c4N21NhYIK
d3ayyF7DtgFK3smTrfWikQM9Vh5RX09pv1d1swF0IPWUALM5XJSY6lrX5VmiSfOK7bmj/t8rPdP+
RTddptQTFYpOhZs0fJj7jJdwWyhNl6MFrdjrzl8Njx3p8kslH/7vDFm/YUyM2DcdB8Nooo7v9EAy
n394jV8SvDKl4Se+2RxoHYNWyT5T0LqjCTN7b7/13i8v/f7/Ce7apHZ1HEeIUW6gapzrj69dwQOm
/8BXPPCbumogEXXiO3fWe8NiXZ6GEG192V+VR/h371J1o6k0ti2VR7wV1BkL1XQOLHN0djrf1aP5
6JGhMCf4EBLcB4la8SQ7iUd5R6dHb0WcTGU51/nRitJuwgFHfx98fcZGihQP+HIUHacSWJakStOV
mM0M/445theShkeoOorclxoR1AAk+Hy+/kBqvYPtvoe6+Uc7qSOUNBSW0tPLeNqvDp5MwoQ0tTpH
psULVzAiRX09UUphXAhb+j+Za+2b937X2QRbjgX857iFYyq4Ln0/efIDAkQ88NCHPKLTTXvOn4SK
lSLPZ13uOrgfXrNBVP7h6+fkb7PVKieXMTcytl2NxyKqpvKGiy4Fq3i3UZJN9okkGLYatL1rIozS
IoaKD2JxHxb/ivT1e9qgVZj482+6zpWD70yCiWpvCvPqFnHSJEEuTyT89APNGjEklo2VE27VK253
xkdnS/V1oz4YV5iUZJdrmFEtjdq02BE0USMB9Lzy3KwbHqdy5aNOuLY8j111pVrw72iYKiD55Rzo
9vy7guCUNd8D2ZIddRzNOA/DJZVrsCk25KAMwh7Ld9fD0BlJID2X0CCtOWnO0UVTqNnqbcSZuVve
Td8uJRtDYiRuaRtPpPoO1Sl81cFCtaWTndfjNBvR2XqpV1NqSDwd7ToUKQ79RE53Xn2x/ArAuZus
xnXytseHJ5G1n6qGuHk+h/BNNMzeragSWHvE21y8LHBm9EXjOfhO+J7YmjY1Dpj4A0R1hv/aafJp
PjVcrtiurjygV+kiRBwL6Y04pCAPaYNIRf977N1cnhEKqhj0P26Zy1HZgAwu2M5C6JKspoTuXguO
wmqAs7i+A9rkHuotFEK/pSVgsNfxoa93AXZQJzwsnbNPFrTARN2gLD2T/qT3c+ve1NEZZYx76Jy4
jsWTXQ3krooizA19LHFOJjJ7EHhgj3vqz9bgls/BgjmebjcK3KKJcBVBqmGcfKpGk/lGy4dsDnqX
We7iCd8vFIZinJQXMbMjBOBt0MS4fT1NQQyJD4vGH/dGEWyu6uRaJtSsmGxzAEltbR56HiE8zpqN
+msgPvH68U7M2NckNudxTm5LRTkjjzFbZJLR7rZ1bE9gXEn3UZIwkWqMoI2BrRDX9XUJYEU+OyLB
YS2M/a/BU7jxPyrVpqo9+6TEUXx0l07FTC4yP2ri4kRLlBrmLXBRMicU+T2WMktJKkEaMNpCdhOi
lF+snLgg0Mxs4NHDmbIPxzdG2MaW6TEHjQT1iXuGD5OhGI71xYHf5tDjadZ9v4DjXDzpVq/5Bun4
Vl8VMBxNwHfTm5y9v5ldQLCa8z4LjPP+3E92SbJi1GRVGGrhvee0h6zlRYBYpmdETR7JSyL9Iw4V
ez1+U5x89OtcegHhFQcj/aKyipRNLsPP50Ww9ESXTOuuW5d49tZUR0AFkSzGnTuX1TWfN8RAGn7K
JahFC3gwX/X9ronEliH5QUneAeEfqYAlwZoIwYq9cR3OOjBuCKTz3a5asOdq3lsRdXf8RJZtlH+P
t/Xj8C+Pqm2UtMIvzTJEVRuwvhsK0C+QugshAqrA+9FsTz6S/DxSRMcV7rb2ZQ3ovttObZ8X/DiP
2/fVZhhu1a5KTtQtgU564TGySlycKMh2XZqzyP1yXiGSc3QTEfmiDhHz8HqPpn2SgCz2v8NOQK9H
mjnat53iCav3kcnuwzPPlHE6jMB/7ISGtvVxYsJqmg13raB2irSdj56g3UMJoeKHlqvGwMHcl8UU
uBQ8qBpDVBIfw3GtIs9/B3ZGZ3+Q1S8jWpEq4q2ARsxthBL+kH6+Wp40SNvuMLgY0CIKm/QTTI1h
1ttfYOHD/feteSN6dmr9xMeLVDIc7aUKMv8uLJczZujRCFsLqX08VkFbIkIIWN6dmYpr+b+Tv5MW
EqfHUb3nCrYAF8SEDPsvg5rTRW+cF677qvpB1kYtIpE0prDq+fYNe6AIOu0wCygTYAjlCtCSUg1E
wD0hOtNFtdTlLkR5Q9bihTTSvxENZYekncwZSv9pMXjZIh0tYqIa8AhVQh/39mseCljQoYRiQ1TN
1+BwNVE0wU7XhAWSjawIiV5GyBFcaBfnL01KZDzngzg1XBWvj2NLE2XlIYmAcWimZemX5FBNxlcp
DopaPNQLWOouYCVtJVylWIDRjhrxp/T/Hy84MROIxM0GeEGPqyKE4bHl2R8mF9rdl/eKDsDos07H
SQF5l6Jp/ZOzrEBtMEvBJZ15Zrs7VsXhJdjhwdgkypYOuXHalgElGP2PumALsW6+ocIMlLEKpiVK
v5napGCKE/uLFiPFkCRv/Rg9y6hxEYwhiY9juWm6eS6W5QY6slAXB8TRi+lVdBcdEk40pQ9T1/ok
olVLDUBSvmstnPngdc7i55eEdbsiqk8OKwbXTDqOBSb7GohPr4QxRGrWSsJksL4Nm43PDavUSDfd
9SVfsj1uThD2jPIq93pJlvikvHa/ObEKiad2sb5wvVRq/UH08Yju7mcm92njgZcpPDDnbQfoPoAY
YBtnqINvxhZVW+6UnqwY1uFFdDpAIfgnwV1QR0okwjkbjmvI3DnSptlUNgl/JuGlitalIU4HTEFj
FYhDhxZqdZT1uM8Hfyt1gdLlpEh+7Qaz0COFPS92QvWnRmcWL6X3eHkgQbvLs616TEwIqYbq4/w9
IZwVgUXkKc4JsXVNVWskvL7B/3yMZspcTEBNzFn+JkMYgr+4hJuljoiHoucWa5E9EAI5JV8estyj
9MOQzO5S9hd4z9dxkvbRec34PR0FNeHRZiNQbmz5xJ1uTQfaCe2FcRMbhOPdmthkeCgnqsxDr/m9
z/13C7VGy7AEfYnOlwVRHq2+jdj2eSRp704hh8EI+syyN7PO1/QSO2sQk75Mf7sYlNhWzNBOndqL
L73IvFcyLHl72ko18mH1QNXsy4gv/xTVcCG89RYP1IJtuNvdHkby1IO45iXUCvhK2FQrdWSWrHLb
w+97zNAU1XAIB7teiNX05HT3EG5GWS+UQOKNyPabBYp5EcWgO3T7yaSf/sEnGcRlebcY2l5E5D8e
pOQeK7kunCR400OfISG6goyy0PXtFe6FzK1V0cdLRMpx7zI6ML9n69b6XdiAzg0PXSn+WYKk4MXR
3tb7KFN32+UumzjsUU4IrQC5VXQxwZosHyguFCm0j0wT80njx6hFWtGyiySe+D/8tuUtB0ChWi3V
KxbCRi+T2QTQer3UmrVQJVk3w6vOFatdkmeJ/TIollLysDJXrI/Eg9jfAN6NRrOq7eoCdFRsGTii
6b76VqjsOY3blRj3xvuYvGKK5mul7LFc7Ks5F6AOviUGGU04WNsX13+DkGJGF69jNnSOhNiNACq6
zl0BdoHCrVQumtRuJhKqNwzvrTjqlXJ9W0pDH/jqp3SYJirTxMeVxoFHC3YEyb4mPaVy4SnjYdhh
JBcPJpdn1caaURdJ77NlhXcciDMgkbs6rfjCRtxMPnYP9zLyxPeVS+PQW06SNXcvjvJGMoyfIT5p
mT5IKKCqBeXm459CZQImo7i0zFOYJsqGAbRg7ChU/S0So85/uuJEIl3rkMQ1IL08PRH0FVuaUQsH
UsQ6PsUvpmZf/iHYDtJA3YWrj33IF6hHQDqlRymoiLhc3byf7CmuEP9719eXi7pjkrklDnbnfsfP
+X6/B07XgkZOGMEUoYvTVAgKRE3fdvv58wV4IHTHwLBQd+ba6tuU2QegljI1y1HWoHj8iQjxX+zV
PMLC5g/mgdpWc/bljwRT2IRsHaF3KyLquPVRYoLnGenjupEdNy7pSCbqIJXbL6Kd2JaGzC2E/A9S
Dm8B0gpqJ9/AN9cqid+u7HuAgxx91y/3hG60aKy0uUO6ZvVJA51VzQKIg0N423vuv7RsYj1aF4fN
fdKSwJAhmkZch7rODCLJZl1pqyJO6Hf2hpNSPbxJ9CgKp6jlnVz7EUMUrN3Avy2K/V4oPPdGf0q0
D250eoyQY/oemu1koFkule4IiuV0WtgXnQyenQg9sSvVkka18mvAjN50ihOWpGHWphSMmK0nkfhO
wyW+i9BWSKDAwLCk2gomeaOLWczumaRRsKqPzOaqC2KRhJoyiITRYdoRw+1znn5RpLC/G2Xf2obc
d6+1K4EX4E0YlwX7yzLYxMOIHo4pXSKF/62B8A5+2y70OQVDbU9kA6kw79Tw6NxDnRelHr/VV/QB
ccyh9eDi1z+o0leecJqj+xaHa1cWEUCgRwlOiTWbGbMT5S3BONtHPh/44/eQ8pcqQ0XqucSCBAzL
LRH3pihb0fc0uh0QlL3AosoeQ20bWmkZItXbnmsQaMwgdVyg5Bd9zaO+1ZxUuqis5BWOQEbJyikN
ngernLtauYCCquZUZxKFji+vibizkQb6MaBpk9IPNWt5FpM9TlalObRySJSgQ9hj9G3PvXZ8K2KS
Vz1ze0h8WxeiEF9aZ1NfIDPrZniD61133be213t31VoQmXBbZhftstsepBRwOZE3JCWOXIeDPCer
X+LgTaUPqpNHPVYCejIJUdFp/UyGv7HgYO+/YSo5KArZGyCOF97W5eeL7XsiruXvauElmKCTpceD
0Cq6b/BGqdo0obHIDcvTJPkoBGp9F4V0G1Y5eiXVdml/MZ9E3fQT9bkKHdULcpHjub4XVJjnQiH/
LMhp2PaIaE9+88aT35/rvqQiM6jmpwRoBfQXVb7O4pw5r+5JeL52Jmrd5PU/ZqrltzP0rNTH2hkp
OGLkP+kTNIk7eqchXqoKEI60zrqqMlMTboK2/ionixQ1cpp1waUS931qdPpsbtCHoDE0W5GDkwLw
TQZrzXuCG77FvTwoZNv+PIR/19dwbtgI/01eFUTj9KidfBR1IIvnYypPtjzkujRBgqCyl0Eos4QO
+RjdQp7Kj58YOap0+aq5TLwwhG/5SBdZfkDTiB57aCkteueva0JIVVvSYE7qu3yT9sJCrj8qFG3i
JUfYX2gEt8CIjXQyfS3q3RBC0hdD2gBU/PzFWeSNnPnnz/WwX2CixNu0dOWscMcogjPn+ziPo/UN
o3QIf8Tpdy+E3Q5X9qGhhcu9HnyKEbY5gpce4j0CwFNABmh0Kp0ofamfIvLcf39ATKET45zygDVs
ZIMfABtI3939upvcelvMUc79YJ2qnnPJAk5RSP784oq8m5br41aDDtt429LiGPG+It0mRTA/lqDw
g8eMrEBdCSoQ+GKPlhW8ueArnniUZdsz7i/798He3VWKEjmpCxjT7ud5XOcguJ7mJKws/gfMLzYb
BSleyM8Jif7fxY224LS10pbn04hif6Jf4OoyRZ314ltO9eNoYJvC8zAplCm5SiDy9i784LFDoocz
py3Ap6fhpVP+0W8yrDsoOB96wiH2EKltS6csuZ4QJhdAdiHBqTcP38a62dsPcMktJGukHAGp48kf
1D8AjndDzkYSqzw8bndI/0TCHF/QHhXBNeujRWKZP8H4/VIPqeRiwqXVwGMYAM9VUIGLQbpFhqsm
uICdBzFAtS/bUWnMP6gqKoq0CBv1uWMiLS9mhJRnnd5toHfY5FtQ6ZUjtjm3HJpR+iNPk5StP9f+
Cht3WEI89ypACtS2HzzNK/WJbQJ3a7Dj2JIJ4uok6tZlUe3zmaeiJF0e8eR4OY10UtQNWeYYupxD
doDyTBuIJcnv+MJKgCr1dSS5lj6t+nlqaz2D0GuBp/D1wgFVfddJPsZh9intXeb0WGOn6eFOwSi8
ePRAaMysH7ZFKdVlJKlZreOrb/w9YpEe6ZBVuweUO3mSnYtxWjwCouKsf9rYnP2zTNsE7aR+dbjH
lXCHFK0PlcOMHlS2T43CIj+JMmUFtWn06FAsPM4WMgwf6w0xP8iJuAaTXhDJaIJrnaAAZESV1HQA
VIfCypYDNYbSZwlcuPB9l6/lrDUVbtuiO3wd6ZMonC6UGEwBKpMNCe2CG4u2D1eMPuwDyYJFxRAh
FVS2kWOHwIsjLqsKE7Ldj0JgoUZuvwVXf+BuVWftT/kP9VYNPLT/s4NuC7a3TWAhyt6PL4H5Y3KO
140Ta9ZTCMPfrMI5M86ouu9VPW397YvOctkM/b51TOkRdZnZdkK4KkqhoUUfm9TUAoRqEIgE35l2
C2PS32ZI2OgUmLMO0XFJocYN4eNb4HDpDudESCs73hDVNaD3duX/bTBPvmREe6HZyxWr/ATtm154
F0HORR6PUvEs60tnzFIeS041VhqUvRg7W2vpEedHgA5VRM+CuS2dEhIshFRdXDB9dTgawMociuZO
+/zEtoi6pA1FEnrmyt7ZSojj21Kqd55mcq5puYvTkYKE5oTLt9b7ouxDS3/fEi9IHbhHxCBM771o
2dpP8YASGtLyJ5XSKO5qIKPnLG+Txgmi8ZR55qE7ZYZpWCS+JvIpX+8R73bmltMhj2YB5SbTvDP+
/ywZYZXLNreOQ6dM/S1em1SZw6aaGmsGVN5OMhJpuRi7oNpMI6jLJ0g8yl9750RaoNaEvvFdIH5/
fPeFnOx4+8syD0ohlfhCyFygYCVwZJmTNbLdIkoQRF8z+BNRp2W3Hc428sdHR/dQ5vdv/HEV1qfq
rXoGrAKMzVCSQh5q1w0df2Dg0qkh69nqfhCPodvrQP+b0Rc1FGZ26sNaon4ifDJGoF4BCgGir6n5
btKVMlweczR01Om2sYANNvBkJIgU6YxN3WP4U1XXc8f8ZqcAePpkHxjKWK5+6fOM3RX40F4mFD/Q
YVb5F5LSqCsvqpDuzEVtm8kqX0fi1km7aYCj1IVQMw59vFDucqYTplpOeFFyPxzbnnUliwfdhLJC
dxND41vmqURTTpWNevsJWJO8DWQVKgXU5d5aVSvOGCtqPGWbWJ1IGE51uXI7TzYcTQVaBNbOfFsu
GTWrCu80q4er8GciYInekYE76bD/X9spsxRU7l8OO3nEuDisckC1a34c9MqCFZtY/gqqiG+Iy/EX
XRmPsfJF5v2+ADN3yaXYrOD9OnDumO16XYy5aT4J9Uo5k5+WALpYt6hEcPKVbqtk3qIAzpDuz4qM
Pkhx7FunmbQNPuzA/PKrsGsNb/2t9l38Prm3X3EaricU8KEuY+NTC1sjG+UK4g3fTmh/jk5x/ZVH
keLczv6J2FzAochXkTQMAvLMQtkZN9PUnGD8Te/OMpfHUcWQjeK+jdQZIKTsxpvt005zaITwwerm
MdUjzd28wGuevbQ6ARWgny2UDR1IdvW5/k9ZgAiiQJk/r47TbsEfsVxTD3Cw11ppmhMJY74WjLl4
zRVj1nVWH0eCNS9IWs/inLoTv3I4KX5o0ojhmuI7fz0GNNI8kGZHXPKv0lqZ3QOESRwp3Nm98RUq
Orrakw63BRYBrLyMMqREalfkUr/nNs0Ylsn7udGg2uDGL8MdxgAnLtuF3bDlqDh4K6ve2+SGC+R0
VfGEQMlgluvm6rChoDWhHG3BC3N8zuiXiqUVbB7AdzmNQGf3QwtZ3ho3sX04dc+p3aYRqgs23bI+
j+rmDrblV+/MiGH9mTrJ4aUDgS5gPso47YuUL9fOfIkUnLGRwdCbyKdcZ98cvIk7lmgCACaAEIbT
qKKKhW7tnk4fZSZOlMCTDangHX7hBKOgUPtesFsPUHEBsysm3O/cnWbqtOwfvGQse8UhXX6a9bhI
+WyM+1nGQ2XQiqVSjH5q2HkD6WIl0o4vHqWkLptOsDtuke3s+tvEwHLuTQBLxH9Wf1znq0sxQUdn
VMc1fv3Lk/IsZOw2+HzWnDWTREHdNTbtH8Lpjjkzom/9SdCNI35d7QLZ+us/L073NS81sb+tLhEP
n+7FjVXZAInQpi7oJbHfNVD5EQd3s2U24AFsqixCbh3Bed4O+Yr6YiPq1WJBSqoi5am72hE0xd0g
AhPo5CKu5fBOaRsCYg1dvfOH0Kp2RpDQEqcawlaYAAJllU1sOlTmfcBbFpSa4kqj4oOAy/85Dwjs
TErg3KodjUbihFcgWV/bL0Ef4nGrIkYt0AFap1QQz1ao04cemKZgzQDs8vpBdjSmGaLB2UOANjty
IbU4kJvgdlUBamEk3Xt2U+PQBwxGNEncGKcItjkWyBDUNovxdNMa4lmTxDQY2w8WeghIETWz2PLl
ZDINKp6q62rU3AvM0cjhFTEzkWaniCA9B84He01DXN/v9hkBHKglTwB6hRzReawYpxXrNrfPgZ6T
Yvd0GLORy0xfM0mcNdFvSFlpNaIO5nl4P50aUT799/cdluopedXFU0uJp4lsbhiqrikeqzdCqBbY
+iX8szhPTeBTb4PAPe9126noJtT9+F0VkoPWAKQPYO5vGV65svhGsNyJsnbg3crJrp6cHOWSJUnj
Ze+cUKALmCwmhKD/9Fdp+72HWJ1FCjcfy6tBLkV016axLiIhHcA5Hzn0Ecgbr7gHt5Tmh5j7NCDB
z/v6K49UVCWCRPIzdbL2dTilaV1zUr/e0t+vT+yM0oauYRVIPHinWWjaMtijgyUU2Jr1gGo310jo
5QZUPY9PXkEIiLuYn9SIZtGYLFa0OIhjrzmptJNlR9VykWeGTMZWKiXNX1+dTpCVRltGNckMtPKB
2Ob0nzvZ9qAn+D9syQN9xhpLijHzbcz6A9atN2ibtoDNrO1/lYM5nm5iU/8APcurYzLOy0I5P9gy
SSOhRBMADNzzgsyjxU1/5uXu8BLB5H7zz2dC+50Rd7CTOVfWZX9i5VDJ06a4SpUsBhpaadMwz1H4
9GlG2qcQPTbwy4q9awvrwEyYca6eRMzNdwKVvZv3I8kvTWd0Le5A3Cn4OgVhF8WlWTeRvTGMQooV
LkrHj5wNXfHf01VjA1hiS6ak7Yg04Y/rz+ITMSNKTGSOeLC+HqSDlhxJmp77/9/mA93IklcZYDrE
qjQj0aMg66MjBTEkDh/NuGXx7rnSdl+TJhyfE4LTslr5sWlBZ2B2ucdAoIugSeflex74JJhhwTDP
AFEbOD8DIWrGOjh8Q31rKhHBitsln1h9qUbvWevvD1EmAh4W9tNn5ABXAHNDAN3Q0m0G/3n1acNx
V+wusgTWshPVbJa/5/SqddnYPYVfDAZMu0xd8LHYGH1vZs8PAUI/TQqCUzc0ccQhhZirI+nnggUC
Dq2WvxE7XqRi3OFb2mkE80IO2LVglWUHBSV9MPV3ke6ZiWsTEOxk0ue5bMLKnAanv5PRrAVbO/Ox
/kD5U0Wp6vuBjxSODnG27P6mm3wPVSQR3CBX07pjHEN2q0IZYgt4ejS+PDNKAE3siiwZs7THF21p
6pQDaFctPgXnG3t5OvES64MtYiv9OSb5/Uj0bz3zZETLW6wOM9PJ29/xxeQ6drlgSpIuvSFlKOot
JYgHap5XtC4US5eSzU9yGot7I00YCMquT6RS5Tr5o0a0RRmSo8k9yUInHk/d3Zs9SJ28i5NBJhXr
H7sBSTcmYMkTzActvBkDxqJAfzkUAEfuwuMiFyQwxD5wU02XgvhQjExvYhhadkFwk+C5iaH6u5sB
XBbmjpgcy30/GVVy5oxqe9qzu08WPV57YfZhhUZboLjJOYzAA8q/waKugn49rQv/tpd8MWQixYYl
d2OJxHt7Jn1bfXoKShsRV5tslhDyzgC02h3jP7CLNzUNedJV7rfy2BTEtUNhwfowdgipkG1i5GYR
GkvTzWk5O6efcuGd7g8El/NzF4K8UFoAyBmYAxa6DuiK831XoI71gHhqTCiMDq4m26QMzwcA0De+
ZaTZZVAn0xHWX+brhskwuxxJUV/M3vo3OjKPQY4DxC2Il+SrB3gdKqh+Avn6j8WnR1ILnfK7TCwd
GOPtcTfV4VgMUXSZ7z0QEHUmWjGWMir4ETOVURSyKII+r4V4hkzEC5xRBi6fat2lx1v9iQqUvuPw
4Srl12Dn7X1UuIMBV/RGWikNokznzzKVqcTm7GetYTtl9N/smvRbS3VglVwBuwvgf/gjMHQl1sCm
7YE3g/bQEv5Cc0N6heLnXngCrQBxCacULd/uyCEtFYfe80YgKhOIjhiF/93KTiWUA6lFfb22nVzV
l6yY/C+SN2HjNHs+Uiwq2AhMNzqkvETEftVaqw4sMClpLbAwmxUsKQ4bI0YFmMHSURzbLJlR447X
Wbw5Jzr2wdgWyCHuKPvypbU3HC3JA+MyBG/2Db3Ixoj5gG8MM09XDwX7nu6mnKtV2EF03GBx6W0j
phTcbjFQREZ8TBLK5s6+Rhx/HmHEQgoQEVYCl5e6KxDqzXVivN3OHbMSMXSjbOoB8rTTpxQSwvCQ
Un/1bComC/7j9QiTRV2kANuSxSW+sZeoZOVJodMMi0364sH8LO6DOhY4WLkJScZBesWY5TXwxuYf
3BXT25QRcs0LA6X5qTSpRSGWiRxXmUS5dOyauzOYL1KjLH9ggqIGPGbhNPCQl5R5RcjyTT27cxy3
H/rjXjAmY+gionpnqTFm2I+VHyB+sZe6Yi+ZSUiY/L1VyfwNIEzPvzy6T2lWJA8T80UlG513Fjt9
0+af5VIVd7I1WKedbBKWdev0hn56AC9Goyf+TTw686S0W0KzeM3OGYqtVdHP/74nlFpIjVRBn/it
6XqoMFA2KLTgzcP1tx/DttqmU24pXS9WXFeWRCWue7mSb+EzfXc1GaojrAibge5agmg6phxiQVJ8
T6tnQ3w5MMZ5EYXiFZjMXcZ2+Rk35MXZhVy4NjgSPL0qSmoJcCCA+McCLEia2Bo//mxW8Dyacijo
4nz0kSalDs2z4GvrLLJQ8IHcH1qf+ST9oSyYRImvicXnW5N1D7ayeLSp2CSimQ6Mrcbq7rPFmlOD
E5p2vL27o+ChLegBAwc4ORUJ0z3Db9YFX+Pci2wmmKONLYjYD10ainO4wLeKaL1P1cv3OfQs7WiQ
9uLkDwo3ufI+KhVrD/tzCJyRb5JTC7YSMRETp2dQrVeSbe5Wo3Kvo5NaM1/tXtbZyZMyC+ghLsA3
EfBHGcbTKqHLXJaaDmBO/am1JH6bupBi1AU38ux0KVWz6RZ0lC7inUFq3g6uPFIlf2F4B6QRptl4
kEsK3ioVJtTgfAAtupW50YPPwGPlRIOwQrVv6uY6ibLEEDTLBl5zr/8F4YGJhWMDM7oIIr6dzrUL
40+IlUc6zmT3ETIJ0poRSNuSnbRCiOLVritw7FGSGFwdw7g4t1SXFleULHM0m+N/kyKCRUSp0sUD
kDpxAAy2Fat4Pc7KQpcFVvrMbUxBoxaSSIC44CcdCsykYIG6cDU4bhpSKQ1Imclt5p8k34x2Iu+3
qY3mlhj6FlSPhNGPTKSAsWeWNYVExQPHMQ6sXznwSFAqPiRkn5LGlcrmlMzJFsYZ/16dF6/W7nfi
VrDQuGmnuzTWfSFLSt1Na+34rQlJ0jBALcptxMpq4JzHneNK2c1Z2SAOyPgDh73DyfAIkAL/yIKl
1n0QtEOqAICQv9fP+p92S+oYSm7Y5JZdBzAnhWYdob/IZWY3XiXR5fLZtmU9jWU04D9MPOLqNv7a
ObYqWPKqgMwhYdIUngTZrHXTI9E5Ci4QIU5K7RJFouuKr01IuvGH4CyHDsIefFGBSdCfF1v878mL
YxAWbEJwYxzN9nhlCnhH9SyayGs/IWS2W6ES99eWfDbfAUIFKaPYv38ON732u5+PBhfi9sf2E5nQ
qlLoYnRgp+hkDbaE9Scxxkc8kQeEUjmfcClOmRxpm5R+YnDz/uNJIxyZzxn5wqtxTRt6QuYmlay5
bNKAAS4UExH5pveNhWWHTKroxI9vpsyXZ9jjVqt0UT1Mh9s1D4GB2WWXvjkdDj4TMiSw/8ucS/KP
IiXJ5E+YB2NHglImzIFupCYGNbi+3VpqaXcCAKrRr8GMrrzGUP6esO3CJFhs5wJdLgz+qh/ef361
ibUJbefyZ0dA8QW+B32SQ2y4myK9W0iUC/pROAnXrbK7q4piG1dmfhUeM/N0LVMMGqomL2PEaZFq
1i0rCven2KfUo7CbxNSGftgc95EehaBMvAIP83QoC8g88ZnWuY2nE+hJGt8lqnIFnROiALJtu9gf
a8VsPSG5ms/W9YpGRiZyqMxuibBPJvh9ks411/zKelnN3lLoT8dN7WFz+ycb8gNqHon2TSnu1luC
jUHqTDfc46dXwmS0RMa83wbpLg6OTNabXhGlxKeT5ZD0EhVfnxPHEg7+nT0GJ6BrrQcSNb1G/yR/
BVqHun1hc3kkxRrzlFZrK+GOFcdjKvwjQe1DXnxOqJsXjqJtcQSIIinZqY0uZNvcHW76hFRvLLiX
U+2VDdMxTQx9pgaxrpbVp6da2H8M4A/HgK6rwg/l6jgGkqNuaI/yo3zkqOV5Yj5VlQZTK8OgvXQy
V9Mjx0eewdrtXsqEixKzXn1D2s5g7rbBQoIg3LmFHV8edG/FCntPmwh6gQVnYLPC45d4Eexr19Gp
i0IfwnA7B1oJToH+g9uW2UTbQw9S26Na0nEcNgOq0QRBpPTk1wdcs6g+kL3KnTvBiK3XdHuj9cLK
IfXt94RZZnfBfBPa3QASwgFdDoJwAPJVl4hqMNCGtKKqUuslmZDDxfisCN/FVY43ERQHjbQMm6Ld
jy8U8yaRDgUQ4XAyNjcUC9bMtccy90harNKj07i1ueOOoXdk+5UFgjq6j5osou96aTwCctYyf3od
LH0TDQeBKazY7ExnC0F2CVEFWJxahbtROrmxXdc1Cp30ksgqa4DbtnQ7M4pBrSRyfm2Rt/+Hbd+r
y6d50USuiaVAfmbTu9UgxpwyU/R8iml6sCtfPvUXilKkNvLLbdYzEw3SEm2eO4FgAyzwwxsfbDRr
D1WggxuSGTDZEPydDr5PpyBVrTVGXxfUq6+Z/thXkQAMvW4QZIDQsK7DuGnD6Pd3HQvcutDFoz25
+p4xbUuChqkBjCoaREss4bW1465VqO7USEywXthaLkudKlPtyItv9kgxVvidXxVNgO+BBLeArP8S
yt96Uf69krQNPG4Wsac3yHPUKE8ztG1+XbUkA+6NesqzylTw+ub04nyYi4vxS58xdPXlVLGN4QnK
FruQUC/HywoPMsCphpysky+0ENTCCZ9Bf/MhY6TfNqvxmlW0S5Aeo4vJpG9EeXedNGeEJ7ktg7Nr
xIbRrVUtstfuxDPJNVlBiRUZJvp2uCIx87s3Snbog2xAqgx4CkMTn5X0uvOcQrDNXL+kq9Tes46V
cn8PNiAu32gfcLHg+F1XDkvVCi+VlilVE8Fe2gEUtY3wDdoWz2Q5I9WyAJvf42heZuG0bhjd8/S3
yDyMKxX8YpLtifJeTd4VwcL/3FySDiKfypMP+BAuF8OccKHsv8GrLrp495Gfuq9GqZ1Z+4kU9Vk8
yyT7NikaA2MvA1Pa9ZvtFG2jlEAc2j6B/qppliC2mdu3l1DP1Sdkxxmitm7R9PATMT1IIdBk5V8V
qAzJbxVxgysIJ21OzCeAfURWAsis+PH79TOAX3dUBtBW0PCE2xN7q6MxZXbuj+Z3XxNvRDjyhbQZ
3UagXvFooRxcdHECOgqcYL6V+THFOGGGTKIw9okcPomOlCl7GiVohvgg/pyGQLRAg/lS6yGndkvc
KQ1W/Ih9dxaFOXlrqyTPd1bp1tH/zRfmouO7Qd/pyE9qgYWYmIM0rKHuQb4eyKueBjJpb21zCRD+
vjRIDWtQqnye231kCD6fzXnqU93v9LhpqzMypI0lNc5G86uhkYJJ8z1BEO+2K9VKJR6zaBgiugEL
UTVz8r4JNNL4DIKKlyGwbEir4nkMfc0GJ7nSgE3RRQX8B/WU9mWs21bHnU0scPBqXMlN++I5kCwX
POyVs7bpuBcL35SwjYKcdiYAD+/9smwObaeID21+yJ6XdwSATbLibmIj4hRBJjq06w4fvefZhlMj
yywl+oJsxtqeaNh/MOnBAq0iWqeub5A+9IxURox4EYQ/aKO6pmNv8Fd/boHMYIbLc4DN+R9u9j6V
gFXLOqAKYCS5yGMJCo4oLvyZDOZRy5Iu3Xh6b9nONXzgXzMp7eMtExMZ/a1AiP06CyMLzvroYCH7
GVYUgy5F4Czq944CQC3YHwNvaUPP0bpTInDtOfExDo8DQMNNMov5Fz+iM6+fVI+JkghzG1xVFAW2
i4wvLcOO9gAUUcunrxagkdVYVaTMFjkWTZ3PM8w8sPQM/BuDGSzppvgGcVEjbH9C3HPJNmogBwb3
lvXNU73IwsO+GP4hLhCDMSHBEvXfQou9BCCn84psgMa31hCrholIc5hvDpECAMa+PcWyuXXf2MIJ
bxaFeW6MlZx/QR6rks6nt1pJQiYjDWkkzLX7tnN+FuiVVyic33Fl3IeuFljCuhkWPz/RoOpAIQww
qkrFvtZkBKQztYyDyQMsOSM49FS4YyhuWr5MK8yGHt7CzSx5ud7xCzXu5PLWWRu5C09UlvhYZ8vv
oJaNURiTfU8ywUOGEtkmcRM+gS1nB2IIyiTlC5IN/3rjkTsII6HnUUvNQMSbJkrTU62w379Zi6K6
RX9VW523BLf6J/6MptVgzo5/+R6zswPKH5LmaIulHMg2jrOYrBNfXKggJd0TWbZG0IV3VgWg8eCu
bFLzbiPFstSG/JhVjlbim579JUsRbWej6GksVsH15DtECsH8d7yCGOEtzW+2WnBeFm2B1eh+bcln
viTQnmgDdM8Pp2THyyoBKjsM0WVIpfPoXwTJEaGWPCvCCGQcX/T+CxTQyvSxRuG3bYRnDW0+6L5z
jKMy3DOoYQUkHgnRs3a0nr7o0NgQgVGZMjI9C8LmL9ySYHTvgIpwasyFegmYHIwd0C6y4U6k0LWD
ij64KQEBbNNBf9Mk4Jpp1m0UVh/W0AVSrPAMgNvPWt5LtWUF71gADjE36m0Dmv2lE0aUIOygcewy
AxGWvQj6UeHHf7wDFcSD6ZpS5oujRd+jq6zvjFSMsS81DJx36Ze3/kVuyvNG6//PERyyAch6FODT
bArJ6a1wB0LNqVFBwY+uXAF4CLmy6Tq7C1c1dgyYA9pgiufNtPAIN67AYmkZBKzCppP+z1QRxQ/1
tOO8KXBnMjLKOODIZkDuul8fGcSyWmDz/uq531bYnF4WWa9Ry64NDVa51vrbs3psdz0YTSa7BTjh
DMbZIUONbj6lw0G1lDlE6sEStI+XeLGF458ng1IZZBzb0gqXpQuDFL+N9aphX8W8TI0sDB4R9csQ
4qSjda5BQY6t7puIaKC5pjLMSi1ySK6xaLYuVbT+j8DMHWEbb2MTcAYw21g1YeorlTdG15f9D0eu
ii0Ei4iEdfJtHpE6HlPO1MRvkBpi4rMSpA4Sy7XjvgIJADax88IH9FID2u95CCT/aPgXYnxXnwUG
4KQI7Y6LC9Q/qSQf5oc2PToGjpi7kVowYkiroX4n9dnswE8uQQdKSB1B3KcAchoo+Tx9leLz0GOJ
Qauc3crYhbC4KIypeY3OBhff5paXTD5ZDB4IkjmUEU5RHq9GQp2uFzU+RTfqnbvP9SmMFvQkUw8d
EokmnEHLri/QA+v8Mvhvq1SdFLRV1pzHhCX5G/BJpYQx9yFengHZYHTwmkE5V+as/Jwyw/juOMv9
AxIFqSRE75IZJYDRu9LS7eVupx73H4Uvdu3esUSrPJs/FcAJoAbWalgJou4mBFMtkAAmVS2aZgnx
WhwCRL5jfEkh1xY1nsF2UjSHWGxSdhV4TZJ/qE7LPhhuu89lE9PWREuQi/17IHMeOa7DEoSL/GDL
OasYCz+DoSAkLT4JbTylLC6h0iyCcfavy8KACU7PygxUO4+l2x85flPAafCghCRu/DsOIsTgzlb9
X/M/WOBZXk8Gf/r6GaYJCNaAibC5dOrzUGqA0+Fd8Yb/nG6V7AIxD63SYsyAIG/5uimwDDRsD5gh
lo/M3DSIkvFJlrp5fbOMxh1r3mpG/A6woptcLp/gdT7wJG8Nc0sdcFGP5D195mIsFSI39dtmQw/V
grnDmhtntDLpmlcFeahzU6laK0sOAAWTi1YjzSOiTUUdpqPsD4zu7Z4dEPho79ICSCrcTQZ9rbeO
BCl63Y2izqNNMsRzV6xaRPxMY/gSMEPNVG5a4k5TEts2Ybdxvrgfo73vajFSF9jmY8bp2RF5y7kr
8Q492mMx1InmgJIRBx5pWG9vqhnd3XesYwb2pCh02EqRxzIGR8xWGv6RW82rzkSlaFyGD26dcGdv
Bhew6gLQa/z52L4MbOtrjfAKGGCAa5gzMIUw7oTgTKoK1AeYMxM3PoYMJgD5VW4wPFJIvcW3SGFh
D4ojgCSEFlLtOdOqh603q0+kfOj92GLE9SDq3kywXl34IV/dZozdUjSIxZWPHaAr9kMdhYNq4EBG
eLS+ADZ8SNnnv0yAvC4Wd1Sw10g/7GdsrnnjTfr+PaExHgk0fP9WV0ERVoZq3zbywIjleFZCFK7k
mPif44cnM2x5hj+AH41UiHruxyln0xxFSucpBHp8k5iTJPUyf23YnZJZl2KktM8Q/6jlxRRJj//e
3APtB7qEIMnWFvSwwIMqtuincqBMEBYpIhUcF8n62ooE6tdibD+ZN80nMostbWvpAhqzfIskx+Aa
13hFTSojPznoe2DmKxRUnixJ2npp1phkBdEFsb2hJUI02rd+2O9EqWU2dPG2rKr8hK5muMo5EyyU
qRP9rN86S1f6fmPi4+sOCnsR83fuQvfvbiI3KQc97xQ6FN+j9KVvAohmJoRgZEW7fq/6M1FKJCVP
OixRWECIp1pJL20D8Fc3Oz1R1Lel37pJW672ygCNpalWo9JeYeoYv4n+virx96U8gUoSzmM/xyRl
dUYQYFBYXItOtl1QEXjzgCnWYa3rpKQV65tgv9GPsVEPchdD30ohyWSJnQkpzGZlP7QaUWbMXBQg
o1SCDNhKknmNzxTPBD6Cc41/RSHhppXu6gaLUAefUnLXKPmpYlB6Zd2CStc/lzijauBqoSYz0n0W
seqmIV3/J4Qq6+xE70z3QOdm2C5brqqIewa1zFBziijwIvQ+dyKT7OTbb5H0/tGoabTUNMz9l7yv
o+iHOdh1b+0gr+elntZoJiAsqW8Sb8tNO7NDNllKJZq01bI/FERers+ctIlvUupO1+OSV4IamIgn
Uvf1/XgKhQYV8HNX5RPWTTjyq+GXAaXJ6sCFPeYu+rw8+qXextWJy0OQxWOuKaDUUIo62URFpQEj
b+koHAdGcY/oXeBBJoM7Mui44bHg3XKFcyyeL9tcG/5yN+NVsPJtxM7BR+Bn9nHqXU++xTdEdxdQ
Ttdr54U/1iOdoAymUe589i3yAISEMLCUm+wA4QRDsUc6v6sJG3/XbQ9bSKucNEalilW0HAepg1HW
v19POss2mNZnP4rLMeOnDdnrf3ASTRkcdV7DeEtg5A7wtuDWPfdCxv45Lrnq3aHF/F6YFq5XR0cK
6yqWEsBXSMtH6WzsQaTJn18FfP3dCiIQ/6jXi8qW65mmXgLPo8Yz6/aJDpRBvecS5i85YDLMjn1N
iUzqhjvG+VoX2bJPjP+i6BbGpfocLn5b5Ikixsmvlx0tAPZc8JGJcoxBM6ZoRXZB0Oje/QGmcyvG
VKrCQk+ZbhjGgIENhZzLXH6YLmv9kBtlqfCNyRGomY/TQxjpN0BSjaLtyfky/lesgiIpEVAqjpVc
87z8TlMkgemVah0nYGPEzLBVMdi5jEwjegP8YkTXzokoEuVodBnQrvDQIOdDF+WE2zDd1wqc2Zxl
BgndRbv1IndtjQIr4wShhF0BZdWBYpAWwDFMTVIwJMiqTg8ZDl3Ztbk2Eotv1Qk1BUwNXLeGKL6t
CB8/1S5V5Hn8s+yZSHPORGOJ8yLjjrzs3O/pYU80JW60VfmWU4KWyIJlgFTr1tuuUPd47jXgFK5B
w5AtBhAXsevzd3+SOwe1einE22tVMXgl72GVquMqhJkqAVy85C/8BxmA9M9+KatViJRLILpKeT6s
cWPsZf2U0eBnyzsBn7rNCkfwVzAhQdaDrZ+/fFAaAr6C3if6iHkZTqNk9J/KzZ6548Gg/CoupYqT
CnmVpmfWgclo6UkfQIWjowBSMAcJDGTowi1Ix6XcomqPblHGoaXJE7+4HmemEG8qi/DeUZ/KBt3B
BFVA8zWlzJXIeWojEk/QCtAnSeJefMSfo/D9vKsUXHdLHDAcTg23DeYBkndLd0Zzpo/ZNvnMD44u
cT3x/XV8L5Jzap4vPyz4PmeJIcQ5UrED7xMfg2Hitg3oi/R37KkVaSeTJuVxfaprsAoRdp9BhgB4
cxqJw1yIi57qqRZJ8tLNO9+6udzbPWghmgtlQyKo9nGvbcRBoi8Vuwf5VOrxPC1TpOyO7PwANSIG
2iXTgxB1ieVCpdPUOH/C7YfYr2lvJnEok8R/NPZ8+M8xnWbDyfO/17uGmh8PwMyPcXthnUjNoniI
xkRGhV5ycl8nkCr34vOiTMQcn8djb+joPmiG0elpShHM2FGcA57hb4fBu3Vt4dzHWrMffLoOB93X
bLZQQuCSmqDPDHsJxS6bf3yxIpxq5HHIy/5OlXHyvzCSk1dTFd2d1FddhO5BfavG1H13aoj7JTKq
3qJGi7C3ZXS4Mg7IeK3ErcavGPDhh+VIg9GPy3APly5jc/7bfhBkh7R2EerVl/USE45Bqz3yC3ZT
DP18WiPXgV9CzeMeALDxQJZfB33rzlam4O+Uv++QhlBdBxKXSKpeuu45JyVpyu8ZKO1GkT9qkdZ2
diGnsn2FAxBLCztUWsa1aEF4anvy0XYndYrpOrSNzE7+2YL57lzuRzU/uOW7+2zLOGqFTbtmFPfB
8d9Irb2gPenzUeTF1yTYayO4/tjm3sPM8p23ge4rU9pIXRSZy6LQ7LtCIw35wwK1G2G6TriJz/LL
6GN320nvPxfvPv/McQZ8627Hcj1kuXJSCebfCErzrO4fjgusNPXReojAVTOQgOIG1LWwKf4JkD4Z
cnI0MqvzXJeuxyWhJXlHcOyoBelO+Hg6OnJ8RFS77pPIMVE3uxWXwnwdWv17facAqN0BHUkpTcQU
vOM1+097OT5CbYmYrGEoTrHfY18JC+OA36NSkGw1SGidwktRkDuzXfqHfyfWqlvEQuWEqJehTNhr
7tPI7CwGsOJj9JNROpkHonSvbYQm4ajuDGjHDVXVQGqrNFEcqT+uTPjaCYOKSlJGSvtq8EzL+ElL
WSidCrCtcdADdUnWpPXml9h1LCJPe9ZMFOgOcSQhXsjBhzQu2JwKx+i7JblgfIskLey5XajMjT3K
NI7QRRr2VkfcR8zd+IFhzPhTmRZzJh7vir8J/Psm3bRiVUT6eWTF9d0qY0AB28ALGjPTO7MOFxqL
LHkKVGyTcsvl/It7SaoxtmSbBcgxH2gi4u7iRI4gQ3Hm9C2lED6+jRQMOoXw075QsmOX/5ZAWszz
vhnDYnR2NPcJMIwWr2K12HbZmirFjSuqVJvX3clMgszOJbyw9Pm+tpcwfSmMWOvC0Rnsv5luCI6f
93LtjmCKB0yi665XZpXz4Zs+ryHk7FkgkxBovm4KCmewd7MiPFSiQrWlEgNUUU8LV/q5DSw5y22v
XM5HkqXfNdEpbXqs+W0CFiYY5qmfABTTFE/QJOnGcZFB2USe6wesJryxDQJJa1r/G+9emw6Twzey
Dy7SbAJxuYs+iOr9ELpOD/xtFgwJ5zaJ7TmcKWthMlZxkmQDf1RfK/JItx2Szc29PQcNgrMUB3x/
b1YqBe3EF6mCMvlsJNKnAWbOVe4Ava6LjUPiXkRmr7aILV6T6nYYBZOAxVNwMdDIFMoXjXmluTol
9ILX4SqfCAaPERp/xlU78PeTw/rW258qRrTUIsJMYjmMJZbQmOTd5P8uaThTzNtd+CRu43Ofl3sw
fsZcrzinP6gFHwCBzJOyb/Vl6duDpaVLUmHggkV+sP3c2R9cEQF5Y00bY09B//h8rO4Sp9ajYyoU
sPIyrgLveveCIOoif1LvNCd2cL/QOpKGhKi8EEzHNbvplc2COY1bSuuDg/gndpU7tpjy7EKm+jHI
c6rrznkMb8OIxUkizVUEKunWh3hq/8BC++TjDpI35FN9VcwyjpGB3OKyWXT6COl2Hb3hJa+KM/Ry
5xFNUqKQcQX7+5n25vTxTEOB2t72yG2tsQXw+Kbky3WKnhRNDUeao/Cv7xk5N6xuBJsFA6gpl6rK
qpyLz20G3pTjd+6M2aUBculEjE2loav6wZC/i22YvruX2SbpzZvL3quVUDu7BSebE19bi7rYJzbU
p70rQCcBJcW8lybxEmEfrFwV8vjvs/A8ztZ/1wzsE7yeWxSuXkOvGSjycbB69ofRP2eaIbdf49ms
vIoun9KKIkHpd9Ojmrl7zOmrDiDtfepu9Gox87d6JWArORJ2aOXfJEM+t01GmbjYOYw+Rqxp6srd
5M6cmGDL9qrj9c4jZi55x0m0nJnYIfLf4i2TeousRBPabC4ZbQ7AC+LxoZOFNd1p2snBRMawjx3R
haAXsTWpnFkwnldqws0Uw7Srg5T9AKCVnkSAWgpe9VhfcCF1qLQE0G71RddEdYnVTDpYay/U8B32
kIpZ3o4OQWiL47LL3d423rS4JOwzrwZT9PuIn2cNuUmVIS2GXjmU2CpSOHWxNblotMUgx5U9f4a5
OV1Yq7AowdDAOAo4K1c8Ve5XAMgVCFWuxNWe6qJiLAxw5FK4Ambfmr2hTG+I+/qmpbRQklNrToHX
MlNQKTxfm+nuPwtSMogaup/HjooZqTNiyDAbKfFgJHcANngmTDtm0CJQAAlJYWcxPCayBLNKdDFG
Cto0PXxNbKBpKHyhI0jDlIgSl17PckoG8MBDCmRgJCC9SddLlpbfOrJnTwYZvhsG5n/90yqi8O5H
DnBDutwHby9Ufq1DktYM9h90yOlPQjY26KbukCtfArU4PPh9e1K1kNXwjFfyP5rH3E+wKD14AaUM
eJLVSSkRiP7OYFAliojGjfLiuayb2pd6PPke1aIBllzcS6hZuLV9JPexHZDKDuE/9IvNyfb3FCQj
6oZfmBjuTboe66nRM9Sbc6sImG+GzIJb9LHAHI+9ja90rperbroASzvg/W+MsPIN9/Vwb8mnzunx
/r2xtrzmE0GRh2qIMyQWJosmYvhdyTIPMqsLbhMbJwVZnlUeF2HOQikHnhn5DrpU3J4qrB3q+8/Q
zmDnKd0OMvEuqDnNmEDbVckUQDmJEdk4woEAeh1XfyLe7WALebh5YYcDfic4NRf+rDnpKvbShqNW
l5+MRur0aNaoxEFGB0IgwNyKsAdWy7bsjZjz8oM9lr/eHPyrCiqywHTm1sgb/98waS8iibXK816K
i5dWZsCrK971cO36/8KbpZ3mD6E6q7KaQ/bcUUJRBQuSKPztNHkuKNIADuiXOvBhy6l786aZRc0j
SbqejlKzMCTTJmSYC/nKpqjTvCYTdd+b63qWo9nffVxg0rSTNKWi0Wfq2hny61VZrrm6rrWL/g/+
SDoCuLcFbbZe//G3Or6B2qGrQgcVYdZ2FRtY+YLX2CO4/mMM6zjQeIFfgBlpiTpNV56/tax80BnN
X13IDQwn99a50JCbAYiD0aMtswuKxEJPsLAzp4G7ARXJY2i8bzBXnfPfm9LARqC9NcZr/qgYW4a4
+5whMnCDZa5+2O3KsSJFoS4VpfbwMDJshOrN9/escEiOfx4R1Ex1JncRd4slpP84b7SuBpEJs6Wi
E3kpDfPVcppMyX1Vri3oAc6UkMO/7QeOKf8PTN4ADznWFA8vQkLw6NKvdOTnMMKJuvT1zuP1OXcz
/KZmER5vS8esJmf5UKreau6uOMAOiTNoq3Df/WC/w85uiWNzcTECrfTOSz6xYH8Y6Ddxi07eW4hE
SChDL1XW3UktVMcp718nsz+drwGlQomQr1ckCyWD4s1jpiQIUW4W1Gx80xBNJ3beKVpf8EOQIrnz
Ysx9pno6a0rPodDNYtmy9PZb06QVIXyzcCbRUvfgcIgrhc+R4sy/eC3vjxevWPcfrbOA6s5P8w2W
Dw7Vl49Ohoq39JbNVH4kYubW3t1zQgsuLUgmKYr5mJTvtvQNpe87F79I6xgmrquCmUJ6hqeHBRQb
CYI/FwWwWevZ43TBftsbDRL+3VHQgqYrcpQups3TKXhJigU1yR+VQDWt3+4U/IgQTFSMfNE4mRXG
OeeoRepP3KkyZp7ZAVJUHc866TVs5hxrCMgwx7O86I7YoXUdfgtms+MQwBqI9IMld3D7RHV40mj2
2fMyWIKKSw6D0soNUR19yQRh+URM1OK1yr0chMtvx/XsKvmtOxAkRAA39rggmnwS9lvUuM8iK3BG
tvpFoxlw1PsfUJboQ8xo0cC0fyNtk0a3Je1QF/03HhEHIAMGMHfKcMLSVkUowv2bfD4iLRtlmGWU
s2wp7wJ2PwaMPh6irnrGvaaurdhfG8YPHmUnrRva9cTLr3eYkKbWSKuN575U5ElasuDw9DXJ9iI/
OZqxBC6bQIZc3XPlDYtjTzrWAO/6lV66Tw5Yo0oI4FQL6eWMt0aDQx9QqEEiopzLw8YPXWFh502c
gmxMdFrRFYcNypt8YjhNYN1WYcU1e/iwB8jpFQNDChof8vIRPsI4hYy0ZAdeI+TnOM3YdnIKRtdo
weSjXLvpnEaR7I/Zoiswipfnxa97AJ3n47H7PDbLL5dUoAJRL6m1pG8Et2J6Wd+8yVzdhmbA9sQH
HH9F/KfeRD3BJnno7IK/yybb/txYgvoiSxoms3YzGYvweYxcgorwLKB7cmnk+Cj6Sy9yJrCBJZlw
5Ids4W6fm2zvSCmXnayD5p4cvTJ/5vHyLdROOXRbPmCzMDYFzELNllEvTBjhMWkHiGsgJzoE69xc
G0URcgad1bLtn+m+Rv1LnWJnomhu2qHa4WKZILyw8K//wuo00Dv4pvO8PyWQ3D8XqahbN9XlCzyH
irlxBplcKTE3nNNNRMzjnacy+l+IkF1qdn4DYnHU4ip+HMj8/vIFuWviA9am4s1mEMkQVIH4O8oT
JMojPwunzspeHrkjJdCXDtRps4i8Ty/L/Io2/fgPuem74G/2bV+9oil2ZU93I+qHNpkCjbqSOjVG
R7Y7cfrE/W7DKdS0seNeQfz6AeMfDuuPi0SM35VyT+GbvRFq/tfh7zYAWoByZ+W+qiPaUjDCCydJ
X7oeNBLWy9iLy0Lt058mMqHnJ84DKKVJIT1NTLtqG/wvMCLdnF9WSfD3PrZ2xz+n1Uj2rS6hgCDE
Zp22/FFoB2TMwg6ICIysXFaa9KpY/urMNEytR+mazLdV5c28SqUZJVPaQpVWjsj677bRO7oVyjKz
TX/y4vM3Jps3S/IXSfKRwmLk728tzPaVNp10flhYnXWyYn5MIoHJ88J1lrMCvqyD+48sLui3sPG/
ySwtXWr/cphn7eJ87MbYZWpxtXXY1XW2rqwSEbQntqoq4ee8HMITv/NZwJ73Qc9zaJWjcgdRQsd7
M4ibnR/tPUnmMf/3HElZ1Rt9IP5MNDT5bI1dfcYyGfuSG7K7JR71aio3YFXoSI32/QEkLy4fycNK
7gNZ8G0owlV1xmImD5mAIdaZ7Mg8WnqEhAIl5R7adNOVPzaqahYeEo5z2PbNazTf6dKmHjYErnBW
WcfwXROnMhlEyQJ3/NdHQv2OTOpjYSNRrrqYZdsZ11Z4sXfqotp1YzL4+nopjJynyfMPYPDniw3J
ZT+g1j4Tv5bnx5Epan3I+lBZDaCtQorOY9B3e+3UfK/dep6DAqwSAPUGf5PmiJL81dKsN/+gW3RJ
+cgQAVxqxGz1AUyFotEigsPgh+LrNGUrgnKLafX5E9F6Jv1wp6F2EkR66RpUwv5rQo5GeIzsSJ9X
lXvvINZ7WU5s+W30FuaJDRAsXlwep2BL6X/KeNzX8OxOBoy/7aGRmsOLsvre2O1iFOq+l+HteE3T
Tk/wnXpRu81vZcciecOr243tO+g703gbt5305m4ZFHnm1SAnKU+w8nV1ZPx6UfnJn8fbtDNiba0Q
rDFUiyiokqBzdaWogVM5Vx9AfzUCoQHimTANOuO7Q4e/iPpHFqLBFm5z+K0eF4U5z9re2XFuFMa5
LSwuFCBttl9VIU3YzjIlk7NCzPdSZ6prMhIrj5kDfG2Pf0nPesyNNCsa/iMkUTd5GRjVS/F2k4YV
uXhGJuqqyynH06KR6t5GrOOlOx5yXdqBeOEb47E78jN9FKKB6OWD1vgPnTo+N0xinS/yXLfVBtff
25yWULAqnicN2LBIncfQ256lg/cXunWB/arnDgpzKMEiC/LsXF4CuLzlKSNkzb+kEUDY8/IwV4vs
vlS93T5CFGbvJhl1Fo4Oteb7/rvJvSDVGKjWm5P3kMnlHDXsMieK6mG5n8LmGw9pXQno+4mg5Yy1
JmfnpjasMviCr2TYLg56xVIj9ciUkk+oVl7Vi8dnYNEogFk0M4o4s92BAwhxlWIuduypoGjWL0pR
yvqbxYu0jrJLm3jSbJUm6x0KmwYTgWbm1xSMGRHNdMyycKJgeNQEcfAWkpQxFNDIIDlmab2HyN9i
EhEw+4mVpikQs0uxHOji8TX3kBP2FZfxxx/rBi6jcacYxl840/NVhH66k81UKuWcl9h/bQ+xAzsC
og4UZKx6Kr8n3W6Le8sJRU+8lPeEwYYn6AZFxKV7mHWi/aHVMwRVA4kg+HtjsIE79PHbdD/mwGR9
X37cSZZjknpSTlKPDUwzNMVQpiSD+bUSfZ8A9a9QmH+6ePDiKLNpo4krhANy38xIBwhhkcvlIvcw
CmUu/E9Evb61ic2Fq6++BVoGebtzPZQ01cD1TkanToETzoyEzrcxKoOm6MiWn2LhQaQzOxzcvgqx
yH3NHExFGYixia1IhTDsVwvMQeKzgBBErv++Kr8js+icocyVpXrzydWCgb5+BKF8A+yVaGsoQ9oG
KeX3Zm4vTf2Jsqw6z4COIHk5c0qA+saWQPn0yYK+Y8WZhGqLVB0ZgjKpvhgvbhzjfpooFeHpnF73
/us6tDsu9T024tDdolBhRDdNBhp9sSnejlqKg0Zzcb5uZSZ0JHA0V6CpdbZHLr87COOF0YRmlNFE
91D9/Bqz5qwfSgjiHf8e+BlQIKwfKkUmESrz4wBi87rVmUAizB2q9iVvHZoBd1aGGGqVDTDvomys
f8hRPxB7/EjMteq+CKLXceGWtxRRZQ4IjTePIXnDQjx3yz37tBpDMbw2vcYqsw5HlimuhA0mcetn
UgwROvHi0QhgIhDQ7pTexXk0XxCq+otXlPsx9d7d2OKpWV43SCI3whOkNoJ+TcE5LiEQnWwCkSeW
t/Z9oFoTBjimgiNjz1eRNFfLbXpSiptWVqQAHYR5dolG08B6pVsBHmbQAMvZdXZ8SE8J2aDfoFh1
f9szqyG/AG7Pe8XYMRPSNDwWvYvY8/wzBgRUoitmhcDcGGyUGglqSX0Tz9K/BTrPWwMAuHvCKuZR
twyPldL3PumfsYI2tRVumuDk+p+cRgrE6MBaOAl09FwuFxCPmjq2ppNbfrKDQujgqTksZgDdi8PQ
L8doGbr/xza4QiKtwRlIMOVurdrB15zdbRbt9RLzSMonxd2jDOTegKprSf27A9uHEpsC6tRDzezA
F7VTRFA/c2vZ/Ik3SrM1c8PHWOcmX1haP3oireokBaibhG2q16fuzb1NHRYJDG3Jn4g0go1bBQlf
t/CRZiZZ29Qh060gdk0/Os01RaZheCEF3q4RhEhvO32XSkf9ZwXnD9ZQLWIdALUNqEjaDkNXYZXx
BhGN3j/E3tvBAklv3t+n64Yq4AAuJWXobyTpN07T5phU8CEynwXqWFRX5H2OGrrsRtbszwruTOTN
Jd9nXd0+xe/zcCwWdr/gP3VZhp8C5FJGfF0+nw1gnFhkNTCo0PemUNPPWgRDFNgBSijMo+nz0P+u
O5X5MOg1Qe5Mix29y33La8M9Yit0ZGYAJkMeTVmGhfx6dvezruWQxX0dn+lrnBLAR2RIzVsS7zrm
ZFL2MXYDj1izbuVz2jon8bDaIwJsa8P7N+M6dNfLwbLxDX2x08i2fyx5eJTSIohGHOHWBl/+8jCy
sT1REyDMRxVvfsrae9/lUoLCmuo87JGJvs5NIVw9H7clTeedV2G8G9B3KGPCxOs+q2NEjlhWC9xk
PgcOv94nwAiITfRWAi10TcrN3xbyvs4eiQ1p9Jx7Ag59tkg/NEUV3dpQXOhsd8JcbSmGonxwCPN6
depUC7CtIdqpAzqI5uIEZFs9rrlV7edBS9zRO6HImXYsHhhovGcNO9Hg03TyxKNxWP4IELUIz06l
uKp3P156aykrHV4Yt37WZp6nsOA4reWBFSg971s5XromnDNc+uAmCYcbtZE0ZY7JbA0cMOf7wHJw
bMVPNCl3oYABskmWdyvIIo7WKTMZ6vic9pqXLm2lppWfsYAOkR+ZZqdvyjrhvk+jZecP5bCV/Prn
VXpYm0n0L6Jv1MW0TESWVjPOduDGN/5p98MqLzflmT2q+aVlXj+eb9Zxg5WJyID57qL+dxAoyQ96
gi+WpZ2fdIzuqD/puDQ4PjjRfVL7iiL+f+fwyug3hcXfs5WHPLNECM+s62XksifL7PVJxdIfvGt5
t2I9RJS6LBH3pwdDx72+6oQK8mhIiAChH2VkjU4bvVYrC/eJ39r4IRKWp1NpMjDal8zXrG96oWqT
rPLWXEqB+oNzVO2Bx9hP9EMjk6Twxi2M1PuqBaOL6ZBgBS5whoQkCNo+/kkkSURl7ySaykZoJaFK
k+V3eJIBQJ5yiukV2n77JMTvRyoerNR1XxW2vucR/KV1+Wv5a1dbeVO9pJX0P9+eWC/AaDPTc+ec
Y+6SEavP6ukSBTukz6vZXl4cDH5n0jH0nPgW9R00JGvlSZjZpncucyg2g48WMFA7Gl2+zwsZ33jl
diZh1WzksE5Gg/prhCFdrc1xDwKRPhCB9WYhQoJOKJs/N+yVVo4m79HbbjKN4FQQEKZK1E6WP75D
KWVmLX0qKY/RpWzzxhF0bw6gKZE/MWDVcaeMiWxRK2RC3zYiBu/APQIL0tiuq2uqn7TkuNf9+reN
Fm0Zn/79EwuaUFlrv9iejkLfoYn3IHiEBSp2AJqEYlY1LgYbFJZtVNPENzYl8m6Wqws9QS1EEPCO
dQcE854rdWvAQh8yVruNxs06jAyZYrmESvltkYiCDWjH+fd/eWpmKeZdk3tKrjnV1eBBkv8owL2H
9Trx0/pjsdBUdF9oKA4y1MVulo5uAvhY+2PCzqGai8UgRdXoS4G7mue3QewZPCF2iqPjGtouVuwf
gTHT3dNMRv/koWF2eMF03HMgwkdTcIwGDd1asCMSK3xXF5NhByP/tfopKEmh1ytBriyT58heykPG
7ckAH8j7ZeMBwqUCOhl+CZT5rk2oCP7Hj8HUTOifitYYHGlAtCsKCmCubPXElZ+z/7emP5RE9k5Z
H9rfAR7utqFtnOxJJHV0uioxXh682VCQBQJIYl4cqBSb2al2YJHWhRs7NToIgrrq3PpnVvF5OXSb
ZPjJUPdv4UkdoGrrfRdE8A2IqYWcyLWV5Q6g0oPJmu/yPdsS/BwKBIpEUJuHga/3oYTMXkf0aqDZ
grdP9Ag2PPzXd653OvOmivyQeWItXfrY0AWVxZr80S/UfKWh+pUKolZCSe7cGaB8AK4fEMKQRzlI
OZPg+7b+gspCk6vlsw9Esd5s3vJny0qz0UjnkPcuMc76MiFDKvXMeNFDRzaa0GaTIFnrZSRb4DSO
/t0rJf/LX6v4JC2dVfzF1QsqanPdpJFYKHM4yvkCyOISCc61Y1Jo0N6UpW/v9inBYiFIq9FQ+uvG
lZD40q7o2dyYGMLLMONVqPw7t8hHz8Zsmkf1m/HgtUwQKjVs01deNpYzM4+tg+wzlBFPwQqzz8PA
polySIxYz4u8zzJAM57Cbkh9Co0inIhzUSnnp0BYGRkcsV9dIm+3l4OfzroXo3H8JQAXdl5PvJd7
Zb8mzILuUqST6VH8UdFlVzX8knoJ/D3wy6eSyo+cNqZm/gnv7jtIEutZKA+XGWznlV3laxaGuXCQ
XP+HezhBMQ6856YTAkFdRcoBz4xXuzQuiP/pFpgML6q8o5TpLalBHIjeA302XuOSleVydYQ6tzWm
MzBv4G/M7x8sWJ1HrxIlEoQvAPuRC6Sr+PB1qM84/KATDJByjQXxmuDS4trR16eFUXqBGgcnNMjb
3KLfkfrFJd/wHSgVSp1P3SXr1pO51uBgdJXk0ZX09iF7yXWeuYFyetGI7MG/NO8YJh4Vk10oiFN2
O6hofsRK+DJ9YW2icMkQHGKVPhOgNaFH6n7IOZRx9eNHaAww/feXv9iPIGvvrbQaATDjBwjQAbKM
bhvjraxk9i/n+lAhtZotD+vWsyVLcMHbjZAHNyg/59LhUO0wfWVe+vUSWOrtaJmvLt4OKr/d+RvD
xVC0feU2ODMdQ/ortbxTKJtojfaVvoZ/Qe3/6e/3l5S+VxVhY81J6ToDZ76LQLN4DLHIVEnFpaEn
GSx4KlhKkKB/BZmRmhbJqhGNGyShtSkU5rBEGLHONnRdUNESfSITWv9uIZoKtedzJV4Qy03zUH0t
hm5wARjMmH4zCwumjFe2Bx7csu9EjBhYZLiQH9+QwleSBXoSd+KBHkVUMoJEKP4PWPkRVuUchfS2
pmJjdJpXl1fqEjk8FXj2eMadWdK2IfkXC0cXnUV34NT0ckjrlIqdNOiKYEx5mVJflKaHzZO/HGVw
+too7d7Jod3UGAPJXSmPrKv+vAze0IXZ9NNIK7hFtFQVbz2+UcooRr+utOp0xiLUG7XQGYEKdQQS
i0C7J61HFKLzzcL4ixbdDwRc83x78FCKRP2FImLZ7Wwl3r5k7VsGFUJ1UHUWNXkGOQZ6103riMnJ
fuwY5V5mJg1HOu/Kn7XKtEWLgOD05PKCua3dzqjj1r25T6mgkY3QgEObtafYNdfwWqpX50s6ouSs
O6iypVabwAXPaMeeTHh8MK3Hxq49ueMixmbD2sTCz9LbcC7KRk2S3eknEe52iL4YWCLFN9l926GJ
jhg1FeTuqNOpQiY48K/pNvG5IQ6W0Px0OMkQK8XdRZEJWzjqC9dwVCHsWxjHxzJk5YxpcSDbwMDd
PYd3g+dmhNVhgPEujGD7beQAqstqSx+Er/P8jE1/K1bU0FJhsBpzJbGMiTInLmUygxTVmYZjXCOE
ci417RMYBBx7FbXEzKWmaH+VGuzlz1zeX9BfTl3YpL89ZFkM00YB74KyMlb9Dg6sw8ynqapwrl7f
ep1lzBG8F9NVw92swL34cNliH2X3eU4Y1iGolWHj3/tOJdpU/bpLpafzfh/SG04GU/5mcVxeKDZ3
J6DvcThHD4SkW5OLdkV/GvoujArjg8JJZlxlhNS2EqtwA9Najoo02WRkEz3kbwkwXU+jdtSsVgC5
n/z1RwxRXSv4ipe3HHhbm5+YydSDLv8z5B7xjQXTG/P0Eq1AVTusaRcUNjjGkzDQLSlZgqlFcexV
sOFpXEhDbDvcXHVB8ItErD2ute/c0pzrCbqhXDiCVdRkrXIMwBKFBxB+jWdYh0uOHyOn2EYE6Fab
8p4PWZIopmzSGJqGPfqAmA6LFQ+FPDBnaJmD9AN/OiHJdlaUYqYjr+ZwjsTcmpnEUX+VMrYqSdE1
qpnKknKQ+GiK37ldpaXghthtXomivGVoDhXlxHdr+DBevZr5prWrYpFtlvBOSvPadzpoh4ZQ+70w
Ki7CWS/aHinN1grfmBlLDZe2XwDr3BiayWKVsnPKq7kwm7VHZ7//YdNFJKQjBt5r7w3CnYkHPSmf
aTzWga3L8vZDEf8PaUmYP5NRKaghoxmJThR8mFBv1BSpP9WbC/5fdnZ7FywSuJ2jAGEjTCNkHi8w
hKL8szQSPtacnsNtzL6u8f9mz6nIyftXUre6D5AyaVzq40CYosHsQmQOf4RiF7YC6Vtg+oeGIk/P
sZxeeGJXqwv5aJolzE6QOYljvdggDVlSPkE907t8x3B4amqq/NszO+hHCM4dNHjLaVuLMJ2J9xq5
3KdoIyY2SJ1Ab5mbhPI10WvOxGd1QRAXsD7AhVNiWp3zt9uttGR1aLd3VKHcEONgn1z28zwnKuTX
xYXNNoCrcZYypOn5JbSl0+HMGKVj7C0XWkniVBnkJng+QcStdxMmBSjLD75sWgxrn7S5vTo05dWm
5as7s8Cz5d/Qbg1JKzZh1c8efon3qOgtd7H638Nu3Up7bofKurmulSQg9f3cR+4STY+OfHpUKmC+
KcMsBlCTLlhlbSNYlUUDcaOg0WDf4Q66loRS9HhOPTSN0qYHqbWkF/3MvmGA19AN6foiQfTsmNnr
YW1v6ngjvrj5KitemxGsdqHtY6eN81m3mV/4Si8JwJ09AgxoaL5RXTnMiBqFN28A5OxZDTubLH8U
3YH2fnH4oPmAKFYFa7Yo0eOaeJ74wVn2e55pIXNB59HXjdW3D+0jRJddHFyRkb+9YuKIjCekTJCy
pBkoXkVnlmjCKwnKsh1QjvdN+gsXl4vqWHtG4XZ0dOIVk9Jzk8SRI0nwNFPEHT/Bd+50JMI+JxOK
EwfHMJe/hda82QLbwBl+OQBqC+ed0fQXYE5NTLRNKnlyVCkz1+2yF+8kp38lDnmz9zVimV0cPh21
CYs6Zz1v0SKtO7M0rtUz7N31uBzMpLlg7IrdL5oDLr/rahuT5IoI77Ht48LDRNB3GqK5EnZw5Cz9
EqLujoY/RPkp3HGAeBOgPqCoe09XtLDdIqMbaNFXz+10tuhkHU1nTX9vrBR4EMi2G9R4TT0PAIhp
y9wbJwOmgz7rs2vljuuGC54nrjE6BYrh1MynJLzgReox3QLj4J6j9e6HzgqmrYRbOh93e9yJuebQ
fLSMuRyRUVmuIatgNrz5v0V7jg5moejJFT5IZw7L8xIl3kqDWelVnK71q5m78xDUwnuc6Wj0j3yA
Zy0gGWC1t7zG3A2hkz7GpmNAhGDq3kDhcbk2v+ejH5FPoihN6/tAXmgBXevxxHPdkdxMQS/7JagG
Vbm3q8KCApe1CMbz/dECmWeIBeQEzN924ZdT7tnHHOAGbXL3NvzaCd3YpwcLuWceITG8Fwzta0hr
LT9Fm+01oYB+IyUzSGrVGtgwZA7SpmWritjBoAluPH4Ayb6FvqyviQz7JytulxQx+BclQhgufxYy
SFub2QrTeRT6IQ700EhKXhQ+kqV1VxBEmx7pqSNmvug+t/9adRtfmp5lLtTU12idswr4Xmlauhb1
0SoYQ57D1ewS03fm8u+4zE8tQ4vPEXdOY4Qmj2w87Wg6ykcZ9NHTmXOMMh+/UuZRaZrHCbVjjyxA
8Aid9GL02WOg+SMLpBAyQJQ5lc7Xvf3kG0/eFVJCPd7gQOPyZTJlu1xQuFawOgDB/BXqXWMEbiqM
s4K6w2rv5sEzC7ZuxTJoAiQBJg7pqNVbMZwQpMmotkKRfawHbLzwYotlBgZDqqoLJvscnlF1bCK8
bt+fQuRXeCjL04u2NRIsTUmmk1kfhPukP3ltXKWozO7ls7A00tHW7M6Sth1YxhNCmpmOvtLjlpj9
fJCvIQaTu1kldojKiuE3gAtyUJw2pJcQloG4qGdBHH+1RMQAlvvC3e0sTPLvFw9S/utIeXcOb1bU
KAHEdkLpvX39xcH7i/TwD1D0Hn0b/dFavxqzOccm5q8FGeuYKYDnHTl/3qVRNBQinAkMN6mNnw3J
28ESMRqU35uQkluMicEDuvjk/CVbUxYVbY3bsnOX/NLtjlftIYtA9Nu4aj5AlnyeL7/qcIw8q2tp
UZMhNS7YoZjC9kAcjF3biNlT1TV1EJSohWA/uZYhI5oOPqPKIW78Ir5QSOPA8wjt2yRub6/b0j0Q
V+Nb3Ic6A3+7FoEYTZ2bkmRh3Jl3TJGzfsK9WOGPhxXiO89p811l/LgI1ydjlKPC5iJkxSEqpEol
iAt9VLbj7R0t+hTxLr1ZJQRF8R/rgA9vRR0pJwYjIQuhyeF0VefP6sCQ5yp0RO6RPWx9fErxSYyp
yLKietT37AGpRLhhiXzGAPIvQW2Uth9njOcKcCDpMX4esBphLaV/XTGSQCwXmVW3SPr0m2LuM99U
yXUPkcaYyJhq4aolccwDDkaGXqphqcDIyXT9yE8rvTxVwGIqyZfGgpi7MHIss9ih+/fxvGzAn7sU
3504L4tbrnuZWD+7TN4qFRaNPDAaiVJE5AXgnN3+CHIGuPy7sR7joOnDGpwrO4FXiPmzgcFlVAy2
B4MxjrzgNjl3egXkiqNFjhYmFilZArQmvemZT30IrB+PDwMQhDLmsk3ZXWOrGybZcB7ac3FgURhs
/uo9CpjiWxh9fuzhmIEiOniNVigFfXRZ6AQZSeLWdO0fTKHbS2ZxMYpoexOOpTViW1ng+p8WPvhc
665peSm/bht10OH5z6YMr1cHKtc5xAn+Y7JA0LPm93hf+FCc6/0VZVY9Cc5X57qTGjEkdlGSS8xy
Yecon1vTryzRMKfbnitZ4tTD2uvarEZhwxfUFCVcjT+uHGvGhkl5SNXkJqBWS5/jy4/KaGFaH9EB
YPp9z6VuH9EgcxOrSA7/0HBXH8YPqi04BlZHaRvx3tJs9drWEzwjuyQpwXsEFYTvEuUmafFSD4/c
cHWmDTS/4oC88SD2zj7XyF+6gIHQ6b3OZNGBkp44EXB10a8zxGiEFDXqt0Po1rNihOUiePKexvy3
9GpaWM0u6dPxFDRJ/1c+uJfch+fv7tcJnqS4eK7F8nnyV0kwZXL2MTVc9I3DdleMXntWRVR7a7vB
44cU6IRDL6dEhVbt1ap6tz9Ux9i1+7ge0b+Vb0VWm3jiiyOQ4Rq/JkL5T+FwAuUB9mtTDKG1sqOQ
FinWZdx1heQ6JMAUuzRbA+CoYUfJWZFdvZPupQE9KzJtigMNY2j8RH/qJwPYCefUnKFAHEHVFYVP
kkMxrqUxetWO61biXoI47D+tbeiuCfvLqfpZiF7lRfLW+i2mZsIbMHe+Q9+OU5UEwP0XESGXEwaN
5TLx4CpA+eelJE5fHEk1TUUbJsp3AhS4w1Ax87QLirKQNv/Ksl1AbR50LRX95k74GDUfN+9nC3f+
m067eHKWgD7AyG4xIycCVHqWhJCZfXbE8WCtjNMZ1dr5Y6IoMay2/b7HGGeImvziUtiGV0kBjJGb
V83Nh3Zca2G1PkY/RMkpGDUI3VlKEK5PuKi2ON/MP4biWNqWB6GTQdk9bpznFqOAorT32TnD+TEi
LWC/xBdJAkoSlTHuDJ2o0bg+udBphXfUIcO6BaEfoxLE0Gnt0RyJQR1mOdEu2lfcoNHFDCI63kha
FvP+R3pofNbdGfV5R7g9+egaoQIsbZFpz0lxpcMc37tQjfjatAdrZ1gNECDcGB+L/M4rqG+4Yt5u
BjVRPj+0q6cNucOcgPS2YjF0Ea/Mxn+4QIK6TZ4tKGI5re4kVqVrwXJjXReeoumKHeF6M01h8o3C
UyZX8F21mQMi3NQEy4hWwJ1fSFj8Ccy0hkBfeR2JLMseV8ZkqYAe3kxXT0BG1l0oQQVYAp1Fv6CI
f0awQodcxD86iAh9XPA1zrESi7MGyZkW0lSj3CbH5SgW2NGUekISF/z0fItuMZXF/fqDr7yW9c/l
HoOUFcAkPrNabOjXIw/7yLwZCR7lOdS+/KRQWA7s9gJ+i22yt3+183yXrUc+BG0g/ulM2SPbf8SR
wIV4TPMsOF+nT80SJz0bqnmTWzEXRdfnlBHhSRm5eYafpVvtz3ZkaRSV02By34mvKsYBToHkBdef
ZXQBGQXDjHVLLg0lKR7tHdvnsRrSYNGPityVWV2+KgEbDUyw3mpD/8R2DmHfPfGFTfk3m0bmOflx
Vy5UCsgtJRG4pm+dlquGs6yEUzZUB6tRHxIDTh1MB5km2QXoYP4L3Dwdu4SIsW1l106kJtUeWYwy
lgo8gq3ZokTqUAC0zC4GhFuOYJDyTpXHYyxMA+aHPxqSbIfpLivd3xB2ndKuSk/Tc/PrM0495+gU
AjleBfLJXZb+BwlP93G8AcBGVk7EhSGSE/SRinw6noz1o/7ZEE+HSLJw0XeCqGGFN0POr6xPyF/Z
pjcYVybzZk5CCMHgK2qhtR3EULOz7W31AMFpED7AXNuug1onNIFaOKjgosjeuP7VkGGhWUVh5sq4
iX0S59xPT2/ho840NhNNRUCfxRLD5Q22g2iT0u7+/pM+9Yx1zaRKE+bPT72ilnAnyRJEAu/2y75u
a4HsRBTPvGlNc1KhUodrOmY9z8XvelE6uFGWu+7dFW9j6rHfUhWvaidkis7ol/HIZXXKgkaBCrrj
3typ9yNt5Q/kV8rUCZJH7mEw2M5mveCFuNMdwJI22bFPDt6MuPNxJbQLRiTuEfu0W2XH/icwRHuj
i7tmjBY8bevXG1uAirzfgjVJP2Zph1hhQwIqPKXeNip7I2B5BSSVs7o8X65xVRQii5xFQKBTnAGq
fUesp/D/I6HzsKh5K4YXoSLM8N3owMAivwaHj9/EQhG+kANmUKGrmWLC4ccM+MMMupS7+DZC6NpH
lg/Jl1PSkxRnL1gx4snsAk+JtGyXw5VsOU4bCHs+JsdQLwCWG8nEoyV8pW1/J1t/cYPPp7ZemILe
ud0Vt+vzT5/EauvCU6Zgf+AIKRPFPX2gRumw3UseyY5aYf8inaZOsVGu2uL3ZidCMf5qE2j085aZ
FSmd6V54SMgFxToKGSTewh0rX6B/I5iNT71awUmHUecL2RQ+fRZvnE0RvpY75OyPOXm9c/4prT1X
1hGNtcgzl4qIjLzUjBQqBXhC6FdLprcP5GvbNg0MQm04YOYwFbo1g0S8Lf5Xm/+1CptIMpbTScG/
AgUyJDg3BxiO++V3LlmnPRXt8t4cj9+E/9/Q2EZGZ80Q6BoYiTmHPQtQKf2112RtBvV6KDy9WFbs
J6GO0gPCkBdln4/Wz9tuS2eda3B+I1Lsby9YQzuMaosaEf98vphs82GoLcdccnizw68tNi4ih/Fu
9rvY0WOwFoStSBVp6OLBOWQTRqnsl3QsFw/4dAvV6qFdTxfMqIT60K9JdDP8iDFNV/22On/0OrzS
QLFqp4sB69hUPcjMWRyiX5gra2HXcYNrW2nUw1BAatjgG7gQ/zfvd1yCMfvAkaYM8CK244dzZIHf
aHp50KleLqEj7wcEkkiMlNjVlbsuHcf8Km9aFZSc2Drthg1MWzfrzsqG1CdqfEGqUadfwq1Ecjoc
or1VwmQBUmygcF+XQV9IWbYBw3UkXIuowMtbaFOxpGxUTYT/Ym9jpfgv3siKH9g1bTZLlOgDmvwk
USFgY+xGg5v0wBNStM2m6jsJk07nn/OJ7LAulYD430penq8z2Rw9vT5w4eBLjWPVXMhsxQRYSUTi
DAH+QVtOaDJijf9D7EFRJI7JAq+jHlsLsxVTqQvEAUzFMmyLz0pk0npqWOajegZi5w+vxgjvIk0I
44DIUR7JlqjqCktULv0y9tp2HAvZz0Dy6x71QITbTBrvfJUSIrGYkupXLMmxZeOGfkWNH+pqj6Rx
Q6dwKHOkantp6enaREvWJ7goC/rAuq/jWBjKhZSxRMkq/fkqzkA67JK2H9V8fjUTI/7GA/hASBd3
oRtX7qoxo0JYTVgOdeD0yglNOdZrr3b0sEgkAvaQWckP6Ni/lcC6rb2Be5KAPi960Y5mfjrn4Y86
IhU2ec7NeTDu2G8Cs5ctYAnKWTR+ZH2h8aAZpeA/9yUMJMXkrhkPgtsYUYWmBEf/3M57c/ylck4O
EuJXlq0wF7AGkWVmnR1cDs92Vad0rVkzyfSNOqWxHsoO+cuXjySOO24tnnRKksjUZVya2fpUXelf
SgU9rKlnK0VVrfzHT0BaaMvQUFVsZwHoCenkRj99+i0f2/ghoVa8jNlBLMzZp0je0Tw8C+hSUthw
m/QSmripv8r0sxWN32Hurdj2VngLtz64R1II5T1vJTXtDdpVADwKjJpH0o7ovfjn2qZ2vinBzrWE
N2PkAE1/yMNxKP2VMoOOYw2Kkm6OlJN1l8IK8XxdoSP91XftOr5A+7HLBZGhUSIvY9arVrRQ1dYw
xUuhAWG4RX+sVWZQ151z5/GgwwP8XiQOZSUFXFcgmqTp+ORxlAxy2dXuB3WUucNun1mKVwsDMWLI
mh1TlPiI1mJBzULu3YAYozBlDaheZELnYuwGBbr0kLQ+vIcqflTtbN41Nv2y2zUdiy3gFwVIr0S6
BMRmFUsEeHpcWd8L8pCWP/Y4DsQQTvMA/ErdE0QaHwdrHcQyyGVXysMljRkaEv0/Liev31mEw124
iO/0J1G0uRPdhAGPRsKPcTuRFWyFZ7X4+LkjrL4yvvdFdCPKp+fFEPj7AixCBjp0VXY1HE0Jfk5W
5jpZbHnXw20gnBlIcYfb+JZUPaMsVpx5rMTyAHAptdD1J1cOQpHqSthNcRvFBmW2aV8V/jyIh08S
EMdjpYX1diROoCxivx6pl9DU21fIz5NtXT0mhh2BrsY6KEAfDRaimgX+3HIwobMo0kjE92ZNrc23
4g093QUKSEbSH9T+Nu2d0qOIiHqIN3xzHNnHnzeCI4orXXZev7q5UawZM7eKPJt1cFMc87L2+vd8
ubAnybY91SkFW87ojUhxx93xLuUNstFasy45MZE6gErV8alxr9254vSSg12ZzxZ3djYNF8h53/BN
eOv1msD3+ammpfpMDcrsbuL/FBKyfYgGOdNmwiF09mJUHgH7cXlHt1w6FT+MfY2rVHOlaVsxvmc5
QY3SOVFXXpZ601q4YeTQ9CZ1t7QFyFDFL2nHTGTGFGnZmfw85pdDQk01dE2zROrhppN2HMYNJ2vM
53pdx4h5ceCzKsTJj2Vs6nX1YcfsAYZhuKVSCwYsx52l3me3s7OYeU+Ki0PpGrboUlWsSohcB7Bn
bIha8cxZvhXgJGgKgSTLD2uMDc1yY1vPs8UYyNIKbPp7nvVDhl86oVxIrpvGNtBP5V1qTe/VOeHk
S5Bf78valxd3350awl7RzFHfaHwGjVMIHKbLB/bdhUbFW9TSg8FWofo4cuMY0pREv8FLX0RaCKJQ
fmyDmUIzP1i9gOSgORk2XezqLP0PXWdaKBIdDTcEvMC8mU9ZqHQEkrLYn6gNwPHSEerKsLWP1bMV
5f36rYPfQg3W0+62YlAiKHfypxJhlXn+fClUx7qePhTDpsZstczqqMPJsRbiE9OLNs7Jxd7HhqB0
E0+70c3PTM9vaQGhGzSL5CuZfNzhIFQEkK/R44odAV+93RBXpNk61WuGOGQuDLFZjUBJsNyk+am5
LZNBeejx0M8pKm94gQbGnkOeG7LTGVEjhDkSsq0BsRA1Ufrl6O968GiCHaq1mhppU0mTcT9rICD5
IfKxQ/4wplihQDp1cGPT9U9I5aj/q4v7Rnu6K4Kcqz8DdtypoWpENgw3TN6jDI0FXvb8SjpBwZgH
esZ2JSv1axkAoHyXEQ/TzVHUVMuXooA1am9UX1vDuv9bCz+l+K+yRDvAhDM9/OquxGJEa3o98KbX
ecjgZN22f9EcfnalmEIDOhVzvOSfa2bSuE9k64X31XQP/4Y2YtqUB5VFCZ1SHbOb7oDE43ioxEyp
ZJ7rbFi6Xz1BANKfcWL1IABx8h+SJEoExLONMJr7Ca4v20Rt2WWrvKZrQ1z/xu4/ombRfkP3yUuO
rFpoNjv5PjEpnPl6dLxZ/8lIfkKGAfH6dMyQBILewu7UmulWfzbuRhoQpTLuzUm+7OzcUy8nm9uV
ga86TE5dBQzjJsSpaZYklGCvodRYfZHy94DZTL454i8zT4ocbN+F7RGYDpOPJYWdEobwdYQlWzNF
uAFnFVzBj0xmVdulPzag5JGUyGPGJILwZn6WwkqoTyBBdJzQ4UOjbHk+SIH9V6Lj9LsVVEjLPiNh
el6d+TIoSpr07VSfq9wOaZMJZiavY3t9B/kXDVtZpZ66T1/Su79ExKYVF9XPBpxh7SUhcRtITixs
tvn5x38HdL6ukFifQkxgI8Ggt+S1Ld7gyUsEfQjdTg+QjNDtRrzAxCwGl8gW15VDZkutnhzz/RiR
hankTFedaAfFSR7TEy1qzHmtlySsjnTFAlXOZuE8Mh0tkoVHgNUsVy3i/pZ/XEMHpdBh3+gsbH7E
0YEgZrKTIlFZY6rQrMmLr9LLiA50fOgngzZGqsMFvFExUsxXDc8vDHSNUD6bOLoY5DbFEWKimq8J
eo6W4xkO/pjwpSfPUG+Cr0daGDtTE+KvkbF3Hol9Yj9XW6UVckjebb6OySh0KKfIBoG2J19ZN5Sl
mRExtESALrRQsBcBctCh8ts/bLY/cEWv8cb1sVzFkUCUzAnMMDl0mvm+iZxKnUwI8zjzPCEbJFJ4
nlSHknfS+EdqrVNZCDRc60JF0WV+cFnJ83433mbsr6qRSE3Bv0QrGlpuioFlfYKHx0WyTnHLu26s
SrevtldiS7UJ/HbzuReT7YpTghJnPYsnpupU1rKqUvb366dtCimHNfpnpEs8a9UY68SDC55sHHyY
O+A1e4x0nyao11kiYx+V1k0kRmpN2fdJy/kqptUSFETxw2EILGld4JN+3cf1Q7Mg83TaZ3BshvMQ
SHvoc2snzZt7IW+QZVCV431uvATiGXFL85RpdL/mFloZ2USfLnnuDlWveN+YQnKuDSm4lNtjpqXA
SeKBqPUY09YkX4aZhVRjcjQJC5mrQd9Em3d6i/mtTUQSTIhWg5w3s5//lwOJY5aHQ57zAT1M95oc
9Pu9Zr+ieUcl8zGWRxVsU3jKpO+Sc1PCH0G78n6TBeh4VZVE93St7SYSiKjmXArPq8eHvJ8xvDmO
2Amui4cxEWi++QtK1IG4JSw2G710DLtjXe/7YPo2fNP9YK10VgsJiKn/Nnz1JnKNcBuyssP8dDMP
ImbRjfhXJyIvkmD7yv4m2mnKuycCKb7GxzwEsDDWINrsVqQdvwVJF5Dk/OeEdk+mIx6N460CuR9I
YWOo6cKXDwY+avoi8M2zemoIQsuNyFtaZA4aLHzox6PeXTmikjOra7hr7o5xMGLwR7DR+KbQiiAz
L/N0hmA7xTGgjDolG1pg8fRjdaddCogXbr3yY4oWScey5rb77h5Swx+OKR/3oAYRw2o6gM7jrYMk
HkamrYke3J6MnPRP6HL3cxWiALvKsAf/7t6i2mIkgDBzu0/oitDD1z1VLTSLvNX4GTqk9/eKE1w8
oU08u595lJ5mXnXCUcoYN26nG0pTnYTsa8eR1BabXghsnslBD+oY6Tjq9PKY8c7ZYw+9vr5InCBe
4naPc/BsmOxyKi38MhYJ2+CnkK0kW1nbtrR50mhmqDyQ7rLj0bPomjLavQuyBoFFk95wTtk0Sfls
k4Ev0I3nb0PM6L19XU9weSIIU1ayDZPXs0m8w2jDWx41AmDybUECS3x1QI7P5OhVNFwd0zmPU2t8
mPUL/3TAnlql4TTUNwoMRo52B2urgGduZrHmQfvgpMzvAppX1OQkFQZsnZRqwPtChflV5JRa2NNR
XyOm+9268sGOk6FwE/j6JFHAelYYDHZw7/vmmwTKSuTzgPUCNYLZvWv4464PpoG+dwxMS5DBZSfP
dCje1CMfftvlnqpd37bi3iJvrEHx8XzaD9TWa1VhqO1P3Y/r0nNPRxSagcml6NnfG7mTHzPVEqh3
22rHcDDTCXw+cX/nY2Epcrudi7wAyY0vvIhAulJabxM71k4grSrYdZeJs3VwuzjvnOC8j86EHlQ6
pdeGT/6PyEbEnsGQCD3ykX4mKTjYdBs1w0Dx4NH6W11EMUC6As7KzhMQ1o33PbK8lWt9/nkKwL8S
aH2r5rRIQFXpqOEppNOq1Wyuh9JLjDMfoyjBbteDJ/112tH3g5aUcmSJfo5up+uJAy3MUn3GE0aV
gqNHhnRQNKqbl2DZSsOSaLE3QAHLkIQkspQkp/bZrvx6snwR/cweMXOZj8WfLrI+blj1fRsvg8FX
f+1U6BBMiMNujnExaL+vG01Aj7qyiksSTfOpA1pbpYNvlHS/0wQEjaLcgerxpmS89hGSuIkHK8sQ
+Wd35cVc4O+O+e2piHCIQ5EOfx4ZtZ5Gybv7NnszwxWeUMkFRlr7CpiBn8VSm4Ri096QyWX//cbq
X3fTZx6JoDPTaaiMxQK7lKwbU13PnNueLXgx+OZ7cKMq/PNRNrjY4t1GdOBChmh8rbpBHl/hFZhh
ROlwvIRWq4TrLLQQdwJdI/QIZpeA3hYYYZE6BIQTYvu4qycuMvShpNK9eCvda63OljADiJVlSeTX
1ebNW63y6d6FCpvgwKRTan/gqMtz/S4t2Smnppe6GPJJ6ThbmGMrUGmkT+CGFC5u1N+kudr79jQg
AKtXbLxRaq6PQ2SYD4M7UavzLB1B9DN3CFNBHSXB9ikp78z+q27DWrbSavblFoNvH4GSQUUxRkmT
+Oy2CZgFnw5Nbqr8dQay59rdZSxyzIZ0fEn8LQVJgq+Z5AJc911mWO48QG17qJWBkCj382ywLf5M
CguYOMdYi44oLjpNtyYAk9ONsx3TLhRKWdnwXngGkVd0hz9lf3JQCsH24UjSm2GbBBlHawsX6LqS
BrazFuJazSfnBkeFk2TFvK725UFnXSy0Dyqf1Ub1oxB9DxluX++kE8ascy6lwycmykzOouw1L5XW
eBOnl2dmguxgYry76IYqLvoHxl9tt87bNIE+gZsQPZpsJzKoVmSyZscFxbsdxPnb/kkXGcE2YWlW
C3ubpffYm/6MW/qXAKgcGugyQSDPV9L/CXRl8HeVMxqP6FDZdmLms/Veo6Y//fy6Pm/3IH45eH2P
PluyNg5SDZIdH0lV69ULgVmH72/xewbGHg/R3u7GJj/7JoDRX9+TDCa4FOLGr28J+PRwwBtymhto
3RGnHVnMU0RgDv+rwYHrDtBarNiVviY3wY7UYI5HK+dXMNm1dIhpGienbITd6ZaAPKxo4RfbM+wC
8FMV4kN2d7C9NP2aKgccxot68OBLAEtpK5688txD/1le1uIY3izQmBMbar3u8BfNbbOMCb4xSv4I
uSHmHg4LC1HXg3SbjzVO4ZBMqssXacbK1xorHUd46qVG6skosY3i8Z9TLgH3QDJDn7AbZxB50PSC
akCyBzHx9isjsTSbnPZ6nUFwuTaDNacitx/YpLxLbDktxk0k2Ha317SEsb46Wq8HTtC27W1hplMa
ISZ10/02eL+Yij3zJJZCWDXeY1CCJalymA2c6ySfPmImEvyM98xA9OK6b1F34vyQZOuxUUwtOCX3
b1wViae9VRfV1mrCd6ArEjiOUUYdbP0U15rMYwrA1a2fXVOnIA4tx3AccpK23Q3GWFZVMH63zpKC
D1YH6at7B+ccgrI6Dw9/G3a3nzkt+gJk53rjsFPoeDTLTB3VoMuzVT4pLY5/P4sUy/WuQDjmv5Go
GOJIPpjw+bTbwUKoKXUhRDygeK9ZLTr5JlKxiELV507FnpKmPj9yeMxMfshORpl400VEyOmIl0Az
y1TMuD0k67vCQXNrWkg2+Kb/xMJbiGh8YTgu3cmoNl9VPDeSXR4rdloYGA2pI6HxnD612NrmWfZc
/rhP6LbML1ZWL7ORDkXLXAoKQONocO44N00dKEnkxakcPkc5rrSPCohhVCxAWcqq+MxIQpV1KoW1
H/ntP3AHmu37iDlXmA7G3JBTNbLlvi69gEwmjS8gTYrBJVOcil732Eg48Iqgd1eBKdc24W0Jd7Ox
l0QyofkXqFmRFo5hdR2d+yEzFmkB9Vg92e/9W72Wybynfp4GqKeAMLqpUK2rmf9Laq1LweNgcXfV
Z+tlXiDxJ+1mZqkDYXpbJQARsVeRjpd0lvnUggkSIun8yvHH7IBMBKN6Hfa33p3e2EEVybeQNcZi
miCWTTfzX4Jq0M4gbzt6fXAqbUT86p8LgG+SU4oK9IEBuWzEQr1fc/g0ZmfSOGMbbjADaUGTHiNl
KSi1wJVcVFBK9Cgy4l5x7lSl6UdIC7cbg3yHp8dfjW/wuRDpOqE6sOAiXNZ8++QF2boYei1IJ53c
OOaFHEkILmmQk6qUzAXVy/sdq6rlBBhpS48DZ30VctFDG41da8ssx70w6F6NZ3yv5el75cSQnKMl
s9QD3gJhSfLwLaJfcGVCLEjH8VKghnMVdPsA872QpbeuW8OZrUQy047Z2bGw0aJhRoupSYWZ3mM4
GDGt5KvQNgKBdJDYCA08UVZcPTjVY9MUxzhop0ZvAjW1i7VYppAhXYtFDcut8GeclW2LbAFCKbP/
JbpimPF0g5RUJzciyEfYGld1n0fI6OdzPKo7Wbwx2ORhQVA7QIK0286jGmHmhPnaqxNnJRGFUTLW
L1NdXYycp62a/i8vsjNQmVaW7RIJYU6B3btwG+YjMEif/RHSEzObHhICA07zsNzkeZzEi99bl15z
xJwPDOaoamc0AanCd1iNyJA1YI2yFBVVnBuIUCpU8Hwgk8BnR56gjlCd7Pb5fsRltH3itnzGVdFk
k4kJKHkWtB9Ezh7jj+aTcrKlA2vfXSTAjEQC78Eajzkz7Xbx1NfvEikjtA1lgvT0EwUO5E6dqn0D
RttzQLNpIaKoPiJmLb8yVqimyHI8NPLZoX6yQ3FCY1T8h3CftYzIEIQ/7/mHPRxUexqcvOF+W6fB
0A0C6BHuLw1MyDmrHrf2tLURZlP0WEsE3ZSJUkewLbFYDzTP9rSZXq7VtI46zuwqEbB/BMGgz9Fp
4rtcJp7ZRFfkjYRuKQSHADGtK7h1vspQ4HwiEXamA7X9UWsUnys+zDhL7j3j0f44FV56e2p4qC7C
Plk2BxRb45BnEGK2Gr3OdgymoU5Y+Z99En6IKQ899BE+jtoP53nZQhuDbseTh1atVydCWtLjMV1N
w1y0Rd+m/+EAMqY/o49rdxTCSTdXUxMeulJd/5K2JN6kNRhhgQ5CAyNCncmGjPhRgaftnvua7r1y
QkkVM1KvZ9IyG8qkQC4S0kDgwDb/xbCpwEzEgdoxpUVfx5OmEeD/Ib/7mXfqzmxefhSNYe/JmMKA
p534naOTKh7azbKO+peoJ8lF2ry0XX7L0AV+nXyxA7dVmYFjgayprZ4a7fb8tmeHlKSACHUHMryL
x+u/34dmoNJ9JCn3AeaNJUVa42Kf+mwnW1HP46f57m7237ogxa+K739+9aMP0WxSgLmaXmDdkO+o
D7thAHht6S+2SeXTJqB5JvD2AFIcpJi35wNr+uiKwHJErAH0GpoEoiksJ677KKsh4ZhnT10aymuW
8OlpZMCcFqVPacWdvy0j2aY+blynbpVW+hTxLBs1Xy6+nvqnh4arZ90bu3a9uJvM+3NL0rdq5v/d
Y3qFFBXEROyi8Qrlaz9v3dTCQBY86t/d19/Jhh5f7jQcEHmgy4kshONBfurbF6J51nPEWhNfFLBr
yXTAHHuVbBzTHNGJ9naJdKJCidCqhBZbyOeAPgAKtIxD/AprsA6M7SDYKrIKpNdl5C2PAkePzl/I
6VuLk2umOTqgecUEK6WFYVdSc+YSIwyd05cLSoZw5KzrXPZ7ZnzcC8vdLRXbSyw1pUE0QCByt5v7
VD/+ySOIcEk6H44riOG3hYi2r9QPJ2Z1vYw/oyzNPh0Y+o61+DQ9lL3zbi4GRqrbF/IKsOBqgP2M
adDOkOp0QMYseJenei7NeqMLUpPZNPqooqFgXrldfc+FZW74Hk4Q+ERmdedQh9N5cZ/+7mKC0Xh9
lh74q9HJkR5Qj6IPOFFhtE+lmkEd51TNc3ZhQAEl7BsbcsyMtd0svmsSQTXRP9Az7RSi3EWx4yI9
B9gDA/pgkxKCIIqInDjPwmeCOUfuMKoU8yFZ7QqRFddK7Oo6ReAiF7onbjWude4gS+/h1Yu+2jWR
MoNKzlcAh6m9IN1wBSFwkMCCRVBBTM2IfjygwoTgqI2PAto6HpBIFbSD1+5DxxQ/wSCYWk+Yp77U
n+fCWkg8Pgk4YP0OVlqM6OP5D9lIiMbSihEc+LgqZrQYcyvlFWGCdK4ceuFNe6MIRRl+AOsx0mu/
gCFIeKh6l++XhIHVdE/piFj7Jascog7GrERLcxpFUsiBsWGjuEDQxRdr+BsCeaHM6EeLvgoMAVLs
AIF9zJkPYPATs4nyc6DmQc7zSw1azGG3uuVUMmQJS68WmoB7EfEDeXmEZx8lgrORA5YCjzbx08bA
Hm2z1knz/mWiZ5vMXYBgSFC9GnkfJvJX4GvpUfcuXZaf25byNu6sRKGjXPTy+sLymHOvwz+YX8Fg
cf7jHoLuFvAeVB8CvyVAkwPeP/r/ZbQM0z2PIYFdZrxqIAY3sezAsjgz2jzd/5qvv9XlV9OxpBk/
mpAwfb//7eZPC9jhcJiBiGeIX7jOjqArQ+GkDFAwm7pRKTtNZC6YD8drYkuCxLJrWehkXuvItEWK
9JjmouctdULgnxjiO99EEVmZaTM0vMUSh7iY3dn8puUaYor3gYdpbbbpMJNG7BWe73Xmqmzu+HHE
+U9qmxAQ2BC5eDym9qjjjKffq1IwQqX2zNrCtK58KfKAyt/Yr9to4AGf6mqZjqN76Ttt0fwR9/T2
0376ic7x08+K9lhwUjz5ac9eV6meSPoO6aLZ1mbFiqf/o5CnB3MDNgk5O8xJWiPfiWF0++6kkA5y
vZCKCSDYrGTDCU1qDyUehurzkBSlWXknMrP8RZjZ973DBPXbVFHlaGbgTy/eISoWfHWNG2Feohl0
wcwnrvg9SkE1/3tgktYrn+v4+Etwytr+KsYxVCfoPl9A5idUwpXt8KOMeeBhwVBAehmrD7zoVIZo
v4oWqamgxORuAqgUNuhN0HHzmNjhTS1SusapuKjTyIGsV0PbOwRc3SbnUPQrKFLy09hg8rudFrim
x3chUlJ3PDbaFIfMXp+sMYw/l64LZq5ATRpPr7k5G2gwyj7ftrrq0Sz+bvjhP5wt6RHb3nGDjIBW
R6O+LyZTHiUTHA3vPhtz882awIJaeT72ujacvKwas/Kt4QpncolACsJ4Ez01Y6eGAyUH5IxdojZT
F7+Y0r2s1srm1d+TFMULLoYIqjBp0J7PiTtLZRUnS5BPqQD2VSyP+PyWWzpgeAEjJkAm9JptY5K4
DLXggFdoJYqEOB2KVV//pP2vp0hllWyPSGbsv796euEco/ywWrXFcxGTtIZlmBgxQtKep1dUMud3
tWo4pzJ4gY7en/JBfcN1ateNLayZlCpo2de1nx5lJ6miB5WCdx0oTxGYMidSOCEPxQk8x5Uv91aT
EkF0+8qX14PUjrtFaTjPp1aX+FPeJo7dY0hZQKvWSuJajg0dNNLQQhQMp6kgyGRBOPdO3fmKdoUn
dyb9kM951cGh5xEyBvikMFrB2eqdT1FHOJJyrkL77s3pNgjSWMJR8GEy472U7oCGiEb5UMW4nIsJ
5i3+QyUk5vE2ilOh76fkR1XvpzTuXO5pg9KDLPjqetM/g3ywIRP3a1P7kAwV9V6EcEqtbXcWltHB
awgffkvspyakm4b5QWmxxSjUuUZeFs3MhMd0FwuOKIhfsQjcmHVU+WQstvJkZbxMySveByj9ew2K
8plJ/0hzWDG8nu7e/mlCX136hjB0JMacJS6H2ROaCLTSzxWxJsKyaSTHeQFBD3azXpyhRtNm0gCW
+aG6Ef4vbwCA/Mrkj11vLrcbdDZ0KgPK2LdVgsC2EJzWSnKjbDm3TXToJjatjY6sUo7/VfMrNNK6
YKJ6AoOOOYNkj8RNRCCBX3Df290yZvrJ1P2U6t5LQ9tGkp8HykW+dhEttmAi4U5C5+yx0a62pbO9
TccIO9uZ7jafp5CD1sNLx2niHRwhiz/Uf4b9FAkB1zjHGr1O61kVCFEQO4ww78KPDDHXsKGLXyxV
ghVqtLq7Tz5hYl6YVPmJD1gN1PnhcZCN3FfjrE9jft2ExsfXsNI7KHxmxw1ZX3zPD8eq7RULsEaZ
nGOAAvYvmTdicr1ySVk9xRp/PaJ0hte+oTrcNfBM9IHsgUU4DQ9GIBTjnNBVuxdW2LLq20lUmeD+
+W1LtTiueDs9gY7yzTepqu/MiPphr+Wx7YFOLqQx+cfWfK26TvsK1/T6Jl25sIBZTKeQtucABEyS
KJPWLMpPKT3V0Jd92yGeR3xXO+sf1IowTrdVCZiGkQALdBPG1qUi6imgYKGt5IheBGRZsN09Eyfl
w1rskHx/wU6G9Mtf7q1rHuv1YzSnbxCCPiX2tcTiY4Y1gtMR7Uw6L4L1SggHORLHJVKsBSTw2OVo
2sNX/wf7atmmoDCw2Px+o0gkL/lnxSMt7nC/YuHdHYvVzKXZwAff+Z5DhqrHeFIfhNuYxjCWR5XV
9X4zeHND/nCEu4aQ2d1fgiB6Ga+8Q4aKPfbgGVda/z2TrMVX6td+STXfvRh981QpEI6f7UO0NCGx
0mcOjeOX5rH0E338++Zuxb0A8QLcYOhVwTYPNe5IvIp05AiK8qM7KMhQodUoJEX2JYdmQ0oSMH37
e/EERNBkb+HeUy9+tbx7J2bzl9rHQNGasuUkJZETg5614MxbVfJ3LJ8NyiMKEK3NbaPuPtzHOPp/
uJYlNGgB6cFmpQfcA+hcGRcTJCyeJUCAfxeOd036DLCDJgO7T0+VDXpccCkxvT2gdO3JufpmHtjX
0IroFJW+3Y/lNMMPaX2B0lXX+cjnFrR0XYtpWrGAzuHrt62NYm3zeVylT3wqUxX8zqhBptWFQX46
p27oJiR6UIsyPq0o+6+O/2hx73GwEkhZHZXKNjBSnJK7goxaPm2zE8hL9K9BiKpIXGj/I62+ZI9j
hHEDp9x5EjEp22jFSTYQdmXBjnZB35gy2lnIuf//WuHn/nWJhVLUH+5oFOEBuFTmp4JqhIseRkNH
WCgmDZHWsfB213fTFumNMT/JfsoIpfDt+OEkw0GnN1Gv6Bn//uSiMau1Z5WlpsjTEYv0C/5NbRsR
MKiiVS2RRFMH5yU3OO33yBnAFK6S6433LoV/R2yQ5hE57ptXwV++m6AqJIXwLSsk2DiAaU4Txr8G
cNjEDEXPJsmOtDssGEVD9xq3Lmk4q5jgj6KN7xTSXKeAR4npb32oWScqmfHW2t5ubwOyu+iuwVRQ
01SfEA0KgjtMXj6X2wb/uQPtf5ojvQRNwfb10SrFf5H1a90cRWxLZMbKHdccgRh14t3Tv3i8uhKn
NhK/UtRFBgqDH5nNLATL8MGp+x5HI1iIhfVfJT8Hk2k45xzZnHfPQX/LZYPfvH6HtgZdvrJF+09k
LG+++4jRIX6WBj7JvCp9ioVGLFM2L4AjpH8exklIgceFpL9wC7iEvCwHDbuRq6Ykk8vL9HrI/W+I
+MApWiyxvdmmrPhyxt0h8Nt1XR/W/scOOJ43ZM8mH99EAm3s04NBi9Kd84OUeNXWbCTIfHOuqpmH
0sdBC6Re5m34m2FRQ2tMtXg+j6ZUjUinx2Lj6nvG4vXuGw8sLmb++5ryidJAgr+Rq7GXnvxRzwkA
Me/4NpWrnKO+DdArddLJZoZ31+pEyv1+BzIA0XTHgtHeT/FnLW3iejEQUuM/9vZJe5i2DHubkey/
o7fg0JBilHU6C3l7f7+XqRzEADpSkAzbJyueVTM9vaENaUKQUPuH/m0YWt5aAncwkHzPP/xHriQf
d/+qzgCwlYTYQ6/r5WqwVgrvukxuonxqZ9AcGKopOkjuwhZgMGl8GdMZfO8wBP9jFDYgiQ4Fv4lv
xlueuyL845+nFAbyWy+QsdMPzsczfL4hzmNFNTWqVUdSMmxet0yqhaBnAQXYTIzRhqpCpjrjnu5v
Z0vU6e+8xAFd00cLYNJaGYApBsGymyBak91HllMbvcPgWSs6SmhLjUrc4qzt8ZTyFz1GxvIlpVm/
4d9+48DAQyDxix6iSqNIpM/TKv/+iS8VA7gl6gWtTH3cTnUvarW0dGcX8iRC8SU73dKK02w65Ugz
f1YJJCyxrtFb0ZXJZvCeHX4JATHHpx46yRK8oHi0X3eGzQosrqo8G8f/95Q1iPBlB4PnLPVwQ7EA
5Wc8Qo+G8AzTpL7o8O16S6s7dwpisBvpg4Y9cFCYvDToRM6ztYLbOF1yLHvsU0JgZlHGfyyCYDiW
ouNyl9AljiwSPR84SKHIeQGXsfLQK5CBKDQ7z66mhAYlsgJkxbVZv7vQqlfJkN/XnQzUynPXfGhE
K5Q9Ka2iThYrTTJu4mNi41RE9Ks79tEz5TmvC6M1hquJ7Nc4eLFwQOSSf91Mjk4hncDbdKi7zclS
EP6AJXNft5qyUWj3LRz1FSCLSrRUieQd3jsrGJ8xRm2nyv8vGZKXXArLCXfd98JHcj57oOutzXER
382yElqWzZe0ADVpcAzpy2JtFfi8iqycG9yrJWr5edoz52Fbqh19+dee4T40pjIffqcsfKyMI158
vyfC02ewKI8EZK/Uy7dPUUdMAuHV6QKz+JpjB/3OcUkidPoGy7RBC99o44f33/+EGd3RdCbeoV3C
5d7KgDdOzWd+qFDu4fPycDJu9JM+D38v0UonsCA1hz7MY4bkXhzNA1J/bloXawKjG9TPSuHsMD+a
nOEr0XTDnOJWHUwei5bMgiUSBkRyisnNduRJ4UTKJmGImRyunxXR7y/U94/jjRFO6F+fNivKUdvx
ZGtaSCdJ5vIlRrtk7sNahGkQteaHS6XcPlQ8XBPLHUAIuJoSU2hp4QHl6FAoFEXvvxkEvDdT/FlV
xyT+m/QSutVPJd0n2thKe5CWnn8Ggyohs9VMDnxpB+aCvm09NF8S+5g9abMbPVAMlIfZjFCTPEmF
Z67YTChLcvx8l2BftwPrUDFs2RRVeARRJepbEURAHiPHnWrbL6dmeQ4pR0256WamGUZ1EzZN5fgs
wc5MmKkoR3AHQ7uOCW1SEzJVnRxrfaeCea3wXxc/fq21czUMLlDTg0VloJGlUjMtL4OqL/ps4d7G
U+Lpgf0PNv3W1CV3Ey+jAnWhE6vlK12n9RSfWL2+JlbXxZHlnoFXdTCX+SG2kdYDAsVajpsj3y12
fwN612peOYFgl8TT9iBgd+8xbRSNRKHDRbc8/C5XbwPn8v4z+i1qEvyyB71+Ks8GlIJUGSqxpuEh
3ktVbTJEGwuU3n8M6Ak5spK65pQj1cD85K+B1HimjrRq3Y2T2+FXHssaMyVyEn3IrxiITpYNMGnA
nmKKpGmvTWxPj8DCuvRFR38YcBLx8XEwGLnNnMXHmrbVbbNfKnpe7QWleNqxHs1Tnwsp6GxQbOBR
1LERgIpaujwkt45c8nbxuAmBw+btVNLLtgi0cjhHrl//QwG2yT199Kbca+2VErOCGfHXjOt0PWpb
PgnbzBOMvbbIbMXPqlhu6x+46mKh30wa7nzmbwBM4m3dlo0qLUwZ7fKrQyKtgiI+m6Ppq1J9cTCo
mjp3rMT8GsXKj3WOBH5tB2Vtmy72CMD1R6Kfo59OHLlEw3ffO3yASr4YuCU0LZWJatBN8O4wtN2f
zBuXbwpGraOYBeJ8pBPv2F6DXpM0tnigzErs5X+fc5TR6cA1K03KQFTADlIS3Locg8WmDVlPGZh9
m9o8o4AzYby86D3X8UspevfxGJoBFISI001XG4+Zd5oGFYweSaQm1H+6+qwtnUGjeoGAPZibDlVO
jtbHZyrfbWTapag4Kp+7T0u0Xz8bfQcmTU4PzPzuaWVo7YxN8zFdvLe9Hw4Bi1aOZN4Jvx5FYYM3
x2XgMBSq1Z2FrI2mWAFED3Zqe3uVBkbV8282JShN2rP6D4f3Wknp/uGvRT2EYFTSxclBg53MQUkt
nGDUQWu+s3cbpNg+k93q5HGGw4JPkFoWPbM/DQtq5BFha9mdm3c1A8dTFyks9DTgl1XVp12F+9d6
QQMZlxyP8a77H+HzINS4W4ZMMUyNbMJh+l55eo+5GWTSAfC/taWeEzCLLeL/YYwgLLJQ9bAVWQXo
/6xxCZ5zDqeXPIlXy5idiAg82q1Ja02YkrR7BCacuFVVUY8IQ+aQoKQYMRTm/RbrEwAdGjIqSHii
2LLqIckThi9LygzrQ2OvqDmZ24WK1sPAy3fXtlVZEvb07ttx6hJRPo0ml07D8RLlvvbovTjSsp1x
9gQE/yGtKnIGuXbMQUJZzepVUt+jhQBZVozc2CGPDxpv/CR3kBs/Kg2qIctQCGUWasaO8Q/tdtfH
MNXysqPWF9661nYSMQfI7euWl4rtHZ3lAUPEoCGMeGnvXX56gHkiiQU7xpPA4VgR2iG38ECePt86
DRUcqf8pYnYViWYkh7TdkSI+lRnx5YEoRH56nZ6c3vmjH2IONR5NoxhfG8KYdDAT77TmY9qNKfD+
rOlXVyTFmxPPlMN2mR1n3zQzqmPPGf0xMOpy5AOaCKNCco3TCFiYGRkRDgPyunU5AWt0OVA0C7at
mSW8NRmDzS/aqbw+8i+tAjRWLbiN4DQcDFHMdyegRWuhkK0fpCqfkm6nNQJJ6SqPmrH7nRo+B7+Z
/6aL9nT68YoF+MEk/buyb8QDDUS+er1hYsJQlwswgwqBowiJ3oi7J7b7nqaIR6sjD95hRthqe8R8
i6ECahT4YhkcCIfTFVQZcMB8BkHL5OS8BMddFpzKeLd9kx/ThI/NIxUIuH8qBgS3/J0vIUl4CCng
SwrS7SEPM/2VkTonm3S5xe46Kt2YpO5B18I4CsbXgkaO4cery4iyxris2hVfEglvwwZKbeQF1e6L
UI/5K2pnkY31wp+I6C0A6TyJ+1Q2h7iX4SqAMTqE9bkx3EzLqMNQmFf26eQJDHkKcL8vbV+Qz4y5
HwZoNyP/0jblOHYQxymJ1zceSxTRiSqZjshn5hIfJQSQfn7kuwKvN0Jjuj63YzYJ2apRJLs+VSIC
d1oicJnxD0c9TRshOeyMSQQxNyLU7aMKT3uvk9c0Kb0F8CZE1Ni/sykCMC2E6xY1VVo8ENn3Ps0O
xE6zSfp777bNjnxMJE7Y9bF+bOCnqUDKUHomBbb11OEFuzZ2VlaG+Ob+F1KU3NFc+eQD4+HRMxg6
UbKum2a5XmusoM4ifQo8mvYo7dQEWpS3nvYzd+r0/lbVNEFilamvJOmkbHUUdE0/UTlBmND16YXE
vtKH9MFLflkF8h7sB+shx1IxtUjH8C01GKN/ZFScPZ2edL35LcveOHCqB0aDQmhDGIlnsrVGDEGl
g2ZivWxBmNSE+U6gBzmCNPRwe//vTOba9OryKZFUw3xkpO/3zPn3FyzHJJ+RVm6+GJr5W3lhT6sG
8Vz6bnArjB7XJPSOaP7GTr/rDm8h7xxqvaJwWz0YAF9P0DWKDhEiTXJhP0gcvaCNQTVadPg7d9OG
XRR0uKWKO3eqay8gDeKaJrIHQnMJYhikjV+I5KWXERUNU47V/oL00CpHIJKxSH9tsqmwY0QJqEg6
9rzWKd46W5L7xu8Lu75Hnrvs5J1A4nxGCRiQxzQHEnZBLp3Zj3hq/PpfphA31SsO6RHzc3euE7fz
4XCbVtCMlAOKQvwM1IA07kqBLVQktE+gvfcs+i/tGVcTwB8Cb3N782ncBmM+pAQNUYQADgncTyN8
QmuJT9IhGdsjvrl61BwS+S2b4o8/xy26c9Bk1Ps7dnepevCKj2b0MbKsprdbdUKU27mqHJcHhn49
Bnycfwv/wSgM0KmQSsz8MwL4V7Vx3K91ZN69YRbrtMqcKOmKYihMc6dRxtLF//0C+TOKfB41rR39
4WNqvq3fnCIbmFmFUfXu0OETs++qc6HCtHspEKg1cOwFlIB3ldF7lvZXvCe15zOVm//280qUTu8v
6DNlSl/3wsTCLGJOARpxskkO2pzSLtQZmBUPvs/kSorRWfwmIxmgx9xHm3CP5i9JuEhTkGULR0o6
QiMGDnpAk3LZ6fIu/i10Ry654WqHRpk+x/wYW+TQ1lqduNSi342pjcDVYbTNuvoQGG/wHAuaFJq9
urEwu86GcGiuqCn75gxGy8X10C1Re+/hnMiLyv1hIT4JjKkPlWWWry7tUuNjJsQU1oAEwgB13wtw
Z4D1bYAXL88ZVorcuzRegJKkF/ZggBe1ZkQ0cV4/f5uwTODS9vXUYQtzIhoujD6PbtlIswbBYqoE
5isFEvwC8qjtuvhVmKzz0seRCEYqJPXqW17pD/gVTrQb5N7OZknOoexddPvvuAtCOHYeYW72Agxm
J3Cy834VgCXfe40HQfo9VmALX1oHBe09zYkLdF7YWr2tdzjYcx/EW+Z28ejWIhQgIbz2beS8IJYc
+d+F0mMlq4hXr0szmW1po6rbVwaEH3E88HUmDaz9W65oX8t06NLQxTMiPrCol30NUB6UyWTHhREc
JgwWz7MDiR+XqC139ed3Z15tTPy/+uGbmKbdHgls59AcD48mqMKIP89MCdP82k2aQew5WMjQVRqo
97F56f6yua/7Bag4IlrzRmqj2WSJfv0ghLDnME+ecK5OTwpOc5yiBL0F0pGh565196eCG2r8vDoK
/pjyjjRS3LpFzViYihWZgnfDudub7ZNOwcV4D23MO5TtOyGpxrMV91bRER0h7Ho0xokGZo4AqmqW
8CiuliE7kuGORD+Swg7eLlpSyBJ4R3UZ5wvMTgsi40rMA2YQfNoQPrQx3IWACREdLGPcyQ7GVNy+
H9nrFam0EjlJDDcB8nMfJZ6Ty43EVvcM1A/J+i2Im+jo3Zf/KQst2Jj8YDYFI0GmgUijgEZcMKWr
dA5NNX2eQqSt3GMkaccFpk4k88EkBOTDKVOeix02OQGuwazHaEnejJ44GZffn/c3oj896rWUjL83
AzbFvo/lvkxjk4UjNosbAEgW0YdEZUIFUFKKfITsbWrIqAmI1UYWdXp7SgkqElpwz46UQmrlnrzc
0LGIZQnKP1GsdEW2u9RjlW4a7I3ZRrOI6SI6utOel0CyghlbHR9tehdvTF+9bRmyHPHVDV7u2K8P
faslKnrQ3vCLPLRbmSEZYhCu0KzjPLih+bg6VIAb5SolqseU1qnJdCxTFpsN3oqc1/xR6uYtsSG9
f3xo79PaImxvLShcFMYslaikdg2yfuNxwUNSWykhS+JlHGLtnSL9842tG0uCRZ8E6V5SYq0ubulp
D8Z7SSTR8QznQQfMb2KqqHMl9Vo2mX/Fgb2j6OBy95y28n9zq6GppVE75pVmsdOUevrkBtR452E9
wXL0z+c8SOvOB2cI5aMkiI533x1pXgG/3jOt9E2evbHGU8N/Uc6kMbFPVo3DfhQHjXL9ux0s0Emy
TIR2bosrSYJMqSjmogwg4j1ZxsVAcm+xseIvrlcyQ0uIxgLh9/EPeS9NrrPsd3+P8ee4vT09PHzy
QHr/V6qmbIjb6yjLoT+ShmlOF9+U+VtZmE3yhnGbfkbCd0RlfKgVWXMCeQdkmbjpuAcCpgYHiVzE
enIvwgMRc8cu4kjvHiLT/1ejgOw3huhi2xv8/vIEhqAgEgtkIcqOHhn+45TXcB3aF+miv9YdiUOR
aSTRl1QTR5BF24EToxrh9zwjXMxUfgNI+On3DS7qyRDwYst3py4NRW7SXXYqqD1oc1WcfpCu/Shn
yk+vUE0ML5EAvy19KMQ51WHfz2pRSiWxpurL2/qorvtaJ3J3YeQIYPK4enRY/G0FvexnpYjfTb+n
7KtAnofcl0YX9ms33z/M+LjsAQTBkc7OiFJImsnfoiy0R+JTWG3FAcsmo6hk9oGOaB+IMuk676hk
gQiupErP0StG+HYhquwIkxqZSUXpK4K/aIwCKrdPSn5HT0439Rzl8wMjq28/NgHJammd3FnBdNz7
aQCg6oM9MhScjDbc3cNjMXrlw1biOuyvEchrgedH8u3W8Wl6ibiTTMUwUIrkvWcWnFS2ePyfPbyv
V4SZYfOPe57w3hdpovqd4nyXDen9eHaKPArylB2XGVhna8rHU9jYyCUXGtKdtwceMsCWRloEy95I
GOppdMuKPLbLo/VDbIgnkb497m4ZC2vhHJpNJav/Hw/UlGa7MNQzIrZtVdoAXRHa9RJXQwJXrsSD
TW24YW4d5Kjk+gkNdRBJ75I92Cn9wl85KqshBWJLl4zm3+hSVrB2/6jQLDD9A6bRefgE5NS+JwFP
d2hNfvccyqLOu/PsP/z8YFs9yDD4aUA+EOnz99+pO4AFglxhGIXtEy5/PZ8I+sjdckgYwsJQsmj7
oFHyG6mWiTgIDVUYKM0ZIm3YoYYsWu09yjeDr465KvWtIA6AqMcDR2V1OEQIjbHeBQhnogDK8pBe
0wGXE3XfcN11SfF5AxR4oW6ydC/J14qr3IG0aEieT7hR4aaFoOcYGtkf+Hvr/yHKRG85DOnbNvA4
o1WYCLEn7QRO5/eg31SdGQ3MO19L3OF/X4MNsmbky+zyxBP4Rouvfc+sJ4M01VPLd2livp7WvDUl
s4HS0vWMq0kgCYLB+j0s7HBAiUGPGZy9UJIvvQW81QtinNrrVvuChVJGokUyaASAeaCmRN2UsOhz
qJSLBWh7D0yTSir2mq4u4YdUT9KAik8KCHbgA+aHEok1HJA23ES0s+02NSf+DmGbbFlsXAsZT9cn
F7X1+4gUUN2Jyyk2j6mBbN2TbDpktAR5N45krQos13aGGYhhaFWNJpfKytqMJObG7MBzXc60A5JF
OHRDGDB4/YviMEMphSAvPTRgCGv+AYPe9j/pTKBpqCYoQmjgmF9jJj4q6sm6Nj6i9Aob88nqQSOj
74x9qJwUqNBERwTLMKTb8l3WsSj/E5dgA73YLRPawusSQpLmBoBtjKwd9BA1IUAooSkYGOgmNTn1
pyoM+7HAPGzSM5lf9bZVq6ytjdKmM+xsn764UyXEkLGFZp5xxZjwJVDeohcCdwf7f1MI/qUgFLpz
smQ+QwXdG9bKMpUqsRq8gJj7uZLTbcbGIIrT5M0cPG/BZ6WdJ5CryNNnW+w6k5rKVIFwX/EzR12I
KUZKQ2vdajMiB0++jKTJ/6R1BfWjTPyB51vv2GC16QVuI6V1+OcLqCtWjOVTW1FzYpx7B5ypn1IJ
+V16Jf6aOyz+iz3LzBKPxLKuVR+uI1dt8+DZmpAULfchnQRYvni3ZLoVYx2F9hHIppFNmzhN9VNS
MDFrgLhzjg+pFWPItUuFzR86qskFBfmYwH+7uOcXooAHo4vyAjiHMkIzKxsoWvmy8t31QeC76MV8
kYj6pPETTRY9y9khRePIQmmiUEWSOAKEuByG76VUYlWDomgByFnvzlbX8M8BE3oNf0jxrU38nQrn
t9YGtPFR9BN7w8lTWd9GyEv3LJZUrqtRGdvoUPLQWhUpsLOcGmNsK5pjMHcKOnR3dHgeijKT8qHV
p6g/RfA3SLRx+unPJPj24w9OhOZP7gA+cShRv9qYbCGR+fBA1ElDTtbgSxhmDXxJwckjYETCxwCy
2pZOugFFw4fmGN36X8wSzcroIu7S4Pwe0+vizaYvZCOfdygPR/RqPJIpHmvaxjxdqxYBsF5ogCDq
H7mSZd1AQbw6FPa5QimtVmTam6/Rvs6xSHiRdZYhbYAn9cXk/xmOuVNrVZoLAEgKH1NyDsHw3zMJ
Tfdbk1IMSYy5fK/OkhjWRfbtbX28uDglOgf74fYEmGirTmCoPA79SBT5wCJCRchBRMaBR9ebSjOz
zWLy4IikH0QzGszL7lYEz7SwYgkubbxpTCc0dnF18JHQKDgshk6ZR5gLqreT7aAAjIt3hhRKYyPF
vsW4+AZoHpTedrBiyYTllcVaGxEtp0h4YSr1O2vzg2zCEtiaivV6VDZxS2ihQyYk1Aww8FxyYkvg
rsW6heRRLZ6f6K918MbTMgsI2uFfdVLmyB6aJCzSAhLkO7M+oP1levWfi8LhZcVlnpM9x/cCnlle
PF8pi5EYsQGOFpYG7eI41zPtJk4zz9e00oh5nBG8vLa2oye2+Cupe/E9vSbKvJ7z6XVOarZ+TIhW
6nR9KrIR08SCAyt0yVKERbWyJQHiRg2CKqiQgCAc8Fz63HAUHousZSqBSsAeMOVPcuP1jJfzDxJG
kAfQn6pAnmv71CDKiTjmktBoH/3z6BctltNb1BQW/zl5zR+tVHAndaDNOM+/u/RRn6ba7dyRjajZ
qXqjT9EUQ7CrB+eMqdFy6UDlNCaqkQLKwI47xh9BcKLVyoQHRK3u8C0Hy4hSKaRppv2ROWHBMo4Z
ORGq8syKRP9SWrw4ORZyTLSDMqNUWoUtHpgWh8JpkD0ud99AK+Ojv2pypYoRgqC437BpUeTTMy8b
iQ2VD+fUYR951iYu9wFX5V81YLONgyDrXXEebq6k4hLnYYKQ/53yE/INNtuJp7Hk1NaPiJLBTTNk
33VIh/7BtngnW55HHIE3gXUnLju2iu05cmYuf7rWZkAJG/mATnDY/MwTY1B/XoLopQNWJg6BHyPL
DIsH4W00mlOPmk8BgNEF+xluc503EodAK5XWFalSWENJk/JatRmLxi+spHVvnYWZfgcL6iCDNH0d
ZWqGdnZ0V0RWLtmCFMzfaU5NKji44M+HpZy9jzxanJoKA3/Y4mquQAtfrcXCbbbqnMZuDh3DCqbV
7i9dkHfpWapg+b4kAQxf7fecoasR01jffpZf0NHE0vwf0lsYrZDJIbtdqwVTJkmD4J/VbwH1MaUs
NuglWpDi/3UwcqvdnNBwVH0P9s+ygrXUzH66NOPEBIYK8e9oktDNrbqZK3aEKar/fuKF9HSSfi4z
5NZWTFIzXUMr4OgeCLC2pY+hldJSZ7fHNhrPrahcrkhwbLUdVNKxdpa2ZeLGf/NSLaxKNNUQ7nKy
o1FzOCJEgeSwG2Y42rnNupK7s8d7JIsZbVwxr6WlQiFn4OKFXyPf9RMk3JNVSD3ODaSYCpz765TO
KIi4RmUDPdJwbS9t07lI7K7a64YaDaEwZwWR89IYaWat4kbcTt8tzfsXL+kRFwEB6vKvisJKoN9K
1HwK0THQeYDh74swDvafFHNP+xakjXR6PR9ylWLzf+aA0bFp5cDM4YrigTtd+NLiHsTQXiJeaUm6
ON/0HDCocOSqiJLV8/EUI+U9XPF/HLM8ggsR2NXA19xlsRcBsxxUOOsLBiS6l96sf9qXmuC5UmRV
JCz0Q+CWrz7AlsLaetu2LpMMoxVNgDa+aYvOq0A2zGGL7QrGrVOhgOig3s+yuZf3ND4b1lQrwOjp
z1R4qY+AxikPC4VOR1GKcJGI2KL+uCL4/a9Ppul5McQMMUs9Luv7GlFuEHfVfh9M1e9U3Gw9rPct
dgtFIOQxwSvwNGg04+sNWAm+bVHGxNtyS7MfC9TAGPxAe/z2/lN+svFr2VYqBpZ3q8E0kBUsVXj3
D/coZxL0/IzdMGM7vwlzJCqFAJ2WIxcK6OlhLx2Nw1qAddkat2X7ymBd57uo6tXIH0KWtVtQ+5js
IaOmHVDDm1vx4N3+QIYrnZcAWGmEROpGTmvWvaS4MR9fbocokX0demW0tsaXNuMgXyGiXp2JY62a
Xa8FDyXAdt40ZP5h6vOh5j7f6tDmK3yyNb5l/PLKkEthLtbUXuPZdIc9oaN/0Vx/zOk/G/Uw74vW
RaqTM5XzhzXQyzYIxXFR181efR7F2o23+lsSUlyTdtkuyMy+tM5SF79sRfcLF82DmLIADSS8/DbT
c7E0u6rEVp4MVGnZSe6ml0+cq59I03izD7Am369k1t1mSqwCIEa1Zvejrnww9O9SunkYSPN9+sov
HiV9zPRB+1Gac8MXJYMWaYp5QfbkrKh3jqY6UbiBXpSdBYiXnzX14dnssHQlV0mLmaq56UeJAjM+
Jkh0Soob9q6rUyvSjnybSsbtkmKOV2e0A8ZmjoHY/UX27vujf8kd7RzDN7kUCFUuNm/8yNjVHAdN
3gy+bKaRXrR+ObyWtHUsMj+yLrEmMPoISCh67Q2jBhn+OQN3QYdpvz9EodJOzSQjjCVRQK83+olW
0V9/aQFjCLu3tzS9c9C5SL6KLXIW6CMC3Px11Q6LNB0bVjp+E98f+wbgUF38nKMdkq3SOOT6SvvM
U5PCa5sDmGWuyOIPKyjHidCMZgASvmFcJH/3LOh0yioxOEgfB51BBBqEGYm94JuZSvIu5XuLiheh
KDBJVIYwggN17GzleimQN7oIYMb+GbPsdI9LiKP5S7g5KoXyzD0CfDi5BYYehDVHgpj7JL3YhK+2
+fMTl7nMNGLQU/c0RBk+YxTRpcxyPB0iWQnJC9TRWnpWcXaFRHQ/6XUZMXSZ6NKlYLSXFQJl8Fie
1eKC68h+V6pe7Ji6rYx7x8BlPdyL+sAkJKnRw0Z9/uws8vkeBs1PZNjBlNWb0FzdsaxBkM5NEyLY
NPdPd/bQ3IArQQtmvFi7dlV56vQM1WpZluiNLH9Ei1Mj5sJBjA+L4l1//b4FYvRqMMKJMEzX54WX
pD/sR5ssKiNgY+7tA7WxyCH2bffnXOi8xqhTwQszS3XTberUnQn11xcOMFCcwZzuqrMvYlw=
`protect end_protected
