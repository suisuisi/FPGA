`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S6shR9DFCbbp1SGmCV87Y1mttswx7ceDhlI0d4p31pfTichOkL14ZRY8LFZLKaQeZ/MboFd1A+aw
X2cwAoHXjw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AfRvJF5cduDMP8kZa4+MW/uvbbUQNKd7hSGvyhQUlFug9FoHKThRHJD6+F9EMM4WYz7R6MJOC1Uv
t6Lvxfat6BvsVo3AQKtUi5HzUXJRXfn71mePuoqz0YdGmikolY9R7uT7heOAN/IOVcXxm0DS2p/G
Pppuuhq4lcChmTXH5bg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IhTaYemNEBY0SIg1gE6YHwimoDa0Fh44zETaYs/Iuvk1tQk47WX4j2X0LelhhiiZZJv9qhFA0XIN
K5N4QtdKZJ0BKEgldXZ58oxjuu7x8WPwzXZ3jEJDnws7zKnSxZbqz8+piYRJ9hYH3cLRrfYhnyWT
9eFAOCxXhStX03bGOhcrcdeQwoRhiSx0vcuaAbBmMXqAiqfxi8P+TmsuAFRNA7sslRFfRQi62T57
dJ0gOOcwciDkjAbpM4A3Q2H6depRkauAEKLJ0dq8ecLh43ImrVSycYVsPubFdERxmq5zMWtUsZd6
JZ6Z5oJF6+EAlCNps4gTJdQc8NyaZ8pPnavpvg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QFydrhpU0g4XMLr5UpljuH7JNVcbvuW1ASbLIjTFdIRtV9gn9zXVjUpSFRx/PWM7cWpV6N2iUhnk
w5zXgs/t+b1plEjottTw9mffwe/65e8PcWCaSsMvps+8/oSFYHfMUrtQiNuXeaRle410mR5deNgq
RHnXXTi8+WYougJAAnBjavUZZu/hu6/r3h534E7OHiKxin2JRvblHVbds2J0gu+Ui4MKelgq8eiu
D9DoEi3HF87cWevYLDXozLFhg+m1CRQLM3pLvtFT9s6nM0rA84TTaDh+3mbdh16k5sKyHelc364e
7RS5vL+qSVSate9zbA+w9CMPBFYZpBzCBr5XTw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dRE+p2EvNpO+WTmcQifWazc4jBomu72qXp59zbjKJjUwEKRP60N1OOp99t/TCe4rAooY6t61K3v/
Oe6qbWKFdyE0YVHWqWtzEFVeomjjfUex5BB9711QlRPnHbTZbrMDMxBJGssFCrYNbrfveabGOcZa
bcdm3V3ALon7exIvUjZN2Cs4sqs+FJ87zUHFbKnwGJkjrOQL2IDDSMO0l58wo/+V8yxCXNNjGYiJ
NTbZUs6X/mNPq8Pr+bG7k2jppt5eiq8Z4maSjBlnpRQmybQimcZg5HgtmSu3SXHBRCTEKpb47iVC
p+FbVqFuOGXT9FVFp2WUd3b1nm+W1eYKz/8m2A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uh+h/anHX/PoPY1TPwW3dfPqSVMMQxsE5oER1bXTzsHIAZV5Bn0JI+gTLW0hSTm7S9QE6+k63ZvK
NGJLNQ2S7Agpqiir7lyeWU1dO1SoOtriMEyl+L74sBUAcWoEHDGB8NRDYn4vmKT3GluPisd+2+wd
TaW6szJZOKn4dYkNO3U=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UkvBIedEbmQJaKsByEar9/GuhQhOtUb2zN2RvLkN4DNW2ZRDkxgb7XlUejcQb23EY75q1QyfWRLe
8UE7yBNo2/h9C7E6HPktM6g07JetMlyj5jFA5ShQtZQKGEJMLDqryi8VkyfuvePC9oQh5PZZui/N
z2zpyUQ1GYGijD5N7xl+R/EXR5fF190HzK+kB8qhKll/z7jcqABBqKEWcdL6tjQ/YRUp1hHZcbxU
kc/THHqKh1hEWiV3m1mWMOo2EMlyIJOEs36vj7lto9+sKaVZbneSZKMyz2EbiPnMsjXTbeydMtuu
2zEmg3ND9Lv5qo/LQDRxta2TucbmS3PqFP8tfw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175296)
`protect data_block
rYFCbWlrML5dA6inoAg1W4uwK1j5iK0NrgO2ZAIUiWNSYmZDllDYnxcGEKfcffwl+bsiFS8BkK0W
vq7juW+7QJ6quHEg/VL/kXLnLsMpYD0dMoKZL8xXY1GDcFnLt0DpjHgk45Qxj2BlOIshmUuyd9Va
9ikMsU94rXvviPi0YUAIgCOPfSOyH1hhLyTB96e47memKzSbLLT5LOH9TEjIT3p4vSOqcYURtjvb
UVdjx2Wp/UAdNp/zgfWgn3/Pl0fEslJyczGSWezQhfu6ZtEeJ9+xKbU7v2dtjD38af5CgFfIcLHv
EtfR7Eo+mScdD/vHzSZU5HsuiUekvMEQHB/12T2Nsjnz+l1813H2cLl0EoQW9lR2lSq2hGav3yBw
/1JdeVbGFHM1CZCZegdmtbRs+UI8sDlKGk0snRei2XQmT2Tm4t2yeW6yqMYc03JskJjl47gWwMRw
wvYwEYH+OQL0yi2DiBT98muIDME/ix2FlUSFb2uKmt5U9kP2eXoBZjrnMQQKub9547vIxyAQS2wr
tBCe+wDFjZJot+qCacdsMJhc68jCzOCZT5ypE4MbgBB37FTdCw3kSDMOvvChJXJa13dyr5atj2/U
CvNhLSMQQeD+j/haKOqKjtPwqebOOyBdJPNNvBGez/kNhTImgYZDQQRxj4GNMTN1FJVdMF18pzgD
qQq/XCziXoJzaTxzSR/3EFKFRFeuWpg0n9n1wNSOOYFf9gn+HlrNmknUGyW1/AoHXWqqOkZAzNDX
hxg4voEvuVxmFKC1aC3BQZxSZ6n/lg8YSe7ODgSvQu1sTu/pjt/worioAlJDgeW5dnAo5R2DG8Rn
gHAiqxd5m5cIA+JKsLOJEb/Pnke/QjASXLpuiIXrLWlyzAircJr+rPkDG/TXHxXfSGg1xIsN3bWq
nqBRFzZn7k4LK/zCu4+LhbauWOivLBv8todKSerCfh7vpvMYaCGfTYSeBsFLHPm3ivvvAAHHnFPc
d4GhTh5Blzb4DvPkGmEfq8xWXlfFXB4FpXDLA0al430WGK+2eXc7/glq84t8TB3EVRwdFAap2dVe
l+x0tdisiDHXyZV4CfAt3iyC1Ngf2F+81ccu/c9Wm+vQPCOaruLLEW5tKpwV97OLpXVImPD1HkwZ
L6y1nrKhRVYraXOWVUAOVUrt8/P4fKe5GMIV02gSpSn+YLPevvkiCqcQ41GDDqbaQRTu62CvpBoi
ewt5FZqVGBKNVmC6faPttZigNF6y0m/dSRoswAn5OK7IG+0Fa+3IGuMdXzsu8Tgo/vl3SRQyIQwz
hnVatm604SQ/9oy5XkcKqkA2bfbg/gQPMmwSb70dw+qbVejkvUxL+ZTHsAi6vxVKTzwmQSW3pcHj
mxuOJjrFhVJv0PdgylD3sYw5zNqSMKCwMW2uRjyNSN7gS7xbtxE16Gtj5oeE4xjXHE6DBPG65jN6
2ziwVmd0S/YAYrgXBU1nhjYXufqf+e45AM8rTP0LE8iO0HMC7b/ayRZCTPvnGPin3Tal6MKEeUbK
tMTHoBmo4cbOo+dgAnZoaOuVj+mWosabaQ3+rce/QqaQdduDJJvmm7hWqLY5gqogyeOJsMgVa4Ht
IDFZPoN2rpC72dXQclXR9SAF7OPUFpeS2vNiAJ+uHq4v6OiJl0hukpYdp9p5Bb+oX//9MbryA14l
n0qH0Npnx9WIPvKfgx9iVPEF9OZSVStDsKNp6P6UKPsyMZ3pkxbvgUCpwANjmFXvEuAnekW65Q0e
RJkmF+GMAxI7Sh43SAlWOoFHnhpE/nKIQojZnytMAYnmQ8ZqsjIoQQAgsMeH8Pcu3ByFJhnECm3n
SXsOxmxCG/XHvzoM/fgOtvhEdJM+4JxmHxzB1J1KmUPOWhM9jzNLqCVTT83AE9GiBv9tYvFWqCM8
Hfwy+RuEsx+HtkLlHCF0fuDFf8O8Eys/c04sGUGw+q53uEzxpaHRyppK8pBaDO3A1Ht0GuuTt5NW
fYu0c727Tk7XCWQUhsPeOGNebVHIKlM+WD074QkTfXmmzclwoFjiNb7iqC8JXMPHA7gbUvBcfLEE
c7eSarbmuP6488B1aZTQXXHgCOyhQwaOO08asC6Cosb2GkmGjwpilVog+2CIHCRNYTaK9WH/22lA
srAiz3HOMcj87P7KpHIRjcFdJKUYOoN4nGQVyiibrQnz4XtL6W1/+L4Ke+0XfggSKKn+gtn7UGrg
odtIh8biU2y8SJEUvdjI6h17x29qgeZ013x3R2nXWtLnn8O+MDoYPVoLKiqVM0/PkQPB13djgmwN
H1xXU+FvEIUBNqOTJlWpg7wHdckwsZEByGqWMFBd48joVZw3HVtJYtOr/ZJE3dfN0NOtUzxV7ipG
TYZDrFwJLHZD0pflhoOrl6NQnNODQf+LbpIjrku2IOFGDzTTRz+AaVRncVZp/fFQZzjtwC8FKSGG
afC73/iXdd7o9ojuVC8WJxP0HSVmeNXHjQIyXHvIPy3y09iS2YtjHhxvBPH+FqwynDHEanGFp0j/
YhT0VgEZEaHMQ0VE0UxbGiPiq8JE1ssAe4pnD7oSOsrwgJULawsC/I0XXdFObCwwz116lpLv7SGW
9iWZRTOZhfo8SsPqQA2HnyWujrTZyELCh+nKL6Ot5/Y8nE1BfYZi0tu8exGAqee6mp0x+UvPBawb
H+XQGCIau0MDYJtWVclIsbF6M5AktS0lHS0Wr2t0CXmClp8+rKN0G4vF6CkRwmcS9mWc9dCVma1J
kKNCwGM67DeLTbWaXksa3RraSClGO+FvlhzHtic+sGJWZzosBGNY2jM3mnY7kvGWbPgYCQWTYsE+
MGvFbW2p6NL/sNvG4HN4BM+mF8NAk8bLjciALC/cF85Ls4yVN5thXJvZCbCadqgV3h+O24ZYyfKI
+MO/U5114F1FkUE5PKyS//J485XEpyB+JMTgVdwtSOqsq8UZzX7G8K3cQrdnQ76ow/DQuu+EFjDu
fPuCHUg4qlpdPVtEd++A4hu5KlN5BD2YbUzQHVw4cbF8Z1I2ppo6g34X+g1UToI/wjQzK57Pvbdh
gs3n63ZXX87lBGH9v4ngicSsa29r6SjF6fzUrq3K7KRSPL5M/8CBehWcMOTOrlYH6hbZu9pNiBJE
T52w+upyxcI3CJLxglvU/3adw9wbrQxRkfDPI5en4GgO7REx5ydJyDvxaZiQGejtFL1M+phPBht3
QIBAdIgccJh13iGBV4qrK8RgJnRWC6XDcz7jVZsl4ygOb+JKzSEV533/BbcQHMeWuUtl3barZDnD
CUwNoIrl2CGqHserw6gGdo/sl1+g1jCqQLYp3ZgtV/UgTRR/mkzHiyYujY0bdrPwQaFWUxu9gDAT
FJ94dYnlEvtd5OY1H2AsnLMLGE84IiNK064WNlcsxKULNoZRCMoe4OsKKVJfS+MgmNEFEu5e/+FK
zW6iS1zgH1ypI2DqRAYRKt2+zOtUpO498EDejfOVQxaJ5nPk+dnclPC2zPF46Xtsy489LzqxVPkL
ap4cMSEEcy0dIPoqvsTnQPjt+KzppqxCo2Wk+fjErg8h2a7ohrJQCqaD4O0nvbvk0UtJYpQMbdWZ
FaS8rL2l8eBC9t0VnPz1oqQN4kDwVxSd4f/CtfKf9BUYrxrdfzbyeG6Mm9welCgKgqPJYoo5fRRG
TgRq0yJmq1wcCwKnRR9UA3C1IsrnYd4d5Bmi3NxeqzC6vE+6JDqx6uVezGm/BsBYosNEt5YBDiJi
B6z3LdDZwPgdRhV07jKDPmtqdKYTVbgvI7skS5qXYHeyW//tvwY2gckrFfIYYFzknBUjy7u3hHng
2csQcPJnisMyL7zgRnoGV2fSfDgHFl0o8FEaK0f/7Ru62nhd/DCqUSfsaNdDzJuCH7kVr1XHt8qU
NEs0l7qv9EeE1Zpfkc7dP5/KCS8WEwQx7DqwdNCYI992CxrQI4UPZJ77oIizanQsRvw8J/uQGuFs
Hl39fq+/+sCO0XlDDcx2VzeB8LYvr65Hpt++PnL/jMeNTBES7n5owE3+9gfyeL01uNVa5gUrxbXZ
ffrTMWXaO3f71+n6xea9sA5pOaEXklhO35uP8zAAqN9X/9JOLJAPq+XTyV4nPTRWFMlNwTAeyjUu
zykfgJ66o28Ce1gGKNQTDjHIqyWLzeZrhBL3JdSO3o9gOIvrfIORYsZq8s7yRkPsoiJ58fyb7XHx
Oj6s365VJRSru3AQ+maEeMvtQKY+xy7LWKIxGw2NmFUj5hVOI9Kan3Z5mwbyW4P1S2wo7kRQh564
HGee1GkVNVYYSkVO1VerSzhgb8x1fSfQ07rPwh2+9AkF0MdGjqrr3QLqo7MmjyyxF0cLWOps8I7n
C/wxMooAGdoE69zTdEfUhS7cwOC1ld6JnqMpnJQ/WZmF1VvgXPGcDM5F59mqANBydhWcteyDWpqf
w70vCs4bWlJW5jozKnIcpnUGFDZqrKKjqPsnNWH5VWSJlqsuSNttuZiLJ8pyv7RwXdN+PNNWqJ27
NOIbsOffu2qQmPqnWEf7aVWlGOEAdJolY62NqRzFapE2A5cFyofGTzy5+jKXKKxU7U5HVxHuKFuu
I5AW+t+jfHToQUQMq0m8UkVhxrynET4TRT3gYpNd2uq6wfO8dzWg0Zm9QC5Ocg+kMpJFoOaZkGPP
BvQHYMAZE81HM195S5O2TYmXPs3bg+5viblZSHmUB9HweejUs3LlNOAUv1k8RW9NXxgLGV/xuP5A
gB8EQ0vm4bnOzurF9NZolE4oZxUx+kWNe9yi/frwtmXOrACy4lsyBcbuwvA9TA08aXwZF6mIKU36
k4oiB+c+92xmCdHx1KsP7VCGCKoRzHRohxw6R+uUuytrRCY262z8GkFHTa67jSIPl/Sp7fWXHsVl
H9YJuk4lKQoH5rBYukCeAzf9C2YG5Dzxjc7YeIJoQ9ozt11VrvYeaMasDdU4p4hsTHHAJDzLG9ln
vMrTfmLjKDgNBGC7OEFsT4AhZjTEGZ1lWIvxv9XhShQ4IT5F891O2XlIHXavXK94wmabAfsBlGIs
sgmjaJxtNTW+FcumUN2EyQQu4YQqdY3oXr1PZVH20X5Xag3Z8YvCCvDHwfJO/63NbPq3iPp5jETE
aWPC43f6RMXkSkv45/vBdf42VUbBduLwPFk4PVQ9dZFYOZHtHh10wFy+9xR61S6+y2AxVrMpiDPa
SDvr+Se/iiWnIyIoTnlFNNA81mGTUbXex35jr2kfKGtcm3H+rJkhzugdbjIDUrMI7Dw5kBapko3G
YYH7vLv+N6R9cWEQVCoaEEx24HRomgi4a4HVQeK6lQH3HCLpPMEDe/ujx/bP7b4xFg0bkiG/Bo4l
Ma8/WOTTBwv734mSCAvhgez+rbMOwg01scSH48kks4yPp5WlZEfSqDgdys1ay52e3Iu258xwy2Lw
JqZ9B2t5y7Q6PsTf60uPYH4r9IUXxHqtWH1mfQ3Hsl81Ij4T0oTgtb9ZvMNhUWT4+B+B35mnm8/Z
NJ/eHs9bclZ25pktu+WATrU5+7w/EhrF7cqPVMi3yld62mi6/O7DThBJ2Mykv6SEvNrBp6GPzmTI
TuWfxKvr4iPl/vUE1u6mgA5/RTHZq4os1NQ9211FxCyxNBGweCNNIASpZStQPvDJbZ8nGHW58qxz
z7OQhe/RpG9mvRAjFUvAKHN9f2Zwm1qbr0hM7HwbKqEFci2Lesb1QOP42NQmrJ8TZ3m7fDsPvcqW
OAqeEVZDS8MqRWY/dySXy1NuhpmFOoOALAbtjBGj6bN1D5Cw0ywjnTLm3LBFTQX7IvjEVvfz/C4X
nBr/ne7xrBgiiC83gmt/KLmom2pwnTI0SprF2SZYE0bYDxQGaKV9MuBArt9I4NOxc0WHhoV9c3kb
ZCOiDD5WR1DyIgq3MmOP2iBwiqfgPD5pOHSF5q1khwADn9BckjLR/+6HhWo1rfPzvEL/TkNDuepL
csJehECa6tEPa6o1emM5OGKa4zlX1c7PRNOal7luJP2j27hint4qpxc5/oJfKVIAH67QuaBBVhab
i6OqTdHSQTRgmIKS3uh1wq7hU0/a4xJ3Dn9te9Gmn9LPnTrJUW2yafWpcxSb2w6LIiylgEDR94NZ
L9d+DZ/cqMbFy8GUu/Zj55iNlGM7LGhCzojSEXX//1H1bsthYWCG2w+2dOqKPxkLnhyNgft52oM8
heuFNZJyiXeN7gGog5d/f0bglBngkXw4wlQkX0lJamkldlCKr0pbHcpEvpTcbfYXN8NsEFq4ICS8
cBK70uR0wfixy6wTE/qgGgsHY2qNXmgvRJKKTXIRCVIaPolqpdjQjSrilUBa4lxp0GkDERLvrkGB
2ljOxgVvfI/zTf8k013L0uv16apqzBOebDVOeQIqYyhFslqmnSUIxq/DIrQPNKpN7soSgkSOdl27
DKIEV2FUIc85XtM6QeK9BWjNCkYPd4JpUaK+2jpdIapi+5hK1BmtBCtBuy0rs2/YGlgzGxvtSIIO
Xv2Yj4SiA/WMYDeFvwq7faCmow7qJHzpw39hlScG7a0+qn4nV1qB47ugV7LLYmdXXwaHidkzeZQ1
LuyabTOrc7yC/35FUqH7PGIm6Kkiav4IjvryRMinY5Y0UMIqARGbkBSFZw69lw+urivwT0TXs1rz
pKuM7AcTZOFnwx11Z7L8ovPzdr+iVeguuOYYF3BWvgR8SmprPQKKuismNn5hcD2xx4YyjjKc8Bd0
VceY20VGbMJSjrvQFibC0RBkIkialbVYeDvbyWwud0AkAVuqyTNcZRRRL1MpVzouoHR2TcHIdSXE
goJGZI7hGMbqscqoGObzk+9T7v4OZHzLbG/ShzaTl9ySs5dj6czbxC+L67yviDlwDBH13dVDs9tg
rkKvSw0ewq8cC8RRXeR1ITtoiWcm0dA9waeXcdrMKOz8qu2j7d+uV8ANn8yFgZGMvQhux1Y6dddG
NISOI7iD2k7iYPnEmM4VQrqgrZPQVVYsKYVUomOSIqPsIvd0MDJR9+cWB60OxzIx6SyppAlHqm5t
mlq7uSKEOy+sYJa8b+VwIVrhalZGQzfm7tcVAKBZX6V4G2QlT9NLNuPEDwudO0Td5js6CKvzzN+j
wgUsTEHNRADhOGKOU70u7NnKlINqKaRvqdOGiFez/dHj5374AHz2ApEsb49ZKHTpTtpfNr1Eb7sc
AffE3dw2hGvpX3731fFQ+dK3EP8quU2/NOggg0zw7zdXeEO0fVbzPT1rsBgGoU8oHv+9U6ejToUv
ytSWDI8GmbwJFhsjjtc+01zAXmtkPxiIk+pHAcGB/f1qFb2iTj4hVKWbzvHtgfx9ceHOCQR+Nm7P
hZqtfftq3FQkInxzFTeiXL4fldVkDvF35wJz4T9WT/rMhU1ax4kgf8mbcSGKw7ASxjKnVklzLmZS
cNEYlVoLJsqY9vJ/TMEAHdktdmoNFg/qvcG1chgQ1R4hTQ9yH6rISGqHOrXgcmCG3Z9hX/cUXtrY
SCRebDBfBpZe5IcGRhgdZnVmkjU/Gh5YVLDWK40uDAsY13OcTDOSHZAPKTIG/FHqphWXldOIRt1K
QXWf5FJCEpPpdwmRaLcSeKU9aIAr8G33AcyxzLL5orNQ/pjV2pDuE0P/qf8SnEZH5NIP7Kp0l9cq
j9L3xftsyeyWIect21UgyNy3EAxK2xM2XFzbQKdUx3v7wFR74haE1KPN6XMyNaBtJYWO0hIyNlJm
E6vthmOu9btDXghkbB7WWZnB0LrsE5/F4A4J6XWhr1teI55kRiqXn737QJi2J2CUZW9ZS8cmsGPx
bOJ6gvDndZbQr+UIOc8Cr/QmX4+PTKPTW6B8nxlxDkn+0cjAVtkCVZxJmhUMRz7HGPztlNy3u+yU
VTGUVGSP75a64HzmcmdsFCqFYsnS3kn7ctXy5LOkAbzejABvvRZAmDXtSh8SECN2jYrZDfiJPUT0
aG534Ks+JMsHNwFssVqePL/F9YTxVv5S0Dj1/tC5gYvWNDvSBHMYgfhRV27/awEflfH/Wl1xIqCV
kMtz1iPUX3GpUOf69OJJqqXLtPmQqblAEh9kDdFx1ryk99LPAd48rW06CObEXl9OaSEkoPTIs0d8
Ty0e2DC+WJSdwuaXz+mujLjh6ddlyzdMAy2t37f2wOwWIWJz6M6bLmZhoa9Bco8+eKDQUBD0TC3+
uzBba4LMe5XQQmDR4NDnvJN6oE6irBvp63K9zmgP7QxybKdJ8tFUS6WsSxkppU8b9W+SCfg7jQ7J
XORgLnKld+XdjlbZETVocC6p1lEyDI/sf3swTqA0xdP4Ls+BjscvyhJpwqz5moMIzbZo55gYcPCy
ZimF7J5rMM7PCaFdXA13eyMipRJ4dXpCcuyMgG8+l+8Gyw0DL1rLHeFlMRmjeQAgoJds4EbQT9Qb
E2qQq+9T1WWRDP9qCZcMDUM58RDu+XFD4J8LE4ikodUIxNJyv6FHx6pubd6f4QEcVAstl8xx2/6L
nwsUdk0IoG36nANjQFZT70tAAARd9XLbQi2bHHV724bhBqcERf36OmHy2pO0DyoyxjeQ0ayuKoj/
aGwMvET+vt/MsEzBzl9EDwu2/rSSOnnxhxiLtYR4WXLigmvSEr78otESjUJBZjkgKVUL0vQd9XH+
bYSHS5bh5aNhiiw3ZcGZfcQcczlHq65EpbbUNuGJA4evbCZBIYUGLj5DLkY8CEvbm1Y6Z1aucDh0
vKQVd7/35bk68GSyObhteQR2hNSFXZtqw0GyAEkkD6anKQKNhF6V+UbmV+5M0ADGWLeXjlwkOmPl
v8ylPYAORBCBzzTnEeQTme4gYi9hj/hLyzOLQ+N6vB51iYoYb++N8Nh4LF8vb12yGSgt+40MDL+a
jcFkoF0ANwbtowTTpvv9BiUuZECxrk/LVzqm2f2yY6Qh5Nh/GPPjIap4oYp/u4ONDhj5kwppu6Lw
8TDPyJbt/H6+HMn5WQXL9X4V0IeoeGS6G8z8QV6BECMA4zUP/JfYVg+P/NTg3K4CBrtxI/zrYKnI
X/ivsK1a/PohGFruI1oRFsFGQ+vglOM1Iyo21bd6aSwWp+2L7E6tGEz+KljPk6o+gU4p9tsebFlE
Iz+IRGSZjw8PWte3bWBB9cn5MOs0hQKgd2LfMT+dglcHzEwg/dHMtEv2LqHBNeixThMAxXM/kKQI
nCDp5fPgrulw4RwszVWuml4buI7lwiH/w9Yd0InW22GqcwSKMufOJv8zojEZ2nhCK2h4oRuIInSS
bLDoGOjCnkxZej2JNPCdPRoxIBFsIcpiM7BlPAbKTejdxPbDTthErIhB6UkE7ADCA/mirCc9ARnE
D4SDVVlfNtxqVcQ837h5UrMBKsTv9lZtChMjRqP3gLX1nkfmP20eXczNoH/l2S7ONapQgyWOhghM
6NSItkXZWj3hq7bdCpE0o81JOy/LYmMFORldZOqtPt4Vs4fd7Q1PvF1KDUNEfwpGcQpPvIeYL3mY
L9x26/PY2VIZxiHYyP90PLeYY3ng01wIhOQiJB3/VUwCGSvRW27RJYmU19tsspqKqINfxz4wTtQy
tZH6DooU7u6cWDevaKgxO3dP9vPQkm0fKY5XCXYEpvStw6GlUfNCEdJ7cURWNsZHEYO2C8vY7N5c
qkVCFchkCxBqYEf0TBCwQJnfySPmtXhrKhZZQvpjIgEbpmSPHp0rhMoMNCV1usVZZjqr91y/CUJp
Gls4/IWi0VtyVn08E/WpXpqOPKhf4xKkWJiPkzDi3DdRk2ogrbmnIsAt831rRvI9YjsljtCWmRYo
gMJeST855jfaxPrRW7ayAK03ZT6ns2FEU7TwVCtFGlkhlCr0Z+AiQ+51EX5DoyS3esQLXV9/uSo5
12LaugEOsk4XG0nZfWHkhxeLju1waOXRmnaklZU5GWCr+2SFFd1zMYe+Qe7F8jGy/DCh3Z5qN8nT
04y8/HNV/edh8CpAKjofKvjDbRm8lEWSzr2WqJooam9iO9DEo0BdDYdsPUwiC1jvj5yVar7LHw5K
AhWz9jgZy60TL8o2d+UNM/iiYYA5KtIo1RiW+LMJE5efeGUlvGk46QnkcTFojUCV+Qzg1a5nNbXD
qpS+JSjGHTyvyZfFS2BA4GiF9tET5AMBlB5yOQBsUe6fEDQeErMPudoF8/OMBAmdbEd2B6/7VPU/
fUNP3FWrbj9R5JdDL4Qq3333o+Q4afI0Jy24JshcjLdosC20enMgeH1bp79MGwqg95bKnn/M3dfF
utGthfutXEcpTpwkYh1jzFWuw9hh1i08KuBGfX7pTD6cHmp15b/QEJVFD5VfmcPkDZqkZ7Jkyhc8
2lcbGjyU/k9E1aEHMq31eWjYelxuSyZiAIgBkcZce9L/f9jHUFALlOG7BWRi9JKeEhKeQc/aR4kO
sWa76d33rNkmfOYoQo0WT7/yZL80IosK55LnVZDp3uK+baOSpG2DxBPHZe02MPIRylK+TQVszdNf
IMcxFtkVrCYOPwq1OjjiCbY0fEHC+F9lPqjA3nIvFyZlvtm/fSYK31kpacqNKxcp/wERj8ZAih3m
YEjeRmBooiAEBpMD1SKrn/wd7AlLaMMgmTagVmhybGfMNwc27TqrzhKZFakOWNH3XYRcvIvPR2ew
jCu294+Gdv5qdd2CSZfpMYreOC8JV83GS10x9x1ULtaAnvC0sV6OTZ4Qs++aZ5tTpoNqh4ap8Yi4
7Cz3Fm6qTqnuP6kxf5C0ZZ/omUsNhvVib89jK9N0O0w99/BtOg6ElHMbMR6o4jVltlO4lj85OJwo
P5vk10wkBePG0B9CknZbNmQvhElyCmDOxF4tZwWTRFk6ITTNekuaVFfaadEOfy84TLLW/fFcMv2s
a8KYGlJ53Mi17c05CgSzwqocul01B+OR5LRt56fhTMQMude183hWbGq1g5g9KIU0Aurrp8z0Q73j
Q9MRfH18BZMWBKVoSkH/Ahvhx4wugPSt/MqQm/E+d6nnxcD4R2XrWgHmldQcCoxJbPnjuxBAo1Ee
Dle7Py75PmhEV8PUV4wX6b2mKpQQLsfHSMoANA1SGUPFLtHVwhqtpcdBtYte7tUu/H4SXkECENsc
Si2l9Pv++aAiX+5irXyVekSlJvizhYpuasOvB/p8+ECbaKG5xkzo0vKqvYtyNl+3+v9tREr340hU
XdItd1BgoQUugxPFwT8ViXKbPj67Okfw3MyzC66dCVXwgIDFpmagl5LvMblrmP53kojcCoCJMNm+
kBpqKGNLp1sgCvifkpSlLOs6kRTQtgqv87458/1FVGP7FnbqQAwm8rJXczUcLadMbEcwZzVbtelH
b+UGh6RWhQznF6v+sSmugafn+LL9XJnjWIPqcCbqMSa30YZ1mH2Zoub73uXBubi8dLYEKh/gIyos
+SW/R3dMDJRk0TAViBmWwOEik0lb4ejbqZDaeUlH7wrS70aYd1ExbDLVHeyBMDIQXVT1qjN6G8eT
xj5oRQq6HLXX6bQrcDbxkWXwBa4PpOcvPCNfnw8lSPRdQ0v7+RjqS0r9C1N1eYqhYTSHS0tiSqph
SDH0CdE8CXqVRidAuK56i5X5vg8T0PaNvH3O8IDbDp9vQreKCj87QijW2Gs3g/i6MOQm3zLg7sdQ
MWgDOtIfIfqCpsfIBB14NrFjQwq6AOgmrubkJjqMv+eDi930ZseF+3bbjlqUJW7JyW5PomVTfrbi
O08CRRf09dDN2pm6iZEeIvTqi5xfa/h9JW377+l9EfMXkEXANtbH3JrdDlnxm6AnsuNkShm8ZhtV
7OPL/Fs2wmFMYjyB9Xq+lZ2/ijegWQt3fXl4rhyFsErgUXaEyIGWHiE1Vz0xBruvGqWPwqOGdwXZ
LIeXu9RPyPQxSErhA7lAPGvgDDKLuMbxvmw+d2eQkeKjW+nHchwZXEHStNAtFxskADt3WUnhiL2R
oYx1aa0perbW3GEZ56vbkOqsOLYeujZw0+sfPOC6ejD1GI12MdRXijcf6NAiCZ0AEddqsboBh9dc
pPizo7WZIZ0wGSy0/cd2a5UDofnx/kBBg3ArPcVBhJFlI9UvY6t4RhiYWGjOcboEKicNqX2QCXq7
XdGYauBv9u3gZhvaQT/2F+8UXLtKQUNno9XF8QQ5axx1N41aKWcBSuSw5VDmYAgEOnqYXpPomu8H
wF+Na1QgWdWeXALkYM6++R1qKQe+XKo0EV4SA/kkQI1nZQH4jOIc+27PvGzZwJUWbk5Yc95NUZKM
qfLjmeScGJ0VUl6i50/m8m+10/KBHYVmtd45FbZOIWW8hqfyfrW4xV8mssJAn2zhvyMuFmuFz/dN
kh4GxrWAVur8/XokfliMj3MiOh+5zKi3wclzY/8rECt2yJiWhaZPzlWWfwo/IQXPAihhTXYHn2QV
7S73qKt4uRGha4nrRyE9QmxwIWNY6ac+cCdEq06J2Z86TkdHsznUcWDI6+W6ebgjgLe5mZbe/wVc
4ieQwD14kc1V+57dYZnnGnjFaDnmBjpYHMgW+WB7zOiCKdgtpWPreqSB/2tvRWSCiycRN/WJpbZ1
jChOkIsT4doATzmTpTIokSfFaJCFPM9WDUO2CeaQT9iebq79tJe++bkJCiIpcv5DrSHWrDCEVDTU
iqR2u4fBNjsa8gZTiCFKRyWvf0Ys8qr0yfpp1Lj7Iub6vQJo8BBaf3vXfWKcY2TAFbIScBNHgfdy
8JZXRKUnbuTRj3YqLCv8ChRutbFqZm8m+iiLKL7bhYDbBcZtlMzm+aK5MguTh7dnnTSYNKXcuJU+
262plY7onawdCg+tafMoVVTjgJmvVFeCuaDSpMs0dwe2NBrvZEn7+RaUzTCZ5lPE+1TUNhreBICH
FC5WNbRj4qW140EwRItVcY2A1m3kI6Lm4O27L3kalLkoEMUXowa4FEB1Gt0Sa7qrT1vmwUguCm7h
4xUmHC2XGLTgB0Kw/6YcJ6M67TtF06LCfXnle5FmRYBrYbKnplk8x/YqTTPKa2a6OW7U9O0QYXkZ
SSWxgJKh8xFY9f6SoN8Icnvo+yU4RLpd8QNld0DFu7bceLG11nkHVLaOrzjrNlOUfnRETr0zFTah
MdLN1YjohCUHA/riF32ozLPXcma9pmTbf5ip7Kc18TDeTY6st7GPbtOX1+9h7hjAj5VFxp2C+yty
52EdVNsOsPBvQ4GorqPQB4NBjz/izefQYgJQXGXBSfGfhPTKEtUeQmE6R2trnxo86LO+0h+soDG3
h6+NjLbjkQVWbuhFUEfi8uSlLWgxDnQdLYj3udWuK8fNdT7w3uaUv0tfflYGIojdxpf/2t3GdkJj
7PdKIiEDyzQ0xX140XCmMmSq7YfJzzPK0v6usNle8EOXuC7Jvr370tw968WmSoQg92fo9sv7O2Za
wqbrdSPoGTRFsqyHBmvHb6bEvoSXcNYCdKqj+o+BMGV5bhQRh7IbwWg/up5F+6FvLbpl1g0LpzpJ
aNFns1BvVfFI3cLrZyN15+zwWwW8/MY9MoVXEEGyxTR9LfbhSPjiJJCGUwO8p4q+T0UvazMMyDxt
iayFrky5HYX6dclaFq7mHUnTW9xq+ya69FAs4mYKJJeh79d/m78XqSvarEtZLREjs1TPS2nR/EM0
+MBVp4KWCkwGgJkEYmv3iCh0F5XwexVdP4bB2xUJgESvb17rh8jctqht8QGLcN9tDCVOFMaSEKvE
EMjLMBBycglfu6Q/XfX+SWiQDaK7XQIVl9YR/ozExsdAimz3LZTf8zMRLDxFUAoXqDztMji7DpR9
IU14g5SnOIy4gIUwWg/iCMGuAS0B1R28dUQqbwSgz8mKjmelv/zAPmT884HdKSP0DAp62fBYQlbz
HR1dAbyozbeTfFSU5g7lZPjrbzZEE4KuUoFazvJg0bz8OIyilAm6UytNl0z7EW6fA8Jgbn+56xA1
oY5uqf4lGNHMpf2dt0Oa+z9cWfXSCsYJs2SnWoycZ6H8O6QE0E4Q4/ppCoKmpACxkHQ/n5oJa4JP
h+kMLgnGJv4fhejFPFhGkYWnOuRwvsgv0/m3VUM2GasDjs9nVpDEVEeXXZsgQiC6g3VE3H/WTysG
Rpb8BG2RO9ZkRiqzOl070Ykau4WIqN48I9Dx6AlwNeecQJi4doYG1L7l1WHYfo7jOAJDn3ylO5h5
YFQBI9+sr+eglEsg/f7bnad/8mE7jItiNsIkoQSZZaULQZI8I8YwE8zvR1A+lKxd2OHvBWKkiY0H
U+//l+ArG+sqRHG2fWkEzN6G4d+n2XKkYro2GZ1+4/hZddedfdHgNcsP7jWV+dyr/n/00eG2Ws8y
TnUiBKCbeReD09Lzww6Cj3IZ5g7OkSoOREVO291E7XtPDwE0PoqbI6rcwCgEyL484J55tRaESMux
u+uoB0r5Uzz8a+ba8sNMoimL3X13zx8Mbha6EVypkjnYeLAupifKJIHsIU4S1HKaQftG3DqNOSpd
sR/TSkEo7w1W/EDGogW8P3jbqEvk5xzxsWRTeEq0ANphQrduN0IbfGmCDRH98cFfqY5x2C6oSdfW
8hoYVhtniett/Ih71V58JFCOjfSi0UYxt8bG+iVSVNM+OAGdWWq0Nb+ezsY4EFnJsATJQIvpHpzH
WFUwjbmWXJtWp1UD4e6kqexIJC3w9smepErFkxlz/c0Y1G6PfMJB/aufaqQJOC+ZteuKHyXZiaUU
i25qNa0WZthz06uGUQYsvpPDj0a2EIMl+zbPWdz6JtAndzwAZZxbg5xx60muUUn3BKc1hNCLUzjY
t7qqyxZx8EX2/m3xdLOVaHbYlkNXjfeTY92QjQUMkz/SIkJ8OvEO09nywOat5L/Z++0BqeKmwgcB
S1tFZEeyQS/gkad01MIAX4oO25Cb8RwHNhr3tgH7tpmb+kgrzE/gFv5mVAHYJYqIe2/fauwqhYJF
JLibdV4IuhoSfctl5ACZGXFgjExrd9cGvY1N9t7azAW5VHsH8UcNbRsVFizRvWEdlYNfpKFUYaDp
UhdXoGfSxH+8grXNaabWUCBgNu2WMPruYc8+zrlMNS2tpUddHef1RcXibw4p71c8HZcHn1LMJuX8
0MmBpWClGCQIsGntb3kTUFo5g889ZRUn+1DDq5gLOH/GiwTEQ3K0Ou9w9UX7kPdAHC65xWzZNFYl
qfFLz0hDLMA3zHtq+jU3317bjLgWuJPUjKFGHWGYsbcsxLepLfBIzZRai+6lwKhodNoeX7psXcxC
n0tZQSLqMqcW1iKZEUb6NPRGrJswsBksn9nHgFoLSz263IJSIqXxo+a3KiEfBUDTJ7/L75uqZLQE
2kGsa8g0JCxHkGTLviL5Um21Y3FNl36RLf7fTwT4EXfes2p+ZvYbrUfic0HxC3uPm6y2ijPrQtH3
C2xBRic0nL8PaRHgHc+gX4BGIeO2iQcgLWqMmPsxVJh7ztS9UqnFUyueDd40DgBIGKSDAv8hCdS/
7q5Z5dYbz0skw+w/awHCuF7IfVb6PoC3dWkm3Gvad4Tw/VLVqY4gSgiTznb2cvxa1yjpmwwj5yoG
U86ZRfR8Ho8scyFbFXdn2TvJ3L6Cbc0Gc5SRCV4Lm+kZrPQOjEW0rDbN8ll+K+5Em6009aR3S9t1
HeTQcyG1tGTh/jgBG/8jKPmInL/BQ8v1UJdMxFvTPqdat4nKd2vvbgaT+cWcppg4n4A3lkTtq/Eb
PT7swJ8b0m4LGJMr5ItHpwN9mQv1CM2RJgypLOfcS8FfzceLFkPaaCXvQa1bcAhy4yXsggYiOSC/
o+ZfeAKvvkf0va+nkVm3IOqKUsLURNPQFWLXWurY9gE/+iL1oo+LlfKsrFiu6UHGu3KmqjIutyej
T7IxapQRnFtE8XZjObrsG9URFFeStao7hs2KZy7cWmkKoWz1kDhoKN+R1Su7ZLxbAPPKOCso07Cb
g5DxNTkKwsZGe3HQ49gASGDdTWKc/7r2w/n9G1zd/p+UK7GyRYwmymFEmJseCEbXM0jDe5ZetfBa
ABbJchwfvp7MIbl1lm9CAYuv5wEojBB1gDjAO/b3Ly3gvclqBLiFvAxrwW9TJcrRhntfpMK6FUrT
rrBwOLyE+X8GSHqZc3y5IDgtdnNnAJ5Q3Rx6AKhSoUOFSngn0JY3b3idv+n2OwT5rF2vo5cKPWx8
n8piGKIJffZB9mg9nO1B5Fr/TrEox9M/WyAZA40joayejVAFTWicFsXTsWSC1GzbDiVqxZXp6KMM
2o0UJbXqZEGUienGesR9/ZxWTc6zuHDI5tohx2LSe7q6RMvTx49Ajc4px+no16iJ4T86RRB5b97O
GFz5qI+q78GTtkEqYv18gDvydk0Fr8OGS7qjuPU/7u+jWG2nxIljz4LiLLkiDryiZYefu1018/mz
b4jg7n77k9KnSHyTAaSyeuQ0AdJ1HuaarJmSHtjU1oWMy6kX8fMNV1OT726DgOb7GSS/cHKj6mUS
hyL2Lv8PDILRBk8L42GSb3cndVsg8MT8sxwX0OCZNEUwB10OfHkEUghraRfdv61oD1Ms2HzixL1q
H4kqsr0SeWSaYeO25KmWJsyKVE5CW0U+DDo/0SXzvWM5L/h46Hcrjnl9Vu8g99LFCfLNcVmKmXiB
sctvd9XDfhXO1ur4IPD4NplyxOi41ssOoqYyWCp6UyiVvpUkxioHrB14gS4iAqrq/wTcNvEaELSC
+PccNxZPgO5XWUR0fD4YDkcajE9yskP4oWbP/ESHBxu5gEk5fn0iugfLgVrjnR8VNsbbIBfAgoxn
cU0R9tq0tAHKu7N79PDrGTX+ER7JppQzjJcz1TBycrpR60Bh3EAEG19m1FMueLBNX/TNi0Vp/mdE
nwHZ9bNB5DmK3ctla0tjUG5sz2IJGpt0VZOZlvt+vaJMCgMY+kiZE5GcO+yRVAsNPzx+w1hCdv9g
CeCJaXHo3lb/nLN3q4tEkyLCkuPWJPGTEUOs49kbbcW6kjZA2VEqehtK+djhgnEAfl0dnhI/905w
T7+7guzmx8PMl5K2Mhmb2LOhZIoEsSm2oVfkNHG2ZqDIlv3Kx1xShEW+Y5WcVg/GFCuLv8yKHuvo
yBb8PVgzNcvEeol7BZlGbyorbn99YViXHIrcaRCC+2jSbTVBVP4dLVjjjMTjIQWos6PRKj5GtDsM
tyjMr5rdpidW0JyLAS4yRO+20mDIBV/Kj28YO9qXdKNb74VoVXAkfCh+dxkcgDSqXAQ7Sj4EIEbN
DvasYtr7nkxdFE+DZ/FXDCUgbMGN0a/qPbqtDwYcNkWgCDMCR4GhEOj4O3KfIe4WIoZymCaxyWoU
f6Qmjg+NxHWGHQbNw3T/d6AUSGhrBtOKgDYRsQKrh4O8idfToSUnd3GOvXXnAAD29moanZVMPK+F
QA6lYa36W/W1G78V6IZYurDuN1bo+JsD2dB+LcYJdmiA6UmDssuV0/m2tdFaiGU56kBVf9a9heeN
Of1eq17VfNH+10XiK+vkEcIOOTA5MCZGEq+TPmeW8XEZdWOdhDmIO2bGCKYgoV86vu+3XZ6As+6M
Y52sQIhEvArlIXYutPM5cRyd7z7bA7ay/8otKYy20kkjSpk1sLKBT5PXXTcvbu6+w8IkhB1M2mvN
fJHBO/76aIgOn9afXIeg55D+/rMZfHoAtUhgKel1Hw5ub5Nbj/KRjwu8hlfLzak09OOc9GQTHs4Y
uGYj3A8kANDlFYsW8ZjWZyCyZkPfoGs4C0G97ExE3LS2YTxw1F4a/9eRj9iHwZdHT/8dD9+86H0n
hjvMyfnMW5f3m3EacVO7DcbLrU6lpcUoW3OcrE8q4dt0MM9i3W39bRe22+chAK8iAwLKf9pHR8B7
v/R9fGg5Q3/Dp8PthosxJHcsRc+VLNmbwU49mrmqVAqfGdPkMV8BPVs4reGl4tQf3DRtpZ/Uo4MO
v88aVKV0rtC5woe48sHn0qbFL2XLNb40bzUNlb2jAB1Yj/LA85MD4wvg7F37c9Uzk0T47AE1ri0b
djqRtkNk5MH6HAzJAwmhhcgCe1lnW+1ZobmT8If7wTqZix6IxWM/VXfEJEkUlCCvlb+1WlnDRY+J
Di7QTbTzEBnMWAFEnR4XQIxu7BTGjkm5iEkID898k4EyEdU4EwiiO2WZMPHKPVIMyErAmdvfDxLj
fwZSI2iUTBGskchRsqKDH8GRA4hzN+tuQgt3Qa1jtJKf9s2g+3BZHNutCYFLoQyhvhvnPTRoH+ME
FwPm1x7MKyr3+NS9u3jQjn3+5VpO4jzK7uEZjwb4/4BPIu6nWQhJz7sNijsWjh28TOhbF8QN/VDm
EDeUSioMn0A34q8Ny72lJtsP1GXYJCx+JaqX7tPn4j6jm7RgS0fgTlMkqe+TP5Dtr8ss5ZvIZrJc
I+MciYQOZhQUM2hWqONjKSaEs+TxbggJ0/OrCsg3dcVkvUWDBoYNv/ASjBZlAlLZQrnCW2yGBUvx
k3+YbkW/C3nsfqmSQiBatAL8rgAprPyQ9oHqmxS//CP24dgBw3y7rjboGAVrOxBrZ6pUBGPBGoNC
Ptbr1ZC9Qpuh8yN3A5jYbFmgd4ydDYGcxkTzveIMbU2+tt/3C3HrywsmofOcCHEo8KzhnaPT+3t6
qtYYrDmFWEgZc6KN8sfKOLyShAE/7i3f6MlqEVhtc45eOvOJJUBFPN2ekeeWn/hZ93QyDBFJLvV3
lA/ZvF6wOl1sdEctWcVDaQn1/8rkwL13/V727e2iEfM28Eq94rdTMy6u5pqe/5w90+phTlqh7GBE
SZ98Wd6D+Q5RqH9HqM/PBUODZ8mbhu7K+No8VTZq0pGb0HuomjaibLtF79lgWgBOJ0b45V18VfXh
GiOzOSbj3rBl/TYqGHfHkYzQ0R64Hup7eBMxNhXflQmlnmkeB4hVE143G+40+Uiqt/190NBXiheZ
xMCs55e2EoKRQ+yTbjU/ynw43KytgoqyCzwrrGY/sCP/LblmsDKO97AVMkLA4YL3MZP4AbymUz4L
dH6DXdOaZOtG1mz65GHaseYOIF6ih9qhHb3mTjuwmtc2D2CeG692SbOMWesmhvs3z23MthLcNHrs
JTda99Or+MrUT1QKxWCJ0Br5y8DfmWVK5sskVEmAaAsAkpKlrK9PI5dm4Wq8YfSQu2cvJDWEZnak
npIym++WQVwPTbM9UMMr7225FHK048+gyUzNI8pj1HUInBQL4Gxt1kTZraOyQp2W4ej4m31npnTR
oc9Zn+bFldrWtQad7k3j5H2bUtlqFWVcldtrXOQ8i3YphOZ6YVglqOvoK3uo1vOaUNyzrQvAncVb
HNM0iaIuneNcMd4vl6gCxwkNPfV+xIXYI0U3SYWvGj2wD9/9PKlIGavYK3AR0kvy8CztKM+ILYzz
S1PZmtcOJEIyGIbHvlI9X7A62yUcIVBIMPVIBJ1DdfoJHwwIP4f4WohfxEsF7y9wiO0Sl3okdTY1
6iomXKK42XRcVhEnWtr6hNRpnDbvqr1nfXXtn2ivtgCipzPwAwVWnYphaCvPAzSKxq661KRmxAHA
PkG8wO44m+VjyLMqSQtlLyJ/lfdz2cWeQ+XtHcAk0x1x759sBHv5CMxJV5Zg0yVATWHSGgjimYjM
6t99BkCstR9BtVap5QmpB5EFnVZ50aFPpGj4c5AusGc+RQL0J0o1CNL/nLBJtF44dCvcakVPTRqk
XXpljbvM/1W0jN1o7/WEY/G+mCyJPx9gHcH4sD7Pr1tlBG/AK04IefAhK8bLjJ64w5726aOXtjdw
hBQ7lBnO7aPY3L02FGECPdzzIqyEySsy/90D2PjAO0WDgDCgqWsUIig9TA2mxNjvoHkzU0oV/YFG
JyiZc0+Qnz7uLvzca7xXgu4+/VTc9KfzQKbEDqRJHAWCwx3BY+gDZ+4uJBKK8MhTdT9W251TC+9q
k26EzIE9YcaSsT+sOc5ku+OscCu04he8v7CDCh/+bVGtfQUZth7qmdB4nlYDsqYX63lvx7gztcia
sOu4X5zfmyxm40JB2J+mutpMOzrEKAI8BrLJ5KloMZrIk35B8XMGwkONl/QsCmMSbNqFdjm5Wi5C
stwaQ203ElB7TaeFcRpUOmITVnx6ph7CNQrXFfHQto8IK7N0Kt1xOc+o1hPWyd9nW0MIpMlBWWct
5ee8LkldlI3RITtUexdC/s7QdJCpNB0d490AnxGQRgpFcDdxA0ewVX8jFc55qlKQs2WuFwlTDvaS
/26uItkUsLFRYFV+s7IXr3GwRjVS6eiywGaMFt60tLRXyofldJnu3TTACDaRl3wtL/iJL/T6u3od
Z05aL7tGjp3s5UpbrdyXmbkkC0d+IDUEbMYLw6zgttSiWsoAw2pmwyj1ewNlPsZx6RNxmi80BqaS
maJAe/kwd8gLFairAziURLlW9Y1shTtpiiSYp/gCAUKXsNXioaU1mDBcG73mJpZOtcuC9DQDdg/u
v3zDnyHJzRA31t22NiZjAp/iRn1kH2hwL4X1QPOmSYlYPfGBOJhpj7LPdAonyLTD4CDuNH/esukf
wle9OLINnbDboTN9KIkceSkv3OLKIMGqfJ4u5uGZgB0FH8b92B0RrLTMZVBHvppbizUYHZkR7tAa
ZjbrCosS96nnGxH3NeeqzPfk2X2wFbkuYpjipBwQN6dDSZ49ZgowNUt3loQzpsncJXMUNEmMRafh
Fy5OqrBDGpF7zJHyZZAvKLZ/vqtBljeGUVOi7N78eXUaOahHxX0XX0sX2BBu6PPnYt8zEVB6Ijgw
3dwC1JPZdfF/tIl5c8WUPF4NyqcspMZuD8iyzpYV7lzSMRx0/pAmkb9x8lPYCWg+FUtZzNt+wKf7
Ue0r/eRRQ+5qf9e5re2QmDCfxFyRbimdEj48QVyCYkXMYgpaGHIUGt8rbbGiGK3ngD5C4OJCzGOc
v08/77pZdpUQbjymZ4oVcQIlZfzApX3UyUfvxCiFxOWwnEO8qQNLtZ1n4yvj9W21GDylWp8UO8DO
4vsahL8KWMImUGHfK+15x4hDPWVeu7PLATrPtD+2jCo3hilJjuejLAUanQ9QjWb+i8OsduD8miiS
5u+QHfzyukYh/Oi3KjJq8Ri/WSNuDvX1djRmWDVs9ARR4cazukLrAdJ+6q7JKBmoi8B1LaV7Asir
0f0HVVLxLI8/OR700Ljo/SazcsWyKAJXYRoYxcl3w3qkZ/Az/YQ4ecYHLSAJmPQPmZ7uD9qbsMxs
fNjd01Ng+afVxG1zf63q/o9Q931gWY2Mj7JeasnOXSQJ0KNwDO++U8D0gKYBUiA0RWDRQgWtXZCE
sIeznwARw7WM1qe4HnGopSiHaZLlY3Px0rchqXXC9l/B+lhivlpDvvEDcWIwo/Jdh31oIwbfP2U9
SP6Ol4thzWTA/OFiCt60PZFtCq6ZUw5Lov16ENdnpH4/fajDRCC85sAgmERCI069J+deGRhy4hEn
lAIC4NKJDIASrN3JNhBcedkK5MyB9R9jNjgRoVRNkboemJiQD+AJldYSbgQI8VaIqW+dSsNPGIoV
RNpg1ZhFjUyIhinrcWIZXcM34iwPkHX3ziugwaYxBzcCPQHpa1TPXIB+i/j+4OGXAYqSOze9kup0
BN32Jkf6JTGUESE5ajxmGUy7fCK+EoNk2tDQ8ZbmgCluOL5ItbKFcaaY6/7kkCTa8ydYRzd5hWrx
lknhU7/VAm670ihEbLDfMuOIuviKIogT9siT875Ihbeia3kVCodBaiincJ/bvYIYYt5k0gBTeoiL
OipV0QaKFd7pZYnRWPS28bTje8Gb/aOv+ms3kGZCMYd7tT2666+jmIx+plpYBEwKb62q21sfRYBa
q6vSx55hJ+WVSS9Uf+f79vpMk0/vVXvbxt3zZncfinXq8JYc9+9g0eV+wqDJ9ReRA6mbGbGKYTtY
LN2NsSlWhGon4V+5yy5YZ1Ga6wSrZlQpyVMkkJz7rJTRcVC5iQp0btFzmujUUJiEhtWDtvG42I5p
4pnwVX3bkuk2VT3YyL3fPXTMoeRMokunmjRJayN2L9CVqbIG8kqTU/3QBJXiLJqOPh06myXR4TH/
YlO/C9gcvGci4OSHz2B2NwYCNdyQGF5E1p5zi04k+qJfniimCaggsE4vGPQkzQxW4SwOhydMp3Tb
waeRE769uHsah9AZnBbBqixL35gPJWlftMOwqmYBtHA4u85Il/kxs80ALpfz096mFb6YU4smeCw3
xwmlMgnV6OjmoW7IyTuBHNrAqziC7ZADBOZgGXRztopZRMZexAZLMsB+F9mH3YkSKBO8mSS6JIK+
heE3uh2EdWJBOePiEqF1OzR5px0nq2VffQ97239QmEP+u/qv+CKq6N+CMDTy7L17VuV29HTdd2/x
AtQQAeROOXeV3Z05sdYodUNznpeRGrBNGFkaInuuf2sObnHWzPzxZqSby2MvUlpK471NGi4YfKYz
u/WC6auMIP3FIsu+MRf1106L5Fhk1Te83zJ2qq7l1Mr0T6Wu67lB6i3pvcTItup4aKdcvdNNpsLb
FzPGrAAHQChjb3UZxEExEGZKzRPseP5QF4RPpwGiAHziWW2HTkj5k7DwUipVGXVrKawl9nIPsvWr
ngelgyw7uQOVmGEL/zeT+X0lhZFBFeIzIYahnxAX/CvGUmXrr/6qNmi/BJhvt8OaU0U56chV+x9C
ztQmbS1ESCobKLmKlPBuzCJfOSHY3EteUxWoJXnMY1OlBioFlDAceGiC+ixrkSEmHzpnK7P34A0q
AE37renqwzbsOQeV4pOLFesrnJWtuYzi1kNJ4Jb+IVGZiW27m5s4tn/TVotcG0RhlWnmrsnxk2Gn
/W/SiAlnaatuTJNCZCSU3Es8OT7nZ/XeUvPQ0mFQcAcm7WraFI7LAw6YhEveizuCWik2khM8g6N2
enGgefo7RtAZ6GzPI/DWYYwp71AeUjCx2pr5R9rduXzut05BIHqO5t+bjGmAp8LZ9U8GJ51J/9Ou
OKn0orrJiIx4FWSvG610hSFq+U3pLUhdqjmr9w+MAdGfZoATE4sSP2CeLpzijTub1N1J0TeKTy96
OJOi5aTfyDxo9l9SXF0OchdAL7/zcfGmU29fol8OsrLsduIQfIKciY7CEKNcqSOwAe528nA+7nO4
51aDZANETPqI8w9CdbBgUqrn7sno7mPmCOO9PkvxNaBE9JLsF3jQ4UlVZvD/wbSChWVrXiWvzD7g
Lg2nrD2AXB7ejG060RQyjqi9tR/Qb9N5A5dTyCL17OoKWWKcltlMaVtY7Wv91YoH+ItyxUqWfIHC
vdjIJ74liuJv126lVCoLTZrVN3zmLvUqt0as5msDt0lxxa/hY8CQFOG37rDcqbQNzYYJVcSgMrNb
9jhXKVCapEwjccoFs8GFh8kFbittL0WEJToWyqGkIAhDjt/MCIqtFdDHhf5wjxJg7RCVuAX8/hkq
EENw1KZ8rfni2LGHBj8QlLb3Vg6D1NbB7YVP09SK08sw1q1QU+ofQoU8pcOYpAs1nBey0uhOLf+J
NQPOKQeDsARsoI85QcAJROSYxD6BL0CfJjb7ga08eqaqNhVntnycjHlqMyZQuvKpTyyEw1DGMf07
E/o7XVejR+0Nr6E6dvMaCD8ZmVFqmZji9BmOaHhCulDD3Bn4zGBFe/Cc1mTYGoEGaJxl5qluj95Q
Qz6rDD9MLNwRqHMSDMe0k9wNV8yedjqqgVJw6W31dQOtl7y0ETdepGow16RDHy1cegYTUkp278+B
5Un8L8ukQjt+sgPiFSXepF6PiS5O18ATgLCw50zejfr0dmlJazRk3EMdZm0SGcKUOjydsItyaa5j
bv0Yx5ChLmK6i4jB5B2n50jU6Uhqa/S+82UiXwu7hJ0md88fFY20E3wCMiaE3QkE2njYMn4AgBVo
YCBqsBXmFLaqvdv9WtfF3OSTTHydLAHFX70TlshYx4iqUQidB+2p1N0J50bNChewm1C+7qPKiv5T
ii+nHlWMPQ2WrKtA8LSsPkgnESPeha1d1yklUR10nMGxGy6BUghRpXPdXHtVsUnCPJQhz0Lt2R9s
PkJ1Sy7PRx2smuhEz7y6mHW2NdfY6rHF0CkK6riXL0wnEumTVOZbsAYueH7oyzq/RGN1RZU0zQsg
DGdtyNvSfrd6wvtLMmWcbATCC0nCQHtTr78s5g5hPB+Tnmg/uy9FHGOy1FAo5tcjev1hFyP15p0z
eRGenERZCAPAzSWVCCFwzxsyOfc5FVa6inTQqnOj6qes0suuLlfk6lVREqhACSOU9accPItnH5pO
nbVQL7/Pxp5f2ZTv6eMuz+rv9tMFqzQvsqaeWun89wV71TEWgYDI5Po6Aoj3Z3rFgFaor9S6bWVP
1bE9XaJujd+HNezSXdfDv9pnH4HCLAKAGk67TvF9S/74TNJOroQT5ENuwN/H99U69600hXWjAYGY
tVzDFT4dwBUen+tjkt8lb/SB3aXpYMLmbo3Rl56yazyGhQD3ci/SJy/69sCSs9kXD0iKmnrYDU5Y
3CWG79NwyjDpz4I2g/okfHpSGQs+OE5Wg6new3kpWJmfPm2vloHNYR0EfFX6PaL5+DHeIrryeB9q
e9r5wXPL/eovwHIhvffk7cCFBIa/paLB3TwiNrG/ZPZa90G/Q/2yUHaGx/4GCBHvP3BNsWiBT29O
NZRQ9K00MjWQ2T9/e+DnCfU2WUyH0Xf/hiC/dODhq7JqFYv29PK6YuI9ytAU5YmReTqs9eIo/g1P
VfSaX5tBCQHcN10HvXQmsfqbdfbUCNm8gyZjEcSOxle/sOSo8UVc4ZZqakXwEvCbogMPXBl8dBBf
2S/159c2NkSZ6W8R8g6dUAyqrF+MsAD3OeVGMBWfeAWVu3FhDpVDpDpePODQ6rOl8Ok9OxkZUZjM
oVCLzsiaTjLG+cPfIOt4bkJtc8pcNbY+RtUUROlwyY1MG6LBYmFqZni/qT9wF1KnLosRm7gMKKJR
z40TD4Eif+Y4DcmdchUQ5dj5urKFrYeUT5SRsoTvgX8/MXr0qgDfiu60st5t+zJg5MMcgzoSLuwJ
rFE9t16koTxPrvgTqhJqXbODI9mAqlHhFG7OrPo+7eG/OS1erpRzirfrAvnvPu7v06GL2I0UdpFm
nlC7PHmzvog5LVLCo8drWvCSJVAJMn1rCub9YCZXpyoV485GJSHfGrYuKQdzGvof+/6O7Xhe1ecv
BbFsF1wTEdVwKcmPTAMYi4dji6cNfvuH02LZ5gZqHLcxeaRSnIZSQAdo09ZD1ZMzqvSx7hEquaw2
O47sILlYxEt8QicvuXIGVZMfLhKPSn9OxOetLKmFwxWlBLIbcG8LETSMv2lvCr4UERElYXQF+6Rx
oTIm1y/Kr5IvzyLDTgwVT6UUZUPm6Zwu0338pSR6BLPhHcVU832hBQRAFDjm+9pq0A4jiAsRg6YQ
E8mEZbySx04zGfwIQUWyOuYKGuJSa1EFDgla5Lh0bpqWFG6XdOm5MGM5/92Tomtvp+m0vFZzffZ7
BDKHPaOGhji+UPVI3+ETA/iN+H1C1bugurjzvkimkCOHG+Vn+V/gadzkjj6AhHCMGoCUOWGdSu9O
cJVhgn3XY4Pvu/nKapgRadcogfovojBURheYsik/+wIrAykgXrIHZDROslMest30648d5PHXPudQ
9kUwPZX+8LrxeYI8HTMckkD0JklWCwCRnKIssm4vYfPvW9lrBPRqdQ5R1Z4y5ipvEatg441JTEpW
kJYCDZ1WvcBqqJ12Gl6cwDKhhhaOamdOMIHwLHyGVS9ULSTGeWmHjmIJeyeOl2p/SiHvPc3eobah
1lwbwfUjjUooGvSBfSTBL4gketMuyV321uvku6FA1FtQPbUTgpxAkAIGbxCamKUXXSNApIwoRWhR
fB7mAHKmnUhtz+XvWNjzpBVoCZObXVUcRAwZgVFq7j6ChdRFFfESuLG3dIMxtoinTD3OEcRC0tA/
0FeWO+BnmKUSYy55KlJj7BqxjdHy0exrBhwb/sx5JBisubk0kK23kznbadp1qx4o0Cb+GpNUftvk
GtRPpnr4BIWyXSmoB9MNZnuErt8OWyCtIEmpiEg+9dHFxRxryAgE4/YJ0Knx4YECp+NIUbQvIlrZ
+Sc3dJaMUbMoMOtKxhzUnCtRd6fi5BewueC+snlXxe7b/iEyhYEPle6I3zBG6Ht3Y7f97AOWFHGz
g1h6kGdH3/2UuQXVQsQbTyI+UaoWaMjELckChpXFRpMr8D6AXbrRcSClMb3r+TCJrbnuYHfTmG+O
l6Z0nK4dQjxfHgvFuG8ZeC27Vh8p6tBwzgFYnxM2HuJB84oLGGz6Ac9ZL2510Z0I0C6Nt/TNLpUX
ufNH2b8MpCvCIkrPUc9iNrRFXiDf3oCqc0c+Gauq1r1+9nDziIOIv8Im0kRbzNo5bVmluJDtg6Or
Rb/riB/596IvDBZ6yFz/JELyJiYUn7RnT7wWLAzAVHG/Tf8UN0Qn7LtnsfFpgs9981ZwFZZtb7iw
G4khcC159VacB4whYCxSujyp6A0eGgym7hu7RPFxdTHwltDveLLsJeRCX9bJE7BhG5jPXcbbgTTq
j4vdn81UbaV3ibnBxIGoyQN4c+sglhiem9gcU33mkvWkGldxI96EEulNqfzMOqbehxzRiZgKyr5T
UzO1YfOs7IQmVzxoIXXLeAbOSHjPevIZiSj7QD4nnxqUix1pQPiOix6r9XEenXnhinRL5gleKd2u
SetYs6Nx/Zw6ukGZ+Gi+JbMZSqiLdRhtFZ1Z4Y4dd0lQ7ijd1W/WSGyrbZ+Q75F4iw5SKl/PSUmB
OBsNXaX6JnXSrYmEfqI5jS6owACApeP0+RIWkV9yjASNIYFPfge68NLebq5xebV6gJ6YzA+hIwBW
PBc1iDa4LkU0pzNzI4kKmLY7Z2b5IYQRnEnYwTvSABgYdaBIMtF2IlvRBzo+GuMkqAFl0XyLzKQM
9YmA/lDwUBnjZmhhq3pDwXKwg5+tlkLMIvJZsZkEVoycfxcU9rXySGicA+2gnzD2Ame0Vux+WGxm
UNjIVZQyno+pLsSfHSa7ghmTluXXnIjCVDFeNjmrgnM4R7CWrnetH2gp+mZgebBZMwJFcVNhmt3u
e23fw5VZ4MZoQCCQORXfk2w8PEoFvhMeatfXivK+abmhhUEUCn+s+jJhbAAFGxjdyUFh3iO9klCr
oLOnzigHfvHJrQKzNctL6NErD42rdoJqlHETIKD6N+fYLoAa5mnqtblQ/TS6h9+dboHT02nqrCbn
6hM3V8jdw4Sy77qb7zro6nwsopRDIuaei8+suFoR4bTWotIUVHsIWKXS8pibFWEe4cgLA8TQdKgu
URfZq/Vrlz+CSHBIsFlXI+gxCxiyq5lWoZhaeGJzUrr/EnfbFK9rfRwXidRRe5a9lrEBPJSbhyJm
YJdYvtcT33+sVgQoqm06Jjb5dzfvoAamwI8Plo7BTL19XdI2RYMJmjAH5YVYlFVJWdLX3BQYzLk/
/DfEvJqCc54MTA01qn7+WCBvCB96Yj6LEHqTHNviK+VOoJHreU2RMBeIpKulyukq1o9DOovG3g26
Kbbdr/kaTy0ivgdVEwd43z4eYR+P3/DpGUjYMEVyJA04q8X8Ob76LcTxefwSsWE80+Rr9guccYsI
KGgDShV24CgAhqSCJejVuUFM9e7r4y5K8uH0iE/AneQWQYzGOvm02M4RL1UeJo9GRaBy5nwimfjF
aoboxHIvrqXpFmTK2Y1q0OF74SGFM3qCAW7e5j5Z1Ec8aBrjOuUZvtx7A1uDKYbr26qZY8GyNMyL
PBPfHVyOrGPhiy/Kna3ppX+VSEYWMPNTd7Z4O8GFHM/8eEGm8XJVzk/VmXzqS+LymI18wwm0Ah1A
AUDA8FUuwng645PG41LhL3J7lN48Ka4nylvRuD87o/Z26DUYp6EIHdiP68gWlWvJHpIQXL8MaGfd
FXCsERFWcSSJfQhXdBUBjkW/aa//VIbBdJckNA6fGxifqdnJ+//kIN/jiGPAPdBCdV+CiTjQHBVF
nl5kRo4U4CvJS7wOxqxbiauz8/aHRfWEK/Zsu/14s+EUFS3F+TRWWvmseR2islEmRaQo5WZHGIs0
otjqRp2q7+QMJe6AN08XEviUVngTy77iIctDHMyiE0ohHjuJplj9Y3gzm5tUNkj+jQ6Fg5/4E+PO
KnwxicsAvHh8MU0e/SHCM9D2LBAsNVhMpQec9RT6+inn9X2XOb3MqktJvIm7IagIwlZFxtRM7V1/
mhOZwvGVBFoCvt8KZoePl165tR6Eec9KEanX0Bv4RQXKPc1dXskkvNjiHYdCFnip4xiJnlWi80v2
ToVgiQYJGBDRh6Dv4KqcLZQB/V7TAiR3Ttw3LQtXGlXR16dj4t3jZc2nBPnmBHBMSEbHq1dFDaMG
XCZ1hNRSNqqiRCW8nTu91Pm/xTpFlRMhAeezOVKHFVlqDIOJrEDu/yzJUtcDoQZb0DIbNZ3xkD4V
y1evjXxbR9cnQ4KJO7OxTn8yDmUBEV+Q70o08Ur/vfKmRisdodJpT1kmMM1rZf4wVJvG8IfFPRzW
e10h22zPxcpM/6sBmfXoTIwhhv4QfziZ7cxJPSf7P2XtDeP/DLH640ZzSkJTtatfGb4gVtH2Coid
eUVzdrJ5tKnsweAy/QQtlHJZbj+bwiqyL2qu45ZrTOXdp6Ba4s6I6Psy4AMMwQzCB2fQnZuROMqS
bq4BJTu8flmLMiVHHdXpnvBK69H7EUtRyIzXsaIty/TBeQe2fz3dMJjyHSXS3qgGgoIKzEdGY5oK
1tzDJox545w67SDdH9Wa8zeT4ePSz961+3y8iGS5QYVYFpSpmgIShBxGwBrpdI4oTqorKp87VZyK
pmRO+FkSF87SVIRumSQJtPeySHk14Hc+kmGGI9U409t+1nw2WhmWLfP9TbkvcYWF7vGF6PzU+GWk
6gDQ/uVkOcv3trPNwiyCVB+rdt2O1mjPZjijgffxs4vip8HcqBqDfyzhlf4L1Uo5eqNnRPFXMfz7
cgyZNsomidOygrzK8XhWDYBS/uaBHM9WPDpGK4a4mYaxX+294FVKJuVlQD9sPRNGK/N0eZJIcbEN
Zb9d+iqViIF5ClShKHnkmqB8LK2FhlM/Lii1XTFypRkZ/qv+x+sl6BHv3+JrcXiobCVEnJ7XI0vg
Qd0iSnFNJVV3OMZk4WKxPPuvcDcvRAOPCni7w2BpNdCW6RUYN71+pNBsB73zVmPv/GrYpeGbgPie
78wLaz93x36S09g0DsmxZXlcF1LpDFPMAUN2rEs3O83o9B4LpnCu6mYSFZBxXzRVOju/ofSGXWyF
QHhXXoIOZRpDatGmX+/4if5MK9PFWXICsMozzGTo2v6QmxFJGBs9/lefTwPO0f+qASgsDRjGr/Sb
TpcPlCoc19VpLVEI7N1mxCUGJFg9LW69Mce46SXeby9tx+RU/Zv7EyBvTVd/E7Mw8L3gL9xYgQCN
EH4ZBuxQ9J/vAa8hIP38mkoGoDWsCmfCxU5JTwZlPR1eGgwwYLbQ1yNcGLYWzszqLF3dCGZQL7UT
0FCa4Ds+qI/3sqWKYdBx/9bf5ZZWyf4p6Zj+/eojfQ4Y5hqdJHucgFQn9YEf0A15pGWhiPnmYWe1
FQVJWa3XwpNbPoVgBc+zuJsuHFzijXvSInj0ZdvfWSFNkLVjHp+ZbGGi1YgDyvnC7w8BctqFDJEb
7BecVYNPduHB6nO3+GpBSVwtZi91s5ew0e6eiE/n/C4Y9yUiai9OBnJz3mvVOQkx42QCa3YB0x38
N0LVJOX9GYfCg35hVn2L4ju7COElLui6gRay+WaXP7imnbyYLB/S2JFXdphCR1duZdr8qlgI/8Gb
VlpRJMKDVBQDAZnoX2meC3pxWy7oReCGvfI+V95vZQmjdcVLkpMCHM4kjxK8IbqmNN3/rKdS1G8h
PGMdqLYM1vtQavSjLVx3aM5RPQMemHFRd2FiNIcBcUPpfEoQZCme3N9CvtmGF0yban87Akm8k7a8
jmXalPayr2b6IJRfB7okZzYbroZr5jNgRYVdscLXkWfoeYVQ+KvL1x1ITV7+op/KObOnqSGoSDDB
GF50SLwwq0cRzVvzxXztvbPFDE4X4ZeTS1ImB7fXHxFtTyMRsV8VrthO0QQXXx6bNBvsm7IN3nil
EM9vjyQpFZgl9udowkMMcM+kCWLv041gqUzkGIuXYOM6MqFp+ObgmvduySdhosZdWLGyu4Kl7F2M
m0MtY/ZP7M2P3S/SmsOYvUdRwthVpBec/Loy0v4kki2Qx4KwLDz7QMy2zVciPR+raLuOwiu34xO6
GLdCMPoMp3g3zrMUrSafbdZZ5TPRotM4bR1oDiJJ5Qcj/YM/kQevk+etKK2lQuSKZse47e6dRBUn
Pcyf/cIal52sKX1F9cuPC53pRLIJjIG8ai7jPGoZrvg55PSqzF1YX8IuKmjua5fi3LpecL29MOTs
Lkgk0e61dHsA6T6eF0sZp5RJ08+H4JktMHKsM29ZnVROl8x1zQQrbTWHqN8AARpj7550bbTbN/kQ
NLcpZszb7MiHddSbSR+6nVWkxQtx+pBPB5e2JZquRcTf6y/lMeWGTw5EGdyxYfoIJsq5+G7OVDpC
99cvfe+pyGEH93dnnVhRxCnFMth5VNikRqWVDlSlWqYADD6h+ysknuKzRSteBTe5a+aZT4rQBBUQ
KIMSfqERCT8by4SexEuMO+W1agqRvY0AdY4LSPfQoPGmhVzPs1bfGO69i/fKZY+lHr8YrL+B+U5P
hzvKtsn4mWAaIaCMbTyL0SAIxuODpwltx1jbPo91MdgmA0xX6UrhgzPOfX93CHJ50HfECa98gfcj
bU8POFXn11hhmbL+Iljg4WML7yHiGKR+81Uk9rMYV2hia0Rk1hwFgF5loGzIQa5QvUExeNEs2JhP
ccTkhaI7/sU+WpKkyxIsGulXAEV/NDQiQM/n5lt0b7rdf+CpOgXXIRs3F3eYTBXdFImICabE6cSr
jSURWsIxmmKcUHWUijWlEqKm34osJVS8Yp4SHVqrDBi/ViN9cwjD8yuk+eKzkOQQ1O0TJ0JbQW/X
iilOITO5ZqrepPht9o5SlQZT0bRnutgJEr3N08vTsxzqgzWtSitxthjye++8G2C0YCDv0fqAnfeQ
5CD0crpKX7f7eXdS7TF4YDR7PrGaXCL6RwEaWvDSYi0Q76Hx8NgAKnNdcitUlb1fEN8+1Snhn26M
NqHdr+TMWsueW70GiR32GIdwyydIHcJJ9w3euy38rG53zaHQVMhLlFwzxT7sYkayNaIfwbgXNsbt
ThCltnwu3oOkcb2x3fySNvV7MWC7b0zEMmrrg+Ta9FTIZtNGYDcsKdJMsrsEGzR9D+HlExkn1ZYb
iAVrbrkGBKBJaDPEj7LCGUTOv1aYpO/1KjkhoHnw/YMd18i4Kn4FaovOWCdwWAA30ikgEkalpfDK
GVitUKOXEbDC1p3BpagRGMUT6lbP0X74kA4T1IVKDRfk72LM2XKivTGa/BCHCcv29/EQBP4tJZ9E
/xU3N8OQP7sR92WhSLiiiVwMe7z3mFGM4NxO1B1HNE9j2/tXRpiufCTSNJeUFGXDBw542u7N2JAM
Sxt0MUY4GqruPSfI7l91STQNlhoANotClTHdEsDnv2j+T6YBdl4b0fYXOUSKThHN8crpby0V4h4G
MXDnRkoYAyf64AoFkSaIPvDSV/ZAMDJktjtx8cJl1lULoCm2GeJbynEeoVgSG5h7LomG9fnfMc2H
ND2o/B8ly74D4fAM2Pinf/4UGjytMAIRj5x/HKsXsG6hfnsvOsz7McGGCRbZuT7eY3TKjMV6WBBC
fn+KuLUsO88+zi7seic38vw6mkf+ZsSziy4VGLkcI05QXYrdpDuMx1BVGP8nKSyG0HcwR+e/Q2F7
ndqLYANXBiOTcNRTDe6FdOpetrcnJC+TtM3L2Snr46/Oj3hgRUo4MdXi6E54sWO8rYU4T6A2diyO
RBw12jKsKKrCjdeGGTSV460gvm1f7eQKX2dPXQWYQBEjlavBl06i+nPbTqlK7LOKlQpnxxY7i8qX
GJ7+V4dCKvQYk3c32Kjh/N4RyR2SAnH/dyj0Rcz55n/NxoU72a2/w1mPzMyR6E2hqV0cio/puIG4
DKFY2Lv4OWrkIgGH60EOvZPqbuZtYFZork8rZXg1SyP/Y3CjTKwbp0Yt6/yajmn8pMFVZxiF5g0W
Sa39h8rFNhRR2coyAgAcsfbji4V2c8TYZ00xaEeh7ZevKzhZX1bFTdoTb3uc/w6SdqyiJK0hhvVm
0md6C33IAzx/JWluMKqJcFbTX6Atet6kg0vZAUL1l2Cb0YipDyUbGd5bdDqsQiAiVvlkjgN6jOG2
jWbvSCxsKvwXvhtcOx+x7wVjsJykjM1Tvr1D+ghbEPSyP4gFVQ6VxU2qshUa7afJvwoMVsoUjVku
/8dxwcksOt2C2mMMZV6rzoOfgIZCTcXKPUdUT9Vaa9YIQQjnOPusMNI72Mzi6YrlFywHIhAlcJlD
3UM1sdXk0/AVx5n64IlDPFVYxtDkUHknIO2DeJ9SuUiyd6R0lXiVAbSofvEobBJ/eQuVopxIXgKf
PMy2s9uWvjEgIzjoU20My28Cv6aJ7BBziMx5Y+yfCauEZrcf/+aVkXmhM/WCJPYNZwje2PCJds8S
eIWtppUko8rdVDqQUwcrQY+m0Ilb+WQXkrivsglU7U272dfbaXjaK4li5qoH9GjKqjWfvSz2p15h
xhjBpMNx5WrZ2CzShkimXX1BeUR6E93Nm2wzNK99xkKfHtvtqX+wHbsA7pu/EHGWFwrVLhggQSYM
UmXPabEsD3c13oEVFFmabrpEYUVyDPdiHDq/7OpsJe2d+g98Y5XUmDvyHarjQZ09IERAy+HAXw+h
oGAoCFP8R0Cvsh4K0SBusVQzPqEw17xpy0OSHpjn4Nm5FwpHocZhYgP7JQIX6jDleP9LzfEUstqd
elkfjWf4A/TH0pByT0ASrc0q7tgBqNfsvu42i8Gtm86j1iM5i2gpRaMYUv9FMT7aWxxPn617yYrb
1lTxD4r2YBsQyc2ce9eVdSTOix8mNl6EzeRvxmIPdtLT34CswvKcQ74GSrzTrIKsDtBuxrYFvtlN
bZ0Ejn6cH0+PIwBL14uHCUaHRfABzhQ9pKUImFKQYH6/gzOIx7u0cQt7kw26JkccnAf7rgE9E6nw
wQbVWKrKRYJi1HMIluTcCUQe062JY0RN5mb0epdRl6EbxMNQ1+AbZAOoVCrXWMaPcaPMrmQtm41E
VnjENvubj8VsHHfHXwES5lBIm3qTxLJadCDLCsayrx2exjl4VSp57g7j67ICOnYwA6upNLYolp7k
X0cxzbiZINQbuLhWYaPJzJgZfU2YStgD6AGJBaKYke5N3dMMEJztCapLSv0Hr9ZOfJ5IRtjsmHaG
0yLTjv8Ocw9PfUxqvO6fJ22b/UQaefejsaJqeBmtLqV0l006y7IjtbQYqMJEmpBL3QCA3vjrIjwN
vdgoEe0mF6QQLZe9F2ysfvTYVb+kBXlQFTjSnRiqTnh778Fo8vt3gCJrqlWZvI+Z0q9ongi0lIG0
V3fCySvaL0j0lSPzoNGOOu2CMykBbuHvM82zPquXsZjyB1OYrlJyqk7cn8wcoLXR5DhctHTCnikH
vY5wWk+Z9DgVgTrVJhtB5R8NPbpKNDNZ90IQ97Cy8xS6FVjVrjVmKDqzSwub6PQrKcuVIMgI+9eC
YKjwYwnRAE2Xre7yW1FwykNgdeTna/85h2Q2cFcYz2OgMgOXEco69olQInLpF4B6M6LexJg4SC/y
2GyhzOzV2O6kZJWHG55CHyV2zVNju0615MgIy+dTuH76nTa8RjWXwXoR88sPw70zEb2SWewKPEYV
B3ThaaDYs4ks+VQtOssrJ91APEm/DvWrvAvA1Q9gumbYoqjEL4iDzF4iWiVXu7Yg1U2QicXhQ9FA
VKyX6qkzM2WC4HnhVRUlnvgbGbnPTKFO1xw0EYWNWhbfC8faxt2qAOTB3/+CyZb3mV5OsB6LWyFk
lmgX2W7IU4z/R7SuTgNex27XSY/PjC2MdCU/0PdVTLjtJVgcfwRMotcThO1symRfOeAHxH9i7zgX
CWAzUjpXAxz8oqx7HhshwFcPUnDtqJssyeHpN7K8OWPKGsriHdmVX5HvP6BRxnk5SUXsKbvVVD1S
NX1L6xRfo0noQt+NvR77h2PUE1NxqteYWU9Fh5DdNhtwdX9ndhA67BAL/IBLQXdaDby3J9/zbEFf
jD+jQtnA/WmHELikUj7geTlKNTxDbecXRNZ4Tw3rqHPGH1yfm8WI/1bUxzC1gm/N1ZsNLs+bG6wC
4bQmE188zZVqu/iMn6ksX1T9CuKXYBCGVVqpCAjwL3IlscyF5s/m/llV0iYvP5JXdK1SLDWh4ULc
nNJjjLXLj3SA2NMo9zJsgcP+wqmZgn7xkRALYHlHzWabH8u5OKrEd0PvAAQRRYtiNh1FW+1zaYXd
0TgF1FmfN8O0YfBZ/EMkw04fqEXknx4wQKlUcuSfpZae7c8+BuB0uxzqdzJ0zfDGJ1ODUjVgHv2F
s26v4u3ZaHp2y36zCDgii/mr8gnlu+DxXsLmKy5sHawXjKTbaltcU/nyJZz58LLv1DxJ+E+XNIT2
hQI7ALXv/vjQNez6kiIMaNJCFNsIZeSFm2ted2Bsmo0y6tdK00lJp7Byplpe0+QxcwtJGyoiOsqu
e1P+nr0DMl6cm6pKhed1H491FrTiIEA+pcGOul9scdKQ8iK8ElhAbzjeYI3UNIHYJiBC/sJDj8jW
4MgNqAd4fDNL0n0tft7XpFUtjm06rLxdQwlSSBJCtHotverTVqmnAQ7H9b9CXxUJ9N7f+yqOGwnN
AbncE2coYBIlBLUgcnJIFi9kh2AFP4wF93cgr6iobO/IsDHedwzU/BVRluh1I0oBK4g83J3WGFz9
wvLPH/7kIeRQ8GMcr/4Z/eEQE+FwCKgGv09oGpc9kaqP0V1ev51YkH+4BDoJWsX0jpum6tz+beIA
it6gC9sU3IWNxPdwsDop2e5cbeF75FyCJKs6nk1J/HQRKhwyYvb82Cj7pMmLqwdFL7WOZ6aiL4OX
jhYPNlcSv5TTwNaOkHEcciovkyuiuQeG/FBMVkl36woW2A//36/G9dapQIjzZySvHI1VDX5JjcDn
leyUwI44+36aVq8YFQ72TbJSvNju2pfTr8fsSowtxy9VHrO5l+KoQPEXr+E4pjoj0oA4h5etTlVD
bh6TRJLv34Kb+moFR9YK7Z3ghvrspueSu0AZuZLia+VN5TeRqmaIHYFM7ZXx8CNFx8P38LnCcenT
2sz137dVB7K7odwdJ3h5ZfyDSht2ES3LASRO/PJpY86SF/aJfavlPJPAmybUpIRCgH1SnkZ02cfp
s1MhMfSj/rwxLxJ9DWO9b1wLyI53O8O7muRcwTY524a2gIUobO6hZDX7Cd161sOxA1aDXEhmYNbo
jEF2EYmye2X8+8c9e0NRbXS1BOykQB3mr/Au205WHM2U4Dxv6ux0EEPtSMlZ3yAdU8O6GZzM/n2l
iallWCK11STyPxSbtGiCcgcEbzs1DYd54LS+gXvTnMlj6uv7wJZ6tuv3ehyzJwP1lqclRNAHoK+T
pvnObOaARpO/AVb1ucRlqwT8O7sVIsUVF4KOfnMwtJIVBCXGDn9ajYMFjBWW8zYLnGEuKynmQH6G
mRWE7Fx340lR2L8lWZuCangmZymrtz7hzyh9QIjM8/0FXEvYgiB3z83lBR40DzIhshmvCrezpEec
PZ46NOtHlcqP5AkosQHLJ/mdYxXLcjqDF7d264uD1jw3cCagDLXY8f1+WMMXZVXscxdhPE3fhbRt
b/0bRxj2DWsIUOLWJgWqIbZ3mf2M79JQ5MeR55O/fb1Gl6aBKHQd7xKgR16daLaiAri++HxGxM2n
5o0I6s/H+Pzih7MtjJNn4c1ObTeMVmq6Lqm/2WwapGzmJ+RbrBfIJLCgTelWm9gokI3ycL4moRA9
CWzZhQjkWwBIev8UxZ2IVEnpxdMTVVmJ/8ynh5l1FFnzIMqNLraeXaPSgKtm13Eh/S8BIaqqaagX
E4JrlGl81C0U8bZ3MOi9B2Hj8SC/VZ9Tm18o/jwssvcmn3DlXhbXS7UTp9DVVXBGcjTlZ2xTuo/G
30yfvUrXchHyJ4BoeK8GsmgLhmncoAix7lKYRT9nNgc3eE198K+Qk65aoPweky/y1bA7P35V20/G
OAI6IQqdNie+JUalKgokQqBZ1+5cigttGVKK+cK/8513SU+HOlvXOgYka66YzF7/Nu7UFQFKXr0I
Dqn/pR5O0inEBYOwAfaOHTpUvdhriFPpzbjfwmC6CUpjBNbFFEj1/t6w1jJ46H5NOF6R0lGAP7/E
rSito98Vd8QWZsNZwLVlUMbHQOFXDmkoSrmROhoOqHl3ecNP5rj6ebTjgSB0RfZ+oPb5NCXNAmGY
taRd70EmUsoyTZz3GwlXJPGe3vQFXzcP3/jASoYjPfASbzkCaHNwbQjcKBAyzjqwvJL+L7T4wTc1
Spa+28fBhg7Vw85fBIwPlX09MqqS0E4ZpnnQihjduG1OJnBPFgjz8GSUuUKMF+PuhudEg4Cd0aDz
IaCXPDxiAsXgY6WhXsWoErFkc0LKKr0tu94KdVASBrwkvPmtZSzUDxf0LqSfQ7DV6MHZgH4johzW
y4g+uQu13ZTB+j37jZXnZU58bk9kDJxzQLcZr3HWfEYu3Dxn2wzsSwTKThHqO4L5OrYy+oNcAVoq
Wsimm+bbB8GIYeyLOk0ILvenNwEuwis117CV/ejiPquVpBbHXsUpa2m12cNr1eav/yUyWcNw+Vv6
p2EG/V1dDa/P3TE/7q1JBluujiIVhrbunk5VomnEsrGXS6vbrXJZDvI11PG0IelbKL6wBp6hy0F0
5iPr/rgOb1ucF/279M6ueA14pY7gvriDF7nG9rdAFZMpNd8cgXW3D8TPrqKv9lz8aERyZN4v63ur
Ts9OhVmugLkghHbPFKJYr0HW92FTcI6AcB6GNkQxW6/3JUrvpFJH9tgCAupQp4qGGA1xq0QdShQ7
wats164+OZ6PUZp8i8tyjubv3iIuAmEygfbM7uYLcD/1gJ5FdB20SDBBxUA+UFxX1xgu1w7PRbVG
2AmjncwQ5qMCrRfRwiGzT/NbNGpcgOxezDjJM1NF//jMEaSwR2DP4Z7Hzdz2IzxsOxetj2o4GQJf
oD2RMhLAocV8k/On3j14YL0Ou7dBLyPL3LmRWzZ4+oTvt6cdKW4atKUZv2nna7tGizgMWruc6ymD
JVc50YUGA3HCq/3iH+LXx19p0M2s4J7/JxT1JkhlhBzrFlXD8KikWyZp87pYFPVqtRX0Lg+0WGsr
/n6xeC1B6/XHmH3dkVdpImgmr21bFyx4kUIG7Ew6hufQbMl8Vxq1IZDoylbuoTNHdyAjDI6HuN8q
aaVtcn9SW8L3LunFuxjvbtlkSfaDG7ExlzS++cuqMtbJMl33UZ/Zpe/eVU428DIVSiOEb1AB/JUl
nwbdO1kaQLZjjKRpWv/kevoSkihY0oTo8x1U9bgNQEMXHew0r1223TT3HumyaqUCY420s61BDNVK
K0U5s11QmOUxQJU4WWtDnHG9MBDvhmH3/EMPFavCMunSmk1tg8lYovaMrCRRkl7uWnn95haPxocv
GwykmlZlKRzGtDndKEJfxLCbK5HxjYS1wK6XgabOOyZ3EDrdXpb6vtlSadMBCF0s1rW+TKotj5gP
YGavASAhyk0GbursXEH5ssL0NOXOS3rj0B2rFX3OoGziLOOAU39mrlfCS7qHJYd9Eg2jkXKwGqy1
Uct1UtXb4RFgx7RhdMAug8yzS3/3xf+UhhcSzOlQgDZFemPMA2PUzvZaDBidaz0puZrxJF1aEQ/n
Tra+ZamjUvIAuuSOYqB+EwXpHqj8IbkV/+xpP+MgCRXtqoNAe3TIzl7FHE17Ae+1Wb7uS3B8VapE
8etiWiuFzn7bKxgHNg7Ih8RfUyB7n6iUxvIp7/t9MygmAXfTH7B7o3E9blJgH4DZ5u1B2CNKYS05
HGunZI79lh4c81iBlxkTt2+xAxEJBME1W8mPYbdwGEFZBtyI6hZCYBmFTS2zgnD1Asm623dVar6J
fOZpY9ehjffHc5j9ivvv75HVrVuIkIRG+HGqBoXxeTJr1GNq/VyXjXchETk4zhGZiznCXko+lc2B
5h6MJLf+vXuZvbR5wp0qg1306wxq92qoiWIXx4KYhaehnZuxXk7DnpMPw237mezI2nHGtehMECxU
wZK0/uJ12m00mS9/+w4taZbIB763BANkEJugiQjBgdTgJ8w0hwQd48FNGVcH90Zc/OBasbL8JFbI
AMqwsVlBR6+quP46lKMAON7DECoRakenyGvwzmpZzQ9CpkLEwO0sM8uUVl4vdKhKmqPdqdPgWbBp
gnYu71hH531XzLOMfN8SppNZZsTv0+GyupugqmwZkbc//TUsM/LoClhfo3Kzpf+4OEVRpFA+wwi2
rli+CJOpcMEM5WVU300x/Fqy0aJ+s6q4Kv8sALlmfmGuBn53nefIcRD6CFR4T6609AAO5nzWS+W/
3sFj0TNhLnyxAnbRwbCV2TOfENNykMC9rIsFE36LFT3muDqNROhYJIp/YVtey+iMCbhnvTHtUbm3
CWijcJoTyUvN7KFmTTTxikeEKDtruYpLpmDwwm7Ba14DyR/gn+XHFK25MB/zSTvyRnOzXikwAtNJ
zzexijfkY3jIF72g+5grcqc39tG5c5+E2G2IsOi3Ci9ONZHnN5UsBGtlLpHDmq/NFrxqHCyjvwiQ
V0B77S1SbmAltEW4eRd9jUugPujo+sMgbctBchgMPLYi058ph9+czN76zDxPINPGpSwArVboHQLJ
vt21dnBB92WpHuu1oDw7ZSCXYWOekakQQNXjhBHp5Z3As5/Vcv/JR2vaaN4MC+C8HqApsnc4FkPa
hIsgApE85qaBOAHzIPpuvBg5NL9qUsIFRyW6s+IA7Ho/dk/VoCOtX3ck00AvuAgXTRyzaqMFr6Do
Np5Dx0X+vTbP8S4HeMg8ISGyF/503kLSpWxTNH8d1yQwGuVxq2w8vr4UiuHVBQVGKbWZBrNJ5g9z
hjGDfxq00dU9YfOMEN99cdESVh9AqlYrGfhmpJG1a/He08swZEB7eCZhWylt4Px4kxYtnix/3y/p
b8Ug5Wa2++28wB8ld1sBghjSbd4lGSqzRURVqKZQXVPLLbR75ReXbhJZ2C1gxiO+YXbLQ48SXEd1
moEoXHHVF+Ft2F6ReVJCP/uhBJTSVB7EEEgSKlfbfBmwWsRLdxlyUXvZIKJOBs10xPNi9Zyn4lYC
XeMOO22xF51dXv4urbxcVDyoj9WBB5UyBwP4lGJyfcRcgRAQrIOXWtnTeaufRcA8AfP9BFIstuHx
YfD7wR6OaUNXkM+x8Fk9L/MVbAK5PkjIpL4Tw+FuaAkSSrGKVT6LdrdvfQW6DcuN/nBlKYAMMbLD
S63rYUR4UVOQTcEdeb2fOKkqFx+LCiYGwd0X4McUKZRDHthZ7LT1C+l7l/g213JmbsryyI6Vopif
SUM6BS/9m8A1hAqIKKFjDBaSUwFG2uslyL2vjXvaAV634H0xqN4Nn2d2Pr6wkarNM52/Fw6+3cu3
V/u0/QwwTJCL3aF66zToE/fNPkMw/jxFviXLuU5L9fq9bLXSY5WOGVIqzmAhyg5jlq54Di1PxNN6
fO9CE3D7+WBC5OE++nCig5YI8QD3BhFL/g+jIK886pUoZgZqHix2SY6ld2rFPlhvFN3kn6XfTUCz
at7G7fxV1EUyNj1ZOlZBGJYrntdHPvRgirc3XnnOVK5LW3P0xwdx3QlxJvGnpsbX3T4+e0xaHFAU
yGDTLXVGyMe103kD9p2ck62dcmuoS8gqXz1XNlTrtIzL+j3H83Ak0k6CWNQBC+kIzJOhGI48nB9n
Mttj8oQwK716v5IcA1B/xll2XXdanoWPdqisvwO4lM6ZLivlSKofRSEIA+scx+JI2QNo8FIXHjOH
CtGl3S1SzdZFeNx5H6n9NaYoaVKgDSdZJrlyxgm+E2B9azfZoYXWeN1ybk+K2DfZ4RvbwAQlu3/b
C8EaupxmEIBL81MUe9r90Wq9STn4g+pPzTm84EdSSww6gXa7LAd7AKHpzNp0CRoQb13KlY22hO4z
VzxJGvoXpxd1qUYkxp8CtvlkaAdA0PiqOQKm8OpK6AT5Pg1PbNGG614IFDRfeDi7m36L+Lr2dQmQ
lVbH2nCxANImzF1ol67+C5ZYZgs5JboQG+31PAGZGs40hvip4kkk7rPzYJ5wQ15hhX7weT65qGOj
XcoLV3A6WjVKvbIrVWacV+Z+lrP+zNrzJP/Y+gI8WU+7ko6gJ+njrGGQz/KjjJ499RA9F1cayv5f
JqtJLWGsnNxAq8jhY7WbYuuYUjJ3WX6dSaOAoLHifxRQm7eNCygYu4DFlwKQ3br5sB4PnujNIRAu
9SdroLKpZJFXTtgRFbjvKuDltRnMXev78Ua7Q59FTV53dXqCl2ZGqVHyzgL9eBgLXponGVgP60Fr
+DuPDbjYJTFiQiWfZRWnN8JVAk2zHkdBLXcMX8UTSID3/6+H4Vx69zB0Y1DJgJEYn7Aebf8o1spV
pT8k1iubpHXiLG15OVuKRfZ++HlQxpXQlXZlCzkN7PCmqEC6MvWfX/V3Uyo5CHcQJvIP9Jj+iX8U
pIRBCdhMpM+UMgNiGE2D6MtWZFbmbWXRVFSlVksD6JwWaM7AZDM/WQGgjTYt5piTNotHoXy8BXmg
9gSY80BFRd4En+EtL5xcXh7qrT3ABlDxtCb6Nj1HAdg6O7dPk5zZriShlyetbfJ5deM1Qjd3ZQ9U
VTjexv0P8HtJiYeJ5Vu58/24i3sL458uEzZQNGaECq1dlg4dTzTouXlvxNi5TfHmLD0NHhKosguf
krpVtGAHzBmfHy+gBmuqEc0zo6YE8dYEzBCG7KikxwCoIRyWelXXxEbtF407LvVwKnTZrrbiPxwN
SLGCP9k38h9/Iny+7FgS/7fE6S7zFcFzBeDAl68VNimagPiNH0S/VzOK1DjxmfzfrYenueXbB8oZ
LOG3cewOEcLQS60DQN3N0QnngCK/RW98ckrZIoKZABh1ObQh/WdDTbb6BlnJ45AIp0LAvv9lS/b6
1p7lAV2ViSyOOx8vD6yBS9YHKFQrpjwMtCEFHBLMb0DyiegMwXcqBwA5XV0zhYvWC66ppBU7P+jB
JHTIRfgm9jbM6rDHh+srizbePdDM1GSLeYVjtUugXhFC1Fu8fd+qFpr1vd3Aac7k2eb+FKy9ur+C
3T0rdLTkF/qHzJUEdypvGicHk9m2Ru1l6HcDMjIt/pUvH32SRbYLHajeqTn8brjWqhPysOdtfDf6
v2U5/eQFDaFXSIVkuxCoLjYdhQAJz6rBWFwR9seFeud77KM5frjI726+P8S/4Qg6jZTX/Me/OUMx
ttHJyXKjetlHszH4bS9k72RcpbekhzQsxp6jPxbWtTVwcQrCLuond7tuTFh0RiQ6HUiA7FDzLNx+
Y+TRDlhVCeWzuZQ1+OU4B0xSrf/1JOKHTJD1AdV2P1eI7bgIObKIjjOM5/vbogHr36HJwhsuE/bw
xUNORLh2M4BJIJ7cMWX8p3R0LgnK1t46jUH5rT3y8dhCDd7/ZHwZtjWEk9lCAdxxSAsNSmCbBONu
cGednqV+ftFRG4gOPLlXf9qeqE0VcRtXCyLtxkgN1Syjx7MvitfkVJD/2SF1phc1Yqiz/9iMcIGy
vrZFQHktw5k3C5Qk1fSou5q9KTkuXkKJjIhMnQ0J+Rz+YHPuE4hIq9oQ36RLcDkH/w2KFxvbzGIh
9J4UxaHK3sv77u194x/ahEzevC3c0FsMh7t9zh9Chj1o9cEMLr07I17MuAZK5sa61DBs6rV22ESu
r1DwLBlsRj+iq2LEeVLGNvB1LU/fzj1VaPAiQw6Gwm/i7RAIYSSoe4WhCsQGkxdUOG6Kdf5mn4KS
5FKK5zGA8DwuRlH9ly3nv9RCrJUvH29b1r8Xo5qn6P6Aydhc7oKLSLKOknqmHkIVDd7X+1sK2e7M
J0pkK9MfT/cTs3Qd7b85+P9ZBT9i7kTe7WCpZiOy/V987VyZQoHGCEwtGekzzZJPs31wSb6R0GDM
17tQB8oSViyqbe9x7W2ieQ7Z8PX6BMBmK5TrjAekUHPY0EV3rZAxwPCgTdfRqPXSpt17Dd78czCU
mugpdq7X8oQc5mO318O68ILeH4rW1nF5DyMyGY4uF6BKUpyPw52xEN9TYlYp1YgBU8AkvrZ/VPsx
C8GppKAM4I3Q+litrEs5kkBoUvrEZrJ6sC2htcFgPYZD6qP1+Vcy2UJe/e/15ARStLGznQUoBtWV
uX15OdU7YdZAu6klgmdyZOMAS3eHxJApDGm5qY6boXawIjkN9VWSFepNT5iGQx8nQs7Q9PMSwOPa
sehP/Ya5NCcmaUuIV/sT9ZlmU/ThOEI/V6DmSBy6V39Tzgdl9GiTSkhahnx16zv4yOP0LohL22F3
9Z8vrKM+4+hTXt1eWqScvp6sD39cemVqoHUaSCck4XSfMkLvnl9bdxj0US/H8gd1FGw9OetZBaCJ
h1Gf0GBupruX6dwMWP6PaGxBWL7VY76aRS5+xItUEXKhDA7zHb78O6fFF85QMUs0WPPgUWLGnStd
w1TrNmI6lIoEj7TV9wF4PeXsHZqPu20+5QkZmSLB9h3lFj7LcfAjMRDBP8y3TjmUD+X5wTs4r7wn
nVT3aK/FkfGT9I0DXa/S78ON0o3wdAP9RogTJHa8cSvVQ42icgroaw3FBhBaGRmYxB8YVzcp3lVQ
k5oUW8xI6vSLfIbw1NPwstvNEyvOomQswnS/WupLCLjOl1ENCiXtXo2lLkCK6+opiJA4dOZ3k26u
l2ONC5cSNKjjoubH7dYQZXRhCFYQDJ52nbv3Hbtyr4gdymlYJZ2QVzou0SR2ofGMivLKAvWRSjjU
1vbBRJiMXYpdTHwQFjxDVgWMKMMduQI5Y4w/SCX7N3/kdFxR3kEeROMcY/V8KhysBUFVEkL7ilFf
LLQK/QTL06DyV5uUCvNQ+o1wm2VonXTTAPRhSQjiXFQjZNJ3XeYkhs9ci7EPs4qNJ+HZknNFcOtE
eyUMzoesGg2Ly/PUXd8aRSSIbfQTeuwqOkf9oBxZ2VhBZYk509nTmApCMIqrrDXnH+SKFsynhbWC
Ykl849ZhlNsdW4eLVIuOcaTXBa64Jf0ST+8p6ZtCKhFspNJMpkGHie95+bpgdAsY2+Xpr343nYQd
3O2Yafrrz+N8K5BFIgf/VA0m/F0CcEPoyqdK1RaR7yV0iKRqyJYkieDMwxWfxrF9tc4De6P2Z6Wc
F+UjIKjV3+OX2ofRIgDN+pelB7pTazlBvrAc7wKH8Dcuc4lc0Hi8eYA+hojVR5eqIud/026WYtYS
2DFmDy56oFHRlDj+I8JwJb1RtRLew7YrxPh09ohmTcKVtLLu9YsFTiG0zaipBjliqZBDNdEVFkD5
g2L8Em7EasOIuz8VsGWIR35VD0u6fLYKa8CUFrMVhD6ZfOGb2lSLuRd3e/u/7RbfqtOP0/0LEmTu
2OylMfDUWZcEGpfsWZ0ibeCqepuHeno/+jp69KBYC2FzyWsePiAXmx7GkCu205EZngIR95emFniG
bT0I+98zMJAVumVgbXBqB5VlmrKFGVW+VP+TbQVP2obuPR5t1/EZ/L4HDdWh/EoZjwYoCCmMbHJu
dYajbm9BW08OrWjM5czU0RBwR/qAcyZ8pDvRAIxVhw8cQ6qa+//QuD9fLvrj0jVSzqzPbC3ZpV8z
0DmCIr7E+4NNBZWNZnYW4AjExPd9xMVf4FAmyvOEWOhbGRBY8saDPHExCOjD5Rgs4RML2gEihjxa
m+ANqRzwAiUdOPvd+vnzuTRMwAmXVCnetdNpAv9JQNiDJCGPQT8o1fR6tnTZo8MtV6LRPgo0VJBh
CCjb2UvjPyMDB0sU6L2Wifc3JxMLwKqWsPfGCRSdrrX5uULm957EDl7xbnJlk9gy4kbLfmvkIS0N
iOIIac3pbb7JBKs0//QJNk9YpcbTsIp7zgeFSXkk7ZFacmrHGWrenrqrSAs9Cz9WuYXd/SSaBFDm
CNWqj7ZAFYL6f0HjgAg1zlTzgn+A+BsCm0p8bnGBEiydEj6VPZyzUSCkj86xb8YwNRcNKl4xtRaT
bIorcJAkVcdvz7r93STBVEbqAYvx8v5mVn65tRECSXFjPFDQcT2WDvnR4b3sFl30dw5nvSlGr/Vz
r7IJqsmkWJGjnCxNxUuPFV4EIIqJ5ENSh2sX4Nggf+3a73L7IbSrPsx9TMaxWNl9dCsbI+xw3awM
bDIeITequxdhHaEsDffCd8aCyi5GwFbf/iI63H41k0btwj5GdWqNJ8b+cl7UzPIyjEmeXP804k6D
mxSGzTJD5YyEepomA9rBnfaqxv9e6fbXARJivPby46hWIfjy4uuPaxI1gXzbdb8NuIMQJiuUpvC+
ijHVJ2HDeGoC56uu6dKOtThT4qKNvKSHY5mWFppZzTsOcSlPpvCs/kGtupiIutc2WnSKYG5ORFOr
z3GfLyxAABg/bfPA5/cEgcwcEGR2m2SBcH5gds9bHvAUvdasNlkXs7uGwx8vQ6FiY2i4uyAOllgQ
a2jboNxRdBXWVLek/jn75IHRTY171l4yS6NAERIaM0etxJnhASRlz20pEVWNIMt3YU8pylxejSSL
8HlcwAzx/SK6dortsmcjdrYgh3aY54ZV06JU1b2XltD8jGEgLKceMo3GvgO2ziokU4RYy90CX7LF
l+tY7u287u87kg5wqLe6+LkpqkhQcaKmPr1QWxmuTswINRXbE5SDTEwPk/KJ4/b2+UGFRHh1/n5L
4N/d2dZg7+pHAl2KOKa0AyTEYneXDcjhlNlvPbpvRC0NZ5+7gUPO9XeIYXscHx5yLcJJXyy8CEYY
GNzJzbYnXGU0BfwwaM8u2pb/rd/HrkUCyFiK0sxhjM8lINEvJlE3xASgfJPeKeozufjVRqwdkCJU
mY5kT1e36Jf+orYSdUaIlpiUQ4euUR+B0AN4Vs5o12Zi7f79AUPg30applVRi01RC4VX8QmfGjpf
ihtilVMpTeTW6JNhBZafGOnnwYzItzwZcgS/vIhMYoVXh5Brxds96i7DqhtggkvM8vTjceeTabAY
5HJwESFIKHKvDP1Fyw1PaZWUpIVAAAMLkYeOVlMq3BvpWT8+nHamcrzo+FmbaT9xTWnmRrjf2iYd
2OdZpODSnpkBROEzKPL2sHJDleChZztRsmWW4TTzO066HgZv4tq8gIpFAVH9y3kAikOv41qRIZsI
ecAzp5IA9R/da2uEq9sU9LZzeS+ZiMfdOBt91f3/mEEAro0myyOpRhcNuQP72XGy1pZMwi77Dc0t
bP33nMixvsCOoR5i1ofTOr1PCYNnDYKQCA2o0iaS0EpwyNE0pa7BeWfUdFfgC/TktEvw19Wtmled
1s+lkhBTX8vUIqzG3otbfLlaT8RBXTRmV7NguaN8y+sCYTIpFRVaTtcCehfQJqYTW21+5kKnzeTH
dDnWjO+hHhEvPJ4FQVhHpPZsP0Tmqsyu7SsqrpgTigmKEAYegVpm5S5IejFM0Ef8wE22jxWGWaPu
yKBl59hGYM/vxtnS+Tg04RV1//KNV5fg1LXY0NA/Oj60NCkApk6b+GnKiMY+wcaccBCQQr6dI1zw
dAppQ34Q8oEitlJtgw/vcYgeTc6OpS2iOl4xA6JruUZGjmo6xVoDQJhoWTxbJsh8Azj7xlWEEV2g
4yoI2TfVAlNXKfXvvVnMjafQwZ7K+EOvJtmbRY2/tkJnMbTd+k7IgiqTV3MDNT63IXSOIKNnjgpf
zp4LdU6nmyH8U7Q02IXx1QE3cZB5Aagoztuk54ZVE3Z2AFHghGMu4XYl/JlDgRRDvp/bidQhyXEq
/NGE59tbyy36WS+EuqD7bkuiyCwcZ1atLY6eAhNpsrUvlTrkwVSAg+yoMvNZuethOGy29sRa2cUn
VX1BdX3FEHZAhchcl9SsIcsy2sI8PKUBdUXzp96KZTcPXPUro+VYt07nnLpvfe7n8avU8F96EvV8
qp8nvfoi2L2Yz2kEN1UX8NSf0+SD5Jxn6QXKKBBW+8XTwupjz13ibfT2k6piviu/Z921MmCZYw0j
WuDfSS2xijPq9GBqziE12VApDw5BoJFonzv01iPY3wWDf0p6j5p/LAzbBJu1IzzmNKPGHhrhpAAM
zoprcSu8lXDv+60q6XIA03lRrr5Xbf40ATWWeMD3PO/D6nhaecYv2gsWGdWTADAp8cpbXSNh4C5w
iHyxce/uI3YGH/osRPTopd1Qidk24ocKEVF24lOj2w9XmTsn8w3AwI9k7g3GCotRplPSqTTapcDL
dbohl0ucrPBNeM+Eb7hn84ZqU7w7xYk/ke9PpVoAOX7WYLg9yxE8/AbsCdNkPzPgGzv8774AKMSj
YdRv2soSuW2imSbFlE0BorfeWyaQFjQk8GDML5Fc22ziDsU09o2SNsu1YFqJqLCK+3E7q/11VGvB
xPOs1xpJ0robVh0KN3yJBIH3is2SDQzO8X+3X8WQVoExMNwf9NvpHDNkMloDVknrRVHGct+dxSyb
/YUU8jQfcbbeOGA+qvYRyESoC2QbirVU0WaL8Ku1NDlL40RK4oPGs0DUPLVyAU+MGC/eKDm1Y4GX
yT3KkZazgt/jnzMDHKRwOaXpj1YiCV2diKnk6Z7vH7qYdlhZIHRJUl9gXGrF7zIsw8KbskBfNR+U
Xpmz75xDWtXwI3PrC1s6LL/zUIlIbbjZcgacufoWGPjlhKo9Pxx1B/5rOUECTYGmx3c6RYXqYx02
NTcb4BtxzIqtqgJjUJMWsCbJH/R2VsRG1ZTyFYv6ikWoo7iNxBeco4yKEZ/ozxQJNW0XsUhBfyhN
E1s7BKjOz0NM1DvQGuGPCq+TF03ptfUk0V0yqv/LN459q5QZ50sPwKc3f8M+l4AzE/PCrytJCC5W
kH+C/SQmKwDpQ6GnTIpKj4gMkVW+WR7+Ozx2w6esV10+5TliN1Xu5Q2o2Y8gBBXFVbLYxN/yw0vt
9fQBXyt8DfFpcFJ22zN/h2yTzfiljFPFNe4Er5mr+eTNaEHK71jdk6nqSkD5heXfw/7Kz2u9PFBU
icx+OBNzx+DWUXdf9L1oJRv7j/8kTwYlvhVWMwUphMLa+iU4Nqr5GAbwEeSVbLLX2l8zH0yN6ARv
C1LevJsEebKcG9H73TY1IGHYtchqEJ66wKuH3oFQSyk/nDYUjqx+Jz4Y80hB8EjWOpb6ClKdD2UZ
0jYqJ8Lmfq6AtAdNelw6cQT+THUvwnRpKHbqXVQnL7AkSOr32rotvt8ZYNl1uvbf9UaWTN3NKvI/
dmqvS8cnmqjHvvVN+tDLielaRlEsUadRTjNWZc0Sg/WVObmetcjxIiBDPdA4+rnCi4E4/szIB5Q/
T5zlsWs9Z455S3hLdWfDKhylb9/BLIm3zfDyDBuU70nrUkapWa0iq4D/BMRI9KvdSm2Xc6m2bzgU
FeJjaeQHBL31u3Cnkzrw4/qaG6DiFLRNqLawkOGTMdMPXoj8l62MDSEmpLlT+/jkVzYv46UfxTV5
taJB5KLeC0rxQ8zE0e1EnPVa76qaPD/JuwJ2tjprDYdpDccu8LgU298KenyCJ/qvnag2//neTnuH
SGXKPmyQ7hL1QwQ38VWSXnZ/PJhoqjCY9z+5J7+woRU04GsST9tZdcuETDiVZEOK3yC/KWPnZgNy
c5WU1LiCgZZt71uh77oMUaTNNlDo+6ce/61/P4KqL50w5m+yY9LCWKSLmyyqU/Vri+sFMzCaviAj
0Ju2Enj3J9Bc2Iyd11gdj9txusl3HmPxHyx07Nz6c12sA8vGt1Mg9GCU9IpKav/oag41muCjL1Zq
Ei4s5OootkUisBH/Vf5WswVWW/qoXEcjFJav+S2ix52WnAx/k9fVf0SHFjRaSqbbHWXb371ppdr2
h1tJzlaN9X0AVG+/MpyUJaORwtjtKtJ5kD9v7GGUf7/Iz3eGsm8LJOVNDV87ahX31yYsMQhaq0V4
ZdPnKdx/wVjTyk3FXUa2teixF4L+zg/moMaEeSzBpzMBe8Ka+tFrKJs7WDf7b6P0XDyJSfpwf7vS
3lAfYBsjzW+KmVWIXafqoVRqNYZKOrsbyV59eft+S0/fh+VGBjn0nxem1vfMThrguxMW3Rl8ewpW
byemCxKOfK7oV4xJ5NeQGO1me9UEaK4OCfBGtMG/D+LBB7ccAl12NmHj/EuQRkcYH7j+/POk6fWb
d1dUHZT7Eih9A2HETCcEuAijY5eZ9fphdVt7KSn99rdMojOm6C43r2uogxji+YQw2jLGhbGVLMqw
jC8tFgnBlnPZhsPcEHlJnVVl7hMHXyDpb67UKqmZwlM+Fazp/1iDSAZ8BOoHVB2x5/7P37yaNKhK
rM1e8twy70gK9RjbfXdCuvMvc80Q1Ajp0nRKHfEfcQova5FE90dZ8bzBWUT5roJDiFIAvA9Rl6mB
FuKu6FiGIX9XLel79Ikwko2IRepI0kPXvTxnvBwBJLLqNKe+cCNe9krdj7ZmO4GZWLLMN5h5iEyl
dbxo3Mi8ZfgvpDRP8WbKtrGd+XICW2m1B2dAjenx5Vw5aOoPAT3HMCffKtRkNkI6K2mYLQI1DKIf
CXM5gS/EPzVxXbQr2MIIkRW0oTsivUJj8gmbs0jqePsz2ohI70qO7MR6GNkGwgxblb1S1zPBYYxS
cgslVHm0Px/UcDrzSB7SJR+mnw9bgHzUq6WWzV9JHlKZ5SN/hB87k/YnUwf2nE8rV40BSqeGs+2N
yZYi8ReHzym3V/fxhexvjeEvswJYFN+0H61KBwTew0G2UOUklsi/rkRx9fwra7aYIf3Q9Fj4dbFu
V7y+STWtD/584gpmKuWZeA8PafEFTUu8QNcRZ8ap4u7Tzwnvp2LfWCFPfej1aLekDjP3RqY2ZWdh
GllscTiXgNDfQi35zoFYmdvIrjJTzXsSUMlba59/Zc/siPVpOpMwDBvo2cvSSF9K9YeKF53dqbDy
ZOByYHSNX49bK85m9OCiWwxbv72SDzmmSj8VW/Vi3ezld7pDsrhLhvv3vmtTz2BvzXx+bMb9T9Jd
qTmr4bwnNLRXyHlQ4YCf9Btfj05f/Dj0cOr3rRRxrR4pKSq2b2Y1O72F5yUKb5kuzHhc3H07VwAA
/BTq7Z1hgmHzZ4APiTfiTltt3yjxyhPku31UnliWYUxV16TAObkm+IkwVBfNDRqfVmUm6ftj6206
WVrlBv5r+B6oDvlB/kCKzAErf7VRliv7SGx0VfNrOlN1ISfkIqCD6OBH9SPPvgibQh1tYcNBv13k
dxovnKUVvBnM1FS0y/C+oubJe7j0WxrCMsxf7sB0Pj/Jl9k6PXaDqwygFDYD8EzVvE9g2b/7v9Eq
H3PYoBDZdBlhmisMR1rJ0YBnJnRH56bR2MtkjKpxKoeqXD/TK6SABc1uDTfzQZRP7zK7wYmFXfEL
hRK02IQl+ELkvBWD1cEvpqMQt1sYcZJq//HNe3kHg7m4dWxNHwkUDiFQyiIk0RaDxqZJ8UR59PKr
ul66uMrU60Twim3inUv+VgsijCDwx6UXzB22hxMYg/WlF13eq8nOEjbMApbmREFmcZFqLlaNKviV
Qq1SUdOFkYBOkEoPrExMim6+VAV9V2GtIQtGiyvlZ34V4ep7NvnvEvl1icZpQSoQ6MoqXwcONyh4
5zcPkHcioGEgcdcxb0YvbWfmy9NnRsF8ZsMYzTCosQtkqJN8Ked+bHfh9ExJUXPU4X0rDG1112Ay
vxLyFn6ETTpwr9kG9F2vrHJaVOa9oq5wgq+g65AflmFUTmls1Wh4jtO09z0GPlY0rNycqOQ15Rvy
AxEELLxwrFVaKRAxt+gpiBP0UEaULIUp+jt0SAQpTdfWlHX3g5zKVjdafx5eHPbgUqZSs4qI59LY
Lu6zMDXibnUPRFd9AIplVzzSZzhkaM3UpHqvrLL5LZJSlA4+H0Q2UPESM8M0+8Mx0E+0UUkTVd+1
bl+35wtyMp+KEJoLrNaek+F7HCZpjULpRq1KIDpnmRykwcWefdK7wzLiJSqbApghCEQATLs3Y9BI
Tj2kf0jwTPyyFXKLnEhOI4g0Wzdun2t2GEi+rlbyEGvIeYCoQXbhBiFPIhw2qiRMLpOoqR2Rffru
rYtznLlQ+B00SMPyzcWFfiqfVpPhbKUtkIhIgA+7ENn5WR7oNlOhzU7DBV1ig6tLjeRF+IYzSraf
2uQ29eMeBq/I3OIykcSfsLMzXP10GJTbUHHKqNu0GmJu8ukPYHISIm0XoumnGcoJcq4u3FNkNmxN
ST+uG4rQSTdgV+UTbT8y5y6bkRyIAxxXveTO38ANVk7zXjScvGEaeFXnEHbMw/q8DJhUR9D2qZI/
M9Vnmcn6db+q6x5DXKxWpzl8hwLjCXZVw2ruXiSHSQ4YAKP+tznDL2ezwJyU72MLu3MJQrNkRTNW
c19N66neIXF5R3+pbhfD/0BVfQyjFS4M0UAOlNG0G7NHy3Auu7c0WTsEM20C82yOpP1WKJ422n/q
cFpdYqNkr/WFMNfwB6Den3RYAzbGYTmy0RO0CIOT+TgXF9c4HlzNqClb5fKKkUHVmshYoeJQ9RWo
lRmBAxixVNWXHyaMJTAIQWYLS2chWykXAGdhXj4JbZYu44Y4iiiAOg8W9D6nLQttlCd96uHdJvBr
6d2UPpvj8kSMVcJjTOWMXU+Uv38g4l8DrQLExOfhe9kq8eGGBVl2fQTa50aQg20dDQzENBPsdPQh
41NTmAgaqvVSBoQlwEBUGQtSs3xIIYOGR6IKr8Cf6WefUfA6Rt5Wc82VHuWybDBU/HzYRLVWmDvI
QdfTw13NqbhO3sZTnyTkWOGMjtQAHii5A2ZrOfsWQlSsWZJBLudaCuL0pfMb8ZUgXFrW7q9+mOhz
32WgHaedWBBO9VpiYBXhsrO7u2zJCyVm4PCU8AcWLaqLm3VhT6uro/Sin3Uyti0RCu7DVx9Bu7i0
OHQhQ4u1iv2qlySs3LNt/KrwyfbtL9j5/1ccLomDIKm5Ru/FRxSrFEw/k9du/XnLRanZmgm3enzP
i1RKuqFwq6iyHLXEG4RCUtml5x+zqUxCiEVxLxlzkBvYaeoONt9YUTKb7XOuTbugjoedN38JBwTC
Jnxsiq/82boXShgQrHfPYSJ14y8NdUSnwFVgiKqNEnFCF0pxxAr8b6+iJEjktz/g2QLMCZNZles9
zvYNP6Sdc45iOaKmyx2QBc+ileR4TEODXtFak0eXi7mi8Qy+6IhA7t32INNYSmsusFL0zJyzbSr/
Iz1/9lKTQXQWnBI/tSCRElob0Z1+SfMk8IbS8gq5qTe+6G7EgF2+PitGfNuPUYsC8N6+O6BJ4LSc
xni2XXATl701E3sYDh2WCf2qLT8fJ2kG5i8qfypcKTV5+G6NAsZS4LHS70Z4CE9PDSNhievgb/aZ
g33PEAr31xmtBIDHGhlyAFAqSL4y19Pu2OLUDlduDGGLz0pPGn6cwvnKwVX1NhIPT4zLMSBTU5DD
JVaDhTmFxnpAYzbmAE11mr39lw+pbUfjl9bgZBeNJcQA5nrPH3O/74om5LvrzXmLMsp4GHar58ng
+8ijVHgMohd7ejD2QOJ8JX8Va4fXzXuDYqM3rWz8c/zH0DVek2k/TtpZ0Fdppi6DlI+vK8IWy68b
XRUEyEumHnN8HkuE4YrDf2wGTw+HqOEMNEUzjzCK6I2hntrwRtL2bMivFyNQ1POCRTx9O8o08G/p
QpEgIbveztSfOuIPM3sVJwJVoqqLw6LsmWqFrmbFKCpF+eHxfxKwd3P+vwvZW8Y/qg5dZSCLMbT4
Peux3waupI2ez1Fv592HiPGorDUMefo0w8lkxigk0RssTugbvGBz+Sb+tP+bixZI5EkACKSwja6F
v4ERlase1nbJkd244ugfJG7NF/xOZpSHbr8dUgAf0ZWI6q3FgiaY7oeuL0M/m4sSCBw5zQqCsW3V
n0dMCENJ4ZbHnDkkQ4mWDKtswWf+UHIrYBvxKdkV+VDmXFXPkXn/5NrVh3YVEx+0JMILmbKdlmjH
dCyfJf3r9FUbNl2qwTfmmma4T8W4VX0IlbseeG9WW/7jWyBFAFccO26QOPZecXh52sh/w/Lhoueo
DYarh+o7u8qnQ+menLv9chu5upmmF5ZvMoG/pFTyF2iH4i6HMnS/JhWcZfgIJkcPA7xqyjPc/B8O
W6g9fg9aSdHY31+5Q3ewGPwRq+PzxM3VKwf21kpDO8MZ9ZGbQaDO2FoEayWuIX4KbYAsMa2s2A5L
Lq462zb/98tvXBaEa8o/DM/phupdi2s6hprfWY8s2ofQN6UtrTULPNIvJJdW5XBx6uPL0sMbLqRH
qZr37Taz9HxtOnbgdZ3MCLiv55Bzxcf1Bm8iBnEms2wwgBGgyG2Q1gVX6maLEryVF/+xfyZ7kTf7
QHYD069wDyv+9fQb/FdA9Z8/fFttf4pe3LtJo/wHDHxsnnFGF5eGzTWNylCii63Vy9STLGWI8No2
s/cbyZaWhVDCWj6xx2jP2oC/S/ZOIFx8kqWrJ+yuiIAGZSXGLAKJU1Desm268tpoAzaeGD/u6Fgx
HbE/sem2+4gJxqUfXvFrJdw5LDZXcIlKzxZwo5IavtaeveNLA6X16WNQ4ISwxwVW0kbRp68FaAcX
sbxj3WgYV8lNqb/eWGStF071yaBYae4Qh3jKYnQrjV69c+vseV4ft/JqqkDsCHTW9Srkgu9ExRHg
CPluxYvXvEr05mXMIBriMZyxRyCPypzQtfkdR6xeNVwORiZ9PjWLrTM77mJfBuOZrper7JUJNu3s
kYkEkdlLVusBV0aYXpuSorpG8n6/acQS6Xjqbm9hyhDZnRFLHUNYAgL+kny3LSOfcno6h4Hzz4MG
vcrSHP2Sa7HeYCypNP2a34mK9amlAKw44nKhlsjwMk+SGdVlEYVFFvcslFLmYBLE71qG7Ft4AWOG
qIQZfS7RtJfBt2Zc88XkUD7mM4E3U6faI1ABM1GQN7HQrR8k5SJf0FrrBYqtopPU4KYHxnbDg9o1
5ujZ0V/hV8KQhomM7T3iULJh5B2/Fk/tS4cdgFvdzu10eTP24IpGAHw+hprokmy1XhbSD10v57y6
LKHjw7qCPP4ptM9ooGb41ywaDgdWwX9u+TMJDeRM+9zItKG8rpq8Mt0W/gpyZ0EvlcFSoFr19VQy
TP/ZmPe8MgOWdGbq9NuKQ5Akmq6YT2L5Rt6AR/BPtk5XG5TyaW52qt3vOOQ+fcam2SJ2GIL4c8LI
J/oDW0FWWq3cTwNEuoV1csgKip7KaROGaXntZHJ/IZNQgBtB0RWHDoYov9Y8nmWAlASTjfPs6/mO
9v2TZjHzSEbr476PrJn7be0uIGE73YLt3rZB3JOxiBHk3Hc2uSueF5+Vv84oWZ7lfXgTI4xYJEdz
46PsNk5DjZcH34lqYoXnO3lgkbWW2XEA6Q6tNXa0SXIh/YL7QDj+elsInLWoU35duLH0Cl94M/xt
nqF2orwrJ6t6N/P3cjgUKCCxtsd1yyKPzaUWM0cvOU9L0KaTgPbUAlQInPUUlh5NXQwLRKAm0RAs
JrBtXRG8fKgpmJIr6fwmTC7kDQ1OSCI+6deFvIyAnMGDzRRgpvoXPepafv0furHG4oxCegw27KF9
7iwbk7umKbTkzXVzie81PUP/21bOVbx5layR6YwiVBqP3sPYvwK888tYP4cDeQJSyRwKX0/TNRbs
WbSdYzAQF4Cf4f2ruSOCpWppiWEV/JGb9xdN6i1olOEk3bq35QWk7Bnj/S56rB2aAZjQsRS60CMo
CMOWQ3r2VleWaD+8cwbmkzk/UJFf+dyFMRFUmFkt3maFPdrsH6IZKcD33OvTZZs0IiFn6U+rM8Hh
RwZxOFnWgWmwiSS/zC9IS6KXed2rd5WotEhcvaqsEGdiWZALa39SUjJujWYopenTb2/7PTAZEV8y
EvWjXxnIO0xaqHIjL1ImbXFOfUdQO1BPjtoicMQu4cyDRHGJQ2OXwwoMXeVThgLdOpsQcEwwQMHt
t6UlAhYqPmYNbxPFQNl4Xu4eScL0a26SyZizkhTS4nwb7la9roMkSHvqQlV014hNo4MTCkh+0hVB
2HmySK7zrhRlEHo4/fpupnEkMgs0oui3u4cEzUIZofq27RY9SqR4cCBIp9vMv1kl1TN2iqkJEys4
vCqymsqRp2hGZ2LS/77PnBRW89LaOCndEYRAHUCFi+Rc+ChPCoGE3X5j1z1MLgcjyym2gZIoGRMH
K6opgrXLmc9NXILGqiXADyViy9r7BAgmkT3F1px3t4R4xTlEvbAfQ6BjHTlBeXJlO4Eq9COLIJ04
AVhXWZavewyzFkYD5PqNA2ZBhDWD6gmLBdbUZtgOSQgSwpuyjOF5byw6bif1/aMKB29AYzEwiZCx
W2qRc7aFMtNIF4+vPgeWxloLcOXVjG7KoxtahgK42s/XWFCij3D/NMBJ/c3bPqPSrdAVFhsOaVqO
59WFq/5ix1Mq+2fvrNrrfFJNG3vUppW7xK0wKRzLX6tx7T1PGRl1Z3HP6D9pWDEWTNNXjS8AZGGF
1olZvJQtIMoZOOsMR2jjEu3VjlKEt0yN4qg9uK9WSqTssALwUyT0MvNSOIsyX9e7RKUwpkxztQA/
RwVYGF3Vl/iMGYg2owp3bAfh6xtFcLms2FOEXbamfpVSnZdAyDSE/ud8fZTgSdLTwcgE0IOSu7Z1
K632JoNGSYQbd08zja6rYNXTUrd/YfbhVxrQ3s+PGf0QPOVfe/Nkt5XhyxlHzWYOakxhB4ubBh9B
COfK5O18njXaQHLeRX5JvNrx4JFYsbS5IZ5ggZALphfTKi/0ugPvepe96EBisCsyZF/2I8V7KJCj
xbmzHBCd2QS4vRX8XzKhZrTLIK/dnWYsGZOrKnbfmVoKx8vLH/VcI49TZs+EtdaZm7BAkkQvp4eD
32tZnKneBzZ2w0k59j5ZytwYMCE6F/FAYQ7qQ40VPVQ3CoFNMqsfHJcLvXm4kqSWIUOCW7Jeo3/K
MrMOjPPL6XtczB/UCfvPJBJjsoV1owBuMGCN1bJfDQD+yZ3FuSmpyRTvNSGnuz3iOIkjGhYcW1W4
Ze86FUurBlLni6+//byIGUSGT5JXHdGXQzu9dzIGcc/mxVb2qBRtAnPSrqE7ljjttzma28wKmSmI
I2SrSKwTaVnrdmdvr6VVTz79wdlksAk+nduDsdybLOkVVeq2RbPz8yCBF5HIeecc4PA0SpnZMUPv
YP9mhPr2Bi5126rWJJiADJ899bA7+q8NHmRoh+FOtIwM9Vj54Y3h51KVDl6MpdpjGowh0li7puPT
RnN3DDvRZVO4YNLQf0Q3TOdOOF3qgma5RV1iC2H7LixnqvDnxMzorew0zM7UyrVFH/9o/Z9h9tzH
C6S6O+bs7cVuaPp5Ln7WQa3SinFXYuUIS9bLeY2We/Pj44iyNu4TMXOPgSSnJnCKb+GWBCoAssOw
IceDl0YgZd5aSCNTnnmClLAg/4LQCHThrFelBuZLh6zMe2UMbVqmMHM4S3Ffh7BJs+OY2+AmFtzB
YmKOf9LH76RzJvX3OVLAC6ee8oQB8aGdfXeiarkjqOpASRt6p3at8vX4vU8kvJUnvQ6nV5ewrLpq
juSVkUXU81ITH3yfNJCgYb2bu02LYcUiYgLse0yLtnF3LSHFxuo1RR8qbRTS9xDAm3SmjDFEeUeW
EDCRIxs/w6f9toD9OV9DybWx8m3rkeziBthLIcoFsvegLz1obz4GgizdkguzlEwpTXX7MLzQga0G
NFV3dRisi42qnRmxZe9Bt50piE9X8OSsDmnEbH+OrQIZuCupE50/sIvMdQBtrJZn56JZhrWogIDW
tU5dYg/m1impD1PBwxc/rXZ1XH2bSUrLZOi6z3J5F8eQSfpUxNjAR5YBync7hk6ZZUJnSFIhcMH0
LnqRefEf5LyhV4L5YiM5qhVosng3ZtjIZFFNBzWN/opUZzHbmAdO2SYDtQdDhyNE1bRQIkrW3Ghg
9LGllxuj+N3sd0cJxLCK5dJnbnw3Lv02FRf0aLVHTwrcQposnru2v6VIgCCoj1z0FimVobNdGGlw
pkzDqYuMtr3DFnd043xC8qHJEYs+cssXYZOo8oOz+kKJCHo2rybWyhGYFO/O/iplF80wEKrPy4Lz
9uxBhqSlJRxHKQNaZIsIx6YlVapygOfPgxhto5Q4iO/P1N8uYZSW/AKC+AGs8XxXoIcXOeOB8X6q
57Yc4WZ6Gi1ojn3j93wgzS2UnaNlTtlZORMjubfe44CuLHYYeK33GaXdBlYZ6MimwzLYHcAK08MK
S6DRDJTKAq7G29tgpEVrd4BhljzVgHiofEKkE94eTiBWHfcBgRwldpa9JUD6H1ByqNhNZN/L8Ywm
K9Yk+Iyw3+QDMKroXVagzztAr/OXieF6k7xpHogcCSC5+f+Kn1iWM9FqwBR2Nt/ZIoWlV1WjaSub
B3SLSJLwuQayvQkDo0oowqK2mjYLfE2IJUPa9c2Xihv1pOC3fKcNKTpxAuv13UZvsxWS+cqQWwJj
aqxGqX9dFJIAgRZqj5xSOXsTWYzHhmyVcl+XA5qVRbQDg6BYxnuma0CMceqiBK7BQ75A5jTXovrX
5SdJoxla7S7DBl2R08LEiPVMu8shgnvKcD38J/4NFmsUClL8+AnwgMPkjZXZE/qhBe6jf1F8lDEe
eOfaM9Rqmy4yqCP2mveDUJmWLz83lEttf7c4zhtLF98f4e6nbw5MD6P+7Ae7EKs4tCwmYMU1Dukr
W7Rvt+KbczxILyLWYOCU48sG8EBONBvgKjkc930XZ3SPtltbm2I1Dbr9ajoyVvjyV2+4EGRLFd0W
Gm8ng/lgE5qZPJrw/c09r4+JQ8DZ5+OTE0UyXKVjy5f+e1eCf/QHbyLhvP66I+wJQBMcymcdiw3b
9dw4JncPJt6Cqw2Rnh9Y+LkTXW30mj1Z3EYD/TiWFgetsDGb+8AT751CdVv4mep8StlJjJehQQjV
5YK2CV64lGM17kPtJ65tQw5HUpQVNyPmbDHBJ+RYtN/uq3AJp3XzlLaIEptIL4bd9rs5u8608IVj
G0/aL6124qafNxrkYMuvr81+mB6zc65LFFrhcOiPHuJzULLdnjiQ0bLji57EbXBub/K5rFL/MBqN
rtD6dubqoDcnLQXHAOM8f4d4Mc7bdAbuMGRMUx4DJjhpmvQb41oqQSzBdiVM/Li06eUXtCaqqg4F
hjeIz++3QDTJSMEgiCnrhtJY8eUsWPfar+bw7pQqNwpm03yRj0SPspwjom1PMSRibVaxbiTR+zCB
IRlFkXCen9163VJowhsKcM2iQJAuEaDRiIqQ1Kg4BetTQcwhQ1XXiUASKSanGcO0QeJjyU4xQHYw
bbU7/3MgbuviJAk9Dp40ccFVL0GSExNqNWDPEKJ1S3yTUKcK2H58YTiYUBSSKjS+bh7DD72zu617
wI2MM2BJLgcYhZcymb5A9J3oEU3HzsbQPJqQXLoCF9sBAWq7iL3BHY0t7mreNic7uiKYDv1omUpe
GAKfkkEsuWLUF6sr5DJ6MycnAurLd60PDi9fT/QWtqu3UGvJXFlTIcKDDvXsO7FDGoZU28uSMEon
xE7jbnP8v8+93T6evexxON4H0mO76bcieqd3jf2qlowUg02BYXiXjc/Gq5ohUdZcWnHhJw8c+h3t
BtlvB685YCumqvEmmVXd8qg4rHOgTFGXk7/zrbjHMtugw1fwqUKdDAuA9l89wyB0ywDJUyMoihBx
dpWc6FR6JqvkYc+k7J/szUAwtaAka3MzR450yCbsLtRR6O9IZNIDkwkAXrXvGQTiN2+mIIYedS5p
hK7BwgZaerEOemqJL6nLlyK5jOQDW07SrKs1bxJ9GaZ1oAUMF7QBB1nKsANqaCwBARrYKNOLrrYS
DIfKQKWctK3xAAvG3eQVGCaACEcPlLe+nRLTqFt89ZPJmdQUSrUnRSB4YyFnjM/cC+M8f2QY8fzF
5rBUgo7bp5bgiU9wW5Pb6b08gYFqeChhBLeULfFvov4hkUFM6oYar6SebrwUJoOKc5In1yZPt278
iCT0+yBwgxpi2e0BSlRWuX8qFI9p+p4GwfcuxqDNAEYeUVWPcFtTiQ+0NeZ23J8jyYOoW77yHsq/
/H++rOeKhB+LgcK6hGUIib6NgxKeCHrGKGavTwVx1S9uqV9RveVnL5c6y58kZwLvJzuaUtUmHcKV
I5HbeZjI0h7L8T7edxf4OTBQrGSshBVmbp0I8weanVvtmCR8KGf48aL16RCXzUx4OCAv6EdWj+1Q
sQGbsyuzWbcS2XYkDD9Jxzl5h5+s2tmnHcHYrEpnglKa+lCDGkHgI3di/tby1jNU2JNnZftM5kyl
Ase3YZb4tgj1TdRKaeKVYf8UZQk8xiZ44RHBX2fBxPIPr8dsgI1VSZcSa4RVPsvRD4CIIKXOmks2
bXQioWCS5fbUrp6U9b0CRW28ytZScYKEp8XBClr+fpyiadLko6cTS9sg1D1GxmWlUvONeaw1X65G
gBRsQmZ6lLmQ/HaXFk2Ue1GXAnBwDMN65VG8V1Okygeiea6AcM9N6s1SWKy93tQOWOdtgcjnCajG
FvH7HcuUqva6pIglbaXRvnD9nJmxQXSkfSiht5ORg9qFVknCUP/gcZih53Jq1NoGb3geGNd85Sux
AAkauPqFar5m1bF5M5U0bCowHY88cjeexZqSz5R9a0RBDvpwhwOqZF0AcPnlgGKT//z9ugn2qqe/
x5J3lekJvHUfSdc5tX80PEJn+TCbV+EVpolPavi3HN3W5A28cFuC6X4TczdF2VX7vA8QkN68LGVO
ZNUBLop+PN4IjVlD66lUsdbmIbui8FXOu8XaQhoOm3ygh9NATfIVwkWUCuWpcNanHTTPSImyyZIp
joA6uWFKeBgFb94yejl5k1CyRwS21e9OaudC1HGWRXZmNoYzYbiXDckpyihuVqLuMIuOty0L4BMe
lV8Ub/ERBTlI/2Fb1PfZ9eT1BTyTTcrbEcxwyOtm1LAiPymrKqwqqgAkeJywIg82xWapVE1VtLM5
tU0NqmPtE1cnqHodIQKIayBPdGn/QTvnMQMUVvmHgxbnGFUvNzf9r3rDNTvpZBUU7qchDrhYy67h
6ObLEdxd4TYRrZueC2tbOJgnoETlkIAsQL1rjTu2GbNxepX8wdpl5S/DuX24f4xgCkG0ymsV6W/E
CRqgeeK5BuQz7wDvPiZvVMMw71dsyUs7A/kpJIywlNqZL5NBeOrvmyCIx/8YzkWfnVC65+TbYlKe
b5Dk8HXYLHKVhyBfLrzH0ip7m4xdhSQAdKoyubXnUtO3fT/9e28bEp+hV3GEWJvXEd+2eGfwgGHe
J0hXOBwwQIPgJpIUBbfY5EP9KIOeZbdjHB5ikrbYbgtuRUvVelYqfdssl3IgfEjqkHaJXp9Ggibz
l/WBiCoUxizsn+A2pWMxa4nAfuQ/E/po1HqDw9HWrx1w/xr7kldhyiqy0w1/UnF/IBVxtxN0RZEc
FFwdaP73EArFN+d7qygtwLiejJUrR65a6NwAIRz9zrvBOE/+F+yqUWkqR1AkEmPUHw09OMG5y0Kh
0CnDrbXb6pGqdjF9MeB8tSmfFDFsI3tY9JTk3EeLb5I3Oklz9sG7oa8pVBzteSd5rcyoEfmW7VQE
pFCJD/MlG/R4nmXJcFSeaLyFgXYvxWATV0IlluZm5R7wIb7rENY+i2y+UeXL2iFLV67bCrYCYIJs
RNOj8zg8Y8ojjn79Lra02wQnTv+YGd4P7936a0IHYmM62W4qccwRnX0GP/yK10jlKtQnUj0V8sHy
1jIQZHyoqYro/P5AjgEJZaLjReT2ETeTF6UCYPyBofrVrsOxRnUy3BXlopfzgHxaQAaYcMEvH99l
83c/lZvBGlKLLsBBYMTEkjvd3ngrqVsvVl4QuE8FokjRKF0mZXu0ynt6yqmuSvNpKdSshPp5/27B
6eSyFSHBmlENtV7NsZGmkqCPKVc2R1CH8y0AmESp1B0ZOy5OaPqoqaspHOM1gUBbNkWZ6XrDw6+T
GkP+xM+ftyxpdN2UPqrvfEq4bJMS6iQQw94mU/lF+hzo6wuXqtU9y1b9/i1bYoGI5L+do4JJI3LS
Xrx4R7XVdor5GNuiqkLmEPRIwNqvYaUwgeabnSo0bj2t4KwupY2JlSoMWEa7tP8QVXMVpTiuv348
RQcRUuRrhBoW7adg29CJFml/z+uop2UVtyCOxU6mmwoATN5Jr8AYUIfCR6I+S8LyNVKPUMU5kkzB
m5scWarSnUTQZKRxtnNybZ+4Yg3TYV0d+XnNTAjjc1ImQ9r8kkA0J5zfqyxZxJQkLbC7EbhYWOz4
WYkdFBle8F5c98AI2p/e5gZZ3utaGDWLH/NbxboxLwjGcAZeJEBX33LKKImrOevWTRnW789o1qHs
gaRLyXCpCzVAeGPOj4kQjFM19pV9bRXpUvN+/RsTu1Y8GoMFWDGWXjv/0HF5Xg4TXct3PBVbRFz6
skL1mfu63xIsmQGcGYC1/U5BvO9tX3JbhBdkkU0JGoHO7v5zkIMWvxdWYu8EPWKDwMqQYHK/R/7P
q8an9o2uj5r6YA0Q1sRMRLUrWt6cLDlXTI8iifq82rAYniROphyB+AFtIrrJanahX26TCS5W9mXr
/oCcBvQfLTQs28pQ6ygTaSBDxzIIS1YYTC3j+x+PPXtsnWC9fMNndlVcVEW76xSm4WHIbxdEmvf6
tEGiQAuqsA62C0jmUMfVQNKc3f4pLg74MlElr4In/8YcfUNthlDAMPv6Oz0V/7c78L1iquqcKKkC
GiothZzYQKYfkcU1lRM2+G7Xhb7aSptC9FGY3Kdqr2uvLpUfzby4bU7cp9dvZN3L+mV20lJlYo15
MRIGRyxaSh8AL90pvopM49rqp8DkH4nI/yv8NGASZtZvwIIjpa1gytuYFJQV9RY06vsJz9RqYljh
ksnh1eJmNya+bydS7x56lIgiKuyi0L26qd1Bc1VS8vTwdYqMzcTRY/1gBzchgpcvkxEp8w3Opms9
IXs7o/ZFEfomA3eNtbmGoh03MNqRk7pK9Jzmcorz41pwTxSRhQHB3LFoYYQ9dTAkrrZ1hdC4tZuQ
kGNEMNGTx/NgzGQN27XrLzkuWu9jNJSXRmWelXmIBqAuvkpb8Ji5NXFXWpOvRVT0594zCNbadkea
SMcYtqrEOlIUi+Nzh3nPpQFpCNdscUiTQUzEC7FgxZLkhFJxidclgqA3pxlJu0WHVZW825FlX1C0
YX92u0nGx2Ijs9aeuwcE7ij0CMZF79Qz8WtyipeHPXx468WszNO4xmQGBUj5kpw+IPWGdl6CwY0Q
edhL2Y86E43aUBvZvOaDvAjomTkTKR9BpsJ8F6wHR+XFt+xW12oau+tQtPB++lqcGnLoZkRJc94S
nOI9NsgSxeVBaifnF1JH/ReSm0CXzjGS1Vp6S9h+tGlnkVosRg+44anP2eAuZEsIOZ700gh2HVua
MF3qdYMhvpUna6cgmWcQbUUHhm6oSEzaiJzPE6n1Ad1snIJ939lnVy2vRdTIbD24wikEOHdpVcpp
a1LTkLUWVlXmxnm9IbaeiwZaPJN4JSpsCiE3LDBqd0/2PWat1GAgnhzN/nFqnzKOkySfJYwzzhY3
8W733bGaZGevpP7Wuv8TgEtbdWg8sr3e8OijresjPpddBda+q5p7bbKXWWTrPWAXzbszQXmDkigv
oxviYb/VInLuQtfStUG+CPUO9Cz6oZrI3sC4fDIEpKEcdjCQOXpJ51TNHAW6iMDXT5Eo1Ku7mGpG
6+rEW5PLpkelKop2MCZOyMwDq9ar81OgemhzNvfymMBnD+Nt/7whbmhXT+z+QJC3qyfraXeMAB+t
ePqVcDlmqkRyWATu+AIi3XdyHg41oS7/bL+S44oJ2dEdtBkW6x4DYk/mAc/frzhkK6qiSReNnv0x
OSudRlQPZlCE3wgXS7V40MzgeIkwiTpGWrVqit9LsiOzYneoHKexnlZ/Arml2gScMi42F1KsDpOn
Bs0YyPnDa5WuqxXpS5Bfw6B3LKnVCeAjJDi0KwbT1Co+nxVAQPYPQAa0Uc68wlWIuVoQYN3L5DST
W75rsLiPIVVsoM0rHGpuwZlwZk4hzjNctQjwxvQpy+ViMYtZLEMkfyhn0NTf9Kz3g+YqHalFvUfQ
hKW+9pYFr3mKdKn3OmCebFMfWbWe+A/1DPwLESVLxfZBgsuX8cksvD0/Fe2C+Bs+y/t3ymMrBspt
gBBJoM8opJ9YwZ4O+Y3kN3t4V82son9gkmKt0DznzR6b/ZrWDJAGmCF2TEHSx6JYOEDkr0I9hy2h
Z01Lz1eDTI2bEPh+yZaox/IdV/V7uOt01Ilg8m/wM/AVrFsFGh+K+oqSBv++7yBPh/ONE1OyTp89
rxf6ImYQoMqmc88936XKbOqZmJ/Yu2D2094qsPy+DfECYDJ9P6eiYgKuEkTaDy0vNolMcZ8h/Ii4
LRQEvdmdnrub2B6lmVqKdpFKXwkZ7zELcJLwccgcV9lRrUVlizwHfc5/lMwE0Uoy0AZ7O+oyYYkk
u2UYwCa5UowoBeLnB/HE8r3dxVGtugWz/CYRh+wKEGpI2PLiA336eIljtlIk+lLuCr7DWLoyhAuf
ld3dmyafmYqzyBG91o3EiDO+NqM2TC3m2j2+Xx4NTrOSvJuBx4BCsP61Fhq86JLub6wA9/iKO7hF
h/821RnphQwGOm+atB9PTlDdcdsegDy8jlrrbQD/SLs/nuaQrdxjxzbncTLU0TGYNcMT3nEm/naY
3tWBpUPZuoe4fc0iT5UvxKFpjJlfh6+OEOfYNOy7vzVQgfQoNNMNUXQo7631hFM4LTBzkwX/h94D
ErED6gonBG1lDtXVviqaZ2A7q38lo/FWWwXPAOdURREKC1JVEg7T2CQ1Mbaz3cb/P2NAVmq+NT1v
ovi81TWjgk5h3WYOgRRKcPwXQ9Me+X1rf7wiv9BYLU1/N4gp0DE6KOLkKwA4EQeeyaO7gJqgONwU
/t36nuPMORrjTC76W/AQjmendM8N4x766d0MXUbfzBjat7bNpDvBcAAcY3e1wxrMCpJW0noJaswg
m0fdQ/FriBtTVcCyaciA5ZHNO9AZC0nvuDvvsqaqTx7cx39p4DI6663p332fF290eg+/4IsQaYYx
FzrN6iC5HeRrdQSz80Xke/N3/h+FiRDcJTutpiEn1axru1EkGnhSl5tsJk2lhUkV1I0JTAu3WfOc
w5L88AedOzf1rP32zJsu33A4xTiuLKpX0cmV3TLXdg+STBQh7eqAZgUGr+X8f8Q75zeg+u/fb6Lf
9nijcts8CNxQGZfV3AsVbiKNCb1oAvXi6s3DqdhXziCGDUpmWGl7VWTEVgQz0cqIMDurn5dA/hzp
Ny8ys0qpONdVs9KQG9zd+1qCH5hkgO7vLmyxOSwCEBXeCtR+OjLeivyB+wdK/WtTTGgbdLhUhzR7
OsSaAfK2Aa5Lrpva5VhPgOt3nyU3zRfSzALHrGujDbNMfc97Tl2gglcd1X9Q4x/31Tyr4zOeXiUM
Qhkwijp5IspWKo7S/2wUt/9k7HuDGg7Jw+soaaayPvBa/8euHxhpdRdbuTJQSI2nRR0dK0qA3aNJ
oLb7ccTEiQBESC6daQdJ/KltQf0koQ57x75w906XwKellox0xNMbz10Ejxn6fxd+2nlpapKpsmgG
iCfLmddNbOWzPkT2PExj/D4wm+iaL9BPaQO5MtzrsJExfv+W4REbzLKJN/L0S+5zH5rLPvAkVhTM
84wC8pEpE7O7SaADlKQf86Pvb2En1o+PwB3tPWmcMrQoFqki4plT0etebzrXJihK8mK0H6m441P/
vo2Pl7O8UJtGYVMsBOXbsY7Oz87Qo/Mq2yCo2Dg7RxF828vV+tc8zaglLfg7hyaVo4gBDndpNe4/
2peNEanl01tTUgGbEhIg3BxWkStmRkN1mAOrvHHlwbyBGO8vRxbIwBphRTxzrYHY4iJ8NI8gLgOq
and+bzbJfvifzVkk9CYPA5REJghGY5D+CZp+D87fbZeDIDakNTennliuWuz7LUEOYF9hl2KAHxC2
hxAhdd+B6pUP3otSCLxGozpUhyhQVeWtqLEqkKQaLpOcHnCU/R+jrgy1GTIVNG6ai/NjbDGIAZGv
GUgduze+c0AhOt1e3yBkA1nQDFwxR+cK7e9UCq14GjP3uATspxnBNm6c6pxQe21DEqRfORqe/XCc
PuJVHjKcQJwdRsLuR6D/ouWX+L98vjf/OXg8/zoGWVTBhoYC7Y8Bxs4luyuzMbY2L1Rd8Pus++Er
eFKjz12OIF0zbg/VKtbT56RlF1AqGNz5TqRRAsB8tHpQFWEgbRmgJlWlB8W9qVO4Xd0iDlhSo3Uv
YzwUxpr3vDPToBBkyOLciFoElTj+8CQPsyZ2m1gf8GcjRFSMk6beJGtNwxAx0uPMGUbuQ8IOmpw3
eElUJixCNmvyvZM4tzuFF3QKLZBx/5EHxdZqqpmry9CYznIk7KBYsX5jtyENiZrLCM2zpCVTwOLV
doVJxWmy7LVccKPkW/Bc2tdFPI5WvaPlNcLXwTSupFJgayiWCHEIziVyapXceG88ViK5oSAWOz3C
vfcL5GDtVRl2vovh9GLasf0VbTnQcq3IoAZeYzqIB6BSgpuuPmk4eI8fnUgFiBZfw45P1/1K5NwG
dlVLqz0PicZ6eKnst+WVruJy4wfSDGY9g34llCKaW/39Z9T3zSPyZ9WBtcUeG11jXjYLynZ/2Inm
M3R9PkJGqd0Nlky68EPyByTElZUXvzf7ihtLXhZQh4/SjEXjXHDtiE5/wR44mk8+sQ4KhhRXPeN+
hofRyhYojnMvKsGWX3uN135DqZ5eteAwx7ufdRunQ7BXHAelK9f7wfMEXh8wQAGdfYWm0amAEWdY
uQv4q0q8hb4RPgDtSNXVZVd1lR3LCVJ36xp4NlCIAlt8wRvHbfMBCZmfw6MM7Ws0glh1lmUpvtLJ
D03zEBYdLIGJDpmC+ZRUhWdyurXNWZm6MTOUvfaoEfpEnvp+mqDyGatsmVNI1M2A9NgfYPvXFgs1
Y6QgOtjW6NCl0M99jIr59siModNMOYqY5nIHsjP5JRkUjUz7PEMrG+X4Vt9RW7A9nWAKmirYZH6O
UgIK3Bd02jMN7KBRtKKxlwGgb0mZa6nWIvbe0WxbJODc+3YQCIKiS/ZAtP2c5XrZ7BlFksLvqctz
i06mM5DX0hDkJIIUH7CDL3bVOI5Kb7ROQWKs6JJlxcECWHpmwPw6fE0Z6x84xzIukuH+KqjranvK
L9ZIpNzYP62NyqjKatkNKVuBY8i1YG51AqeWlSXwrUGTN3A2XI1LkhMErUEAKEUMYeFOgssU9Vo8
cFC2JCIhO4sFzTgqykJtr1BQMyZSl3fhpH4jwr8NaymOnxfyJTv+DZR0zuy/kbPkC4zqLzGE3s+I
Ld/wa1GW00aXbxhpPt5r81NwleDO7d97jP+gAFcD9fV1SG6MxxI3Fb5LcuTZcxvkH3GDY3nt86bj
AqqTvoCrE+UWdfhw/ueuI2sDXvRSEA99s/YOWEpXAy9CR/ALiwOLXkCGVWmhkVdiInOGAPU0vhPU
Ske4LOX498MbWiLrkzMo6R1uVC1y/FIkTKueW4I61oa5tXZdp+rPCnXiRtmD8khWMhE3YSfeKWlJ
2Y08N+TyrYFFPbfn/J3YEHDdLN/eRC5gjRFk4IEwzkXXzXDJlxVkECaCY+A4544K14aUWYlXl1Ql
oaaPybRxnT06CE16Pg6SxOBkAFeQxipncO7sQUQaEIa81yTL/9wB1JuLIQ3MZow0+4Wcnk4ZMyvM
0kLXjk5P3+yNe1Wo7jb21qTGpP9z7MNfW8Glzz/vX5XAuKDOJk9ISmnquTPqbNvZJ40/deg0P8Dm
Wv6bouEhF+YOszfgBQ/ebugsD7yAYqH+4mT16j2QZO+oTKFaYrNQSbtLkb8ht9DqlsiTvlVHbJFD
UuT9b02fm/e8UTsZVSYPAiLnP2zmu5Jd8DxEGMeNirrs8CcpBMuz9V0t44DzO5QC4uIIZumJpySW
D8itCULVT2FwUU/xKUBXM48GZvVfPG4AekSSBInxvcaWfX90phvXwNquxboubFBBo5/en1sHk7Vt
AnzzS0wmWrUkkqgpTj0VB1hFoAfqdtdTcZvRhrUm8kzyByvGkGwg8WlNLd9RVZXHEWEV6gN6NdeF
5qkwzOqow7S6Es1I/qkstOTbt2OpjGyqpmEkGS9uAKIuV62Y2O658bV59lhuZeNWjCDh4BhM3YC6
ntH5bMdd7jJtw1BKpBT3+drf1sbfJOyGj93wJYfWSNj2PEwEnG5nZ2RfiJgFZQdjb/vhZg8Rjdkq
Mkqtmv8iqPnUBXVjdwMAPG9YwaGDvjXdbP+4YyhvyusopY17rv2emmyWyNj2rEAYTW4GfiGfyRWq
1j0QFoYGVbzGvRzG9xhU9krGCtFSjbBW4t0vASCahvwA2jvzq6VoJcvOEMcqoUCLQBsgmdOz4krn
uwJH52xKaftFNCJmrKBOmfwZ83A7Tg8LdWxdSikIdS60ze9/9g4IZCBcqq8y8Z9cigraCIWJZE8O
s4lUrBVngb78gfiEaZgd/ywFrs7C8HQetSp2FbnnNhO+MCcbIwacHlPXKb+YRxh1xtnnlsoVoL5i
z8w6PdGp9Ugc5O3DdKyJ635fE+vc3s9W8SeSs6qe/TT/bpUWpNT0njyDc0A3nANsqJoBydy+ysUM
2LR6LvHZeVXcbYyUiqhgTFu45pIQC3vrfgQk7SdGFSWCXKJOEezuMpmyPWm6nuzvMELq6EJ77vJh
EusulNUTbQOivL5XtdqK6qPIgNQE4AOAr1uLSvYaJUIlHvDoaD5qHKTSNmnQuLRpbzmCpVdamDLr
Zoe49jsKRTAgddbkr0qOFwVc0BN3lkrdevgo58UNO/mO6nL5qikJWCt0mor0yi1OSfXlgrvvXYGB
B9zC/vK/rqfs/MXw++rwhLcNPdN4M4bEolh9a+C6ZyMJjv/LSog7ri0Z0UPp8IYNI8hD1c4T5Vuo
pwMpEVIcgqmTLrYJcrGf8w4eIKLUWv1RygCByFpZtpHf5dr9ILVNFOFsoMut2HeBeWHZf+gTHcIT
vu3Ycd7r0o7q8USiUy/m73bpKjdSV+nHd128Aq7KHgftWQG9jR6+KGsZM186u/CeRjJwN4uj6RwC
+t0Z4CxgTxRzg6Vmdjff2z8N0FI1pLCXk2T0fPQjxexvQsIRO4smRIMGNNEAIbAWuM9+dardZSGF
AS2FC67WJM5ADZ8JAYoVuDsB3k6eKBOGwSW50jnoTRiE/5qiLG8B0rl12phjYtBQDIQtkRTsKGlj
9mijKFZMvxKwk78NAPJoNg7hsXsVQOafvxXvCHtweX6Z9v3X2eYiVjjMpbt9cEPMEMBrvohIRnv2
x+tLx5x60j5GNhuX4TJSqgnUaLwLV3K1JhHugmKb8nvQkejoBzAJPfp/o7FmVefmzfQ9AQts7y+G
a6ddj+MkzO/RmnKG8ePkoozZAfDg+KNfS2+FLnf8qDGJ04XhBMYKydiYvcr8T8KxqQ1gCRg6OEc0
KkP+bK4RadAeucfS+9x8zvGiAMMun8/qjMqlQg65eyAibTCbqODqkNt/UiLa+U9bNpPXLavIdB7D
cBpIrjBnJ2yvH8C6zGS09o3glErgiKd7NCl3SqxdOTvWAOLEaL+vkZ+rxnTdRAJg3Ygj7AA74os8
3mLHED9wTAF0uWWJTyye83It02hkrI4sqmTP5Fe8zSDx0rD7+9dkBsJ4q1X30OmjbPkza+yZv6LS
UJzXXRoz+jkICtvAz92L/B3F7vDgg+ykH9TWgp2AAu/j/b8nlwzG7sruJISfcmgymifZQctDwmQQ
sqqymXAmWNzEd7/Cq7x6MIqfKCVleMx+ONfw9kCAfmBUPewHMHCPjDxsFwDlHNEfW9KQNMbOFyd7
UobU0hyqifqEEcSRmXhpnSQWoT83SSinNCC4YdpU2lFCXGHLVYEtHPCStplKRClDK+pm8xeoGMoS
+5HmQmoG9xo+J+9XY+pdUGV1QTyjN7qYJ8PlQ7v4KuNCZctItbPL97CLnHvUmdBTwEl1jbAJeZu6
YrP/1ZDO/uDIRhQUr4iKyQ0ho+zDHmH/+wxiYEjA6NFrQrrQlbejFPJp0j270ylGE1zB7GJhIJxO
pLy6t6i/5NR83YgTdoO3Wx1wcu0tqu6BAEfOiwFer8P6l8+FZjqni5UThO7uhfTjomx+mflG0Gia
C8IF9lkPeEFdS/Wh99/2D8HiXuaalvz+8otFVDQQhmtSbEsJ3P2KYNlhI/7CQIFROluPK/wTlMfk
iNY6yB54fR7UEitjphxWJ0WxpnfK54nGeljmAa8R4Uy+7alI4pZ9o7eL7RBfplA76fu4NaifQTGS
Jrig7/IG5vM8ZvnxfCom5Kv3EHLuv+Kl1G/4UaNnNNMcAWnx6U2U9i4koBfHy1cD1VUHWaUHjIpr
N2Wv2VJGldfe4kurcgmyqtSTxyebJf4XrnUP77k/f9KV/1Eato4UtqGYBI3sN4pVApx0XCEEN4BV
9S5qwRKtYqbY/ajaE49uXKi8Mfg/oLpsp2PlyUbnSdT0VhXCAv6u6+d757Za3aEttl+wJgXUFy5x
e7Mlw5WADakzQTfKSFkeNTjVu4tA0Ym6ARCTnCgriiXc/igWfuHlyyHe8O0izTMS84fpjW6qv+uE
5UTiPW1GoDtlyMLnNG/aWtQsEyb8GuLWlpvf/7TRUJw3oG85xFXdBKXirBh5X+MXdIA28c0+nyJ0
SJkE7gE0HAAQz6T98AqnRxo+cJWsIUzKXkwC3rsNKcFDMzLTew+VpgDqrONdRytiN1hHM8EIo9eH
huhOQyJJlWWKvfnibtS43AEiu2l23V4pSjrxsVVmK9dEuKJy9ulVR4uDppmOnlSsN/+Rl5P+G31b
AuOIHoC+1rlQFguSOB9iqPr4TccBPi8ZMEaABqWSDqfqRBrC1iFDKZAfNb6Dn4RPSablRP4uI6jV
iKb75bNzjTKCHdCVqlLcpUHGwPnee9Ta5IioV34Ffe3WQPq7Xe5zAhsBI+16uywg7atyy1+JHcqc
MpuKudkWmKqEG3dtiCBmq8AsFSRfU8SO+h32ezrSj/yficErPorUMM3cEaDGerOSB772W7JFPHqT
4u4/54ky4fkJI7rxaiUb1Z37XPJqWhBpzFQxO3/x51HbrXeMrgWTt0En2XSroG0U1c81q7JYpqgD
iSbuMQcpw+U7WqqEd1qyoAP/N8m68tcdhLI1dZQz4SLSD32cnzU4ZMWiu1/RDf2kjyh/tpn+X2rK
zVyQOuxgL+F2CLipIEwlDKVbVFN22QkPf59W/TbaTg5exuTSrO+lmjR6cisq2oT/E08zk6AJZbJv
WpS5/dK8b/3hTKwzc+ybWfyuB43VBLL7ReJ2IfH4WwGsSQQYdmPt1GsMC1f6WEP13b0Y7l1g5FRu
z0kDCO5Y/MzFoZXaZmLlD7HFmRos6L9n6nzzeU5oN4lhF3RIOs2xx28iBCLHIo0xeuc0sKHgE2KR
zZZdzd2v10CLJCwjRsMrkHa7ecBhSbPfEsk3nJcu1j9chBDBZk8MwKlwItEEkGI7IGO4Fn/GkYAh
rxD6f1/6Gm8vHRd1GJAzvCZdtMXpnXquIHzWbsyJbpJOiZAbOUCeijuS50ZB40j6nx16rblNzeGW
PnnAoUD6iuVoQR60HmCk1V0CSVdDACBYXrD+2kfk5cDHk10ZYej/22+cDCVNKedt/hqx7SPWUGkq
XR9eSj1cRwmtCj1jC/Oc7PwcyG6WjDPUvkIwAvKUnBFXVX3bqKQo/YLqiykh0LVCtOdUP/oFnOco
6QOxOzN9A9KShOF35We0S+UzAc/HqJnzAA5PjozHrjFtPHKS9GlVqmgxUk5dc6IvPFglB4+p/xy1
iEK83/GJ6YOuiHlBh7pJEVEbNSD8+pH2fzuilN/I4KonamCd3mnZkCWMzudQxHSXhYA6Rg8Kwi8d
Ga9rDuJVJjkNjcBnAkpMm47yliXLbfagHdEwVw4Gd1FBkPTnMawovuYzDKNAhrxwlK/CN+pZ7PZC
lElDL7lRoZsWtuoIgzCesPCTPtn8Z7oqoLD8syQsMLLYHsgsGdQXotF3C+XSm+4ZEWjmPzHmZ3w8
w/3x5WP1rwiS6lwlVQzPhONThoJa0I6v/QmXGkCQecmnn77FhqaOFW7iCHlQFgrv7B9T6bL9pIe/
kno7qzwhJibUP0ASnHEOe159Bd0CgdeEiIIwviyGqJU42u5jv8pd0NxsF1gM6Z1+VA+1KMIEcD+9
YS9VWsVsVeHKQLlb9vgkuTleacqYVqae1d7leuyQMqtP8bgZK9k5438m8e+nkt+0NYMSy1mBDY2V
4P2h0hYhT6aHvcJf2At7r/2+x4gCP8SCWfvkkbUVTKbcAd0+7IqLL7h0qzUvWz4c8yrLn3n5/FBi
I+0aUBG2acW3OPzwUmgRLBertFU+RhkixqAJ296T8kzTdf4bA0vNO+BBNCw7WXQeKFOu0XkCFx7C
zluZYBnCZBJGzVFMJ9vlWutR+6YfSEKQiQIx6TMBgxbf+fxxhaDVyD+NTB+t0youEemvf+asTlR2
5hs59wiqJD3Cgk2KqNlvTMeZxpBPj5Dzez7Y88Rf7JqsrtXcOswjg7s5QSr5dyM8+A+v+KbLPuFG
1tfhwLiS4hoGEwYoJ62Wm9+lHRmcF+UF9pM0B5Xcy1SC8PXtHqRqwYyFUHWqK0X80/tE4/Je14DC
KgLh5s9262i7rYDCd/S5DH4IzACXu5xzgGI27I7B1k3I8Fe5ZOe17r6fhMobJEF5TUmSLAy5pZF7
/7T47LXHo1eNmYccMBCYmlCVrgjGzSruLCM/29GqGtaM1ByWK/4g48mmPp/y/q2o7AQAy+36b6Ct
efYSZx7I/oRWKHaLXHWZw9y9B1GChsPhsJzKb84FDpet+jR2Cr7B0Te8TtaFZyOuTMt2ZNA1KioD
dBPC+BkW/CjD5W8lVQERyheue5Yt5JWV2OsiCRxnc/cpYWrU9PIJhhwIA4xmdK3rFCl2iz2Nek57
riZh8Ety7g5uSEkGzugh8O2AK7JNRNOTo0004yVS3jXEMiXGKIM9WXHxBJQGJOcp/mWOomuMP2mD
ARKBuq6MrWV+sBrZMEj2n8LVaf+LASgair2r8Os0Jpg5iFlphCGN6lLzEdVcLvieRsvG5+nhDrVi
5MHFNk9/Av2rXt6NuP+jeg6DIWWcB6eqo/Ft4ghSlfpI/3/wrJaokC4OeP2PZ6gBzCQK+qxK7tmb
TvrJ5dwKnU3Psl12wlrP6NzfXaDdchI19e84Wdqexbb4CsEHqSDtuYJRfYMQFhu9zEo8iMCujdCl
tloI2eJMv+WuTqif32plwN4+mMvfQGECLdPEmn71Fo7Izuxl8EybGFLhoW0uiHxRGgXEwbLNn5b1
TN0ojcKhX+udc+gElDDeK1pNw7KlHdukn/MmJWOiKpOZ4xjiooEDFJsVrK5mM87TeLCVHV2LwgWm
PVG5jM2FHsKROw1a5THHKgNiSznmS6AuxxVf1623Vh39dDMzTfmKWbNagppuZxYqwRiSfCLd61e6
dyJakotXJ7lV9O/0n4clOsjzLQSQ7KiFbJduUAXKA4uBTrXYNER20ZK4V1oshQ9oLj+0DFqw1Fxs
KR3RgMrRe2GwBJ1NtMk8ZE/+I+ZuM1iTBPkSHQwvdHQ6Y17y+izIVyhQy8u2EhogfF38DjHb7wfE
UWBAbG8R20Du0+UcJTWPZ6HPH0w4/P9oO35+09VcFGJMCctEfkIG23muJESINgcGj+Q6c1c4OHdv
wxbjYv6q8DLfq4gib0krCE0SktlsHartQ9d2wxfb+T+4Ov3Rr4FChsS/ejP47PeWJ0qw2k0sA3s1
J6l20wu6RM2GoccJV6adBPHkG0uYArFfxpD57YZ2A+gsEF2NSPct8HziJaVkJOHEBKXKBLkZHDKQ
xfCfXdCAG03WNziK2sQ5wRIou3BhTZMIG9b03BhowcnUGdOfYgII9lCXKC44DDzo5JVIp7wvJgpL
NN5XGTsN9Mi9t2NGO6eEYItdYg/tirbGEnww2JO2rMWPEeqxqoTMlljA1DZxErLPlQf1+BDzy7g0
rl73V2USRdugTeY8pnN9uXJ18eABEAevRVDbw9Jj++6HJzEyLQPlIIzwgQNk39v+Er0V55sBViqK
qoc4K/US+7jhWjvpghmo98rSZ4AJrt9/XiD6cukPjgE8/qF3R0XI+G+H8b6iVOapmTtxsVxA/s8t
1XF7H1cy9byzGq6JNUFsS+I7bjyEPo7sCusLq3dphyeOJiDOGkjfpTiMDfr9dkbyNA7TANUknan1
0kIaC7WquPcjiYAmnQpj0HJJKFYlijf2llAGJZ2FYDxXuqrjiFltpvc4MXLwZ2RCfYy/PKCh7bpB
88O+MZTqvU/vnhAWuQRUfNplI8yp4tGMicSWopE3AjhlaqZ9xNtuMRitig29X6sD6IoBvjs/XSD/
hQIUl4VvbcNjABmprnnlbwfP0qoHR3WHvXwK2+7z/sgpHAyXWVunWdpGY6kCkGC+hmQuieWuTUtY
Co2pYSa8cyR814RTAYzTsY4WZcPj6t/4cEZcyZqNiCuwOQ0eTxCJ975ARd2wo3JALRzKGvHFi+YU
p2u8g8JwE150nolnYcGPpFeRgKXp4ljqm2HPdz1x+17HQjHq9zh/Ddttfy/PVzRe8zXpyFaGr1x9
NPMpTmVB4y38TwOvGAsp1dIeE+12MCFuimMQYeQskqXR0QDyJN0kzqc/vDjU5NIouf5RcTXnS+cb
W1/0psLf1lHrJf+vXan88UiZFbX5s9gO8qUlG1ANPLAyGRPEBgGjqRnHXO2irIppAqyBI5Fa+oiq
Drx4eZAZwCiBYaaqI+Ma3dRH4TdeeTRcvNB06VE096DHOa/NS6FaITIcyA8dZmlHeENEzmuyI+Hg
eq7qqGw/Ajf9mT8F05fJZR7rmrM2lCQOhAfGldyhCGdfL9XzMatcTJcTpkZO13MdpX3rIUJZ1CZ+
JQz5zSPs0Dex+EJe3GVM0VOaGGCTdgBWMzTjaCYQjwzi0VDPapuGKP3OFq2OkifDTuxkW8zMgQOZ
rLmiRaVLIVmU3iAhZbL3A+p/0SgzKz7pL7tMM1LYS2aM3qR+4GYhkCJhDGuMqanx4zamMqOHL2jD
ie88VuXDM3E8fSWF9YxE0C1FvtmWMidsBonH2ctVVDVlA3si3DK3y934AjuIfJqzB6l9T4/0LmBq
/M9jlQKAQ0RsEldUt/Epz+QRRf2sXrTx1cvGfz2FeSGpBHBX8oPoQB0qPmZPVugEUUb9GB8G2hML
ag8b0HSpjtpXVh9pgUM3EQ5J+NJrzvVlgzJmZsqzZW2qwG6/dxTbJ7FonCds6++aH7X6LbsUEdzQ
dLi591HkNWqmj1QGbU1qYH/C84cT0w56KzHvF7KmB3CIfytSdhMEePm3/kHByfMGorG/utC6pGMG
ZU3Rs5cGbHG2XswyOwATBe/eaEs5+OWoN5+ffjNRBOc6hfPGGiLQQ6jpKVc20ItB5JEBMpU/uXV9
orsBMapAbFYtC8bSYHMZoquqiytIs9vw52LW2op+0aCu0Hya7EF0UUNpNeWKXd3RYPTpcL1XJfJC
MOXfh9h/mEZ2VGZwL4bt76fTFRTPNMzvWEizZ6mWbpgCvyEVL8/0c4LpmDc1UmrPh08RaCwbiw2w
0xsQP/5LZVzWmiKqcoGs9OFnjIXjgoFglImE2whFL7ZPV2q8I3d4DG+7UcpEa7igHkbAXbrC+DfS
DjqltFsKF/SNS/sgKesZp9/XzrRJeGGuM5Lc3/JdmKhje3Wu6ine6xlWvG97AjFu1VW9z5Bv5Lxh
vjr07QMwCiwLSSuZRbR9oxCKcaJdIplIi44QCsmLHL4LKSrSrgoMh2Yg85Z0TXpdxDh9GSJjiJYH
i7qjuQRPvCOwD4sGkzL6G2xYtSOLLIX2yiW27MkoZj1WDYrPpf1WjL1PJFBJjd8TTA+SpvPXgxph
Pjmslm6o8xYTt8fTgnURMzfWKn+aFvzLvSB4U1DsQn5RnnWhQGIYHHzx/N5wMihacjeYQA5uPBcV
4YdUBXH01oJansSEM5nlZgtCj1AVafiI/0EuRlzFSYLxTsMbRYbOtr8Gw4oMmcj4xwqeEnapuJ9a
hNebTkTu4/eNyeyOibIcLGptg0+H5/7hDiLfLBkDWDgxDhz9xbQQoPKgJHjgJ65+6JqhUDEnc4g3
zcp5PRz1NcSvX1nxUcKnRXzuUNGeSunNWY6prdS4Y+DSq5HuVUmK35DOyH4xli78S6snz+QmBlpQ
WEBzQDJ+mvVWFw9Kwj56cSlop8OiQNgvEcsHuGieOcOJXICNVqq9GJvM5lJv7uIlVfBlD+WoUTHf
9Dn9BZRVqiWoPNuUKftR8A4+V19iXsLq169gWugepDV7cPyDKnUMxdi20aPJOkthaCwS+IT26HVF
kpXSrfCYKyDEQv/gRPDh30MtBmDlizY0DLnVMtWGj4fWCMuELz+6MqaUD1l1kHILVqsXANHJx0TZ
KQKeAdAnlXETvK8VlxQ35dicdTf721vKO58eiBca/uY1g4OyAu3JGgkLRsVJw9VWniFiGfUrgfNY
0Br9At6VsGEoQ0wO1ASSXO67CpsHPc+RnOoWoQsWJna1mdTsnFkU4Y19T7nppHakBS3cYWN/lw4j
orlz9b0WQC7+O6IYv7Bojma3UMK4q/tornH0lyyyzhPAGoa0ZqdzPf9AHE5yTpVP4KVEganvHfGw
WtjXjcQSoLklRTPQ/ux7YQR0ZLEh8B0inGztVendjMd4xw5ZZ6/Hrz7aAmpTX8TJNMuNM0CfSro5
NIK3BbSXDn9iJ1YWeNaYbmjJOoDoeyPjfup/PoxeE6fHOGuUnvDQWZCBvXoDbrQPTYvDWX1/XcJr
HlLf3HJrhrO99pxLH4FFGVjAOcLf1ilRcIBaMkKIhDSldGqJ2h4DuerV//iduneN176ASXvICC8J
xBTjcOMRajmi84K/twz7yXOoLt/nZnJqs5aiiphaztHIXmrAkosdxGgMKN2+olSKqKzHcIZx9p4e
0vJxjaPFAp+NLZXAumR6Q+Ni7F50qM02lzAwhM4/EYxbOGZSZIc3TNxw9FAEc9fF88AasOlQJuLs
t2O7vzHiTK7/1Gz+8JRFzcXn121hl6L+y2B/YxWK9PYj0wVrqc6KX6xmnw+oGG86NuFHZCYq6Gkc
1O+09xRYFWqyB4nH08XAvIYl28uT9qjvMPUzKe5bz59NKb54A45v2vnyeWvKIzpokMfVIviImL3p
PT34XnyQ8eLphgezOjW/+CoLUzUcDuKGIKuDwAtNkn9ESJPyh3b79eId2gSTE+uh2k72argx8m/g
k6YxfYzcCx/9P5CSz7/Bc+4nlmHWz67ydfyDPCRw+eM+7h5P7w+aFhuF5xyH5I1eZbNo02GA9F3I
M2/Loxq13o056l9R9MzRj2Qwa/v0ry6OkgUY+teTPnmhn/7ZQV35aA/FBnMo7rAtWoUEmuwlJW0I
FOTtCXlozuFBBMgXYWWTHjMWAlmTL14m/kVJKR0XsmXoAXF8BPLWm6vMf9+AEvC+Zb/X4MKUlTFo
ogR0cfJTYDVcTROn5lKQf5wPYrZtror4SDJ/6QCLSCgloWsw1j9wW1OSTUdCESc4+Eg5Zn3kzCGu
5tUpqqt90PPmRAIp03d3vlyUXWDNLwWREkUBN/TmVPHZFpmRJhgV+GP/4fEc7hO3WaL6OiP5I0gt
dNbHKGoS5LWQ/vMT/jAi+/4wNZQqsgg+IV81/jTg0H0m0q7xgFHn0TI1vWwGxMNn+MMfgm22tYq6
m0bAX7Boh4Oa7XETMF9pKIkuxEAODMacQnb5CHsH2/MbTkYKOC8oFmq7PZ4kNttQn9C6Zp/ve/41
5+EUdei4Oup1fBCubSW2mJrJIqfiAeUiw067xHBc+T9QSRqN5jAvsdgEVMery/JvlaLK7vHDev2l
uDoXk6us7qCZ/nQ+iC8Dir1zaHQ06Nm+SmeVzzEzhKHj2DmXdZMxgaIrQowXK5sNNRCA0XLP1/Hu
/La6jjzJ9jVzPOB8uIcrWxsVeCn3uVvdTWcE5d5Q5Dhjt7QSNBtMca3aVSRBkIEgEy3BXfS7Ubtg
RPXwC2+IzvAO7DWWjvFBxst4ZZ1XIG4+MHbZjH2d0/uE8O2+aIochur7y2d0qrUOKneIMzKtsFCq
gXSwAli/qle+lyGBWy4oq93OnFRnV6OrpuVlbXDbXZNpIKughF7M2ocQvGsvMv/Av+WepAScJcbz
Gd1d0wbXbQAutgmcWmiBpb9+9rzKXGAEHhcmf/zkzAwn8PSrwDJDeNeS5vSZfF8ZT3v3zVaPYy8P
ueRqBcKxp7USXnnvXeuFrVnO7TW+PW6p17A/KzBrjvXhl6Cn7pGudDSy1kwjxLzpNvrzqM3V8Xci
CsowVZoV90O01Up9msm5aurxrk1YROjLVTZ+ludHXzXeLovQSxuvNS48tHNjruHNL6v9BDGpzvEK
ylLw4W9hLmoa4qBqEdl7lyhbEBBzZO4CDdUfwE2a8i266vNX7TvBggagjunFhHhCJkzk0dE5NCFE
G2dAv8De+HpSf8PwdKFFHmPWbQwYmeAGMqOKXwJtMoqqKgZlN5whmAO5YQ3ZAOdIBLuFReiNDYsR
m6OAVMS/3SaTulbnw8MSvooBNjsQGXSra+Z6Q9Z8+vps4rjqxJJuL46ukzd7ua1urG0IK65QpKc8
kDp5ruLYzolJ+MEsJ0xClajGHZ0voTstVAPJ9NHDwnkSeb3ti3pXZAiAKwnfjmcg2T+nUkX4K/59
33Dq6Xiv50e26RYIR23g4Oy2pD47Aw3/Rwj3neqRmsKsySylzZbKDqZt0hafoePDzK4WEbXGo/Ee
VCkFlAYB1y3uCyK1WCYVTuyLjD/ysigD+tOLwUF2MGqPU9OFYv8ClGiZhz7z3AkcSPje4ArOyunW
+vwDYjk7rq2Di8bV/ryMYGGvdtEEXPzknlkjyQflAG9AClelPyMpuK6piqD7JiWLzfk6gqySsFsn
t9DUbKFdnEqSbvi2mhaZcU/bLDiVcI+Hv9f1dNSZ0KbbfKResIxwN7xWJbY6wFOq1T9VwVbx6HGb
V7sQ0FS9kjOCD34t617p1pGb7ov8HH8k98xNhNsH8mdleFEWvwHE9zISplNGyptkPaf66vpuKVGU
CDMpOzL2X/CFXwTN2a24891WR7jW+x59DhSMYnZp+hqsMRN0ZOqrBFvnb01shR4mAvXahqHAWy8E
8H20NaEQzQZPLrx2Ey5jaOqJtysgfk4gUjo892urfuvtoXXwcUtObP0JCdwmEqPt3R4VWbwsSTsB
kh0Bv/jbp+oApqep6pQva4DyXg1/o8EkPrM3bsmBhMHwLTEZu0IFPm9URYRUX0tq6OlRM1uIBeYD
yuXpFJc2xBz5H8YMnO5Xt9+N4458rzkb35gge1NkNEM78UiQVtIHmrhMwV0QqvGuLwdx9cdXVmiw
K1UeybyllkiUsaO9H3k+IpSvtw2p/gkgIfA0QxEsPKgLxKA0SOvMSAHBozn1s92AKZHIdE98IUhQ
SxMUD/Wt1IM7l1wRGwWg6BSZXhmNGXRe4HSayWER7OVLVmOcsXTTV0HRKnMVruEhTRw+k+ZK/f8b
lNb29TJJr4sDgRDRb/cul5+1m+ggk5NKnGovz3vjHtkgbYqLIoBjhcTEuOvnTNuy54hr86hXy3Jj
0lxCJlSwX+mGgQ0YqaOuyDSU7LtWm1oawwJ3AXtxO72XefTHGqiC8de9NWZOkdX6Q/ExzNp/WLhl
FMUWedBo/RXhcbXc/NwxwOtjoL9ssM8P+lKpheH6ETtL9H77Y5HjZlDjkgnfkTmSpSzcBXx5Vd9B
NslGTi1eWprv4vHQACc7bylYIQ4iGk5gR65Po/oBxwVKs16ztzM4xz0GKrJUPSYPL7l8piApiVmV
SVs2xLTmbgK6WmTgWcGJIib1A7l82wyd1b0AiXYzYtpjRNgkjvsBmxkgr1iQ+dzfK2ggJWzWTb0s
phrh2BeLxVbYdMyybMxtX4+zCXYM+kK4po+qLnhKhEmDzoLZLUtb60lXmoTdhWkQzEvwGtn5QNxj
oKXxFfCfARPlrckCAAgaagfvLLjAYtxhuv80Xwmf2EUTYpPz9UB5N4e0DSZAWn6B5nUSUWo85VjP
CM+ge6tVHQlevflspweAPir9oJJL1263tMfYRuIgzJPgbS9Ctczk9Dlx2MMH0ALvyoKEp+D/OZD6
y9s00LGDuJasAG9HN97GpqP+zIuM9h+xSnlqGiIY2n0CUewTzBhvZNf2pmlFue7+DUyedrfHqx2R
nfea0e/pJju1VIA6YDKAPYv83LnmI0tah3/4CJqF6QCjkU/a9oqNtq5zcWohQfcT+u8CcGsPCQL5
gq/ogtKIQmjuu5xN9kuhwGY2svoOTT5DNL9G6tYURkAv7mRfBlUWIWkG2FNJfdO0gsXJo7tgFr9Y
1C7ib4qQlbZ6MSAQCGzCAHAF3b4fTfrw0MaVRhfkSg/gsnqMDfA8X7vmQS/PdF78nQesdgBujLJD
BSj5klBmke7BX/5o15bKWwtJUfH47rzjt83DPYlzVDSpx47aq+VQ7pOaTou1n79khQah9kPwmfDr
IBWXUS0ChyfvvSNHNZ6E2UrtYvaKRhiuBudS6awxBAw8E+Y8rAhixgB09ckpkaey2HV4cZC3rzQF
odp1FxZwOuYugb7NUCWeSk+2isBgRO0yzpneLp8S5JfbBCP3R7EwDb3jX/qwra+AEE48Pe3GDJAT
z5Ufkj5Ga5l2on09DfPoJPC1DFiPkW/epqZoMhiDuduyZV2sAE/k1ODtUdACo4XuDEG47xIchSh/
o17pLYgZuc6o9lXXGhedUIJDkbBmgNRnDBzNNmlyZIopO1E/YYJF+b2lUFwwt2d7CJaG2sI55U9/
U8GBWUYtZyvTGJtg8TuhslFVSxh4TdOIASY/eeNCaiZ+i/Ah2zqs3V2ZVSosZNku6h7oeY8qREfW
OlSPDukjENiwoJ7L12XudcTm4zxKy4yA7VmvA0F9vLebxoxET2jV44+CWnhf4uG1G4AoP1IhHQ5S
KSaN3xlWziQZLDPgBeaFgZkhEhVR5x4jqOBpe5ct4WvvHRO1vlaw+1nrwD73yK+6X2r4je0f68Jh
FJXv05VgrMb8V/MFbRtTibI8hayaw1dnLhPDmHnAAYbxq5EGm2dSvej8LXUqmKaJZ01o3n8s2mIc
BJK/kdWXdQppCPGrPiTesqSPLgx4m3Y72jHDNHT0f14GWs1l5PsOUB1ycv0ucZcYu28vKDy9bgBI
DeCAqNCX1/EI9hT7RCRTj1qgBEkSTCrmVGMOpjgW08tq8Xwa/IRwLX3YpP8Aqkdvn11U4DLZVtks
3bqclciU4ui+982oGruiFiHB6qdUu1NwZIIgBn41Yls2+YVDJ08YNQv2RdeTa/5WZPHwpOlA463t
d5IPrK60HyUjs/KpiD82g7QaLAERBep3iae+O0HK87o8w9jpmZe+LOEXljfd1Uc0cgN04wZY8Bl/
THHQx12wXNTikFQfFCkBAnP1EmyBFXQPkUsEJCYgfX9fqefDajcwyTIOvRryMZxwoixzPlI550iO
us18ZyBHx23lrcuEli4I85KJRUMz1tUW3YvfCS5qVcL/4nNcVXB8eu32pc1SlgV+TCdSYshbAUBY
TvgJYFnD8uwoUCpwnpliELxSHohL8f5YWrR7fk9CyoX0IQTNYxiXZHrcWMDCxDPT19pVlKXpi7hh
p/3ix6VrTyY2/x89EI2LJnwb3q9QnWhT9FSwba9lRpt4xwIJoA/QPlWdHYDmZD98fZWRmU+b5Yev
mID59/2154v7yhqw3LDhjqy7mDtqARn7KUCXV+4PmIPFe3g1xSwoWSBJ7RSyB8uzeUTbQlhM6L7n
Bt+et3/VjD+aQs6ecouGTuACeg9H/4GoOfq6YCB1zxOLMsb0DfNIvl3Ifm5/2fZUYRposrzDTUyX
LBuPAVrihoukr8wnGDaSORfpEQWoI3RFVr2mYnPmlbK+yxGTuWRxKmVwgp7Vg/mZFZWu7mvP273M
ut6QCzrkj7oDTcGN/B9yLjczbVL+cf1F+Lt/x9yrNMlqAjPqshgRLqehttKNxrKgJIVw/LiG/Tih
fTLM3mCako6Vk5CbMees2YqE3Jsc84tBBzz420h1/Fvcbiz7duH0ZeWewXcq05XRka2948ssuerw
JiXihHBT43aEBzSGx205Wb1FJNu4wF+/pSpOfyRnwvsiFCAnluQdgUrOPgAkD+CkVRte4Tk5HnWg
D+iSoeNqX3tlxmWdXQ/xvGncupNO8AGim3D/5eAqDcc0oGGH6BJU8TTNaOhxI5MZ+q2iaYKXIB1s
r0cPQ6NZqODQu8XvGCpkDm2AcwKywl5NIH9fmImXbkhq/JUeeToslOSRXCRB2g+w3n3HtqvlPnxz
O6i3DifAsnjP8NCAjJAiFrdwfGBL43on8iJMdyPy5gOJmvIlC3mJEYKYKaxdFaOZUTxB5V/1TUiG
la3hyo662I4hvqTd1wIH5EmYSSLJtKFJ7cv8lC5ULKnDNn/XnIXgdrN7DdJbSYQqchzZow5ZGb2c
Ga5BE1dPKlFkDC/eCSBtNejBMrc1JvpFxEmXL0eclqscI4HntWwU3At3rcqNcS57/bJ2IJqJmLPV
8qKH56oxaOMl109HOny5UiF3ULqlcBnMtZ3oXVS8/njSWJPtKpgtVeMWi5ZBp1hkwWA0yAT63RvK
aX+wOAUmJ/aL1r6ZyoujzH2TictCgKkrYDnnhXWbCZpx1BpMG8HIeKph6LPP07CF0VhDgl9yhugj
YU6Ob1kjfKoa6uaxZzZZQ8JloDyA9ioC/KxgV43hnOpiN5CuOubsiZ2JgxvT8iKhI3HrDk7vg/nJ
dOh32tYpqW694+B/h394qOoq8XHkqnpcmwVymbJbI6QFUBFbF10c6He41Z16SayK6itYjEY8huDp
mX2Boy2v2PiUf5VJiywVhgM2eEh94cRUDu1kwc9fQ1rooDkOSMfcKCxpK6/xCf3H4a+Wk+VheMxP
L1NqLad+tRSO/hDk6JwLJ8K5D5o9PyNNhL8EHy72PGdwgv7XtDq0XTtZWg/Y9xD3b3NO+qIfP9y7
6AA9nz6nVsKEF8GQYPaPwNA4dM2SORT+N0k4fE03pQ3TGu2P25v4HH0GnGHP8yrh6iFiwT3+9kTy
HloiTCGiNaJMJTwNVHnBeybd7h98yGbvp0IvmZHWFgkh+EQR2sMWEtBb9ts+AvRAhkyDygBjgB/L
PwSjTtvbuVesOeI/Jy8hUkj/4eq1XsiaHXm8nZjmper68UeqhIQ1ycUd0V2xyvhYj/dU1wSKVZqX
luubQWEk2eRXCvvV7wOc61gqQBHHiSF8N+8lturPDSrqAlpqZuFUOf7Kpw3WR5apal9KXttiHGdI
/1HDpOfMANXKhIMwDos0LtzxRmz+um/qVuCDaC4r4jFA4appw0PxTARCgiSsI5gGnmtG9EcZ02mD
MbijuIPTQwz7qN74r/Ehv2GYGmux4hyh/vB3Y05KI1RanvFysAijbLlqStTTYssMicPSALX4pZB3
fEwuVGxtPrYhxNbZ7L8Cpo7ycfNWwgQMjqiHTVYLeN2EDwLTIfRfK8a0ugiJ4IMztu2LwjUtn6dc
j7ztWKeNeWYz+1FPpepuQuiFfc6k3ucdOmmpYBoMpbLx0DZ8zRKEIzGz0Eop8zJnpYCOhnBI6nBg
RfZgLP/va3bm6Bgl8zXV4E4NHrNjrsqAlAa3r68lJSU6Rjg+YP5jfqdNT5wXIQ6N4ioA8eOz4Z7l
QuO0wTZvaldf5bU/HFZnDR/gRVVvqWskI7sEtJyR3rVLdd9IPsJRcYWkrDx9We9ls6fXnIbA3PsK
P5b90LvBDDN2GOvWZPxxfc/M415Td4Ic/iRETuuP5l9f6M1N7S4fZDGsd+pcF4vgjjeWzhVYrZy0
B4X9tWVjkxnSiFEsB2eXVJ7K8/Ic6r+qcP3U7aV5+h/Bw055eRBKbWBx2zuG18T1v5bquC/CRXQZ
2VSriHJPldSnmUgXPbfexMUG1r4S4ImAarcBkep9N6/YcE03Q13CzKRzkzvnAMQPhSy2tg4pm/5q
rUhjsfsl1JkeOQ918US5/4FXPP1mVA053cr+2BWaI62bBBlKEWC0Fjwr+R+MFwXrT0oKguhGtWTY
q20K4rTaD1NiHywYmtb2jBYpvrZnbHdE+CY1gDcqsPy/YOtUfw4pRorlKfCKL/o8DQFGQ5fsXdag
sc1Kt9SW6kYnlXrT8Fsf1qEFDURMW3ZKWoandCbHj16SQwwiX9Dl1tXJDlPQOFMZTeaIx5WsFh7B
F80XAIDkpP7TommN5amADdTs6swnK3sf/pso08zav/f4T4aJDrK5eYB2AzL0TkicnCBmqWDi7YIb
fFH1Dsj+tYZ00pspOmp4pxNiiI+U3UhU61UfQtLaPDMJ7FX/xKh6XXIOh3PaXnDmXfBmn8k0TeML
TC3GTKiEfY1608GGAMFuTFcTTemRPcQNnlu3qAXFQLu0Njc/LaSGcPm9ZJibRaG8sAqZFrDbSKvi
0n4N34b6JjHFhM1ng1Upuipv7O3dTWxmLpZF/mrQ4kCJc3byawt1zdpQLjTRMBGjnCZ4nCL4gVDW
Q7B9MDAne3tBIBi3BffJZpy06grE2uzoBHQuMQIF+GSaJO2WELfQ2IcCdSy/aVrEhAmqo2E0GMlx
PwKsD37+CRjpixp1mA2Aup0Q73Kp6vX+PHD78ZEuikLSRt+mRie5PsbUyQ0Ncx1oo6ZegjmgLz+C
CdJJmbCEseROPOqQvrothc0pZNXWrK0HITC0+AFE22eSdG8DyiXfb8oENbpzGM9gfwZvQaVOtl3T
SBNLt+NWNcQ5l/N/4tu4n1FKTcbxqmNflyf6HxGWuxnKI1Zp1FNVFaDh+9pIjff/SzO12vJflN3y
bnCexo2GaZ00uOtE63UKcPyHRFyeExnUyIYzbE5XSvcaMMfv2UztfFP5vgRduGD8d4ptxs1wJQnx
yrVkfFkp1WPNB920zglHxZI9Cs5RtklI8qJLkjPko6JzetdgqGkSsTltp6s0usJVzoSeXOLQfUJ8
bHk4dxEY3s1bN7DReKXseWg1Rw+BnEVD0Na6V3VYu8pxHjvptxfxemD2xXcgARuf1Q13ntFXyZsH
yJGKrhHmC2ves7/jZXwGFcwTRk/pGQ1XwSy28+E3S2H319U/YARZKEU6eVgRxa6T0AU4WsAkJrLe
haBTpYoJCj4ro25tSym8F/N1hcyIiae2yETfVd64ESAmuh5bSOmtEE/CvLwNTHOWk1iQOuCRwwvH
q9745x5c3AFIG8dQf1qtVziWqv6P030mDiuc9FRdqkmgE2VzpSceaCQurBcqnOyAy24+a/ub6yXX
Bv/AJMhe533QDE6Leoj7elkb4MbT0biZZqKtLDeFckMJT0unsyj3+8RDia/60DwNnHF6vNl40Y72
d8fvrs7ZAZKZEFwAipqqnfOizel2aTY8Hy+hgG2rCVRed0lbfSLraJx7JrooVYkr3bEEAysINgvs
BadgWB2CBpiE/0AxQYthB/Je/+vc9u6ZjlZOG0NM9nDbZjCoz+K8NleOTT4xtqme1fyMYCBCLfO3
3b36jhVL/YTN82ZqorloX+7StIW4quTLYrtRyqd946Kduk6VJL7Afoy8ysjx7k/yfgKGecbX3Jt7
o4NmAPGZ4PMmbjqEtj3ZpA6fPvzJeK1DA9XCjLKVTBiCxNaIB80MhMJYnwz+pO+TGd2eVsuFGf3E
NC9zX1YUdeCxxbS1kB5WpB4k4B7zphb8ZXy2ASbj+TP5+RveNR6IQr2uERiRIIaNbOkahEQB2JB6
Lo9c8rZp5qugbrIeQ9rqy5nghZitTgTaIAMS0EB1e8pvuGdeePkOYPNJ5Quq+WnjDIyU+IYsr4rw
gJsC//pJGsXoy2g9rXDL5fzJ8JahySRvQzg0o3e42vxlBjPOV6zoXxP9zEzhGTv4iKLExrif796a
IQ3y5/xGnAOEd0J3jp91XzmRkfdbD/sVQSggo/LEGxfrjlTm7bMSttbqiWVx77hcDh5B9EOzgUHf
krSihH2yiFE+yJmMMgzfAydl0U6FcNL4yycmS1VTZit+zTjouSOnChmUCsUllz7lyZCoLdTJ3osY
tqYXQMg+ZmX0pu/cEjX2faLVbcZKBKixN5FtDXLDcn3kMPpug/HjpsqvirzULGQVQG2tz53hV4bN
k89MmES4OUOHqsxvFH5vAvG1U/j5oWTAEFIbrCPUzMks3DfeVVq3LsRFMnd3/q5SxK2sadI2v2Lq
o8x+dzxVh5sUDY09mJfnvKozzMQyu+ZDbpyQMKsgqAuJMCwlhZg+RqAkEuEieaYRI5TIJOGAwVW0
KCs1GinNvID8HhSdRY0nYmIUjY2Qx5LKy8/6/gw5TOSbN6gyJ3FPT0+xewO5/ENLLeXQuK1GMshL
m0bpE92yZDYN5SXSGDynnbnqiSegBxYuNqtMNE8qb58uc6GS7ltnRaE57cY0ePVDz9tQTrYKxr7W
VchtZp3x8TpoSNeBIvEr2zjClGiEU7iCtIYUY89REIerWRu2ME8gdQLKH18Vs722GzeQ8S/X3rVp
Rnk325q5io0GFVpYz1NeakWLo1tzBxr3b6l+NzkL9AWbnE5uI+DdhPPVKOwmfukvQ1dmxFBnqyHk
Bg03frdo8AC2oCxQDpsPi+YCSVHToKFxOFUkMeToaf2sfWjYFvtoyJpHV7GI1fbYLxjYxZQzZ/7l
uDxMFr4cVQoT6mEJqW0fO7rXAD7P72uQ466YUoZYPnLvBSx4YGTNyEgPJ0h/M23V1Tp9Ou0JALAp
J4VMRZ0K1T1j989ms8w21sHZ0lX/bRctHxpndRv4+ZJoDVg+yRsPe9z1Qr7ahBSLngFFa90qmHlm
CfONGVmQWa2+EH3BgniaVcrHHZYpCVbW7Hm6MVryExQetIm58y8nsxtCqYpGzLQqAtCtpf4BJbMW
W77goJ0zvZFL3F0sC0LfKP1tbaZPNepcm5k2Csd6Hk7pj00GgOtC2LFVrPnNPLIdLF8aPu1OLJf2
jRDoJNNZMFUG1YKb5cauiMJHzAQn1yHpMwn+4Iro4wsrFX3KX94VxjX4annTScZMTzOJapzNZHRn
ABZ3yVr8SyBSop6ujIoKvYDrxD2PIKp9dXiBTvG4SrLNE5bDv+xeJfAcAIjSIjQqdF45AamV0007
lfXvLLfNzGRsu7WhtyChu0LJ824mqYKGWSyVtrayezstNiYKX6hEZLTn28b3ZBl0/vlgMRJKiy7H
tQwmB9g3a4PNqJnUSDcQODdlOfnJSMnGJOTyCfyC+djYaA8udYJfgSvEzNQPgqTg/PAoBvku+95A
1tfCBdpMVTXkRsDNFFz/LK23hLH7PKdV7X2Pr5z7hyoa804eJDBpULWkKHUjj09FH6IznoTh9dYg
vab8l+Dmq3QM/jvJck+LkDes91SFnfGZj60u8gfHiRa0Ykb1r6G6ddUDuxwhsVrmYYLzzbxX6i55
38F/b6bFN/ioXBWkfGb0XBcSb0A1tcSORlGvZBSLnVZqKaWi7euS2swXCRGroZ5BDV3w34wgKg0e
+bp3bpwByE0kf2jVrHrFiueYZoVBhbwm6qIZwMdpgoXeYJzHVMLfyFG7pvixp4674AHSibaTJyI0
tWIdOhLY/1r6WGrPq5Mcvf9a32RY161gkEZQCAe6dmaSrUqrVpnCtt+qnMBLZEYHMR5C6FQEeqlr
keFvie9Z7dMunNvjDTz9OkZYMZCnL9f/+hhoRlZNNJ/Qx0SDNcnQ2/N9KewWp97/4UxbFFsFUppw
ABMCkOjQOj+ewtCAEEhwSOaaw1oUuudu8kh2EbQfKoZU/28AYJB4c0a+GvVYZ6du7MLMblBM+YON
WFRG63iIKkeSyZJPn+eNab2kYveBMBUqHJF1OSiFXOWoyq4qTJ8aiq1p6D0emnFwuf/iB9fpPXIo
bWHewxkLSaG1R/CvwXIr+PwgH1+zs8nN7ffS6K81wl5jg/pKRBYyTL4rEJaA2r9vpun/zA81mQ0A
vaNW48oohBqzkxGwztZF5BzX0EVBvxqvKiYFeG1kKP3Mwu9GP/yc/3+6utGsnfzS8mMGtwITAvhR
v1UY9OX84pu4XajgIDiCzl4AG5eVosrezQtUr3Ob2rzt8ZJJafh8yADRue0ceOyzB0OrH2BuBN5B
hYsvt+wxWoDh1JolEl8s+O1EnvNrMLHtjkJ5ef0psOBEaH9VgwVnjC+UG2XJTbLn7UcXKsC5W0DM
xi3TYfwPz0at+4tZZh1NCa8DGwHxk1Vp9/PbF8uN+NceG/7259Gyc0djjjahPXlx6pSUUPS9pSAi
30UKV4XAG+7lpqoSxXY9+R32ciaKboPkq5h6w0up3sT02k8/pfwtitdfaPc53NqWEo6ozTndKFKL
Ij+/2qEsTaE4KzNL4mZ0iz732+0YP8mK7gyGYINfFlhCVbqgk4LbPjjHxNYqwge8sJTtLrokjN1n
CvmC/7VeloqZV6fkZs74/ZZT/hWefEobz9x++soRfaIx9lGaylkFZGHeekyf/aFLd4wgfW3VNIDh
5aX6se9IyRSEFLBFcZGmPRHjmXHU0fJJtDPieO0Sf9YpKMZPecgflFIOu+8sowgZjNZjGWcETqMG
i7P23L4IWEz95JRtirtinlZz2I2DwV9eh+gYEoTcESMdqA07A4FT++skC6cNtOg44Ng3GurDXRdY
AMDDRoGuEYsF8I/kMYpQkcCRUljGZL2XgayDF/P3fLUw2101YqPEG7vS+lP3wfYtd3BxB4XrrWMT
I7WJwAsdYSqid+yG/siXSYkkFJUgWy1BjEyE3LP6dae1jThg/bdI1BU1ZpwRKqrWItRKb//bpq1M
YfGYpgeGVTW7wcQV0UTII1jnfAs0PnbeqDFzYvDKoYAs1wp6ZKk0ZI1FMCCNLUmBF525jjtvlU8B
KgKjYdV4qX9AW9FsojRQm+HCDDeCz43jOHC6pxOBVJgjQs5xmHfXVvjWsBD1YhDsGnep8z00T1QW
/F8AKWexzV295Nd4kpU83ZBHRAUjrL+zi5bbtsC5zH4Fmdt2h8hz9Zi4Pzj6iKSSN8pdNc98fEmM
7dzcr14L4K3eRu+L3mFAVtH+DrzjT6D76/5WTmHx/JY7+QR/bXCVGf1T1aad1MMHbtlk7ZafGCss
9Mun4IPqED8SPTnAdA/kKxb1hixkveitUk68FQ5IbeWzLUrwsFlztRRnq3WftU3vlR6p84/HTX62
E6FQqiIemS7H3GRmvAXLwnXtVZpcaktEFW84SCMA+6ClooinEOMUZpentsyLM+Tsn/5CfnGQoSHf
y4Z+/TQ4eaO5nPxR9h2tLFeFBKm1LTbkCyZfytYu5UoqtRCU+SOuVGFKpZI7pBP1goNx66l67Tki
g5CPdUXvUe3seSP4YQbw5rpol8HiCqBZyL8pE9meGy7r7Mr2Ne5fLiCJbG9QVZE8hJ6pDo3L1kbb
eNdKMuV0XBmmFYdEhLyG49Jqi9OyvS2r/Jm9WmeYJlqziFZz7c255sm4COJZBZfGUMmaSRL5wunq
QoQyeuAX0HN0ep+sr6xLOj9UKrlQgNm8iItUF2Zy0vBti3wD8Ciu7WIXkMfcQHJavlLJTMudcwSB
Z6BpoTGINq4AJgrnu2ZmCxPlfO+Zpn9zXLCF/1tZUWBgjGDhk5MX+yOBX1uvswFuXVSif9MX6U9t
Tcb7WjIcI8WQmJXMXfyxX4B0axtofGPizl2Dao9KHjegjxzGfaWYnxMKJuUE+V/nafpLHuEVP8Nc
d8CXwpWGwbx4CX14VA2BAOSzVoLgjU1ca0O8Nq41q7X/XEZisXruteVIgwb2gScb91HUvMXDxEJG
Krj1ck6g3b540E/kgSutbFI4y1uk0yPBe5Q8cRAgRQKla5nHjxjfLXhcY0HzE7q7VsjJgWeLDJhk
nut7BD720QCLnuv/VXVfOPAcCEDINpyN9O1ATOzXQ7JiCTB6uIrgAkPiQ4pMr8IQ3+ncpov5NWrh
FoWIZa9mViiRfvyNzKEk85J+9nRK8NhjEa4FSCe3ySE6FEk4jDqLh/00qNdhQZHbVmGLvjkylKDR
hpKFpCjMIG1SDdhzdpsMHeLdMtt0DjX7oxQpSVfj3mohKjpx12zfz1ChdWKkUm+wLxNpZRk4YGhE
KRU2eUljycLf2JVgpN8GmX9HImy5/qUHNMYEOH2gRInRUrA2Imi4zqFBcZaT69O9XKJ85UuC7hxh
axAx2Gynb9TOKkkhQY9o3LpYH61bmBqe2Jbvd/ihc6ITgJI8xcrAZxjeX6acgkbjZKTsIvrdUDBo
Fk9XBAuxpg3NR6GLWvkjR6gMxBhfkKkBAV+kKPs2tQzxKY1aXGelDQSjuglxK1/fbECrPMeLl+2h
3ArZWFw08+QrLv+bZK21omvYZdfvKR4qUNSnsL+XcP3AtY+T3AUO+tMdr7RLul8ZCWFizUwwRndf
7mgKB0Qbutd/uQXrc4FlO1K7+tDa5U5McUTv3wtC3vYxE0I1QSAyc6MEyrx/dAQxT08K2GIe10AE
odXpGUBhUqeOExN7qo5TPUYcEMO0KdUtFqi9aVV749SL4/MJc8jn4nBc/oMssfaNjTFlH8Fcljx0
jH28wO72edor4wAYxVFL2pWARb3oBlnlynv5UTfIFsqXiHUjw4FG3lHzc4K49elbIV6uvatIiGgQ
hgV7rspqKJhPtMG9xnOO1gpA8g+1YFzw7RPQU60Ho1WWXduwn42ZMxr7d+sDHd1NXXMsQA9PKzYH
/vHXf54zOBB52WOU1gK+Rf+rAeG98Mn6kslWZ7w3QiA13WjmABRYfpeCuXbP7cQ7HtZXgHvQqKsd
fSXgOW4EB8bgYMosfT1ZzrLBcJYM2+wqLpUPctiQ1Elutt8JTU5m+6FAX5Vm5SWZyR7nqpj7NTd9
G9Uq1KpH7W1ip1xbnemwYE99q0Q+75EUF2TJBhkW0O5Vtfz3ynektAXD82zqvYRL1qk7hWK30Wpx
s1n9AsvCWEY6aNooDmmEJKc7Z04BF/7vDNEZ3osX6fn5xSxWahfF8vIK2ANO4iNOfl0udZbf1AKu
Avg94W16zuNgsLTUVvkxHPpp0h9U9SRJ6m4JhqBdxNAZV/+wxGpDStH1M2JXtpcY2wj9XmBcJUjb
rQKmAHA5hp12ZdBy3+Yu9a+4hdEJ1xcZP62YZIzsONZhnkiwqr2Yl1AVjOfJeT83E1vASKMcVuMf
p+Jo2ev8/1mw+HoRUnSE4A33tw2t++8cQE8Jqaict7kZkTOHdfLUcqDsw33DGlziw3zlGR/UOH+q
mE/OvfeSHFAzph1DYyEdqIaBTtdxgNvU3aI4UNeXnjOwmVvh9a2xLCtygWHAerzsb9dSGXO7pEuz
mCfi1jYcZUJl6evQpx5UkHVlyR6ObgHO80UH8yiG9YlPsqdQL02+NPymzRspKgowVAHSoxRPkVGM
Rfv1Yggktk8g3gKEFs1Y2HktjY/I2F4Tmtq+BLUakeZgg6dKaiA0nUskj67X6NRyuhVXYyF9gAXu
EpD0ObyCMC0elThylgXnO70+Svk4lrsvO/7ZTdZe/krPC5K72BwcdSV7VZMl1XnRG6fQ+NXHSKim
t9WcjnpjgxBxxVpsR+4YBBB6KltPTsDNYVC0FNl8nlm55NUH/PpUZasX+96112rEmOhyJSynjprx
jxBAHM4ZTBgguKrwnM2HUqch6KQfBM0cubz0N8Q1txuuMlo3+8srMXjYlRZesUIRi9eIFrWgC1NI
4xgfpLgKOkHB63AQityS4WSQPO5h8n7G3OSvkaTXu8SIJxF9EcKdj/P1Nk0afY9+av7hy78ig8CA
9Us2N1WZL+onOxrDeRLSNGq3VjxPk6vNiPN/vs5KZsWr/qy1nmiRzqamGpoHWzx7VoBWGlX+BvpZ
5fLZtry8ex1jzjxWDCZFzjKrZdztkloDhEduhYKoR3A+JreNaWcCJXiG9qChstc3uW3TiDpTr13B
OxUVR2PhUaK6tXW5+ZiZzA296e3inoGkvPn23eCctilBRkwLFFRQWFkfyEWGe03WU+PML4Sbc1i3
BcT03OYb/OMjpbEgLgrq4IUS9dATloTM06RDF2I2Yn2v5ggwEcVnoZq6VwNC5V0tIS2gT312e3Uw
ZpHug9rtIFaQMb2lSQmbDacq0wUrhFNuvnTxAi0dCr3E3OXRcoO94su/1f9d59TiZDXdXFtqepOh
KF4OUnAa8RLBnbliKDgljhQ3neJ/9MpfqFF+MtaUfMURLIcDagD51upgMoP7ysd/EqgTnrMkhJNW
NLkUr8PgrwdNXiMnhYHTUJgp5aXF6WNixcevFgeQQRwVs5lgJiK3A/KcUYNM9Vxc434gF0C9gKVj
tqTPSAhezr9hoEyIAjcTw6PpjtEh9laYeS+1gegAAZKYs3g2LZwWFd9fZE6FHy8LllrBp+APhbRO
/gcYDdkHW763YS05OjwY9Y7VrMeTGrpGuarhNmHcd0KtBboGl+RcNFL4LkTh7FKmLgcrS5NExb1a
LPJI03EnVJ73QjpWY4s73cB3Omxs6R+Gr55+CD5jSFHjsHJBaa5M9NapLRqLWyMDiTa0827lAdWE
ELrMX4USOEWSr7/qqu8EHzIAeOPUPMIig//yTkoLHZzno4H1Taieh2R54YQsal0ltCq1iRrIKTbF
AGbFHAQ8rFuCvcCANKTv6drfgDFS0402leGwE1gXdEZv6N56eCoI9tfcxgm8NY2ewYxlSGjlSw3V
SgIT2UOxhWgTbZV4Dobi8OXtl7YVxSqnL0bNGJBsSUecCOvjNZ7CfIjDwPx6Sl8xXXrqycokBvex
f+qX9buyKNPdBMuzDA0TGHRScbFui0omKs2WmPYJEzitAeKOdW1wejs1zT/GhMThFHs1m+PwHdFA
fk7m7tUuMe3dC8rORji8eFIjU7EkaIthWWC4MdHjIGPhAd93L0bzFx3iaUP0pP7EfjTo6NdPJeKJ
UJ5wIvnJBznUJbvgfbDEapv99qqJfGtD3RKDOoXohOeLuy+YRMJjZpgv72fOxsVmUEvITGndPH2A
3K7G3HT2UJ2pu56WUB8pE2dBmcnq6noP1/TYN3aMxBskmnd/T+jcd2u2Racuj7v5HvoDStbI9qRQ
VZwZoXLNKACXGKMVdQNlYhvUSB95ppZa74i1LFUd91bHtTWGalp0rfnwGrPaWfx2TpxI5eY5T6bT
mSMgmDvhsDSqMS3RmuSAcQXn4Z9K+naX6GuNcna1CDQKfnvZsug7XUSJNMgZ/UhSepHy4VVu2Hl0
kD2W8Yf4To2NZYlfk2j+bctFAgWFx5XcgOCsFrJB2RbX7vpfjIuQizQYPKdlLlcgj4lwx1OS9d0P
hwdin0BfyAGNRB9fHVgw6m/fZJYKdsms7X+CpfYKMJh6hRY1hTdVXgVawq9PPHIVyqyYgs7urNt7
R2M6FZGWeptGJhCnd4T+Dkyfhil8MfW8fpn3KBaxgrj7RW2qZNa27dX7RQ6l8u+wmZSgk1eoO3kv
TYXxaiiiO62RnGwe+q50NdHq4RCd/UMPfRodXCb9vSlEVbD5o4USDa0ZpOFuRjhje3RUcTpejXNq
Nw76q+sgy4C4ckSsgPaR86GJjk3XqUfEP5kG212CihYSTXb8SYp8+Kzh789CnmuYbJ5XXMqB3X3/
B4Kze9hJhxUi8a81Ge0ss70UdXUBAZ9NjeteMXXaTPa/bm+EBisgHKWM7icKGImUTYUPkR9vyRa7
4XW91DgtRJUU8S7EbUjtbGRSLfCY1jtOr7En7rGLjInSKCnKqHz7YRDrZuudUaQXpd6JfRttrLNg
XIEORLifEtuIr+0p964cJM4pbkC9CIHgU2W4OERadW11ylCFuHrg6eOsTONgYQtwMQ/XmDrwQNPf
pWgu9pQVsgxaZ5A4Jda8ArxR46YTwQKnKZiywl1s2s0Oa0eGqQKTMlDinPOM2IKWdI4lo9k2sT0/
oITHSPpPUHjqP8myOzbq+Cn+ogBkGoReV1/HdeHYPI0wYIYGxBbCv58YmEpEkIJasKNXdVw5HX1D
yiI5YqR+23IkZkN5B+OiP9IkLbY/4herwTW/H9d0WHyxzmh7nHeI4p3ABsOBPqLAXnSTvK5S8yG8
MF1xcI6gN6ipPAxN8g43XPPUUs85PSV5BW4BnKwg/b965mdR7W0mlQduZREUcOf549jPIUuNmTi/
iZ/gwsgToQBjcqGByj+/zHEdIKZ75vaAFsZcv2gJKEBw29B//06xGVDMpsOeCM4sc1FEz6up6bBm
NwuCTF1AWg9tgUYBDECxnXwT6VXMZWOfmkWTMNsBsjs6w73RqppZ0dfqs1ZOeqejOFIEzUfZEYoU
SWGWK58cxwiJvCn3oAQkE5HMyKrpfW/A4pUUCVxQ8qdXC2J8blR39Do5+eUDDyncRz7S8XXg/Xkk
RNzlXKSDM+Gi5itOrsyTY9zS7geZr+7UwBujrlWng+E+u70Cz/qpvJ9shpAW/ea39DqMVTJuvJLv
U9UFqGRPaAU6Rox/tV3eZbmYCkklloRByyC4HK6kw0ss2W1Q5H7C0O0+8AhskheL8Y3SG8CAExKy
qvz3V6WAa20mvm/BEQosLEUQ3SIyYl+6qyNdTeMijFHC5nXi96BsCDAddLvkDHcW8hZWdEcJNIxn
jEbJyttHy5wklBHG362DmFzMFFVKnb13praL/N4BzvGOHHt/hjR3qWk8rFKV6vxFyGQYiJlRBRmR
m7ttMMsHML1VofNqFeCzU84fYWIkUy+1GKqeLHDSe6nzuMv8S5smXfPU1slF1hX8q73TUIZ8bIl2
5iQjdEXky3CnTs85tzIcekR+6rjkYuBsYpWuejfpQiJya6zRKYHAN/cCWqtoB9qyBTvHC8h4t2Nt
GKMOme8LrVOS8+mfMBeSwsm0PAe56bX/PP1WuDrIw9dsrePsXYHO8zT+A2lTilN7sUKz9eG7OAG9
3GZRltOAduIVY6DyQaNfkKT38OUThgpVLBYrjUn4SU9FC2i1dVH/u/YQfWvQvdUhgBlvIO2p0JkL
P9shzBG6unQ9Cvg+w0uCmPt44VPa1PkTXHhEBgFf0twjw+GsQ857gsygWTZZ74zjgMZ1ttdr5YX1
i02lAAQ/LCJT5GctneglLFv1sRtQAQpqeRvBAR66WdfMOPy4gb9XoYj+uUbLZpZuHs/rgvpytsaS
t/exkdxpFjdNgy9YLZcrgx4VbcbvC5Ahg7bJM4U0UKl31HYtxar7BRlNXwd23G0ieZpRP5SGwR6k
9UlJLNj1iP4DWaHA7PL9n4xQs+Lj8py8gUPDnpieqOKWIGiRCiQFZMJ9zOtfyft0tkHnUAoVU39V
geSLNOijcKSkwVsQoYS6jG6V+xR4LcSGZqtpr4AmgUkOwT0dqSX9Yrz9O2EJ/RPRY5zo1MDRqBiW
0e9koo6kt2LQUn/DaGqEB/qCcKvRnG5rUeu9UHKMet3bN1EPb5m+Cz9blpI0HH/KB8gv5sSwRUbC
qpnlZhNJ7IZZMt98cqJshzIAJKJBCX+ZHLKmLQXNkKKim+N08uSADG7DAwgMyoO1UNCpekABzqck
NqCw6QVPWXH8xKX/2L+BvOdMuK6fJx8IKok3yjw2OaoMLQ3CutCXIgAYUsV7zQm9aWlqBZRnngBh
Oc0eS2pNfu049gc5e3YrF8L4XqN+023bK4INrUjBlO16uPFUANpVAN/ZISc6pGmeID4GMGNch6Bw
/Sq/T3mb+6ucPk+swFy7mGGbyhwVyCGrJMo1SKY3ACc4fgj7Jm5bu6vH0T0+FGRajmbnL7/Rmx0S
x0M94EYrUPTMhITzGF9mkvjg78UUGBYM/eScS+LxxY2NuDIdNzik4yxv2DufALr252SEaftmxrjQ
yXAkLOlzwt6wyNxrIc4iDN2SCxRvplAxUNs3VZS3VLbSPRJ3fjZAJ1KWW1zH9crQZ50xZCPzJr6A
AXrz4CzbP2yBqCGn+I/e61FhakGXEUTchSO3v2MXEV/vsTEphAc0YzI+aLb6/7QUqbgN3eRmAIZ/
k9ahb3OPqkEX5bKPW6FOSXpayfz0DxYQu2vu+rQ/tE1oBveTkZbkRKl19bPAZ2nMBZo/gSQu7fu3
wnfYMwxlJ0n9ZytOATdnr+bOBRlxu3xbK1u797abqFOMMrwFOxQCwppzevCs4ggWYp62+KgGNl1J
XmdVAE5w4lQkj9AGTkNms9PB2mtnqYqJy4HZm/RkNTp/fXlnkUkC/kIu3ped61hsY/42edDleQfu
BchazV3SCPrtNPoij106HE4Wv8Y0EHeWO2y4OEIwxBhLOxY/Y9fnr1RMhoD0GDT2l89qylFDJq+f
6zcqieyiSyw4EbcAR6QK/kWmu7ZNSzk7/v9A9RctqZaAiuWWisxbYX4gY1QN2su00yWYxvKsqRHn
+Re1mOm6nJPzNR7uTzYDZoPIQ8UOj6Hff2rtq19EF18/28quCA3Jaqhm032xDV+Djzw9GAn843NH
XvQYgHfmQrPybf74IB/RCXGSCWCy8/2uh8Wq7PHpWwSgAXOM19x0kTgCHP+lBjp/RyUwPHszmavV
oDbilQFe25D0at4k4TBRkBNLUpZTdCQEe9bRNiCmfYmIOzDzmPUeXbZe7pnEExQy0kxcJ93zRPO+
HTV6udtieAeXpC7SR/rmz8lv269P7O8lrqLLLps20umk5pm7Jb8SwWegC5dgsmkKqlQjtFCnqvab
/yC5YSk9z6H6IY9uFkUGw40wMr8wmncV4Qp66YQnmlDpsaF+yyDT0BRR4UFdmgNqoZdAUq8U7KJ6
CCliuB+uqOl5dL1xvERfYbugjXzMKd+qiTyQKfpOA/QEQZBS/6S/jVERlrOWmwTLoDanu4ZC97Ca
xTalXNtX43eXFgSQWZlG5+zYN+lFWO54TZphHQJj7d7fOhXO3G2XFczVWJ9o5LYFPgiGtWiTAZyO
zwpl07qeCrEpIbet42Ql7QeCz5RAykP7wpSBaLF4i9EF1mIh3ptG6paB4adkzCmvUfCoa6n5Xs9B
rUWM/pUeytn3hd6EnKuhxcw6oJ2gyi/RWGRSABqsRPbpPBbn3ldsfmiM7qgjecZ7oEMLdVZy62c8
qeNRbY4i7SoTfsmKMdlvL4FyJuDqtARcdzcR6hZmrP3dO2Td8ozkfdkG+9vHDiXY++zSRIbzm8SF
1qzRfRRCasTm4c+M1LwwnfptWP0eck3ci6juCXFPg1Din8K0L2Ry04AGPHNA41AmPrb91LVEjTLc
bMKiCTSOWN/8DKB1Z1sveBNga4sNQ91kqlalg5fzmCAzyNKReoufq1hQEu08QkDoSDHAKlFYiKRH
VcpHbK4at9pGu0Z79uN0kKhbLoEevdzFPALqK7He4v0XFPn/UI3aMqzCwWoi1OjubIaoHimdkRKr
UTGqqnLGIqy+oKy+U3iu87nK6dFiVzZMOxwGlvvL/MJpaiWQyIHd5Dy0scVde39bZXkXKcVM1mgf
8SkHMtu/49zSMbfip5RyA/j7a4f3UIg9pDMf07x+tO3OfiVXjxd/iDPTTT/F61erKQvRyhmqey00
Xz/pY4OzZEcTPMdfrUeds4II7HDAZjLPeXcV7JTxAO9ihk1J5tB0vViQw29i0g7WKrJwLkb/2zTm
g9LvzvL5/FF6WjpOasUqxnxpswXq17m9Ysh7vGkraTX77kRyZcfUNfNqIJ8nnTQRTTgx/iYpwelf
Jfvqo3xux56avRJ83MI84x8tBIyUxNc1WSSacIFVOzIWJSmuNVu3x5lh4HC0VZ3yzUOnGvRPFJBR
rYCTfA208FoAvcqsjESkJGvzBxxHXg1rh7hp/3af1Lk3P73hHrDdXXiLLFniuOeQ444ZRPcEoTDs
BEZEik7tlLAVUI+jG5wpeuAJbSEFuseDyI8/iewEOg1GCOqWsHV5ssLR3e01h6+M8RZB9LLlCin+
CHP9yanumzIMgUiAbmu39CqDTmBjaeAnAxyau//RyWyWn5kwfxgTv9FipcLlGFOsY9xexYCicPG0
LEFlNm27PeJ7XITrMhucwltZkn2DcFE2JpiR045XhijEiwgWw/Kb8FJbsFKQTgaC5OKbCQM8DyqI
aiKaxhlFIWXhVtlJx003yacHfX0t6ONeHmo/Gh9evaWUg3YL/9yzIFoiV1yF9HCACq4EXRU+TVpC
q2illlb7FGpEwxbceObq5lgNehqctrqtqtHSz0VOudP5267/UFLEoZXObIwI2L0QDT1WTpUe1tH6
whKsHGCTeO5Yhp2MoC71IXprNx7cGKVjPzoTFST45WixpeJY75R/sSb0qEmf8xHtiEDmYoCbDpaS
4JxGnBlDUJYpYjPxji9cGwiCv2lu15H++Tcc/jo5pG5iOrSVsJQyB4hMgk6OTAKHiDJtMN9oWs9B
mPS3SPtPTvAkeAImIN60OEo7qMUPzd4IYWwssskBSY/53m0SU3130pgxQBEzu5I+Cb+e8r1UZmHa
soODw4dGKilHOnkeV8vmMwPJMPRjfXD/OSc/smVrSLyAvBbIEdtodwmHYHQoU6sJvHrcM4VHevPb
XY0RYFwbyxswoEcQmxXZ+X+XRCaO4AgOXcSh0usSPkv6JjQfGBbjgrG2SLI8K3J0Zj8hURYeW+Xq
iXDN6H36MGEKead804ZRja8nMXhwbV7ypocE4AhG4ANsRB1j967RQkwS7DM5PiHknU3iG+gXo6TL
PJxgQmLjMHnjb3JSpJLBbdX2DDpc+J+Ij7O2QfvJ0IfWO1Ks4G/BdPB4aqL8SG4+drlaahtW2qfJ
sXzefZOm1rsxgZGorCb9UKq350hvPlE4cPT64HOBwImSVr5Jd0p1TgyyCeI+iNw0g4Gkk++Kxhny
/NtlGtzZJASYA07KhJKrhZ6FwXtwHjKsCXngfnh/N2iXGmmDiBOOBXZlgVC+uZfk6Na5V0jZWaxE
JryYiAHJfJMf48sVrB0fvaQT1wTXD+WEf7BnXAQTIbKXSAbqI4B+POmaZNSBV4o7rOJrhbAumsLW
XUI7+tIUXkiEW9byAcb8rZ0rfJKXR1Cjma1hN9xJ6Y425Qepbf9roryzDSqJrLAA/ZZou0oI7JeI
Z1S8PBoef58raKTukIvWHsJ8ECraBWfOx2IVe85nCiY4aMBvGEdnTzzwOTAiKt9rdX9A57Ya4n7I
/LL4gDVytVUlMHMqfK1rbi2PobreGvQj9KExgA1o706yNrxcGXyOE1uHZ9eIPs/K0R3v4Cfca+mb
BmO/LZ4jVYcVgsLvwikDQrh+NRFSYX2mjvJjs7R5Noa4IDEnAuzCh23Z+Mh2rwO/7363YrP3CO6k
wDnILTJYGvwT3napts+XBWuQ61t9mryyKTYCz3CaYBExylEInWZB01nH+yV6+2MH77SqtXDhdULX
VPvt2htOsnxHSkXigPMTz8U4xpLfxuO/ubqBlULWaXOUtIY4hsdDdj986n1lsuIpMOeGkUPSNt+R
GbKObbO4yqJyZ0LZq1Era5RUbiT66rA2q2J7nlkJTPPDGbUwNY7HUsnFiCEFbq7W2Uxv9/dgwbVa
W+Qv0fvZNrmtrWYY9rporJLjwadjNlPblNBwoQRR0mY5TzO2ZYzdJsTjQI2qi4XKim8MA/IZi5ED
mbx48CM0GQJm4h/bWnC9s2VhRDM6254h9tDM8WTd3qypQtCdhS4qV3Yhq8JpuRrMI4Ii/3bTf9lB
vmtYD0LZ/DWqxmVokZSrL/E0ejCEAL+MjhI5cuR5v+EDGmGYijXper3lhIovn267CUojmkqmowgq
w8MqdJFO9Ej1RKcaRM6yzM/GyZS3vFYNSm/25RFs+If++3YDuIWMvpx/zxb4JP2J9Spp33P3yaFs
mI7YBK61X0fUEDtARSgaxZrkWI7U54Wl+OtSVu0WetIJplYkSj235cAYCIxEXxEJiNDEZa7t/JSC
lVfQt79oWEo5F0qRhiXCwZOgNqAK7eZ7510AkxxzyIQ5EBX18XVeLhCQFv0gCIrE5J9sUogN0THd
RoR+pktxQ81P1/5wRX4wuX5w0/RwwCf/kKOPw22QJN97GZD0e+WZwCW05lSfxVqs1Hy+q/0WLQpg
W0pR5z1U0ob+7Z/jk/ZiHln/pC4QupM68FIhX08J28x6KqGMpSD1KhWr9mc59eNgW1PGtaAtFjni
b01cnT5wDSykoqCyIn5RR7yUmQb4SHOdD2TcXZlR8ES4wfcx1959LNQXVNelE+kZxcuuKxvtMFTi
rcj7yWOPtLBei+iOJtjAzcbtEMT4ku9QEJcpXy5MyaQspPBmpZVZT7RJcG+59Er6j24YctzfCv0j
57oDCKfN+rE0C5hFTpTiHSL7v+XGtfrdw+1DmS9nM9UGlxLBcil1TmHCZ3EK3uBSb1VrCI2TgWul
Llx0SFBAlelPIsy8rkuVu2VrXgLdIRv2SynDfyY0wklu6hb8tvg1Qt6ob3jAwyf+ys3794EDoWSi
+Z8oNbvZnwCkjtLmABVfSD6KuTeUTtBFvyUsjPboRS8sv5O7ueUK1kI6Qvk493CRFyL9hjc1ZgXw
vNXa9MzeEb7JNWiARzYn9hwEzflupJJyPgFB7WqzQQlG+Hd4BSFyKP5hLP8xWvQo+C+5ZvEnx9iq
Evk6yrHW4JTy7ebQT7s8Qo3kc6MnFSKaLc/BdLR5yX2gR2/l7TvR8PEhQbGNBLqA3YZ3AnSaOadH
cDAHmUgYq/c9t3dyOoH0JpIrparOj8ZAkELB/9I7CjWLft/S8qsQmd2aS18F/vjSdMcEpO5MVAgO
rfzV1Sn0DEjUZiigonGaHDERLClLDAOLCf7+p778gvdF5HIejris9twnJMtg+/JVMeOYqg/d4oJc
p6GfST2pg9JEdspzSeMW8CQ4P9t4CbC0Hnxh1dX6IZyPBA2vbjo3GmgAU2u1VS9DEs0kLSKAKmij
C5593ySaUYV7/06uwtkqzW8ogV9RJf+2XcjmdZjQIyiWw6dqEQwKxcEhU/mShmFu156RadcBuWoA
/CUEYW3fYhl1uhCjg4oigDYs/E32Q0lOG7FP6TUqCjzQywaEpxmH6cpncyJAAe9xvDH6gLPIj5NI
pTxw5MvVF57MKqDfDrlfJRIp6IPdx+G+ddfgNBhQB9wvyH/wcxUyPA8lnm6tH3sZGgUJ02NpvqMr
lxTAnHY+Ji72pnABEja3o6e6XpZYza6OW5jAyZixIwdultGqx1mosXtsQiBEjFXDFg7acpR1hY+0
RYLPCdrj9Gq7PBvtyvBhlrF5rHr/dUyGeQSBezv8RbTduow3mXFoxm3aOemPovRJFUcNTlBM4PVB
EPlHLMAK5QW9NgMWn4X7vXOWCG1ocJn1vjxls4CzXOFfkTaa7zg7NwWoK7H6Wlws35ejb3K8NkSo
2LLbXOAf4XhtJ1BuvzYBc+s1CQK6CVt1bUvCLinXLjJ3E8XpgCtONGFZFAIf3Gd7pUGfqQCu2cOq
b/ZZYIxUKUwjoi6iSS+9ka+sqFMHzA8MJsIpG+9QOaTB5V4RaVJ8yoA+wd7edTNUBfjAGr9QCbGf
Dky+fWtRomtmxeieaVUt/CGFoZg617j+8q7pgn2BGLdrTkVoQY8jjMHN6liqHhg7a+7DYfYhDUCU
AQ7BsBoxT/vxEgLyHMRwpV/NpwIfK5MvZIA030MyTW7Q5E3OMqYoXGQ+F5emFdQpdkVl1uf8k0oM
v8tpTZllZ4R5YSs9nrWmIR3uQPAlliynYuc0YDS0p5nVlSbLxnCT81Rrw4O37K+xlMygMgpWvrqu
TVGFwRo/RrgN6qOSUz8UrOKafn/WsUumhTV4fB18jXxEZ6uu6197AKHWNki78GdnYyRAYllUZqej
vrl8yFo6aM1E0eablkuQasFYtY3a3wLfOw2tYVVCiCapgqIh/tGDujA+O7s2fU23pxADsumJFTrL
K2jwg3eaFxL4TgARIygz3Hdki4o57u/7WBeiOEZbaY4vveybaaY53/yRSw+iUixmkfjHMH5zx048
80JrzHz1qNURd93G6YdcSFbfFq/+hWEg2ZWljCJlxSPFjz7nI9TcYbvVyY6lDrbTbEltH6ZH+cuP
UsGd404fsq1jURYCo3nhKyEYR7ryT5mQd82HZ9bdxI3bnGeB+UQQ8Hiy1lL4qOurwoGnNX7qA6TD
cOouUL/8G5UbWJxtxL/BZJ7JnZiPVR98/w6scdbrtlq+dxgLhawlyLtgz6JdIP2+4A/kNnRNtBuY
W6iye5zxsX7KcJj0WTj7A8mUsTb/tlWLM7H2CCTvinmgMuzY81hQatn5HA+vHtkVG6WLY7rTlsBM
KLGf2tsBPdOlxxLzUD3DJaVkTSwAeHzwXr9RTv3bYLdioaYiw22R4mPm75fWoLKV0cjWpBocczXH
+xR2ckBVBc5i/M3Dxpop2Chv80o1cuH5Jpy0M0B+O4nZIU40AyrI/ujOMEVrQQfXVxNwT9R8WzNF
ngakWsdp4FXeZD8clkSzxA2SMyZeQXAYbRYv/MxBGFel9uCjLZid/XCYPOutjtp/8mm4UPueo2gu
A34GU41dr9CxOA8tN2Ssq8tv1Jd7m6rPkCB45u0EqJP8ScihjXlWPBDEfW4blkfnPfZldbg9RZYu
XJqDqPyh7SrYK+QCVWLLZ5bbbQdJvIt+4LXUnL7jZvSqvwt5dswSfeze6tfX6ouXF454Ppor/w7u
q6Ajq5drQtQBCUD87ipbJdz+1vyiyWNS1uP1iPiSDkqvXUzrLgrX3edGgnlF4zW8b71sbkGZ+9y1
h36WS/wrLrFzUcr9pqVR3/r17JzUYBM0xHjZd5UHq45eZsmPOnvC3B0Dq0cbAhveWxVmOQTUVyt8
FmS8DznOiAmLChWVx1/Z65tQH45n2Mv9/WxdCNsSTJrHVzCpJzRQFB8cSn3BrnVbekUCKHSTitgk
DoHGxnGmM97mBqZ/W2hutiPC1nAsHUuKBSgnHqQWXxpeWOGGQALmMy9v+8ktgCCE8GxNDAi+jCf5
C6xiqyv4qL5zrCRMlzMSsdKYcRTmiK4XIYQMczNbGP1sqX/FwQkW/yKtQL/hc3hMTt3TZyKsO+KP
RYqepffIQ6q/lxeJwpxxzETb3Rrm+IWWKG4D3oPpONqygb1POpyGxiWr7+q+TH2+M5nDG6/QxHHX
YDqWrDaFt9e3psZfYrb4/5sFHp5BYJSpeKCkKmZ+56SvcUEofouQS5tpZ94Bj0ND2CQb8+OjPvlT
fLfcRv2UyCCP9CCdILeA7flULgLO/dA7QRpVw5ohfd2AKt7LfL0H6PTlPVUoYc95Enqs5hCjuQV1
RZepxSl2IZiqGWxcJCHVX1PkrERPCZSK1WRgrIKshfNnUwJD+cbbWSHrsFnw73JARIxdDJElhFs5
3+5BadWB8HYFQCwugNZAZOigEWzJNYzCi4xCDHDATMC3O52crO6eJB9V8v2WUtDjF8eHct1VbnAJ
xhABv2ZbsN1vEwy8bcUQ/NSQ4yfT1tyI8VK7ltfwSMVJ7e5FvM8ywLrtRsE/jFHEYli1H451j5sy
Lf/qsHMWEpdxsFx5FZ9Ruc5+f55SsxWJTEnrA/lbZfYFVGb87TsC3uLfX6h2oPkE/MvjCrz+4QAW
50+nrscUfL9kPLmxAv9JlWoU5XMJE5KtPg/HDcpjLzqntMzUzS+UP5WQTYlnQBtQDeqIffg1SRpQ
YX5MugywvF83NeH1gjm/48nvg4iUjXdlGXoAT6eX4YcSPmzbQKTvsZMbNSW10VdiyiZDqdRxnS98
kt2DzbOHcrNIsfbKlEg6OBbQ+W+RHIhK8zRXryCqExkJ3PgXDTjrcjUK4aP4tPgEeSO2qaExBJah
CamChmwOgRIjeNvI1dKovEUQkb+Xc33yERwDT8EDamoxqTSIl2Q8anFNlNzkrd8SgrEkoNfnOFWN
Hi0PJuBAzYSWOGsp6ihwLWKkMzeLvlF+K9dwP1je+7LomKucrF8g7mtFLLp3Y7IKELODO7qhk3LG
dUmmhiGJK90cAoXlppHJtxD4Z03Z5pOvIVXWalrNPCENvsiVv7pE6DdaXByLJLpTrKo56EUCDezf
ELAx1TAHkAeFeF8tqZNRY21JRAOOcoIMIVZorFvMX6aHbccsGCDgQsvuaSIQhOhnrmw7QRhljhgQ
hp/dyhYCyN+Gk67Ezve+Inp9NyNGMnvv6q5WE9sSTdAXEnoh3IU1jigO00zLIdrBvRMq2VPBQfyz
gEYdq8iWOdL3LFdqKI1+yd6xbvO1y2dC6saprEDLKb5V+6Amd8P70fcRu3/bR2SRCvOER7A5Pdha
0TvHOGUVEVzwqxknGiq4+MqVN3f2ICwjkwNTC5DnIs3ZVVsjaCBIPLR7hZ3rEuF+ME19Rv5ZY0f+
mQyBt4lQm2Zbk2TXM2Ed6aj4onkgkznFoL/CgYryHOpAke6bcco8ANNABK79wrGHmo/pzEKCFBZe
0R7oyc+W8KSiUQBmcv1FKaS+39HDdZx4iNrsTGu7JVGL3SJD5DCnZSdgM1I+WIy7lZwrCLkSQTbX
CYxEHo3MleYppvA94BRZf9kkh347lxVpfMkiE95XkOjXQnWtn0P3x8RYazdo7MgH73EMtZJIieDs
X+z/7iqzrMajCKdvlEXEvCgIkT8TSQNKU1Z8cuhcdHDKuvW+iWQJMZWFLNmOufKqztEsdJc63LU+
oai9tGLXyZHpAwrZXya7BFWsIZfEbBX7atgb/Obn2ib3Gh1nlc74yEUTNVu+YOLyfvjbY8mECABk
KuZDer/lUZDHeD9qVhgEOoBixH/OU9M9z2L6W7yNPDelnP/YUr329cGvFGSnjxqh9v2K9gQ6WumD
/aLyyBdc/XxyQ2d9LxvnUUjHYQHYW5VFyemqNaRCJIggslk/oZjn7nwo6lZlu7O50LZD+bt2kv/+
n87ph+17dT2WQCjwHTw6WZm1ZnUHMsWI93ib65QrjpvSnPmlHKcMMRqqoeSrO5pGf1Wm2dqRDkp+
hUIDMSBG+G2ePThK57Frdrqe/3YhfRZvx7DKSyZqv5INJ2UKA9XI7YNHX6pGTrtI0Irwa5lLpYHg
mxGUnBGQ0D9/UndCY/WrEyfatAX/lyTsv5wMwr2KCiFKfcLBVpI/4zT7toqHnLyDt3AJZXzpgoIW
aqFzkk516OjrksWygfzCkTdnySt+G4RMY3d1DL3+f0FHw2rG9phdUN4nshelnxAGwBGtVvp0ENE2
5fObBdP6n3u1/aVQWHgd22n9cHPGLvFhDCftvrMiDqRWJjgB9qtDTc6B4zWHK0jdlp7vbgAofMvp
PluBzaCl44NkIU90saGFYi0FpLFbUekTEIQQn+xlb/3oSoKU5x/qWGmgNUs3E8wXuOWu49RbTMst
9PoBQ4xuuQlxfeRbcTv+5Pnl+ZwI/yqGPDo5Ey5XUHSPi4yNaz3zESs4cLac0aukr+2qCfBezkvz
7MWJMB6KaJm5vMRdW2K2a66uf+jS06D+JmoSINozUxFPsdfGgJ5Vcqh0HLnDyGqBy6PkiklLjYYJ
r8FlrdNvFTVTE6W8Te1PM2rDJJ2eiXwY9H0dasNB+RYSy4X0SdNSeAVHMropmNLXgrn0/j9eaZOF
LLq7bzizbT4BNw9zIT0C7IK+8R28eErYjA/xqmos+xoL9I8Yqxmpwl83hTpVsLMkfdBl8EQRwQtJ
BeslHGHpDipBvPf0j+ZVUSJ9//o4lMt9Y5tdf0mR2p8MfI/tIDW6GuwFw9YHM1KVo5e0E5rithhC
iRkxRV9UJ+f3withqH/Y/EcMlSomgLRaibQgPH7sduk8G9OdFi6ra49bXEq/lAkaOCgeu4vDVStH
mxOCh9OfF2nlmWiACTGkJl/4jz7eh5fggn6IoaL9fL8p3eNEesyjSN447J7Ja8SePGIcC3141lIa
LSMA+ySELy6g255/ABy5hWVpxyuBAh3URC7eMEZiyPiW2bs8cS/qxwg/Tk1Itl9qkc1ITlKTRK4H
a27SIcfFzMscn6BiIXQQo5SOKWQtrYwZOtY/ylzW7MfDGBldItLNbKvpTHajyU5OkMMbmVLRjj9I
mwxM4ESkV4EXTWe0ltBwyiFpjJorEn1FqYqvGXcoFJ4ue1CJ7duHYB5MMMFl2ZcPbzed40HLRYSp
LwazFCmFNeMVWT6VcB/g8Y+PEdHNzCd6wXJx7OEn/IGo/ixNP3KA1Fv8lXuD+d92Zv72XnYV8FoD
CVFmV410ZsPlTwu5wV1znbf1SxFuvDpUxcCQvgTLTaXRudywCraMuBBzDYhWmxV5Tdt0CVFTe8gw
66zSqbXk9DN3rzLFNQ8fPrqn3Z5d8ySOklFa0by8LSIZ6SX9fkeawWQUv1cRQsa894WmYhM6fIEj
YlOEYWYgiRSapOnN3lKsFzqZkYClqAMSqW9biKmvbBjwGMLa6y60hedIZfk+10u7BXDe2+UKFQ7b
IAyxeGLpZ4DLRwhNGGVOGB/32Zd5GbfM7hMinBh/IsbnkN0gj2iTTnl1xh8G7r115iX+CTnT0WVX
jCElBH5iWTH5LG3gGBZaNy4i7z9H9x+LImcljE66qIZ/G3g5IkgPQHviFKdsQh7PHvIVEvPY7cuj
LkmHQuCrNxkXc8U7BonQj3/dN51BDl4rfsMoToxfEAHsv2qs2a2HBjf4SQjQ3YkhPZjp1dJuZE3U
PrLioUwHX8SsQdl/rX/xeKx6XJXdnFw0G6SdJr12qLVSd4O8Nm7a8CYJQGZJxr0Y0IX0cUTT9FyR
aH8Ux5JjLYYKTtwE8xMeaCYZvhv6zPRd7HP/QcxBPMRUmtSDZG1aEHaoAfdFvvICeDjqvtI9NwC0
G93+ckoo1za8r2VUQCRiiHsPQOh0Oqrh9V7NVjSaY8UPdLjg7Tcum448QPIJ/O7S2EZ5wbTxDszx
GxMBfQFn3ZotnurmasnfbrtYB8cCmFrTs3il9t+z4XBV0Z4pnkLAFtn7d9hMRbicskCtzz8ns5/x
aWVDYOuirkV3LB7ta7aInnPERk0wbKTY3omyAKJ0QShvITMX1+EtmwGzaJsZ6C+6B56Rzcq8nRTw
UngobRrM3/FU2A3fQpbq8aHwIp+8dT5wtxz4mfMcoa++Nw5NJwMqVLjmkEmgxWE3sVg8SSmMD3LX
ETZOYRyvtdUYoVw02hvY5MLVO767ee/NTWMj8bcCskw5gcZEcGH8Fgy1uwmhRw23XxlnA0w0KXTe
BTRdkqBewOXlKV8qmVkagb5HaOEGu+606myUlORfoZlb5C1rSGO1i02uP7ZW5mZ/Hth5T27xl2KF
sTT81AgX13CmKbDKDQs/gxtV4uzCIeIxJkI160cREIeb8MNeyeIZwR5GyTQXw10R280EFhsXB92s
uE/x6PAQoFVmw03voON9afQXjM6pfA29zHzprhEc38orAcVHkB52u33wSXuDfnowSieLt27t1Nu0
Xje67gKa3p8hKLM6iAtXGgV9A+wptAnxUYohQGCUZL/9k46h6xICf/pMbh8I+CX1SrIrzOxTz1Iq
0TG51lkm1MYESpJrUPAQxaHFHs/mAJYGB2FqJVq8OVI43itA5ytBISHzeWjJ8xsPOigOHqkcEApW
ALLBeJkJH/s6/+XeuG1kV/V+jG8NzfCcSJO72uJ7ueeOry9ellkirE61SBCIi7SRCnFG9OnkPK0U
k2aO3AXhWdlcAiog87hXf0/+h/9sttyPLeH4lonCVZ194QBcvcWxztrSfeI4xrFLGZ8CGuc1uBLo
3MqsOnVkKhBnkTrDqdDGl0uf/LD6eyHsIOkY4sKYeSTqJCZFsgcoPtJK8yJihhxtEv/Daks7ZGu6
np8E37hYA137WljCjNeL934TeQBif7eMHO+glFZOxVklp7AY6HTgXgrvaow2bHNz+IGcxs384sYb
gKJaV963oe7jm/3mcSjs1P9nFO5MLWPGSyUCa2KOLwOqMQBymH1AmVpHjYegvFB3Gbtc3Ojkt619
uHROBcSlN6bfQdZzpL6UxzH01neX2jEIEs9oaHI+zwT8Dci4Ut+t07FiSu5rnNBNsXR0bcZRiw/V
0JLK9dXG1+5Zx6j8s2NNwIDvZ8R8wqM6b4wYa5Mlh//IDUdEWURUBoIKxUOP/x4C7J+gC+6Nk8ld
OrIEZAVuz9IyW7zyol9M9GD2BH1OBGNvZTDzmAE3DRwLgunQ22TIs7BME0878yIrCJXVy8wXouZR
dfrikDYwBNOaM5MfygFeF0ulY3ZhLFrxqnrCv/xEnjVc2lKV6OVPOjoJNVUi+hLVEpI8vO3Zhkxb
ncmMPr6HMj+MiIu4YOCLuVFYr/J8mL7/X7rAV8UglToZFidaPBGRYWOkgA0nM0rZy+Ep8oh7MXz/
ypKYz+WFptNhrL7q2XWJSnZtO28PqkDtgkxwqvDHZ3DvB/zmP6RxNkb47mv7cgRYrCLdiqgWNQ8I
OBIDbbK6W+HLztVnpvREnse0nZT7pYJ+MUvjNh1HHx1uIz4aszoTzIx+FOuABcLZvDGjR+r439Bz
BHjQy5uCYfvOIwRFOrQvGDe7Wk3t0UqP+h6Bag+U0oaGPYOJaRazn2lwPkLMvLxfAprdwJgAdcAg
dwn9xjcP9UnywFJ8FwFd0grrfNcyE5t+0YyX4YKyYf3EqUxZqlgJ6FZCyi7noUJZefI09xBpxS64
QoLGtrak7lcIgk3EQYUzX3Ua74Djp1/NKPOc43UdIGTgyVncdLPBOh4xeDvi2Hx2SRQDfGjNLlP+
f+jb6BlV7Qc6M70M8iGNmBMTMgcsYsmL0/1Dm9ljyM+WGJUKsEBMC674eD6++k/zXIJ9A4Qu/+ZU
XA2WIn+p15WWg4FV175HFAMf65vQCrY3JIzAGHkbl3N/Inclu0l1mPKgENLMSesFDzM6wXaLvF0V
QFwQjYlgNkiwC/jFWHS0TxsVbZEqjPOkfOfPw3UC7sJo/hY6LPAm1GINvubA9JFhw2zoq7Sh8m9X
6T2EI6yaob/dKrLQOdr0jzrmyV/3t6IAvmuuqhUK8OA0aVNBVDPEmkOi+DA/LVMClFG4F2rsTT4K
SGR5XPpclSkgQCaS8bCepTRk7n6le4NHbFdedJ7d1S6ccENfHglCZWENJdeDMBWkl1GpMNEm/hBn
6gQOiX8ya4qVTYVtTRq72XzfP4cLSme5frxyUTi0ShiEe7quk6Rkg3k2JpklH1cKsMvDHT0Ar+SU
T8iKHRcOhEWWZ+Y3k9xKp/HVVSs62DonfJBQlIXFQKTH/EXYcQuujW6PGvdpysVICK7/B/aP9GlP
5Pge3YPvO0rizYicskwUAuLQGO6ojbaYbu8WpFp7QqAPxf1vgy26CbU74oD3aNuWFwjGHZPIdeI7
SKkrAVQPDBLPulFGmdNLH7ka6DRGDP3GjZ4g5cp6OBAwi1kd5oPoEeSd+Na9LWRpugBkPIDcQpow
Dakhmz5V3PrWbqJEA2ZbatgdIqtwUYIJGvDeLKNyjsSEYc/lBRw0GPjU/9NqcGiIrSyJPkAXl03U
CtEJMbAod7SbdRSkZUsmiZ42fSOupLSGcJJNn6DcTpCnykk6LCnEMwKACzpMqbkWTTawO5H3HejC
JYWUY1dv4tlDC4FKXfBwsOB/CV0p0CZqmh83SDwId7kN5Z/TdPooh0UDosP9b3iygPuBNP5tpwxZ
mjguet2d3BH8SEdd9+91uD3Mk3bgzLfrZl5aYaGcukktyNafJ8Ox6iPsRyEt6zsSBNC/FtShxEy1
/QXI38JyyacxcX+7iMJXH0DNMElk1ly1B5XaIpIyQ5o9VQytkPEnN3wcxmLrkO+SCbZ5M60jDM+n
w+F6/zL83BtDqasrV29bz/GGo5eowiT2hT5kfZsQUztZj+pjbH1rKPe6f9/4EDbq/1cYLLnacxTm
2O4/byitPDQBthw2uqI9CNEE7r8XFVtcx1anHcC3A04AVs8y/f9rtrdafRozu5XV0qUrgizluxHl
46xw6puRuPZNLGVfck3dQ6eAcTBDKkSzZhG6jApTwI+p1MLW7Q5Plwjeq+MIkYsIXw4AeDmwn+6/
huB0rqHNtfj7FyZF5I0YYZniAii6OAOgYAAECg60DcgxlJTHp5COUCt54VqhOAV4B3I3/Gn47Amr
Lu196ShHyMGNWavtURCJRj7MqGGm2marXIgZjnLGS9/F6qarJeosJSUCHi8rqaWVaUD1LnPc9cLf
oZ0crIcA3xhbMm6zYmDtJXKwUgrP1rEGu0TSuhjMq5IngRMF4/snblqedaMltEWgxkQDmNtT2bqZ
OMXqG+iIWIh3goF4u8M/ldwei9k6xgSd5TvlzgH+rPbymjPklnVMAkmjcjACS0jwlnf2RVIwY80W
salEuvLqg+LdASwpBK3aUXf9fm/Urjh31aL7Wrv62YSwmSX6Z37dS+++xLlh1MUNg0x/dCBYv2/n
xxuEgp/dHXcKkG1/58h7vXtLSU9n3OruMppLvpwKnnRUvJ/WfAVeoUfCQpdj8q6lKDDSnER1zorx
rAqyYBzmndpRKivGmgI0ipQx5fYTWQpK2FCqunHwPvJjEilbzTpFwMBy8s9F4FClpkN3ZFu1iILT
QwFRLxak068nIza7hB4wKLpInkqRnalsDITvwHGp1c1mFGX4Ipc3pfWNSp5DvyqZVbKjvJz1Tmoi
mg1NUejHPvxOwiPa8EyE6dSfU1St35qhqqPl5Ox0MZrvecn0e2ZCdYOZlxHAMdtZ8pBo/hRupH+j
xKnPIS+LbygJm2UgTjd08nvl97DGgj02uP9bb2truPYhlsKhwy3uu4cuITCUgOqdk7MBAYNx4hFZ
RCo4o7MiGilupcO/iKuD3UdTg2NxRiVMANPEEOPEoppUtHTi3GahZd/tAwTC2ZuTZoKAmRRXsuuw
feuqw7pCSCmKNP4xoejF25wEPF0HHndfgutLXhaRbX7ukEJWaoOQ1eV7b1buuZpCCQ3EG/K0KtUe
mjjlAsf0A2orFOoSaRco3g3b7EYDz0AjvfQzNY22jbb7Rs6uD9eQeRmIBRTpC0x4IGdpnAvn/YQu
sQgtpkDwmzzFx0K2W+e3bGesnK/64Xbqm7nHPvzrxLNZMqIOGuoocqCe/SV6BBMe4PbU9f7HdB+Y
cdEtK+mmy5Q/NWHIapkUy23LpOaR8fPDltdV4PSNq9AqN2d99qTXc1lm8HUVLur4H39tku70meh0
5f0ANWhedryzEcfPYdv22KsXD0RLqMWc0l6j3aarh4fQ16td6nsOI1dWVTlrOxXDJDh5HAXRPZJO
NIztjyu8vX97MfOTCV5N0QmJBdO3GJWWxpyQ6g53HYAPGN9jx3pTL66J6uFEcgPliCGjA7mr28aN
BB6D5j726DJRJbwTKyuQoc8iRFPJ/3gKWPSbAXOQNJuvu/bk40+xO5DxRKRjd53MVPrlGFHyJ6Hg
6ZIf9BthPK/gKiXK4llGnYysuMP7uJ4ad/t42ONmOB2SwnhvVoQOqt4hVkBRJfuKRlwQ9iFFtsk6
Hp+UdrAeul1ZaVhlOCqeykCJiXb6cPmBlHdIdRv0/pvhv3ekiRWo1AMynhOqvz75BxtOpFPsDAVT
ZjpEdjcmtj/D3WkUQfxl4U9b/pswVoxfDSYP8ucAtyJ/bn5h55OuE5un76bgsLUsPRlt/QKcWM1+
FTdbaAYtQxjSTR7h0LmnUKgrIBAqiCmCEIt/a5Lh833EVOaMP9rRI40NdHdK+99GqE9Qqns0JDZg
mbR2t/Z9V0Gbm74lq4Wgoiv1dC0jU4gecVUB/1cty7tpP84dG5YESXery5GJCgTUbIEBIAZL8zst
xbPdv2lFBPLIQY+oVYQoBFbZRsMM1abhzqz0w9qfXtp6wH1kmAMbZJcDggdHiZ30xukdCgTqRUuk
zCafi5bBr71cDyYqudf1/8Bmp6Cmp+WKqLG7SZlKBcZojjKjjXXEGovysec440GeVMAcDsrcGMIM
cUIYxq7h/rmU/yIwDOp3NiZiDlJKZMWerJgsrgfB0eYonYz95wJkgKLtvfvhGtmJp4hLFIn4cXma
5Pj8X9NlTVC7dHwqAI9gwfZI1HCjwpkf1gGcKZlFV5vZsSi+R9PDbhTAZgOZXg/kBmzPT0B44UQg
afNiQtSFBasxbhZNyB6ygFS3IQiF7YXkQhv9ae5Er9tO+BBi4ncRowle+Ec7+Ali6VZShZW2TZq8
6F2gIHi2wHwC967JVjjcID5cXRrAIlLHzXSVJTE7zrKJbQd5WdWFe0gxxVzQfpxeWJN3z0paGyYk
Kp4oVhQ+BcLddWyNCGZd7Ue1jTgFlbtg7UYi3CAxI2dLEYgzuBndz99rXV0teDgjxTvK+GYAf9AL
TitGei2R5+PMR5ZFOColNY+yAw/h6mCpCV8tLQzI4ZnMujt5WQbqJtgmUe+xRlSXNkOaohV4e8iS
yMIJ6e0RCLYQwIg2j1L73V8JXMxKC3J0351YeSQKmfYzWkw85S/xSpC55MDkm/wkwCqOx93JB/qi
Op9lS82rlHrD+emgpjdd+nclCBGHlbhqfAyuoCcJ1fKnDImPVNoZwuJCvQJ6k042ZWdfYK89kwTn
mjF4TtnrYtYpesBunPjwWHx+z5D3CfsWeTFQOpkcA+nLcLBldZP7L2l/ZfE8Vc59SYg6Rj/q+Hqr
5kTaiQiVlAi4VUHsI6O9/sdv10HwwGEoROBxoU8HrN34Jz8P89lmd0wKD3IL222MKqMeDNVw13B+
prTNZmV0/RIk707rwon8XglZZvo+JenboZLjKO69yl+gaYJHmEDULW62tZ6ESYJUjbnMOG0v/NNY
6l7EW2tcO9Yctz24xOy+XTukYAie4Hm2AYvjeAWcT5bfTXIXFHdyleOAvrgi3arx10oo5DqB4k+o
fdtxK+/xDbc0Ey6zAWSj7jZHs32ZsvWTOcwuBLcUZKNhb2tHDCOlP5IIpUXhPs9Za2CalEvWjMON
0i39Trnd//Ud+LB7SrrmHvx2rAZLxcAgw9AOFVjsvPcHMKZr5uKH3gIoLqHuiRhHcLu3gdDgDkXM
MLwWd+faoatpTn24NanZjkvS9p8+fnqAvrh9YX3A5b3vZKTqxgDng33ozvxupLOpcQFkQ/wiuGQ+
5wzWk8zROZEavgqzW4KdkHk9iji6bE8ye5qfUvYjUlf7XRZbm7+eJLNReZ1ie9lomgzpFtWsYK2A
qNfcuMfDHj2ImwWarlGJ6AHUrFBDBzFSRkn4CAWE+UkIPrADJ3MVhbFOs+EsFr6BQNWbUUKNmInK
E+gZws7reFJY+Q1xoddpjKUvLY/201eryCD+oV2MRn75oHN6FfTu1XWhG/VbJROR79zhKha8MAML
UMc6Zi/FYfrv7bjF5p8Z139cIDOsyT+iJFqMnDM/xwLidtoqFjauQ9cdj/QetOsLdBc7TCJFSHOW
FKFhxnczd/hOSQaZbm1vxgSG1+5mgnQm9iiCrGMDFPEiDBunXGAYlmewN+mHgGc4GppuTS/sU46t
HX6WbBzD4Kzl8VBWvr1dPMDZ6jipgscpHdruGTRmUJrz7QLM7OmlkPADaWpV4XPID0ieGSPPt94s
XFArHyelLE4oGexhqRawrwLggn9cLmbsL97Tg5nt4sgYSZ0e+ryP5wTymZOXhyqed+8hX0P2sfn5
7d8EU3rkECY+moO/RsyJHQwJzSbdT7k2UiEEssboC880qgxMJyxSQXarqt/LaF+TZgggReozi8+q
dvOx8LNk7y9z4dVLgvFU/VheYK+No4Bp/OIX6zJbrjlYpcegTnU3guZw0AXXibRblhqFQyu1rMkM
Fpe0sCKmiNgZXpJ/HxnPSovM6V+uk2foWEvkYRM2E3CxOQib1GiF3DunlqpCNMmQg9MAVruyweue
B6dCpsc+QWUyTrWa4zc0HRn8Rhk4tTzS+be8hno6x8C0e6fHm46CgRTCR58YXWteo2MplmqUUVbt
VugqZHXJPMxrp1RTPDmLT5zPDMcRMBvTvWEcxayGxcd9hoXWlpo9W2BLke+WxDxVJWxrwjq8wMEm
TApgSU7dGT9aqyJF6TLfuAeXe5/U/dSHjnR8cFIWKdmHVIQ2PtiyW6fsyHylOGAE8H+xTGPGnRuP
7O7saHwhuZhDJQcomAoB1zlUVoW8sGReLypIlcNDyJ0TIbIBmVuv6e3ym3VSQKuzyuLN3uLYIbFO
XFUnrOe9fkZkGbKMPtQxJ8W5ntXsSrryK8TiAU59NMDA/SXCxl9/Jc5cql/VjX4bwcHu53WtYXNp
0XRKlnNbFuxNVoDgIw9YYOKx8LXgP6F+lYrpOFluEzEHhh9zsnoDRnm51LszAxbhBxu3nogmYSEm
VtMGPN2jplfnpZwgpXoeJ3CRy8ZpOziu+V8bpOljZRyIBVQtwmKbcGGBpkn/tdinqRhzT3RBq2v2
wdW5CXyCUT/cltIOyV9HFNXwS7B0pJFIIfQLag9y6wVK0k0QMBRI3livv8UiiiawISbGfKaO47OK
v+odNu70omdnfXe9Tf6OKRxgHJ4QtO6IUONyp4v37ln0Vc9LvZRG1cIrNK5/kcNSHBuGFjeWSUcg
iR7wQIxN1O/LVtkiF6TZCCxs7Y+BFNTU76i9A+GERDwR9fVlhTxDUUQzbWKERSdtyi6BWh8AAfXk
e7Q/m1272D9+6ArU94FSweY5IVTqUbkRWJ4wdt+Z4Tv+z344AP8kWBZJE22FofxHDwEm4HBKyvRI
rpJy8ztgZ7PrF1OU8Vwvk88Y9mXgNjq1n0B2/tqVMfXhqFr4OPc9Tw6vxsWrzP7z4x+hrYCI7/UT
oofDYtUp6NKFIDAFRr8CQG2Pu8zvX57jfbV3VDt2fO5rzuxd/EXaqimNqun9C6N6P6kyzezfNEcH
pwBaKSugikQYW33COsTpV7KTO0c1QGvLFvAlcrvrRvy9HgEVO3n9A2fxuXXH6M+QkuVmAOEz2U3X
IwC5bgHDdA5cdW4FMugWjhA9ndDbRlA2WTkkLvTsOwpVAvLVvgnyMkENMXqiA8tfqLx3/0qdzjzy
P82WyhZ3m2KcTP5nimdQVzRe6Cu/yO3lFkisMBEkLyaUR2ozAgJu+l6TO1EnQO/BpiWsubabReY7
SbbTGKLt//WXt1d9beZlmGzSJi7qrZEklaYAh8isQCzqJFEbEUug8sSV1L6AYWE9gZLtlIbEkSLk
gQhbiGAc1sZ2kQ6LlQaf1S6xDN/CDC+/D34reV6cvx5AWMhzTdCroQcAWAi1ZAaYHZtVNwSwK7MI
3Q6KhuVLZyH6x2RO4UQe/kpTrUU/CiwD+8fDtQKDVHmUD/NHsZcikxkRQM46fJRSVN6TX6F1A15V
+UzDzAArE7nARN5es0lA7ytyo5WyMz+oZMuAks0ZERPQiyN7xlnWXe7D2UaFGeVxQw0QoN36shcH
sMaXDSe0pBOJpv9QvB6BRrTNqdl21mUZB3ftpKWRvAd7YvJq9jNBRP+Qc5NcJ6whRSIj31d4POY0
g/jL6fRBY5536I8s5D/3I4Pc1wIp5tbYVsPIst1LberHZc3/DNYqdunAfgFnyMY7PR5waJkHokOU
lbS4izFG1zBM1aZcD9R87u6X3/WsKFI21lIMnGd2Z7pv1WdxAlOKxoxeNDinWUhnsXeyXsL33a1F
F829to/CZZPvicAr4+60M7dMTOkG5Sk09Q6YT/6xICPQsV7fU3DVno+PP2AIizWLw6E2J1DTYFcp
RuOshZmG1WiM0CZQ6BtFCt5bdKWszXAHMklCYtXR9Ga0WD2CbbNmLc2wTznv2i905Kb8dVfa21gX
Wdka28Tszmr0vL/Ltg0kCE3dFnUG1Mx4ol8b/y8n7syGL7QP0el4nWq9Y1ziBa2QgkClpYE/siRZ
TGfGEk3zB5717LlFFM6nRHFczEGv/K1ML0bPcJC+qP8q/LdbtTr8YLAg/wkJpD9CozPprVHNnwk0
tYdd5fb+BJnsy0NPY2ml0gl1OxkLSkFg7iywcFYkQ55XMNuZ9K8CZXtazDhSdHerfSr1DnQW/f1J
ROszOHE7sG1fDK69nsmMDbBrGKvrUllOfrStjFYoDKSgAD6dgqy/2AkfJ7epSbPA3l8YIJvtVm8q
m1dK+xmVyOpgVp5v9c+EZRCmGwpc6phXFxBv4NZI0fCUZLas1PYnweWaxr0on7rzJxWzBp2KqE7J
efI4g7Vt8NB5wA//fJPnWGq4Bx9VC4fme9R38cwQ3/tL9/g9rQqrZRS3xMQlgezXO91tiqlO9U/N
/bHy7uWCCk67gfGvya7CKWD7w3ij+gvxTKdqPKmWIBjXT6KtZooUW2mWxirBnlDe5KeWm5Q+nNx3
fJ1bKTlEHAefKYzq4SPyj4LtUKTWebye3cGpavgP1TPTCJixLDQ2OFyf87jyrgwabOpa2pl+DjyJ
GuI7aUlvkin4v5haToRP+/kyjPliduop7JVDQqGS4/DjwBonn2kC8EYufxsha5EVKy1Q2f6qiGh4
BVPDlim68Cbe9xfmoO/8GwqutEvYBm1Ho+1hTjPSfq9SspYbPCKRqDdqVw1w0wZmw8qFBkPHFaBx
4oeacwswRbnTBupnecvbsma2++ZM78yQ2TMhJRqc6xPC5rH5Kax4326VGiNaHVd1sODFK1Bs9RBf
RS+9g4NvT27e1U9nz0H2o9zScfnIW5eh836MVhb0lIaqpFwk5nIRgY+nAgtWEmdXsnd1tQFcfhLv
G/KvQ8Uh49HXLeFyiVEda5bBAuJCqNQr/jG+In16tMX5m9UIeD95eqcOif3qryFvB3Q/cyvumGTd
Gky3zdj1FpeHZaZOrMRR4QFBN0K0bxcGpfzSz64UjZ1TZxPMif7KS/5yS0zTpM+BPKhy9wKIRp73
n8P78GidNHKkd06qrayoRti/74I9LT2CZPquTPdeP22Bj55qJDMIy39j4leV1NcVSdnSby476vdv
9ttwVBPRSdfaOs9Ivc7PnJ7v/48HrZVYC+hl+9xymNBRmiuitKjEieJN4uinR5yhrrHp6Z4aUzUX
6Qel5wNeZHdHDdnFZOubQzOQqX8f4hWbhqD8Nv2Ozcci7X793hP2XtzAsBkualkaUUBhnJUP+4kE
rmJO97UVb74FRRZcTRNf49Lg/R+NmRaeTKmqnredkPW87wi1WpVLuJgbEgEiYBOAyiaQV8uYO+oH
7gCmIffjTTT6kfvnusl7ylGnFSEzv3jFZO5Lf+jHLMss8cn6jv0edbpS2xuDW61HWEwbO+84ZDaz
+B6e+PzgXbEX6MlpzUiDFCWfOR8GVG13qDMauQlbJS+Vr8fZATcmi270xt/RqfSyPAnLyCP2LBjy
WprGH5Yx5rYP1vJZeB2qYfup9aRBcNCXDhwoK8YmSewn1nztW/l6G/Dy8SbqfVnxSEKEqv2Kam14
wuVZIWVMkTZXR64FTPM8sawbvcTwCyv2+IA/zeEPPD/wCpRTj9WIOfVGvyAtE1Ow5OKaC92L0giG
+jmoL3y/2uT8/4l6j2IVX42AlFC9rvks3zgvp3xdHWVPqfTvLuO9QTerD5MMR7jnqRosGlygAHzY
PZc1xV/qMVmBk5Bn4Ge8Fc8ODPwEsl3sK14ICRf3H8NACp6y+EQqheskUqT910073va67oqIfnEd
kPcyMlGNnvNFkMegqui0OtLhOXTRwGuqsQocPmMt/IxlTZ8vTyoKIv0niAkFWWEUGpHYnT3av5pz
SyJbm7OuUUVpU/MF5bjtvclabh67R8cntqf8pRehhbedR5SQc48H/HgfTTlJSM5cIMexL6f+SVUp
3t328chl8vKwgET7eh3SYmkDImQ8IBnxzER3oMZr96bvpXUqvzZrTiG5u0netdK0tzLmYlluCK5e
Nv/IBZmuAdGYt8dCxzaksbz2s1eLHWrDVbEab6VeJJSZwcaFYbITwErEaOM2ju9ESUHhBUtQ+zBr
Y478VCwdjOLEcGpDQ/GN/BkrKrKWj3DOvwZmdNqsmGZpQJuMmhIZdDNAx6nEQCRiZb947a5xO7Vt
xrhimhn4tOw4QONdcp0dOLOqF+Lq0upRjOor+c3Qr/HNZN+KctqkY6v1MZ1JJgpsd2wD9o/6t1WS
mMN6msDIFZla6wflMui/HOv67P0omhOP0IYk+7EAyyxvRbujzpYpJjraguzzqOvXk9IFZzNb3LCU
5PRMJLdzpY4gekxYErGxoWBkMjYgGcv13e6Jk4xw96ESYRmJlr/JHUI5G5rGCRHdCe9yJqfBx9He
A18/cUWszFociwVGj8vT6bs1CMULHnjMjhI3eqvEkkZoZ3B35LKiX+U7ZjRkER6shOGLFH+YxWdw
ltIuO0L/OjkX59ba4VjBy+m8Gkr66SKX0Bgb7MoKwlNb0SnhIEGsh5xt1M9vTxjF7s4kxwQcGnZG
96GxEd0oRXwLyQaDtP7zvnxMQnH5a7ZqKXzOt3umRgG9HynLC8JiNwEtAGmHGR1ixH2qy4UtqCNw
DsV9yTQXQ0dBNY1XXmNM/+/n/sVfRC7ByrrmBVgUbPjov3gf2Ai5TE0D7Yw+JiJ2PvQzuccvxlyb
hgHWGw66yCO0xWsmtPgWZkC9FNsB3OzoIi+fz74WGkzQVu4HdaeqT6bppGuLPHwuQ5oS1pN3rDwt
KuhatmQ26UnpRXBps/sNIMoA9KeWdYPFXBG8xOJJJJDcXD+i8lZbkzUuwr39lPUz4jMh0BMn3zuS
B3DNAkFiH7aegU894k08DeE4bkLcDE9bsuehtyGQ4c+QMGW5cq4Kixz80+aVIbvEMGDhuDfgPXqn
/LqMh/cgGvwK3w9p1JJq01SvECgODXhXKRsGefK1e7wnVXAINHc1j864wxMeWQdjFKjLsQ9cN7e4
+UKQa7jenp8KyBaQoMYGYmNJ8WSjpftqAlp/+oT/fFyuA4LgD4TzaEj4qWSJKKTzD2MxwFGISRFV
jL8D9oEuM5eUEODeP8VKqYs9BM7pKi2yCDqdg6GUZRLLrWNgpWGq69uRGaTku3EE2zH1UuDkoKHb
eq/POSnSAI6vk3xJeLeorAqY+dPptNpJUgUO38ObdmN2OkaopxtdlmLS/dCJ++7VjOWwUJsHY76x
t0JfpU+lKe/g4pkOlsLrMRWJJa5XlSaKetTENCUo9aY3e1g0uobymful3Wp0vL2mJQlG3naFuXck
7pPt6e3PGqMf/tFt+JL5lcNpi1h7G3SQ1gs3scr2YdUf49HakHWESRvg890equ2dgDv5nXemelQU
eYz6DXKvU7gALyRTBSfB3s3YpNS6VY43ajSOrlyRkAjNrRCscp4JAUfcTWHTTIlnQZmbxlfXTXO6
lItof2IAKQFG0H0ZqamRJC7ey5y+zSeU+biJ3ydPuvLvvykN7BIR+R3e8IGR3VZQgNGHb6hd+zEO
sbDF2/9X4XKtdeE0tVNqIEtiaonp4B68kchaoBPnrqNpaELscWfj19FB/pSWNG5oHIORq8cg0Zjn
Q07QbFjKgpVCqWb1mwdE6pGqk9/knS4CTmAQMZ91XJo92/jY61DPTbHshmyrAwDKUOaD9SEq69hU
Ql8qJ7Unh+pb8coaXkh4rUVMbNPnqnzu06TLgE/kU7yGDhaChzV9a6/puFC4JNd67jdbiSpvnhLL
9zhF7S4fdYOL/uYU+podgLuAfTvFK0wj3CUuhTT93rHjhuUVM1/1iNB1xJLHtBr2kuERYnostfKB
Dd+mnMTn+tBQTKs4w0p/cMTngiE54RIvoxXKnd5yuC9bsxl2huEQPJxAso5EX9FPFw719lFB6kIo
6vSsfD97u5mKUh1M2i5OzTQmInHOB75CeQfPraMS8bTcQTNUXp0zfXHXw/4/kfh7OtqnwT05HfAA
nF710yoVp/5jvWdHyAEdd2XfZULGUTsEdWezwObLrsODSN4ppd1rVG7fOUhfW+Fc7WmQBDIJ8C45
rTATQH7JSbEZOQpWT3JK5TtUewITZ6a8DRt7CWF0zZinx4nevyYzqXrnBhwZrF9nw/OZGrfhzqBN
pufvQogN+ZNaXP1GUAbYVyImVEswS9cql2mB0+dyeq+Y1NNDnVOkLxuGTeWm2apVFw7seAkpzXmr
OwKnvp4uxN5EU2r9ZqcIj9iaFCtd1vcKOhUdCH6JDSIxDS0S/o8WFmbHhu/eghV+KAS3xkmxxlKQ
8TvNk7mmf7ZNd23SmW/HdYHJR1YZ09NOiFfUoFo83zEdJCfqePudx6Cize6w88O3G2pfCDmne7oY
blirQV97jbTbAl1Cc82GFGvoYkLqanRZqIc+bJB5cybcDwJw4RvQfG0VZ1s01MnjK7xJaG75kE6G
y7fmSxVn3lSDWU51FVEZLibvUI/YiS2apEDI0YabqEsTCuN1bWBfYNsW79sUA0Gisi4p2BZQsyws
OkypDLRb0iwPw3L8+gDsHEwSFctr4ssqJev/V8ME2QkPWMtd+RktLqywzN+z8tKKoervzPyOPspr
e+XdmZ4/xKd6n4k9Y6VSFIkfIZhnLUA0E3xOyg0kfImsN/ozKcRMGPlpwLoziGOeUElGxCuk4+Hp
GgW3KyVFGUn46YApDyIsqdCNFEXsALt+om4LJjeBofCtvG0RzEphCGRjOMeDIx56lS73yzfyOYuz
rXSz/2O1AM/T2g8FzkE0xkHJC4+TXz/2FtttCNxS66f984HonkMR/iI4Cb3e+gebTKIPGDFkvuiX
KSi4ISOIlLO+Wxnj3wFfg5N3NXtBjBXPV3NR+0DUo9cmoy6Rm/VMol3Xa0lJG0LVFOM372Pzhqfx
Fx0ZbeXdlELvwgatIJjUomvTebwwbj7dCgQFpGcm8/wM8UyDHlnl/5pXSacUfSolD/WHKrZe2kc+
adq2z8rH3kB39Qcl7xxx0d3RH+3OVMVPLhGEccqUKjdEMq1JcnlamMFFga7o4THTuxVray8WS2oT
PAKCczDdbnDuHZTRUnLt/zlBpgqi8rmStSHWTEJLe7o24BuWCJ2YlhbDuF1HWRdnOPcIoBhaKSVw
C36ELq11CdYxKBHSxtuRqmJVN0jOfpnDk2/fO2+zr4YpMm3X+P89fwO/t0cTq8bPExVG7UbD5Af7
TcvoOmBql4R/4vNhIAw6toWbTKkJEOzKQvmiRQU+/k2UeVFU/smMo4NImu4kkMchgBJFGjtota08
MGI5D8GnBf2CNC2Ku7I0bHOpX732Z8F2S5d4i+VjDiARcHtozJ/BFU81BNvT8AVaSw69Jttb24n5
4VOPcF9CVxh3rb80IiymOkbhEebItnx1H0m+znzfLN1OdabsTPZD+B5L+87APPXQw4BsPL7svNu/
VElg6zKHHo9wbqTjzi6f11wwEVGVSLMkLZgHaB1ZcvYZKhI68nWfFTz4vX3H7OJfvx6zbrutIfUm
mrqosIZC3h/Hf2/069ZCORs67xAVuYOuWjQwW0rkvUusAhnIZAnZI+2dNYWrEFW+/k01v1tZ4uc/
gXMNsZ4HkYSRcC6WeeJ2458M/M0y2FG+Q1nKZGg2xf5JsJMfUGGt5e7On0KxMOQBOusPQfeF8HBt
QmuCIUxSPxvlT1C3HkMoqI3mRBgo4sjoEontpWHaafxhuRAwo9ngidFEJAZ88NiC6kAOyhCuZTxF
hEo8LILDmwnHlBNnaYO0yOCT8mHCgZB8oRRbIso6syEOuboREGyICyNi2iAV/MWkaPRLw+xI4BRA
o/LuuD3uyzqOCa4hnkc2hgQ2ltmuzfNw5l8O9mvz4x5iwhcdqmbBgDI+HsyK6lvIDp9TBVVXcjRu
KVcZXh68BeoIQoQe6d4/SzuXDhxClDbkqJhY/vICOdiTF9YTzlOEbcuAikpeJud4ECeTj6fvI7Hq
v3AMKcVc3ustRy2ivp9gKzP875niDp/G93b+TNKX6KT17jH0v2cyfgOjUVSXGc3PFy47ELTpVQrg
5q2c7+kx6bdVgGCpqfkdL+c+aMJwLIqz6eGxt5NzoB8YRMZ+od+5hmHzrzFsakX7ljWx9CA3C3aW
z42R2215mYZj/m+U5+Wb7yu5CkaZuJy9FoHLRujhhNTirVmJnbz+y5TgxTzVnw/QQLYsBj9Pum6h
/xezzObBdPe+ucIiTnCAjNvqAZjueYvzaKj28OwrMx05JLKZyExZx0XFm5iwvce5g4AyhKr4Hwkq
nfxO/vxF3cVwq7/X7CguPh4TCk8Fktr7eqneUoqaDP8Jv9+jjDe8n44aTkZgIz2ACZmhMVlhw3/8
PRxkkcE0cEKjTnEWAZzrqn+ij4gBzlOE/bJt1fsQi0feDx8MCnZqSTUZSDx0csU7YGg6q8APfqUU
RYCNz6iZ4Q0bDCAw9DiJEDa/iGNAIiN6QK3RrMJ9L+1PqspvTof67H60xlh6AeCQdzqsXw4EIlis
YkvuM4io+eXukV1H3p4TPAlBBHm93ubBQzXwWsVRy7LAOA6e77anJf6tC5CxZHYdn2UpEjHtmoE3
pO0T/kbP+p7l/kVJHBY0HAogAj4ZcdeuLud3sejUgs+nGEwCF6i9jnA3aQFFoHVkq5MqqvD+XZHR
TJ964hEztpSNO/EmWtNVDaC1wAn91lftxJuY6FAcwzsDKVmn5SJd+pvQ/veYMTRluF89yBpdkQRl
uVjEixFBGOng7igZGlnDWEx3v2LQGjb708Mnl695fRYpBaX+n1MNufeRS8iJIHdCb/uehVai4Bew
VmRUfyoGEa1CFWUsvjGWNbt93ygUw7pdepG8Y+eyoxnxf6XAlgbNljHEQge7BiSwvYr6ETLaeHgL
vRqGFFMmLAJlV+nNoHj23xXuswNxV5WUgajgO6iQ/KyiI3gP23TM1RVJHdjB6i134QZwHXreV5DT
r9oZ3NnKziIrWl/uM28lbVh/gf0eXWLRoKgpWl0lyL2W4xSHmvt/uggQzVNjvDjOd4OPoAccOZLc
RRfZHbrES2n/qp4a+JZYZStf6ORRMg9kuLgC+GOiS5F9tW4CrQNy2gy33ns6VuBIuFHGF9DjAmOR
nZSiqkyrg1Mv74+lLoO70lyirglE5Bt/0+N39RNETccgGdiZ3pxgeWrECK2VIkMdjJzgcFzWPC5r
0Npuq907IqZnkJwCPOzGfEG8zlVpiSKllX+KBDpYig4ZTa1XgzPDMD6MUPH9HY2dxRmBUEMJkioF
7Q4r6y0gIADlyapntrYbVADvnmWa6+pDEtAPfEFpidggHjRCLB2+jJtFUhdbODJ9+RLYR+zJgaHS
GCSLOJe+ESPBf0KRgPet+6Fzy3O/czkhAKGjvRRExydEDkJ/PJt0bct6hTsgdpIj8Kz5tLvfTKgX
RkWToqM1BBgue2nBlTu+b66RuqN+4yNxON382Mk0u1Ys6mPEoSNQ1F9IHQxNIZMdkZbTO/8DT/VI
Etg4wWckWJewpVp80RoOSQp9YyoykFPzLQFT59dE38zUKLKMsE6XPFavzXWFFOnb/phX512dGBqE
27mMyFnKcMVySiIMO99SPbjTdYaF8xoe32mLQ9unYRWr/LfVmtxsoBG/8dqYkzQ4lSskYfeGRD/q
XVayur4H0IJd6HBybxv2elML+VYTTuRoECx0bDsngcS2mKGmrmYa9bTgaWagnodZW3iQoS/ulQ3J
0MJuFfx2SStqMeS9/zO7A+DnjQkwb83NMGesp7tkD5mdR9PufMHAhV/nJIZyXfCeOWTXxlYLBAh2
pKUVN43c5cLPW5fP05rg2sj9tsShWEcKjfIS0lJSImkw+neOUtekWICQBHhiYaGoeObqsa5Kv+J0
96QCx7CNS6vzUf2Ybq5VADgdL9lUeF+YKJfChv0iD2TUJJPs6pw8MOydUpTAtR1e+3LVxI8tvTnl
Crv1kuJ8fW/u7asn5AhCBCtOefueXCol5dMZNXBvuv/oj05hctQufAz6qvVoPSuygxtkOeWeNjtb
WOGg1YL/drWBejl59udqaCki/f8Hp/+ObETuOeWTNVROV4B25AhyII4Tlnr9OUfdk3erTi77lHK1
q+z32hKyCI4UU/mcwdkKuQpG1EId9BOL4CC2C0N4Oyl1Hom81Y8wQ9JfVPgK2Ozp5Rv445tnFZJJ
JQ4u8SRuuBWDIHVZ1vhO7jZLaSpbiAJeGPozLd8EWuBAeNK28kATGV0lGM2kr0L/UFsVMxoQKd0t
k8jg45/473ZByzdAcZtVNvJ4/+yzicvCN0UCAEdQPgBfhpLWjw4A9/Ca3wzAM25EHeLfGI67oDW4
VswqTHSBR9diEoCIPA2m4eiK9XOsW4IYVm8t2r0MYWWFsnXsvr8LjjNucrf3nxbaYKFYzBOGGUvQ
xnAle9+iREL5nPWngwYnESFlN9HiRwoRkH+chlg7QV7rgtYKT5RbErAF7aIZUTO/Ziq6uFCqmygD
UOrlAY8pde75CTiMxgEGJmp5FgamzjsxKAT9bmc8gZB0acF+Xp4HGmyUclDKxJmeyGf8wofMYnRv
r5gmpmffV4GInD8NYxZ0R7uVzEy81Lxt9fMMPWIyWVbjiWXqXeq6tI68RTwinhUJVvuJMvNaG/fT
/ufkG62ETWS8MHUkgeektC7nIiTetZEL592l8PDCeI70K6PsqVVzB8zoKBYHszeM04pXb/RobCCj
GKAVq6rb2v+4co6w72IpQ41Dpeiy8AJ4Z4ojIMP+RGogJhfCF3qtp9ubOCsYNz02gHh60GzxCRTf
FKaWHfsytu47103z5WUu8e4CVJgyekW8UEfJZHgM1dCupEPWYVjoKyfIM+jdby1CCleuJHpbUdFT
oKoVdLUcrFKY4PEqSujhUY5Tpao5SPf683IVM9tcd1LwbUD3fL2qrUIH2kXI5ebyvAY3U+JEwZw7
FxkR3x95qV3CzYcieOIw1MDfnRkOfAnihedt8dEzxkYN9snk9MzI4Wg1oRrVtUEtJ0mgoPY5FRF7
xTLswopg0RWXIogIyLNEyBbeJxMf3lP9cMvGTvFvRW4P8hQuoT04o3gEW4JUHVeQ/c3MrML5gnWf
8Q89Ky0sLpZyifObMQXsncOh23Eiat4eObn4uMX5c4d9CTfYWlZKVQdOSp+ccEiZuj5ir/vX/lG2
1wd7EqfCEHOxi6rsTy9/Tk/4g2XlhLn2Hc282exhIXLK7bAU4/8Lc1cad/X8k3O1uFuLxDJtLsNx
8dpKie7A7QGu6/npVVQhtHZ8IhMotJl6S1G4Q3aBcguGPMr0dCmS6r0nlH5LxYPAatAHILvGvzwy
iE/GwNBHFj7WJe1mkZ5kKIMRHBlW/oRmbJb6ThODm6L+2o1ZdkVLaZYVQG3HVL0eVl144F+68gFN
kl44ZGrIVfFbs9eosY/02Xm/k3DqU8vY+ZwlzOXBDdTIysDMKf1U2NrVb7pMPB2j8BDBxyb+anz4
DKIZl0fjxPJXxrrkOln1hjD0+3uy09YcSRAWpa5p+ipJj0IsA3Jza67tinn2n8FEiQJom6kN4z1j
T0ixOUxfeCEWWmAyjgGJZEGBcsWGMIM3CcyQ4V2cVQG+x5EGczeHx4Dc0UkKZIQl43o66DXsZCMZ
mgEotdkEb1nunsM/24dSPq8d3AP7Kq106xL4EnlGPoMuP5qQ2aABKEiGuf/A05l5zQfODPxumWa7
tAS1vA8W2faLZJInbtZ6yzMSsogHwQRv4JnHQfVf48GF4LcUGhnuWqU9nU2sVU4zoJ5p2ZPJp2mS
QmFB8iD4SeIDV47q35vTLKsKEbAk1c4S25A0tJ8lZJdzqeGGOYyV5I2Qa0wApL8d+remfye0q//H
8L5fmO+xlqESsM3vnKAZpA9QjLqjdWO+MjwAi6iuox+bMyANkTNBk0piwY+9iHopzs0QnM9f/1SU
LGefIzAm88O+xSgepFqXlUfQU7V6v9BThAdbKpYPrrTUKYFeJdBOl75O04KYtk2jKlPrPcEVxwwN
vq/tR6UTjuA1x2HNID/Y0Z/GnzzBqUm1VM9gbCbmf8W4wjjPmcPZjeBQi3vpIfKcKIstd/Q5j2HP
5NcmUP42PHrlrgmMxAKAwDcHDfkeQ6OC2dZlamiyolXAT2VOd8hefTzahRsJhyuxRVXeOxr0qK5k
2JYVzBt9ydY+l6dVignYb1qeUVgQfBlBz97aPoZHVkwoFdCuhASTUdmzdbdePjXv3TVSnYGi2DS+
lm9EDo7FH8DYrsyfAYIBOI05yWk+bwBM5gxiV76IJCk457taYA54OPFUYFiaHWnxmuQFVtvOrI91
cS9GKiL/dQi4QbDUOZBMwMJhBvUhtNE7JX5L1tSyWosNskXxZoQLQga4VAbR9O090wp3XIWyl+5K
4sudPhJ4J7nq5cXm9s/n9oxp+vh6igKwGCXFeIZuZQlv6AgkNNgAAIR33GUol6O+e2XE4c5FU7OX
nGfJevqtMgoQMReTuhAAXcdgXenxUvgM5FwNOH0eI4kCfzbdx7ZUWwNXfZuSjUwEf2UN34m1xp7A
M0lTo7NX7qX3qI4Rwg2pI8YajJGMIddw8sKaMiCC+0ow5oAnpKYT1ZtHEmZjmLbSlvDw29I4nKoQ
NFa2bqAZnBfxsUASykr2W7SbZw4Dc+X8oVPIK2qhZqfW/f4ynu9iZHHMJh/vATOIPh83r3DLg4ne
LFrTNs0hQt6N/pi0rMyhXE4QYD6lfJPX64Qx50M/46unC4dWgarZFNjKa2yQTjjuZHUpOPUAVV7u
AOihb3hlZiv5AlWoLzX4XwKZP0SXrcM6AmUwk2C13KbvTgFKk1jhMpmQxPx0JpF9m6Jsw2g71YJs
9UmAO+AvJCftZDe8/2B/3MkUax/LWPlm8J9PlLiH2pBffa93VtkEcfUubFR2fZe7RVYRHfkZVU9F
10OsxcstwPaz2lB/K3HD0l98aWG7dqVHCg0EMbZcwyCaQPw9HtqylJyt0Q5v+zrfxObX3W7qAoBx
f2NweGwbk4g1NqYq1KJHtRScIEpJCLR3PT/DTFbBS4M8Lk/ECNTjQwUgYMD1HWhqWkna6HQN640M
MO8qIh6Mcvva+ND0P/UIHg/8KWp99aJUcWOMutiCNg6iPsUedzYKDetnXuC0Yd/qDxmLJqGlIGRP
gPGMvNW+VHrD9K2H+ug+6d3lw04VZ/D05ARLlQYyApcbm/48Q829QnZl4VY99YcADvIbR4z9FBgk
s6jUu6rpN+azaSbn8cWVHRwvuwVazJpyE4tEM2/0SS7PjctxbmEEp48wpXYocq5xnFiixGHlOn0V
8O0oWY04PnchHWaKUoHNX/8wEL4AAHj3wxhlc4uSQsovYoCHDGR1/Nv+Z7KBJvv/tSg1A7/7hCqn
f+fabxJmpmo+BqGvdP6lsI0K2s3y5I02wWiytXzAFYIUIicO7CHxRSefkZ/iiecgX8qhmWO2WkYK
ooIQ2bnNHmTsGNuSsgwSlz3XNArFxxPgdQs4mOnsNbhKrE5FLoI+CZNFJit9jvaR/InMJmZirjT3
KT7uADGZ9xCzJUoYWAlQa1/ehiICHuuxeCKSeQ2vNKVkJ1whKHOxdRnvup068CscY1bNSGslpEqL
lSXl05osW/oNzS2ptjYPOiY2cRVUpWTo8//QW28ArH8LsqzbEDSPBF+zFlIRCmmZBo7TS4SerjV2
cp6S4w3PkUCjkRZnSXfOjKR8Lgr9G8eMJVa6CnhhQpSZlPuZN9DkiU3ENvUnolLUgL9T/Aw5q+1q
pGNl1h0wxqhnILowmfh2wdf0ditPdAK9gBmly2ZMXMgNDTM5riDKouiZqZR8nxvuemAS1EeVFcX9
0twj5GOfa1D2xvrWinEp8fP2vdIBB4d1zvtrq12UNEjBUmMdvNPPDXS9/xG+YAJCii0g6VSyezNs
LgBa28CZNuBW/KcwhiJs2mcubUvRcYgFHo5k/PyL/XU8+G07llhgMPt6QhJLyfkiyE3vqWpZlCRw
pEQoeVxbEZih4TekM1So0lhss7rtTqZmklvWuuEoai8nZZPHlQ+RbFA3xf9Rl+Ao3V4P+YiuoXSu
sTORd6Cb/4q3+ZJQE9h1zzqARMuhMDdypyVrb56JpdLyCw5T7LVnxSJd9YRloDKVjOapH8jzieEr
bP1leSVEdJUd7hWS0JuJoxW2V4IylsUdWpQpDk4SL/8y51UPyqtG7tCRAIbwEtQ4PFhIwmw4KNwG
8h6ZUdHa+a4hke4JwT59UtfGvZK7htfs0OsBGWK/23qj228BJJdyvtXEhpEXI5R6gN4jmsOfvYmp
e+L4v7QFD08dpNrPq7y9twfFG3kXH+M0j6B3GjiGZN3MGySABvi4j3RTpgLeZBsu9az4CM2J5LfZ
MveoWaN299BbyZqz5hcgFjJDDFVRlK5NQ0vK+LilG1O7NaSoorX7Xc7K//F3zhibbOXy/ckm2/FP
v9Jif1R5DG1cvS5N+FyX6wsGP17GJyZTPysEoIB2SejqWyropyTn/h8otlqdj8m9E5qv/9Pt8Qq9
pjVD/+Wzn+9NW1j13WznnzB48ZkHY7dfIfD+zlOPHoPObeLPJCfFR1THOiBuabwLioRmYzchE0e0
GMjpkyQp+8vRICBVHkPqAwCFywW7gu7fAFZ0+a4p1PGynFj77LZBcvruax+NGnHu7j6GL9KEnlhU
7BJvZxWgtOIqJ9RpdwshaWkyuKmnIgMdGNRVYErRNCLS6d6cKaObuSforRc+Fiitrfd0KVSl/bgB
Z4CAifMNEM/Fl8gY6jYk71rOzVTU7v6E3zJ0zpMlODZQ6WhvX31OasaqcVQmexp+YsxMHqSb5PBF
d9YWxHcEulpLxadu0DhKXWydks/VQoKSR1+HTzyIvMqQTi7QSMoDl55jN3PfMgdA/sb0y9wPjvvG
piHbXSEbDLlpj70zYhhlIOSB4EjUkXHLST8OOWQIGu19FcaEfpAoFwTee2CvPk9XukrECQMLst0+
VYVT/pKfFuZ4CAmFZmmcgHH++fYVALt/uZfa8wYYtVNF6Nqh5dqLJjM/FSjRCjlimiejHW7Z1ZkF
FFoZOIv7X50SwvlgnrVauO2SbD7c+Sum6OvZra17Y+bCqd73G/CyZTKp3NQdq47PHhW9iFByAfuG
Pt2ahVth8+cPFyyYoIzZava5wi2+dyrGV/W7rjWmjApICJYzcfP/FHLFxpDjLSetQFXaJSwHAZKb
mfY5rY7/73BGNDLCXHlBK/lb+Er1rxdBDpfaISmzFCLPHib5WsAjwp/dQ2LRnMYQUuW5gTOVzE60
/0HS0ZDMjVlbJWzX+s62hmlrzN6y2QNFAQdcDP312N67SnzZtUOF3YX3gMesWnI5chfkw/b5qADX
4H9inS4NmbZn8KzsvR9WZhZc7TH/9tvxTFmj/5RQbPUeAYY1AQH3nLE/+UQVJBSMhXuIZGYma+Bb
HS9a0/ihXrbONED7kpCylGZGjtQKCpYT6olYp78fGPYayDSVMGoixQIDnm3vtg65AuHYSj5Hdcc5
e1Hh/2+kTLObiR2QB1b3xxbSwK06xxwkzYinaKOuNP3fIX3eI1IL0JpU8SOZ/tm+WjdBIqSi9b1+
Ed4zZGgWfR3Z3AFIcs6W9rzohWTI00UiIx9YmsUEw/qy2nkX1zbq1VFz6WrSo4pzinuhGf/XrMaD
3jYKhFgMWaoyNmi4OqVGjHDrHv+72/gA/36IusBgibpWF+kx+Jcat8NtJcfWlu1J5TGMNC7q6F0V
AfgxWlwdr79H8lZF3RZXPQW4U3hvdqdAReOZ6tB5bMAPT9JuqhHKe8rQCTOV37WiTV6iigYs1c6e
s2xxdHp85cq1d4MJZhsJdjoG5RnCPV+4UXB2htzvVOSTRbm79esCsIdXZ0m7cq/HICtkZBZqS00w
hVDnrBzZTSk+eVlEyKwQcM9i9qo2RfaeGZJ062cihHLBhM56CRq3ENcDwM/k/vxgbAZXHiyeSp5O
nH1scqaRLWtrNlYkbmA8zdgEbI9RYwdAIgmGemLv3HLeqPzFEvnPncDwCjq+NBQd+sKGQYTSfv24
jUlRZMpAL6/Lw/fGuSclykNjsKl+/Ghq1jwXLMRflmHe5X9g/JzwZxYYp+qVMsRYLRuFKh4bVc1K
kCAyrccjgts10wABVJzZiwRzMU2jkkIwIgwzTu7sCJGHJMXJpcwhMw6NOmsP5/KJVVCwufYcgF8t
t6uHrZ/z76644jXDxZfBonGarC9ADqC2x0a4jE4uu7Z6PC70t57qHApYekxzQZ+w4o9uBTslYQQ5
uzCD15IdnK/UyT/PctCimOZ8ujjhc/UrmZkEGdyl/QvuEr9Hn1G64ftSMrxZalGVLDXbSSDs9BSy
KzbCqRescKBVB/qoDA88veir0fuZ8p9Oht4um9Ajb+DDywqW4WF202tZ6crKw1Avy+EYHOySBJCJ
GU3sGOTDke9pJTLlGl5A78SbwYk26FweJGmVHmBklimmQgQpitWMiaTkGMtgnRAfBjOpUsn80DwK
VrEz/VQb4kIah3EU6oy3JqtsqG5attTFfqdQi8tmqWnGqHBMeWYhMmKYdK3ppaVi1rzMin31w9g1
STBVXp2nPrlA1/PW3sw9h7mVxx9XLybRA+VfDlVjFhfzPFxsjfwHI2W42xTUNpz638bOOn0qJZHR
mwBbTgE3JFoFspBWIroV8N871tPoJpuHqCaSkMbWJ/lmzUf30NZd5zSJfFmy8RUILYsx1Ob066Ce
Nw6n+3EJT5t1KMwwXLnyFnttb89ii3gf3nwQsDVIz1LpRDJMDgGfl2EGqUCUvtIcsaro114I/TrU
+PXtU2Iz17uvv7GImLI2oDfhtr97vqwl75eI5EHJbxkeH/ljoUFjyWIj6BKJO76wAOwWJgTR6qjj
qakCEdSU8a0GT5fhiIn7Tk3enqXOJ5TMcqtzwJ6EODCvwy0Ahz5RtnKDeI1nRKmzQOX8cINeZtpg
vhAXSn5q9FtFWfXYpOnhqCT2h1VUINsxQKlM7kB2Jz9hsclii65D2dY4BZ1dl4puOt+SSz2WsJxQ
pQO4I6OI7csJ9PadtA5TocUWjWb9bIOy71IgP0p2NtMikNqytgZsFjXiUy/OPUl6xQifFOZ1sGO4
kd1Lx9hF6NXwhXI21VpmruuD8tHKm0pa2IFsUZapPIh2sXHnnGn05NCPHDL9dXgdDUrekOnZ+9yu
uQFl7pN6FH+1jIt+tqv+BfxQ+84cleYg2kVvcjfc5TIkAjjEIXuS4N5E/stLEghtyP2uNxizeQ4j
Z9I97+08YeteNaKGinYDmimlw6OBe+sXNOAS26g1eMB+fbr4ItqsgLvudfU+BrjfDCBcdM6mtMKc
dShnKoVqvnRpcvQOsU5+YkM8O/na6KLRx8VNWQBFb5ObEM251m8eFM44Q4AXeWuCdNdsmnlNPBkx
5ELMtw8fgWqy7GyLInenchFwi6b704D3n4KIASQ+RJxwVAoAvN0681cyV18QFlQMMtf7xZtqTaPb
yXjs2Vy804LsYMa5WM7IjlYRn7WmmF879YrGK5pRqzaoJpb/hSFMhOkLHIvgb7JTe0HWrFLfHruR
I3pJ0iOgIvpni4cXYpt5bzk8o1iysydi1qM0kytlRRpKAE/hoLsjTMm5aYf/SM7tsiw2Ji6H7KnD
FdjLohhlUk2n7J4oUy/BO0B2hzt2ImmrWywGkBOBaehLXp5QMSKx5Oao9W3J6XB/uS/bGhfjMqDo
bWykxtSWVH71gzdQOyrlgKlDl8CPUzq9Nryjeg2xnW0IDlqk6hRKM5/z5qcTEiSTSZh5DiCt7urJ
N4/pvO5lPQ1UK/+b0X1XiBGClS3CikswfPeHIY+vBB5RllT4DjIT7JF4FoDcNrOi0vnyhiqhRPNA
U1lIDQan8++y/45WysgSgPAyC8+PfD1rJ2WG/859DNALBUgXM5j9IJFrDtI5WJFLb9VGxxfOCP0g
gUu+bYREurgkvDwpuygrYNz7Msf3TifMwBlyFnm4oqYhBKbTBcSviTScHD16fPzVBgGFDeCXk5aP
355Nv0AxhvqygjnWgPpNH3TyPBfpuHZCUkV2Aj1/DQZ9CCbUYLcBgB0APVwmDL2gd6RSQSBG5LeD
kZ2O9RvFmOLDY4wpr+s8tl4H3ejQZ5qKr/FSPD3JUrRIQ1KjokBNy+MZhWVg/mXspl4OyLSfWDxD
X5/UlfH4xmZsXZiZ7A73Dohu4ZraAnzLSDu3y7twoNgNsBqJcFAP2TUTWzk+VfTS/IE5BUMGLGFy
/rypcc/g8BC5X6Sg+I5fC135OU0sVvzBNjKxk7un+fXD9RzVnHeMVUTx1wyelueMv7Z6UM6+gawJ
0BNt6Ptqaerxh18CSF57ov4dkUWcE1dn8aQEItUuS9yjGOOak8zbf434VrjcIllWkYzJLzkQaax+
sEm2hr9R++O6tT8Jy7BMmLNuenr65lxlWyj5OwJDehf/FAC6CXCUG99yq2zfNi149JC05xemVyyf
GK5m8RqDKUQbYYFzs7/eHm9+x7LCqsuE/WwWTX/aHAWkUkLHBFXQhoKpeZIIctsNfGVZBCXdsyOJ
6l7XNgpFJQNchWchpJgGSXzz5ajGPNVy2zghEj++R0hthC8HiI6XNkTb6JJqu7uaLR87yrct66b6
dai8M7ZSfsaDaQ68BwSyp20Bfk1CgZCd8bQtBcfPNtb78g7Ye2WQRWEC2Fhxh3fgTvVXc37w/CcI
dbK1BtXdrbSl2L2DksgZm4MKpmbUPfLyFYaEUO4BSv3S/U7maDrOJEZ20nVaL9LCwp63XJt9VAQM
Eb7ISlcK5yhbAqVS5GQ/COFXlDx3aPyZTZ+z0+Gd0VxtegZBA71zKy2u8LPyzRtw4dh+aflAz0gp
ygx8Hwl/DrZXS3HVMkfs7eWO58xso/QNPDbxUomTd9AYWwK166JzO5dBStKuIIJyeAPvBJUHE3Hf
0CC9jeMZET4x9yaFKUfSpLrDv8gP35g0W8r88vV9FWr2nxXuhuCBRiXMQVvu9i+UJviKvW1juxD4
Jtf/vU1btQVkD1exSgdj94PjjMGW29nEYUYa+0SZgWXBhNZxMl9ba/T4KqaduqtWFZb073pWCK6J
SnXeNRoZNon6HuOLZDmjnlpvVrC0LqVaT+6Be3S20wykzNAilK8u2Ti4z9e+5idPYKhf7Xj1rcEN
u5l351yiTT8lPiPH1HxFBhr7a1h7opBlZbYCUP/pZyFQEzLEdqVa2vDhZ9n9R7yUe1XL032v2XRj
QjO0RGninrUjPfGaI6HXagvzcHd1WP4bwdp58GWH1XMivAZyJ4vI0N6v0cvmqIe76RFryCWVksLG
71bGFMymurEiWQa5Bh0wrhMpdp0KsNHSKJ/H6vn3jTqhthR1Urf0yMSMmJbt8UtbE1P+tbYqBrQ1
5NCiHjEzq5YFFMY8saFjCUpshLhEyX22A41M++HEWoN4HapYHqmqUm973yw285ecr3HepFWm+07T
KfPY5jrQ1ABxxUCV8Tdyp6vJQ9LCKnnEHcXpTgtZVhU47xnCmmQNKA5CjlmfvK5HiUtxRMEytXRn
xAsNVCrUQf51nUl7exBN9npCKBsHTtRHKQOFBDBD5fpI8XuVWJHppHzP+TvjVXPBrWTWz21qAq58
QPEcyihgS1xjHfiCCsD6ff4k+2gynJWp+lWsvkj0hzivvVzrpzvuShw9ko6Vt3wjk4nsvvS7KUkB
mtNyWkekRaMoJyUICiUbvu2YSH+p7rC61AzDNx+zosoL7jFngQRPFcBHt/g1UELU6CdG1BMahelV
Cpr+xR533l2Eyu+xKD9W0/s6fMrmuu3wgYmrnS656TOaQvACy75hkfTOlgh5MjRWOMnbt4+HI64n
ZwyDHc1TQh+vS1/raOcUUhVzxuLwnpZSAMndFnnil9HuQln8IpzuTimxKtdm8xVm8kZrLRFtxOV0
iTq1XwGXaM9kIkWqmkP+93EpOPZ7lr5GtkN9z97mB0QbsGT9dwd2C/hr3UPGdhYS5E8pWN4yFRDQ
UkaRMUMfh0p7EkSON2zHYAgPeYoOaEZH6NUA6imLkxzvq4RPIDVc3vOCDDNI/vzbDUXxcZdN8R8k
W4mzUZi3gJ4dnRaLznt4TD+Kh/99OecmufbY3VsCvIFWVMJ5uYD5wOCg2dcxbpmowFu3fSnFYZsr
smQjlnElmPdLB/RRAgHXREv2mJmBKRNqI93MM8ahRBWy/mUg1V2fblLfLFh+UgPs+IKSP7XCeXo9
SD0JMIEcJ6f6Adrgw5SBQlzAKlslMbQaNPzQuE0SstmGIulZj1Tu6XDLL8ScEg0vZJI8F897lUu3
RhdNbeXX4SNbvcLymBSeA9QkQAZ5IcG84RvILr+lCOmQVUwS6aB9N7Rf95hE89GxCmmSrJOLwwf3
IFApExcp9kR8juj0e8F7jRe24nkdpRKQmi+7Mz/nvo5bFWYpbAL+vys4XJ+B+IXIvs0CxSpOlMnf
qIThiWL6pVi7MbkL2Ubwva1n09oRr3WqkMuCwJrCfyqbZgTzd+dvcOd3nEyqd0OyWmtpSKwhHN5e
wV6HxExeEqqE8YhkUsTL/QITtYrpz2xUBW7ExHgkynnBHLJcXf3a9SXCskyLal3ygU79qcoG2qTT
VC/V+Zu+SRyFX99wYLR/x3kLV+RfxztXYrkHuGA/cnItBWs1aqpEwGtPt4KUZ4YSfeHY4SKI2E+m
ABv6JSps2THFEIHsw1I0l+7lCTVQlcZ3RN5U1dA8PsS94T9RuanvupL1iuH1rMcrCGXnh9oK6YTT
phUMCb9zn5SJ51m7vgwHzrRbzCl2S8yhbp9mwx8JVjPliTGoKAL08id/W4SUBBLZTKJmhzGkEXyB
rPS4O/9Rf8h3Rn/Aa6tWDwqF8GDtYHmuBctsMzSylaaR4Cn8sLv/A/TcHnEiJhSZmaJuvyDcs0TZ
36MVL5RGomHcLN1l3QgcrDR7s84MPt1MKAedgvWr8kbIX6ERGhfSY3rgWAcnAcsoX5jQ6TTMJP0T
RnZ7t0WsVzsttAuJ2oXyIzKvkiXjX8t6H12+pl5uj9SWrqTnkB+a3+ljZOJHDk47zM4Q7Wk/VS6/
dmK6U27uO2GqEtjDDzoSEzU/YtLA9eHZe26FrISI5TkGbfCJfM62ucO8ezClxahzp5uiOebRQMvY
R4sO9mf274DFvUxSwKZ34/srTpKi8FQCYLlKuF129xj5PGMNqoD1uomM82NTJ8KVLqpTrClj0FpY
dRECSBFesGOnQR5Cwv6S+lx5EWrB0XJtUci6xG+/xegnvqk/WsjJcHCY+Xy9yLYR/ZPmND0f/wqg
UU/u0QgLFHl3oZEpt1y2R4q9kKOpUJcghoQGQuTCqxQvlqd0w3kPKzipTGZAjkJL5Gi0N0/njYYU
2QCrXMvfn4pQyLovgHZyEZo+kl4FScNmQbIqoolDB1JHjQBEuAG3kBL5J7gsUC2Mx0svBSqWqRU3
RD+O0833BaimJ2LPudSFDyfK5xel44bhvY/+gnZm1/zznl7bAWggye1t6D8N2ZC37j3zh257d4ve
mcFP0aUg8LOvAtQWe1NwKHd4leGTxFRwCLQ4pOBx23JdhIUJqiu00qr522VSRf6KIZPnwGxvhII1
kNcXqd8Dfb5qwIaWRTcAm15WbXRI0bNoAZgeQrMIQOycqJD8Fz57qU0/CrJReoV8Jf4B7SiFbhIt
yvNDfl6huOhKoeieJXcCljn3ckdtaZFMcfDcoXCe1dT9vrZw8bpL6IRnM5tsOOPr9ERmCoOg7TsK
XFhWEmpl/woLnLRjhtRRy22kquDt16viCF6cY+5znF0Spg8dD06fonykJo3/6L+HwEZqRSnda/3N
sI/nolhN4HWWCzkr0Ux2+ZRaUz7zrZgP9A/BHsEUvtnR75Ym7PXwD/7b+cccHD920mfLR78RKATF
M/r0sLkhN7zQy6EpAqHQhS8xECwuUEZNB7mLt/TAxmDK7sR2VEZYEcS+S/3MR1MCrQXJEyyzW0LE
iPbGVx4aorEnHCLx8z1owygDjhOzt7cy84yDxVbYKchqKOw0+1ByiGIhaofuZ80TS+7vacT6JoOK
NqMAYsQtBf2tsAQR8l/35OsvyoMFWbPR43gogfP+8HSaSGHEDhxJf0+3VbG7PRzw5RMK/muO9dsK
TdW1B0YQHBJtA9cZQwwcgMY5eZeSdT3Y4YtVi1h1oss8PwP4CVEBq08f+MaVv6kjlvxkEGdL0Xbz
czTgVupL52VjfJeXcZoUmbLMlHsG1FnODyVoO5qo0VI2jw+55q6aLGuZsIAn7GeSIQnzqKrOYLkV
4y/jbS4oOt7R3kRBpN1dray0KneP+2Bzz+s3LkGmDUv+ZigI5rVXh1l/ZvtZNt4bDWNQuQWZiwO4
n9iE1rHxR8uIT2J5CZ8omvQ6J6DcNOTibdi95UNaeyZbH4dYiQn4hOOMRc8pvYUoyoHTAkp6T2jV
gyEyaT8g1j62JvmHijpd0X+rwiUJyzkY5NcjAq4B3yqttYvj9Do4oAkIODaRTOPKrAOwl8dHGtH0
uu/CpokWLJq4Jtk2QNgPflxAwuhiK0y7v0W4A/JXsJBPh8Go+lYDieddm57ACdUUfZmYBKZ+yao5
hBpA/ZZnqW62Nleab+ABXh0fBmo/gv19FisULFiruU5JBFvd/Kh7rYcJxvpKSLI2+ARKgAeB2zam
XzuiiVjuQEi+x7ZOijv1LtqkdhyM6wh9tGv75J7KhaEiuhOa33urA3yTWxfYiJwljyPITEK0NCLY
sBirAbMbtrwECxuseETf+XTW1+ysVz+uL7iXPR5M3olx5IdBer7AOJWg1qN9YdUNbjTHKT4WlZnj
ZSHIwWYBCEem8kVoIGuPNc/srPIH7l753MerhAldYRhvtIxScaMwObZcMkKT5Mt/tKCiGmjCxY7Z
MFo0MLN3GwInRLp/WjuA6h0L3urmD7CpQBpBMXLctze/oVq7ZZ7B9KyKeaCN1uipcXt/Uiy9Kkjd
IKp0lSGT7jykEueGCrJBhvLaEDX6AXzjheN+o0UE8AQCz+lU4xc5wQXRIUtv73sMEjoYKAtLAG/c
4fhLaQYrmgeOZBCTDiN3tDlkIJfLyZPgy/pHbHeB/O8QVdoU0qVIyP01Rub+AJ5oB1IFUKoyv4tS
W+cL1UmXC6QT/IINmQ2vLapgkvgaf8l+Cx6x6bmrB51ik+xzR5jJVa7GdzLxq6H752BN7gRa7SdU
JKTddC1p/H0gHdhZECOvfHCLIuvRg3DfftUco5a50dRCkDjI32l3yTfXeQBpDqjpqfn7J7abvQw4
qaF5M7TrZjx3+HTXc0p8sNc64JYCW08HDKxjaZ7nxqkqPrfnhNyVoWFjzpXVfC/DEew0vra63uwF
DJFYW/da0v5Xim3aX9pZwmWTdC21psMsdC/R5ujeu+4uPjhapqpSGzeng2lRvPTAQcaGmlrQhu73
5ptRtJnvU/FG10uVGGAYzfwzEIbw3RkSPUp3k6DAuOy8+/j/0aAWtLufg367LfQ89Vn/DqKjlKJZ
HGKujOyl8269zgeB8iiXHGzqe/AeoQlGFl4bwfkojyuTFw6LD+gicm1WJ+F4EW4Frk5nBKQn36b7
dqoVoSaJkN4ldgBT+IyyA4UiEU8j6soGT0rsY58CSksCSrAbOaNbnojWWRAjDZDKilkwqoSQvFwQ
ixEhdbiEiXvCF8Mw0TIIjsqwkEX4yukUIAV1FPMgxNbuZfOthOI5IggWMMGcVGp6BkxhWmf6NLDJ
4+754nyuIGWsTfMw3/9Hy4+Pd9HsIuTegNNxo+mVO2ra0LYDmdbOQzkamXq6o/C5wq6Y2/VGWMmn
IFD/UcalT2X5Fhn/FU5q1fNv3ECMmTD8XafUVBpKyLDLY7e/pDtgWK0in3BdP2eFdkuZCTjAtv4H
765QGuy+z8HzjIiFr7/A16l9AZAScRwRlvbKXoDV4BFzzqm6Aui6friNFjeyR0zVGB5UrEnbg4ts
lS5g9aYEXzPb6r9pOSFoZtxwpBE9HX6GJED6BRmjCnF2pndkn2qs9lr0vD4tcqKlBSDmY7QtHCob
9n6zzMz9dexUWQH75KtO6V7ToZTOSYXE4VqlF7MgRpG/wjUVGWWVHk9ubVJ8XT8CZMb2+A1ZNMry
mqJA27UviGAAvJo0Myk6TYJBX2Tu/v5+S44fFQw8bMwPRbCTW50gnM/2WbWhbRTrTHHHubmeIXqH
SCM9CKInlxUgCEU0xaK+MwS4HOr7XajkNnh14BUk8q1bTESYoCygmWhKuGw1KYiEmHnU0yH7lnmf
+bL3VOlY0tyq61js1tFx1blc0PAwI9lZOJABh3c8rIYtoE9kJMY9KZKqYZJbwSxq276ov3n/Veyl
hJU5N1vTTntMKLJp4/xSHo1/R0b+qZWZgaFHgd+341OxwcJ5wVP3TyL2WL76s1pkxjtQlu6lAxLI
hbuSSgzibuOcTmDoiEp1WrwjROByspXH3cdYfMoCVPKuYiATPShvPhouqXfIjBXwlyOoG1CCQO8y
PstSEqkwhMxokDijlz8gEFF1je3ibs+bjShhmiW8+FHjmVVEgumLhJL/UBWqfoeXwwYyv7/Wt/s9
b8xEEIR+j4gLJPUXROj6pfuBi21bYImmfrafG9os+VP7YOubOs2K6npYn6c5IJuW/Ax+M5us2GGB
KBo1WcSi27VR7LG0tC8ameWmtDkCMUaHKwOZ4nzLFXtmGAwXUsOth984f1OiJy0h2Qp8shhK2tpb
Qp5Q+W2327Wbf0tAHq9A7G2Ml/ocmSssGhmW0/4LEuDrBOt1qphryaOaJygIFtnuTaR9cGwjnFVr
uZPcy3V08SIVa6f/vvRoBZUCp6JmHwGzdMBw2LDt39q8Pze79eK6ClfYT/3O9on4IUHLi+b/zBX+
A5rbyGKDxg1QZKRew4LmNn9BgRu4e0WilIjsZfoL1UU6FSc2gaf7FyxYnBUAiT9sTF/lgap7X+wu
770TNvY5gWXmzHTqxSmMVoXqHE96WRgaXhak+TdvWWzbzCWuOdlL0wKwDpvHA/oxYctHOkrHAOb6
883w57bz6k0QW2u7izcCkRLgtCP51TujDfR5JCrZBGEXYgpeCFaHbkD3bulR08xcNCYKYpLvGfmS
hIlSSdmHCrOXjV+ylcbjsA21igvi6Ks0dGt1WZQpgXS8VF7KA0XIuu0nWDlsDzXLMgThFOSI1ETv
MNP6wXA4loRvT84lbujnWrt5A6+rfnS3n2I0jf3/Ruc+OtPSrJ/TZUue3rl+25J6PQzYT6q8Hc9a
ncdTR7XvenzFRP1LuK4u2Pd7J9cJ9ZoRgYRlFLOc81M3aspo6f4xJBo9Q6q/q2L3hWa/c1FRvpsN
HTpzF67n1+LwQ4SAuFgOk5ujq12zXZt/Q5Bycn9lZheHf+DX4hxVF+ywsRcKPDfESFkIutlzCRz3
9s211Tyzd3L6oQOxr5IdI3OJWrBXL3ACTRao3jWIFM0tvCsPCd6I98BgvCeV59P7tz7RLWtyar38
kcc3VW6MPRfrzlidhgsDPQ2eSOaMyYfcuyDDhYTIgJugDIgEZikS8trxfZe+yicJ4y7XRTZrkFXo
1vlWjXY/oTTEK4Ntz64llJfw7DK75QZYqiRTfDG75sioGlw+nkpPOX+RkLF5SiytNKtqE4Li8USl
GDmJ+JxZAZCn5r6Qt1K3OerAs8rOyGU+ghFGzr/ZCRWgoMZnHuTMph5GD1qHEO70lDKRyaRyzWs9
fb2QyzgO0ElwKGRz8Bu+Q0mq5VIBlhHmpFApDycfz/KdQMYx6ZKuEnhiED2SSQ2feabeFdITWAlq
8tz9+uK47XIAZvRJwc3cUYUsrjuk/GtFVq8sguc9wdpF/Umr5wzxd4Ga7BHUNmFFBZJmkAnh0kxp
uG3/OpcNQ6pjH5t5zWwf+U4HpqI5wiDnrXiHgb1uYIMzK4tLDFG5p5rakUNBPGL7teQ6VCBrGqpa
mCZWiZ/DFlDJm2kmM8sMRENJ8OaqSsNJn7rJmBlWZggC267R7hHRsdZXbHLjbjQ9S46QLIjS5Q7M
VoHo+KlJ6WTrhcqSsL+C2V7FHsbq31U7jXX1VC8EXQkR5PwuPTNfOXdDgmAnvIESKky+S7d7S+1x
0OUt4MXN+8W8RURhF0OOoHRRolUi26xfHjdYsIKT34dSwlkSNcfc15q3RFKOQoC1usfDOAcU9TpE
RWl86CCJGbKhrqsQyLE5GxbbkRnF5cJGoTFuGIH99f/QC+Z8cdqjR2k1PKcGpoIejSOdCc2KBYep
w/bqYKR8JL+/cwTkZBzs4fKR9dSeU/YksVWHj4urulxhwwQsJsglRfhEZR89bypw4Gt8VZ64McPm
HKAkK+z8Uy41pyt7cfZcIpnVhlJ/KqZQc5ONCXegXrGTv/4d44vr8TISFhEYfO27/yplnGWc0OY1
USLR0b9GjccSJwMVk0XBWDFFjN/j1aD/vDrsHGGNjJOsMhG9g6Li5HmcF+/1CVsoTVWcZpwZVKai
PHzKGCCJ7mGfvALnnJhpxcFuHuBWHJQpkjdQWyZ0OGt85Q4C8RKeVEuX5DKIRzuhwjuRPUD9G6/F
w1XJVtjzShJMFqR4mq6h4O7P2PcwK6Z40nzrVwmybprUGEzox14TdWocSu/CnZY9lb4ahSRlnZep
7h+EX1UGz1x+CQy3Ans69fQWzK1fOk6AhNlmyHzZ8q6CeOQZ0moAeC8sNWJBNeYzZDCcmf24397A
M+e/cgZYIbhQvZKVFTtGLhob/07ujA3fEzLen/GEGzP8tHhjmk9pnx5C34oJ6XldEdZbx1EZBR/a
+luppG+vHS9F72eCmiLiMTroASz/SxBnjB/ytGmALOHQ0AZ7kVTWaCm1+Qo6a2Pf1KYm2hysDX1N
3/gmFW9FVvCB0EWm/YvM/TexzKnWng5uI/PXFI/Kl8Ga5yDynqAe6mdqgklOcPEFm0zhXdRoPKoy
DW2LI1diAaLm3hbgVGQ7D8RThyzPUhYVxLsGn27heMzjY+MZXRZaHIOqMie6VB8neTcEJSxRnGJ+
uq/Y+xIfRnF6RuupQ3R190XlWcoqEckUEbnpQ5P2IPWA6FpYvSTkpaB268LNuhUmm6dvqJr7LjPu
HUWiBoN15EHltX5zehK2Zn5Bkrgfd+ZD+ylXv+sWjqn9kl1qF6bV24Bf+NXn7oc6n132gXIdcm/V
P6EOV8qYYBA+zHPyyYJe0L380+vj3luyNEswrnLbO8p6YNQdfvnNJeHH+Rv4U3ViV+zozcgU6DxX
gb+lmH3kVe6pw81fJNhQnl9qUtl6LMpVa9JnWvyqlKEa4yPyT16czN0fWvXHo64CdHx59zBr7r6k
FF+0N/LX+WKAa8DPpaLY/dwFkH1CM9KTwZbV0BZaFKv2VFY6eL3f5Es0MJ+NHrfqCIbvYZ/KINQV
o1SSEJALz6ywYahx4Nt/9/9XP2m1UqCkOxV1SBSrfT+FH/zjvPGHXCPeR7rJprdA+r3MP+ovf0J2
A9mDzBqIbMkSDVjRrWAOwrJw4GYRnLHLwN6y+rT32mxfEEjSkSTe+brWCIQiKiZ7Z97xl+zYEYbe
ztUkBnnVcPQUIM2Qts3uUsGS/EsE2UJiyo5EbsABG7kdCtqVRYmvy75KPUgW2P0ga1JGMF2ABb7U
mlwezJfhR/L2aREu8NnekZG0f/0FYq/ZUhZgzpdUDegMD6pW/Oi4zyZxmN3NoDFbR8eUVTWNYWQj
DHCz7U2IIYSFabi9fiEmEF/PVjwFFUsYa/UbJtIIyFmrMT12znEYNZ2ez4ToHXgnt0oq3xZKjONV
BZGKCKkqMFl0gi36lJUIujzPKCGFvR9RFTt+TqXX2PTSek1C7Wt/4Xhn40T018BPUof8qOtnbfdR
j8wErSHIbYQuXZjJbXaUDdNpl8lIRmSzt8RGwFFdBuClvLT6zrJi7l2nbe2cO9OocJumGHp6iku8
04bYDc+M3Z3yKGPqebZawH97PsB6dk8BH9/W27uqzP7kSB5xq3aa639yVEv0b7Ux9W128h8ItoUZ
tRKBEJeJUXweuHUQG9byf/VljyBQpORFWIwoaO+W+Ny4MlxePZ+nniABmHYoIa7RmDyRKlOyeJfr
UeJBpdPH83qIK9BGm+RN1D8maz1apGh/iELVFsvcApod0cfl315JJ37882vW5pR4eOp5UTr3NuLp
7exCE9U4jJm8KdJxCgejpcoBWanoEZvKNlBTDUd2nwxU9BtbqOtmaEmgNAxaY42U0JD9V27QB5IL
P722ou9zQpvxCMXX5NV1fJGEI2s/vOlhQrF8eWGm9bRXZ8RsNuc1LEWRlGhBRc0RorOzbHe8cx80
aZdXHRmc9MkNzJr1D8lf0vb31VSCOmw7+LuIT7iGvhmyLwN91DW2Iw3R4YURTnDUtk1KBxpKpEYQ
Xa1m078ymXFy3Hh4r/cvxt4nuoJ8Oj0QLBLHVPDQ778jes6cSbzaRYUQhkBat0YUJRHX6dd6Um7D
hOxYrE6CI4Hg6+4Fc8EWoHzBwnH3+nZU7FqD4iJM+Q1lsxbGk7Q/cL5ydJe3BWnuSc2XLr8a5Ufl
+4Hkka9uEs8SimOw7gIxjAwvnCfOqB7OxXyAvSa9t51GAnieC2MOBIyxwHyoNtF60Y9BOhFCFFF4
KIBTBgyJXUJbIJS9NpmcD/DKBL5sV0CjndiLO1fabhEcSyJMfQFQaObWjlUZwOQwr7GwF2E2zQt2
zaMqKfcyDQp0HXpz+NO3VW9HtbNU8WldosTXRBKfcOOzPCdVdCbBEEAfEZmiprzzS59ei5fTX8ts
hfSKOtiAKMDdR+XSroI0hpC+9d1F30UazhJOVDy7Lnd66SBNin4IvGW5HbXOgMVLBDX8qLUiK4Qe
KfjkBcTgp+m8+S9BXVrWPBcnJ3HjpS+syIovNR2ieGr6wu/bbzTnosVQH3FnQfLundQpHsI7q3HW
kOWWcpr4I2sPODqpLzhT2LR5F3Qy3gq/ZuCcmeA6ay/Qm4tZPYL6Q2p1Dfeptk8hSiPqFrFtc997
Ka1k2lDPzGso74ke07lM5NnJlcb+cfGiG94ldEWSn5dacNeC+8R477MjOlDIbFz4pFRLr+kwPFvA
c72pJj/tq1lAUHEbDPxMIV1bmiqvRg1Io3x+3oifDSFOKcUmFGrKnpxGLZKrm924It1dvPYDpW5b
uOrLRG+c6vx7JTBJXwopDD35B175UUpwYNskvlpwBUy/CWRusBgBjy8VsscO8M2SJECJHq2XbESO
K8HSVfJD+FNlPRikO/LsEb4Sz2/EfI16xFPEwgYWuxeiRT9xIX1YTp2biUyJtF1UNQs5r/A/bY8s
jQRft0YGFBpoBWk4jgHvb7BX+LyqMgH1wlqD8lTTt3qgRYUf2D2hOgALI4YLo5Ebz1k9Ku/+cNkj
iKkkTllX+hUhmJ7jKY2jnVaeqrqBbpOvQ2HWeLRBNSjXWiBNj8+kw0Gz9zo4bncyXV1faAuiCcr7
efFlk2erNyI/xVn6E/2oAO+e2Bt2ig+D6v/q9kDkCoI4nu6LwXKAk+xUl8FbfqJOWbBuBemtS+15
A1hQhLRqJ5e7v7ROkg+iXSpS1obp74YAHTXUNctSvzQGNpO+03sJjYZ3mzH9qOl5G1fELEsJR+oq
wIlJFP5WIqY91lgsc/4xUbNUaYSOHHp4tJYposZwQu8He612YLso9cM5Y7eBJFZC0Up4SltGnPf9
+AIzAS1QoAxxVt4Wxvy2+vDX13wbIUySactlBhEKOXUx42O1YIfoxgFTPiGtKrcOsMf3vv4wOuwC
97hlzlUO3Wl/2T2N74bRczRKRCnRwfB8qsqb32AI90bYXbwCkBWkRlffuickjiDP/mmwtLXKuGUe
oMKcRa1KXimSS82jc2803muFE6iMlxk2179/e5QdNF8UjKHnvQqYQ92WZdhYzDmVpAsNQTRhBkAl
pihl46Z/WW9zos5Hb5rP9JB9R50R6xdYBjSXyoqlPXSIypM496qqOGnk/jaF/Igw25lNLGm6FW3C
Xuz0Zf9GpBUhdPXYM+fLjHrQM090gd4GlRddFAl8VrFLbTMvDpWizZmtbHqO1JjUCWqDTR4/vI01
V38ZvwTrgbm+c+B6f67gYXI35rf5iaBZkDlWnJ5CYWuLdiqdIOcem5YHXcscdxYRURVTHfFN7xFF
E+au24FsZtnUWCa8psRRoFA9qSylqF3IlcFnLV562vsP3ye6hVHaKBKEJtNmG4RBBnrnpLMMV27r
8AHe1XigABDfG1xwRHUtBDYimxsmOFrYV6vWqMoWH+XH1mw2HppUUQYAQWYkNxJv0nb3/OjDfRTN
nzL/EZsNeYU1xC09wF0tm9GARMwyStNxdnBHL18qfsATIX6km+1rpaTaovEAXXjCJRgnbOWSV0VV
F1F8SZDgS0ETv+68zYrC5Shy0ZRKjcnPSKlozUF0bb5fbBpkp8Xw90BKMg0TTdzW9AkJcsw20O1K
/zuV8MH1fpJAepy45+Z9mwacZHM6oEiVWy+8EgxeasDpcmbhJnREcABXDY5QK4w5Vw144GeJjhTk
swxOZRj52De2zKZz+4oPow491omEMz3ITTm8Ac0HjDljQr/qSQZ30Ekpg85S200zWzqI6eNiUz9q
au3uQY0cV6gGSMcn/Tktb2sP7RekhT3tVTOPD4rTtLgFDMCMwUdCgW0WSqqKMeQImOeMKOtEzGF8
1PWIXJ4k8xx7C4k0hDHy/Ggcjvx6xKigmPm8uSVoL/pJp41t5rny2movRqRkJvPMnRE8uoJhH411
xhReUV+EvXUHCFK9+EHiP7Ul78Sv64WFhdZaBcHs3o3cwTj7D1tgVieQHGeaP7A0ZTi4g/DfwJhW
1iweRaKC95wuELKcFPVn9tPbzXKTImLJOK1+PnhNr06osPN1nkFgxp8SwV7u+1p9aDA/yoGZby2F
y5kZ1H2tAXjFFFctnE52E/3DGuqDySnPZlocqep4NXymbmJvBJw0UWJzz3ITs+c9MGQHnu1L8ogO
XTzM1F4wj+N0F9mxKj0bvPcZg0DvWxk6xrP7EDl2Yq1L9GQN/obUgh9KwZOzH7CU2txhjRHeoxDB
gFNv0/co1eURirZ5ljW8De926PNKMDscTy4I6G+naee3KS5VskqgDF5rMH9QgxCjo9rVTbw9WcCg
5KQZ63jN53ge7BuAX1zSFXOJiJgyK7LrhVCoEbkzv2ljLaSbIkFfp7c1OwE0T3M5KvQUr9+Yirnz
eJmSvq/JrRULnDHmCJp6/XaehST+OQBtCwL5iA4zApjwUl7rhgHFbjb3DmBsaLrf/bl8jYzRGmVn
8fNiH1cwWFObWllIW9Yzu3F9uD6uEXYVN4ng/Gad2TtmUseQowiOq5F7zr27+0kRB7iQbOV6526R
l2eaKLp+vilW8M3IC+NQRpxBK2+vsxumoZZrlCrQ4+rhDq1HbgjlxSDHHr3EMYQETOrqQNYpzeAr
LZN7s6FObi7P2M7+k+yDr/4iqxg9sS49BrZxVecRqrmxmm3vypT6G9QD/LhyYrSoiLf4eu1oQ3W8
y9qPo4lLq4YG8yEcJMiG4rtUtUg6hv6AE26oi0Zopjp3DkV06wBzCvdOBv4EkCQE6Wey55QChqPT
lfHq8hPU8NFjXu8q5dQGNEBYe/FAM59LJt3ThyEOTrUSIVtOaF4jTJf2zOaNV2o8vihcmpYF29CN
pxWLV1xo41q7BDZ8ziCr7j197qI6cfsOllvqF3pcGlr91lLtsUG0ubzwGp1cGZwhP5UqGZrlXJCY
bHKqc1lIRiGTIZdwjMVRpIEeLkPnC4o3ah4xl5HFF+56Zj/ePCDqkoDPveVr/AmNS/kZgSQIQ8Tj
DAr6YM4tYnPBJ07fItEwslKJibzyCIMZZIfhpTXLdYm97EQ8BkXChfc+QNVNUGD4x0fLjlcP63P5
2COXGcNpO7Fd5Y7spY4MDeZEG0jQ59RclFrqTSLyYBf3Qn2eL4/VDkgxC4KTcjXN5fOrpBLUdMGg
AKD2TZl4q5lH9otbdvnRNc265U2S1gnD/5xpqDz87zcNx4rb45B4BvpZ8X3fJKGZNjkuomPT+qXp
Sn3ZOOr8Ax6OY7aDFQ+njHsr08GVfxKjDXpEh/i7iVggwumVY8e8rdyVdowBnwPcAZvxANuYuv1y
FRYHYqBkFsJmROvjPSP8Uodx4cvKymIZ0foE0nNYS8nUms9ry+TWP2jwWZ8JYpvitziLDwu7trNo
y7GxPlVKW+i632hIGtg8lXaNAagGSbUGCAhqhvACGB3tIgGF12MDTEDA0XyJ9vRiN3sM1QKAJeRT
554mfITzTZpug6+TLV7vwpgqa4NRDp40J0LXc3viGfivGP1xh2nVHnriNZD7IVrZ9yGJXOOly6be
fk4VD5QIYnwVC55kSzH2rsI9zesi+/G9qxA93q9SFV9rRHt+KYneNUvEe4GTvuoL7c/vv6Xj2rT6
mOVLYItp28ky//9pgQl7HRC633TDcFzr5TuwMZY3gFDomBL6FWhsKAYb9fdTu/2UdepQXi53LaW7
on5Ig/1bfj7Ex9NTztfCg+z0IW5YJTBY7NSdOmm2Y249mbelgrFqTvF/wQ6R5qtjYwymNu79zN7M
c45hvISvGklScdxhhhLNwjjlHXPV5KGYULyrHHBnJkKkpufOP/zHMu2LJgGPZYVeL0koOg8Fqb8b
xEC1rqpsLjRhJVJJUQLuqWs3wd0AvGVDgmTHwyjwAW4Qq79Ld5OPicuDS2dXnbtKgWpg5vTmlLNt
PfvB8f+rxrkS4uqMFyWwIjjFjHu3U61Q8N0V5RQuzP7uIv40YmrN3PQQZmTbLleyjiIEHsRC96PU
Xn414uvx3gQTuJcG+vNpdMGKZn8cARcf3JqUhIaNubNn1WHG56Ed+xWQoHwFs7a3Rd5XrnUDBUpZ
Z0yGuwdmxLTRr+qA1ZykYdctO4qV4/qD5klDGN+4mi+8a+bxkvpFaUcuouZpzz8EKDILZcHOg53z
YPEPUI0wQhlPYEj4Cgcmva7yyn3H4b/SitR1BWr40oYu4Zuh2eRHSwe4Qlu/13/ddoNELmOZx9Jk
/hnPhDocymLnJw8y0ud/skUfOixp52Csz5wnsMyqeXExua5abOW3TAZ6fc9bEqHLSa0ucXgIsZZ6
7i+YX6NdH20kq2RDq9CFOee/v4ftRYzRyvVQ/mMoGoLrbANWiXkVCRudFetNBM+yEArSIOZvI2F+
IxbqCUON88P4MdT5R43GfpkCZoIVDtfDnNHMqQnSAE4gbXKWWefceR8eHh7ze0S6sfSbUTjAk+Vm
DQK9Aj7WP1aMDYZCXh+AmZUHrzponfL2RdgJ6AWJIZQo3dSVFeHU37aQxIHQCbpZxwtFHWho2stf
Y+jxm6PFrRukc5O7ZCBX+jvyngkqIC46CJM0cNYbH0ZnptIJpE6y0N95+SGPOnBLEvLi7yEj776M
QsP2Cc8hFIEaQANq3vHA9ZAaiPpxf+UZNXxtexyQtnS1izAHv2AQhu55zIw5B+S7Q/F1dlY8XDgb
IhUlwTjfXZrFLz2uF7v0TOkQGkhvq8f+vznkjOGwKtQLR4ok8Z65ZCtO4RU2Opsln+omWWG/rVIU
BNCCS5T+/XVq95jFNscD6KN4chKouGvmjFSmXiFf8NDoHDVan9tXfMRKmA91cx/xxToPojgATyaB
oiUmXzSUiD556Mo6VPSS8ucViGLbt7REUCi7zIMENpLDHOVRYzAaHr+hWSjoZdFW+aNYzJTFvkNG
o94aalD6DRvoJ8fZtP/rB92kBPN7ufCFsiNJ8M+Y9P8uh0v04B4t82I3pImyPHkREwDufC9eAo3h
EnHpyL31LSwz6BGWbHq4b4c7W5q2RnsojL0DZhZDrbPY/QtYzzhkENnGDX7Rp6K9xhCCvmQBhN95
ZelPtjBB9/iBnLhiPqpGwwjNs2zzG1j458e2CLzIp/Wo2A8gkUbKQ0ZwGwzsSeAvBVMS+VNbLFtD
VoCVGjRHJJpDr8lLlWoiW8gWwGCBqn8TsxpiLgEU7OdeLSE31yoft7AXdhPYLxz0q0Zi7sfxvI9l
VzPTZklJWQ8KxLX8gUKCwkJTxoFqAhhPXrrnPM9NROQHnpYCLsBdSfu4mjzWDkfro6fshGudhLI3
xPeeHjDTxT8rp/LzhQm39ZF8LYMusFjq6gdgb/ncVm1zaEHJ2EVyc9TDx5agjcamRDUf7h4tl7F7
2LGE69hwhh2v2Nk7E4l+fiAkk+c4XaZKE6uQduruLkT60IyOGHKU+X91qUOsi/ULz8ARWbNd4HIs
TSNskUfiq8+RymWuUkd8EqO93fg5bviaWHpHIMACk6VMAa0p9QlcH8j4ucxvpy6XOXR3sH2woowx
bmPXmzB1JlJ6In70ANhsC1Br0RBsYvGY4/LO+rexYFruGEhlnn1TVJz6k3CingxrMK4j3To5fCI/
uvM6QJmCEi0BDy2eFpliioXaSYHLHwRMoShGhrsC3k4adtGr4Xdb0Tn6BvnDL846G+COIIqw5jFN
ZBoFPpKksDcHBDDHc9zYBBVuCv0ba7mL97vghUpY+hd5fqeXDEMWHdf+lZdzAZ2ik2mtif62HQpo
fYrIbWA+mdC8uZ2AzsBO7osoqWQVqicS2HzrVNlm62Xu7hAhmIOnsDY2FnIBSz7kVfAdse0Alw2A
6Iah92aBmRUZx7W7pfgjoEBVxNl/8q+kWZoOKt9HRRar8Kqi1cLHpGM4MRagpsGgyN0h/t7k6SYN
DkrFCyR8I34aHkUhobhEgHJIFaWLStvpYOb6v6sXkmbftPes0RA+7PiBvBMGL5M2b6sQv2aqLk54
UX/qImHZ0RsJQvrIHrvkdNONQN9x2lMEEQszCWvAG+MSZiyjnRwRuPZBnnNJDoyPyjoykf8US+Bc
H9aQQpEdNELGK144f6oEtwEYuJEcZUMwW4jziTahHopTYqVytmVSqALqKopCpgHSYk6NtPnk9blX
vQMor3Iw+KkXjfL9vRhT0pBRhjhz5pzz9RfUU1ZE0IzaKK393w7tSpzb0I2SdutwmxDbW++T5bWG
BO8v4lUwMyolJoS/eYHPe7RtOO/mZwlIMpBcaC5qZVBU55L8gcVKCjprx1EUwp3lBddglMQSPqVZ
Qw/8Fh438Zgfjg5vynPd4zJRaJ0FaIhbAgom8inwANID/ujpU16F2rR7bgOs4yu2wg7cZY8AVLka
pCCH9qMfEp/qEi3onaIJdKI3n7KwTq83qhJgmcCq/0bG2dAZggNV541NjA1Fqb6EfmQtM14QiJSZ
EPLhabEsQ+q+lXh53XpGFrxnlKz9AzjxHAsGBAtDv3Hb5JZU5JJuaXyv1ryH3SX//OTDexGVDxdq
zehU1T8+FYsRv4QN8vSai5sho+MtyT40Pxu5/fXgGGkAzgxiBO7PZDwv3w2m0AAE1RsNq4sFFnkD
OMEEheFnHojowIQ7pzI+ZE+DZNnRFXR5pjSawBOeZxTpoW33ES4JzLt+CEkSJOiOsFOSl/jCJxNv
0+PNfkRcNd8nF5EDtPLs3ZF2xfFaeCw8QQ66m0iUdicm+3YHwuIpNw9szCwjPc9ZuhZ4Yt2C60JF
cH+JXsjz7ZsK7dRrB5d9m6hsvxesnvdUyPQFXiA3E0P+Sw7bhI6W2FoyVm4hbKP7TRaqwoS9iaiB
LelAgfiWAC1HVwGHKm8K9bCh/NgIM/oXU3HE7GRtAdK9jy4Hcc5n0oHU+FAk/jay4hmKeu+2xgMh
CTr4MUwmJu2kmoFi9eqBuYZ6gaayvvBMy3HHd0GczSs/QxLbXdEwTKEWvM11fIAlBCSZvT/9rX/d
jFpS7EmMCHQ6UB1rlkrVQdCMyX16SeA1MUcAKFhlkCL09jzOtNUH06iNWMGAR7uVQdW5uQFxCLgX
5RjiKJLkBoyd4VeMEANL2tt78LnL/oMfxq4stmFOz5fof8OICK18hWCPPqZkCYIz+bnW5Vyy4mae
iWc5Vx9FITBY5w8LYwQPe8dlOiXMRpu2x5JxB0L1XeROjn2Q/DuKkPjC4irLRVAChqyl8Q9bVC9O
u72q5r4UKTnaTuhkiaDn0xROmqNvEVnDc4+gmDIAKre+3E62y08fkjVXGhr5GY15xSE2YzAXmQe9
lo3GsbrR+4ZXZPHT7Fc8Pg+B/QknUGyvDxt8Ekuy4k+hnOwOZxurncF1D+kCRqHsNJusf695ELZV
HWWYqPaqvFX2kTO+I2gfDvcuFroXznqJDe9iFvZ7ATNi0Wmh+S5DHtOoM4zuuQdrf2daoltEGK44
jepbrtUnUQJewPKfVxCZsKMmr1wPnvHuckt9c5pq9N+4Is8Bwhc0Yi/GTffz2LJNkS8+5bqCuu7n
VuC5+BcRpGJg0iDSH6keaEgzFXGvIkgP7X/J0WV5cRUFk1MG+jSA9XBUFjW48erlzE9wE4h/W2Yl
Vc0klBFpk6YAeugsK7eaDU6d43orpRK7O2Ug0gqeinOj2OLvYHBASjZnws680Y2F9KowWB5phg3f
3glAlazRxC7MLxhIBngub9pYIvJMAo+iPhxKCvX1wqWOh/Bdm1CaRfdE3W9TctgIGgSfX6eAvQ2z
9GKieYjdEUCHIOZZYwhHllWO2ytacFO6YF5VapFsBJFRvj6KOp7JhQD47kyAusuiHPdIbZJMRxyQ
YhFGMAkKKbQwLTSonitgu0GhXiQWDqm59Q3jn5t+gCgxPUOJi4qW88Bur7FEa/y03XVRByXXc0hc
4O6A2pgyWk47LNFpj6iQGi3nkYb38WnLG+BWzdMDqG156r4qUzfikSJITfzGJ1XEoi4jEFvT0CYF
dGzie5DVMSMzp3RNn8NAFlKCKiltfXf5XXH4prHkaV8aJt98Isu8RY1Fx7Uhy2IRYTqJj+kErfIO
2pCxGWKObQVVd5cSnChOclyHr9QqU8nSAc7wPDG6fsxazj/5aF4Is0pvlq1+x5IC9CqcVmMEoiCc
vVsiP6dssv/ONwyFxQKmN8+FHtZPd7ytxAkTghBCeONCfAljE+kUT2RA0J3m6994FnqvNylNPpt5
F9tnQY4ZZ9RoERvaupziFmDrF6zm6ebfercHkkdQpLJMWg6yCOgvPzGJguyuWDhv672LpDwgM6WB
34IZdHF39NXEu4fhDqMOI+i/6hnJnvpCW46M7N8/gfbhA6xzh0Bo8IonmtM6LyU/QCTmYer1Dz/k
U/X/qujDfZLNZFIUn2FRRe9RJZXHOfCcd8Zd0TjV50Jsuq/d8z97lFs7QM1i7XStrKa1fEatg624
vw8Z+xEsLLP/MXTLrl4jclNzYkf0k+d//uIlQOT13/EZVV45NGw3Y4y58rmD3xRt/mO5HwHy7jnT
EdtDYXiwj0BbW2IsUd2+SWv3ShNcjULe3q/ngv0V7ven5oWEj/WQLktWEVZ5BdZtw7m9za5ctntL
DgjxsFSTYetM0fe4GeOBQPKQO9Ky8SSN4NhR9FT3EaC++jJfHjySyNCsDrF6EDS5TY8rMRBiOYhX
t1C2MGuvNmqpB3nbYcIg5gSXCxNsODcvX+zhVnwkhphEpiFw2rNhqCbbWP+fWoZTiMyAXbZXoUIp
an+i6q4OmuxAEiHWxqLfbYvPyVbiKQW3XF4lTH/pRAZg5mCrbezoeLSmxk5PhEg4TK4gd8xo9Xum
bYhqe8+s/ZGEFRysotSI54LaU8F5qVQZjhedqCwH8wUbgMF3iYLZPEesF3O5shqw8aatj/GbvLcg
A5uarS/5n10kY6YZOUGyrvYimIniuftlN1cykyYQTSOa+rH2b8aIggqjgVD1llK6ULEAbANMVC/F
k4lhIFraLVdWk+gJdAOX8XvskJrRX5DIro1MPuH+mLUxsrZUfQfYPVPdEvEGtV4fPlvxZmKSNF0d
tf6FpxoV2td0qen/M2CFwjMbefQ47NzrJZ3PVJXD5C/TJkyL9k6xeKigPXqpEmw1W6JvoBvi+GYj
zcFHlqlfGrWdNz7pPDJZJjS9ZuIhfd55VUg4Q9wE6MczG7nsNjTsOiZA4G7hCXHy8wKI0efyBEs/
VkYbNCvsfjZ1ggnQjH+xpsUKOvv/MvqilKu8RG4fLI8z8ecmwJCOfRFG4VExXwsFGUMG+OliiBPB
vwhp7nOtpjLSRrUmMihoFsCh5joTR8dqmBpw3KhbdSf6+L9F/RG6EVS0YD8DELneXth+JC10hXsG
sNEbweu0v0AoBeBig23fWvj6DjeVuobIPXQ0rRQY80e4dueuA8NGUHzetFcAQLE6GebjKQMe0LeH
qy7Y9AJHeZ7JbbphQFKDzKlQUhyXtGkqFnMxG1NGOw5tkQDMIljtiag4/t847tpd8x7rIyMU68pt
8I3Nw+EemX2uhiSUH7pHpNH+JPOXLpWpfNEfzYJ0F2B4gmkIzBqOvZbaVkNChKViodIP+Gm+cBV4
AoTvK4PEKgp17MfIB83FfgPv9v6keOU1EZhE9ffmgYfiTgzkUzlLHl1Ufq2uSO8jqb+kxeLCQrwo
NVnCFCqYagmWfRl20wgtQKcghuVUBlYRSE6p8gjxeWgTd6VHYRZdpLF6FkD4wnC206tOydhgwJh4
YJ37sUQ2KjrFZj+lRf0ntR1iIxKLAN8jL0hxz9kFEgmLno4mvIArOOx7BvNhappL/tK+jFgwp767
0EpWpmKi9hZZ9+BjAFu/sRmiMHY/7nSqyllGspCMkiXdAP0WgRyZBqyBl3q4cW62iU7fPcm221TR
E4XdX/CSKu5D8By7aqUQ7C7e6nGOaIsMs5xcPYqdvKhX7I9l3UQFbbOar0yMHSy1bW+QRT3ZhvAE
OZVvFfnqX+Ns/Weap4DhCygkgsy6xibQEhPPjW9p7A8JMKKMjxSiVrJ9heyzoZK0gkIaKYbGbupV
dxI9aYNFOWenBTAzJMmugJ+N7/nHjwENQXLQrJLyYU96moc9e7sORsp9ytvrTAcKHRuu/mglhByN
yr0hA7zXjmvZ0VXGwlHgJj4P9+Ry7bRJkSaDbmG9B+sM0Nt8xVR4F3eqlMxKKyJYSxMAJdqUyy7C
rIUHe1hIoO5kK/+ZIrqujTnftktvLeuR8ZZzc8usHW8Eqhn9tSO70+5o+gUBlGlOARvP0lNn84rm
hBj6nlT5Oy1gvXbvBcp8K293JBLg6TA9zKPR/gGz8Czwfepi44W94XNyv4QTBojAt2FPcVeN7qI1
wkn9/qW+cgAP3oAQKFalXrh54H3DEwaI4ZlE1aDwcOU58kEWktE7sHyMx6xJzHPwewK5swmD7bX1
+MlFsgKI520dg0rNdUUbWbJ+2KX9PeDKpMZ0XwRMbVkCsgaRAolet9TbS8D9juMVg9DXiII3AL5o
HW4p/c/0CdUjvKfJnkHE6AA9lurxV9fOTlkwDUzeNGoNAOtTF4QsZTiRS/3I8iqKis82eqz39e67
VDoJw8jbnJFJ9irUuxN+cWVqDHucA9gcGo8kPPHD/dOKWCvpOGQ7lJvd0ol8gwr+gGXwengkNe52
q7ArulxpraHQlGLNQdB+lzMnXUUpb2kqOGMnf21C008TVLRC/TYDkHF9aKAANd2ukH8nJGFPw7Hp
dIsvA3gKd1SQOrfKAfVTWAkLAVD74HYW6DZHvh92dxaKWONlUvzL4FT9eX3Ty83EZJoY9lnZtc9W
3tKtRLvg10Sb3xOiNQS1OrCDdiZOT0UBKOPes1HNkIGAMpj6tdgpZfW66c6G4zPuKTLYrpO6zWGG
yRQ5LnQy+/BeTjcLPt/Mh/TffVNl15B2R89JjvsLH2QeAUH/z+4lWBkqDZ48+AawkLsoxDOzsZzo
g+r5NNqd1IJ8f0jmnW1kVwvWt3GyosQd68wsSRe9Ygw9Vu+H1Z0O/s08OenwIQ8S6t+Zde+3xiOV
7A3AZvTpffTTH/C3dYKhZU8mzVa4hALN3dog6tNj6yZASiEuMJOdeXt0gqyMpOjtANeff6A2V46v
RMsZ3UwaQFLiSSkk9f+mDmkA4jdtl1H6pUpiqjXJTYGigD1/OCUlEDf1edUbOdPS4mjJ7JJZKM2X
XMSXV/ZZ3fBbbhvQ/+dFX9yiOueEj7QIRzEcHcgXExnvCrIdrjLIn8ObpkmQH4BhF6rF1QdXWkyn
gwx4iQ+X/DhJkSNuiAKxPWcasxX8QLc5KMlUcw7uuco7D8NvoY3rEPnUmX53KdXbh7ygxIi2MMFu
t+EOe8n2Ti4owHaV01pd2sXFXun0bj4hjpUfawck71krsAekcNUr3O3VM9zsKqrus/lzpUsuIOqr
+mC6qg1SsPNvf8vgVMLbome5Ui5O775YfutIzX7sLKGJCnTmzYKatvf2PKfIDqBZLBjXUJ1c2Ey0
IqXMGYWnOpj9q+y6iYT21RegE0WBGVtTorMHyHnbn4rWprYW7WpIWNFzY6uLJVFbLUIjH8V1Sfbm
eW9lZ5z3gCq9AB3DLPU0mbxyOOX8V1nyW46T5ijSK5djiRyt3Pal0GBGlvMub9YzoRovDbalSvy7
I00auQOGh/efix8yhID40uCWpNk60x5CsHNog1a+WEsLZgd56i9QNQARyz6MI4NkeFeNjSAbk98M
apZP0aAEGA1VIcUQ5e95iLNAk8zNhMoF1i6XnDzmpOVNwH2LKwBZ9efxWjI8ps1khHe0psxSRrdH
K0WBljI6LDOQJqnl6POvqiVn+rjp/UrrZ5v7tGe/OA5ThTRTCM7CA1qh3fr5kg2zzh0n5taofQ4g
7xfqOOkgIbdnGxeiKT+5hjWxnLzbg1S//m0SQiQdpzTwTT8hUyuJTl7QlZKLB98zj58U2tuatKE/
4RTqIGt+PJdH1zZrNyQr5iMTDGyLOQMHZeDPSY8EU5qVVoPJCVJAtQYAXwv1DK6tKmheBXR6lTER
ip45X/Oho/0X1g26rhUDt3Zuv8wu6hAIV0xdaB3o2Fmwl/rYmxdirlC4kyQn6AJ1F2Yj6cbBk/eE
p7Kp5LsZHvs3IKzux/30va6A5WiKAYigUIleMmpL3QX86YHRfLlzObAR6IqF6AetClO88WtroKaF
N08ncisxA9hvNBpE1JOi1Y9iDT9slELLBoSrbThnnQL7/f85w7kpN8MSjjKJe8hOfhcOoKfP2rj/
u2PJomwk6TN+iDV29FrwxsZ9t94Z9YOZdXOpD6sU5i4PU2KedVa1cxJd+E9V1nl6Lzur/0Nz4GMg
t6B7o/4awCBgkS3WYhjKmpC3b8HqitKTRLjBzBYZ39lAl0tUhhhz7BaeeHbWimyHeW+Xt9+Zs5LB
geczYgr7Fcxe2dIQ8cQGAbPojX+OUR3mkA8lFpXJ7x3BAxU45IdhOoeHAd1qE7x9WK00hc1SmCL7
gAnuyUzuEogS/HWh7ReKfmv1mDRFWhjmYNkvsY3ex4IN1rctDZDic3oIi+As8QoU8YUEHK7dMwIa
KSLAoK3c3+/nvFX0qqQdR73UWg3t94D4HbuGzM0kCb6kyRcyU0jQf+4kCHD6C3BqTDwVDoazx68O
rVyia0r5xmtcKYtJJgB+t691YifWg2FT4kMV/1ke2+ZgI/6bVDs8fWVNdpvpaq4/PoB0V2Fk17sd
cvr0J1g1IRCC2sgsAjMehSDU2Mn9GL6p96+bBXADhVHlruj5YJxM2+qz5gl6RmWQwyvHRlTO0X7/
KuIBQa7PkpflULEjGi4I7Q5zb1rIyjWZyKnbueX4PwJOMxsfJTRFssCXuPOD7Kv1AbaLyg3NImKY
3k2cD8JVaVMey3cuW4Yi9INwdrQSZGOwnWdAWilFXF+ch9Il3lpCEB3v5m4dyEILkbj8lUj4ZaJR
Qxf9bbp8qEoqs3pEst3sLqp4cD1Y/7VlA3G5mkHBUVVy3fyDK0SL/xiGD/69isTJCg6VMq7oNj28
eoSrbj+aJ+0pe/n7XlGK4FZJFVlpY+w4tXsS64dfmE+szKTdnb4l7tb6WL+i2PDKY9kJ2agrHOps
+ljcRloVx7ZNp83va6YfwSGhkcB0B1yHqmyGellsgEtoR63LzaE/TiMe+1A+S9Nfv2WVdrsmeKtW
z+YPG+hU9e+18h/r/GTbsU5RIhye6lZxt2Pjsl4M9YG6G69z1H9mkTsvYhmsy0k74ltAYwkTEhJS
G4OoujMkqW9qzXUD6J2l5OaXq8i1fvl3IpHn7VQxZmaCCRa7W7zPC2742lsIG9cviU+l+6rjaLU5
FlRltlFuvu+iHissI0U+zTst9xlfR6RP1sNlKU9YKx7Ne2tE34ilt9rM2Q24/Urgz33Sct0IExO0
BAex9L9go5LF0EzuB2nYb28cVsJrOC4V8uQ0url6bH1bM7ISr+NvjKoaQIbm8A7e7pCjclETJOJh
lY6fuAYBD+kKR2yaY5L52v/64Pxi/4aKylQm2IJRd/rmqLNoLI1UZK6X+ydAB+kfSAZFpker1Pcz
I7oGltWIFm1xn8zjo1I6reS3S8Q5rvn2bCHD2A6TLd2UN5xR5kUHCaH1418e8oP1+9Tdv9aoBH/v
hux6OnACQvtUngSfnSUiuRa6Eodc59nycJf0FcGzRBhTEs2kABZUBIv/k4FfH/h4xjv71aZzbmLy
l7gn+r4/kFkE1oWPjgletS/36Wh7nRspY94hD2yWcXTfPswWC7eVs6B1b6wKrGPMS3hRsdepZDsT
lE17HQyi9feye7YkHK8ZgmUdv4s5HQqcclXXnpHX9s/NGlNvrHfji+FJWU3HchQAMgI6KpprIlJL
PK0bWtVvEbDnt9Z6iZobCH/mAZ8lPrvyXMia6YBTpPOsa3qUNvr+KUMUIeG803/sr79q+2Ieu796
+FwskoiKUPvoO+3S4burfiurzuU2rIAG7+bMF80uVFMgMOMjkK3FF3SbaSROPo1uXkYzuJ7dxiNm
o+Wpz6rcheSUR45jY6EBpl4yi87tCoWNnFHTR1IH0iVUbFfhCeGQtWu25bpGLXIDDCQ6iZ/rHsjf
iZn8cM1PVkTIg7UiCwdX8U+VXDJ51F5P1z30/ycqshjzYcbtaZHVwzykVXdBDIQICy0HUV9IcpBy
YI5CM+UKViaBNBIDT4wX6cAMRbNHUiVVZ71G7MvLCv400gQDxF+Ii5XUCNnZXUAhUyMGo/s9pHn1
QV84NUlhFA3l+rDaavBw+TqsIrR+Vz/4528AAKqACy28HZ7dBjrmAVI9hoDG+adT8KIVfPqZnTPI
AKKCfZVMhT9Pq1YuMDrKexniQRDWlUIA1hdNNgIORlyokfI1rRydHgGxXgjqBhb/op4GyeLeZPM5
vhjSVEhNRStkOQyn+WaK/XqtKyb8ilmBatbboQRzvgfHnlYwc/MKSsABz1hAQ/ThHpHY20h8j2W0
WUr11ZBhE17cJX7Xi+tYG/9NMigSTGSDpjELtV6nktT6cpzQdluz05ke6UMSOdCpvJXPblpqJfFV
3W70NA3EilkV7nKS8r1UfbAjkP6tB2ZsfEPiVBrC9vJwcqls/SUIbiA729VNmUYO0adaMG2TvfCG
4s+uYyPEyXL9tFE8zCEhyyJizNOVBL09AeDth6MRO9N5d1p+Vog0nTjLE1x04Kev/6phiOaCZbfk
CagDrkd5CkA/fjzUqqkE8bEAel84OeWQ4MTARJaw7B6kF7N7O90oM/6Ot+ctJawdwNxwzPlcGnZu
xj8tbG5DgnqPOQo6a7pECcVBsKHJLmI4ThZs0pqDc1A0xURvfCa+2ctCVmtE3pVUjel0DlIhVjg4
2DG4xrPq1OnwNh15qnYXQruQxSDHU4ioP8i7PUQuggrKlF/zhEhZg6QdnfHP0s7eqBVg5NlCeCWx
z7dv/gUmzDy7W/kAMa253yCRj13/N1vrYFk0wAs3wOj5EfJYEui2rkoL9myFC10BwUg2tckewZFX
1iFITrasC9gvpGo75x0nKMOdqcBimx6pmGvMEqiz8kdWbI+xKzcZeLlgJGeNPY08m3euCgx1I+x6
hGC5e3CKBQHKeOikM5AtrwiZG+Fg9CYkcTTEKQbFEc6ixu5Kj1hQDKP27op4pdgb0Nunam1TzQQN
eA3KSR7fHW6OiIa30A+NuCyTkI05I4FhalWnrPySNssEV+/ZI2xzNn+AMVHTJSsnSKUjhB9355s2
ygqphM9/n81EVD9ptvqOseCrak9qfLhNUJoT0cdNfhKcT3luSTYI3KDv3kJs+VefgsMqR9O6/hsV
6E6LBawa8f350W4zmm20Ew/0sbRSrEBPDWKMccJJWkf/dEKmqONF7dCckfABD9JEiZABClKq/qWA
OfqAJWC0GG7wI1+X3+J4VOmIMY0B5d4MnN07B/DDS7z9lC2pWlGQvaV61hpMUWt3UaK7gITO3FnG
90eMQkslP68GfsznG9bXDrY3ZVMwh5SGU7cfGETcTx2FqwdV5hzYL2oVxA1cYMbJJlE3I3uR5Y2G
b0diycb3Ax/VSgvsLKajyy12r40HfIjX5klF3hXx1ArU7PKUH3RKnkahzqoUjRHGRB2qpc9XPhzF
ud4nlBSJeGL2Ydv2q2Qm5RFAuGMNFCtuQG6TjsCjzfQZZJR17deaPRbxztZrHpGHk5tW8hvNpY5i
6VmJXD2UaQxtScg4RupqXEqrSG94TxwAL24R4O2wYSubYGzSRSnaQYWevpGnVEYxKTj/IoQvDNx/
gvyX5Iq6FmsWLxHGGaeVTonBdB39/ofxdmqLC/4BTsj+ozY52ermieWx/eN/N2zp+nDKju8gELyD
lGRrYij8m9CuF0duwplXuWSXUZPQgxRypGubu9rklvPf/y8K9V0J4x9XA0/Q+hsfMULUdOhMEU7M
27uyO0kd6LcKXYg8IcKGDsDAd5h4si2Gxec8PD6aQriW8VPBpnP96tOPFCc88ERnV6MVtFZjjoyy
943DQpg2qlND9ipBSrGjA2c9C6jS8aHTICOyPXdT9IIqO6pivFleuwXFSignKBg/Xo6BKvplglyv
PW+aA+/03jnAnqs6bGslLP8EyZgVyuup+l29cY+oO0+Lfha4syTtzBq5MIRFOBf+KTXIAln1rVFo
+WuuWmw76cRjqrhEE28Tk/4FBEQpDDX1NxhwkRlmCHmru/tS4q8WCwkXumXCo+e510FIfg3vVpKG
W6O7dKzCxEfkAucRVL/g3gPifzTBN8M5cAaVnMrlq8b7NxO/uZBN2Fu9iSsRXdjGePgsgJHsbpwI
R54/0WeyLc1FpRZR8qiUhtUArY7jUoR8ZhEeR5Yj/O28EcCY6tDLtxpgmrHeUVrBKS+vJ7ZNAW7F
L2LUv23ljda5yqPamfAF0eY3oaFJe6Yobkt0tviGHr6Xu6XgHHdbg8Af1AH87WrHW+TH09dPAtR2
d6dXni8IIzoRGeLa1Mh+Jjd6CU7EKFPLVivAM8EDDkSngY7ptVxMxr0Q/nNOnvILfqAQl8euMoco
0vdnolaJ6IJm9dj0sw6mgXcrAY72JpiTkfLizUjUysIDccBlVhZxA8Y3ymRRNOKDm08deqi75WVx
glBdlxbUlJUPG9qIQIb8mcIgXeXiTuKx2gbzjx2ape8UtSdxSG9PJfkjYY73ZdSgeZVCioNXSfF6
LwQo+Go3rGilbWieCe+d7OP398YEa4K1XnGdf9IbGQPafYDQZjCGyIfhPKWcVUOSmm4QFqWno5so
w4EahRdPTVXx3c6tara/KyvADlVY3NXlQARLiqV3ynm1bpqpmu/HqlLMtHoUM7rpmGShWbdM8FBv
locgKYgjMx1H8CB6GrjqMURsZdV8Eczhay9Ouqwjcb+ncAKhMZ2YRWl3Lgt1mrsJdIWp2uBS6gys
9kOek/wRW5sTCzAtNoixqTn/ORWD6QrJX8rZdQ3jJ9urK3iDvWiMeuFdXrxj3+U2hOP98gMWF6dx
3QZve4bC7i65a3S7SfWf1jlHaCd4IGwkuTfx1jx3z63BEs4k0F0bgCdfcYked1/NdGyT0XJNo6sY
mJMccSwjYXYUWUkt/e1SdlqVaOFxQBF0p0ICJA1OzTuYI0hF681VbbY7+XcdGtdwb2SfZk0vUMDS
tzXh1NQCtuXK9vnq7To+Orr053UM4BwwOUFIK/uA7Rl0JAiHLB+h5X8d1UrEq3Gucuk9MTg1JxLW
ziQ14Tt5HSk5Nwc9146YO1vo85GojHxyOjw1JNHksqQ3zvhU6jmTXfSBdTcSWJ8j0f7NMh+xmbX2
6tvAkvoyar1AzV/iYiDkzP6MBpbvqLasrM4Nvp+Ytc7WMRXpnjWmFiAqxXRn4wt3aBfvHfwryKYj
J7ziz5LdBlgQXqPjtoGRX8RY78TP3wfk1pcQ6G43tAg9GeNwhdqIYjxueBGJEThRnYjdPkY96ykE
CK5uXVIzq1NUEfu3+EqrYFQPRKgTSORHuieD/YPk/osKpPpxbxDGSvJPZ2lJCmyyKUXtASOaiygC
jGU8owgKFieQC53ugbHPShdAHFtmJ95Ufc7i8lnRrtHe1WPoWh3k3CURCCNLzqpQcdMKcM3i1Jpu
HLZjxBXJda7RdmNf5GoziSGfOQf6MYwhibZ4Ux2jojcT+ECA/mNLP1O1Z7ISqWcfPBf41NfezwUz
ciV0YY2+JcjKCogqZ1tYGpTAXAwnYCsTgK5DNrpFfy9DaCPBz4cWoZkOp4WMf3R5Q5nCdHSVnFv+
QC1a6hLez7WE0nDqihFbGeyfZ77tVBzOUoNojOtOFx4PsUubfJN56BOf1RPO4XrcP7cgoN9o1GEv
VlvGlChffsJ1zkK69XMUaNnrc4XCXa0Xgp31neBD8s8fhvWMMjO+Jz03VwbmnpEChu/qDBahmEiZ
BEib12zAhH2K8AAKwJTIxG49Jfv7PXgVUpIsvEfnDMVJlU6aUZMMSkXnkvgmEH0ZsMYqjxewaJtZ
aWecFMa5g6zqMmz5l/U0UTbXtvQpTY3z22Yfpim17h4oUePpdRrvxG7i0WFMpQzajhUleiwhUnlc
Y0WYq5j0h515Piy0jW3RE+Id+9QKGdgPZNmoZ6sA49W3Ytk7kwNy+o+BeZdy2XrI/6mrMq3reovW
TzR1TBc5Qfn1WXCWftZo9ppyIoIh/8m++aKBmbd9QnkWCkI6qux9y+t1/avpc9/qe67EkKXG3sMO
FPuHNL7rjEr1n21ob8CgJ35kQLn3/i3LRoRMx+Wz43TMdhue5/TlxbL6VwoqsB8v+EAMOMcSKa9h
gxxuVDWDh2BINXq1pN/itc8mTiEOnwIAC8U81bqT/CWwuDNQiGtxe2Fw2431fubYwIPpo9mMU2Eg
KlnFw6bWhr3flaNZTjgdxDNl5uoxGAG0kVLxeMw7FvLFeaJ0RuECerjeaiqkIPRGhmkAksn4czAU
TCx+uNGwzBxPc7OutYH4qoaNFV+SyIqecyLY8zzYQowQfe6shhqeQKBqlhHOhgUmMO5ag5fUPRLE
4ADXM6MRbROZf8zgmM/3PYOookD1kw/I9RL8s2Wrbi6xy76a+B+M1mvwfK09RpKuQGmHnUsMSuN7
ZrMqH8MyQ8vrpqQxQbMAkqPTS5kXsAUP0+GPbxqx+Ghh+pUqgKbO+tvalIFpu80EU6xLnBIsKRx6
wjrnClFYCttsZ3BZ4phJLC+IhJgPg2kRmlla3/EVTyvvvCA2G1EwiZ2D3P3ZWj6mhpt7bZ4X0CvS
PL7++F6Di7p9Mxw4ElIuNG2qZ+r3e9PjCPZ0CCOsuPCyBSxV/QgY2Rt+iHRP79nn9IlV2PKrrYg2
xepa2BRdGg3ESIQiCV6jvXIkdnKqhKgalzI2TdlPv3j/4ysh8FAeOZ+aGmxKN5he97GfXdghAUHf
UWw4NWz4+Q7JeiAoe0xt73ZZF1ZR/SwQpkABUB+pIT96lEMp4Yya9wQOYsfqTSM7FTd7SvEeVI1z
FscRGH5ryk9ewQd66O4jjsTW0LOn+rpJOZU2C5i6DDx4S8jY3/stbnVCJcVRKKf65lReEg/3pDlZ
qzTXtwXiNWUwY6gjPNWOdeg8F7utjcmyCHaQqObsHduejV3FfJvLp/kPuzolGzps1o41yLGU1J8Q
5qDV3oO7YUp5bq5tvrVJuLR2q8ORIdJ81qMp5ZQuFMtQ+qbe+6W0vBHhCTx2keK7aGUAOi3vVUwe
OMopx7vFu2OJ4FCqsmx5f2hDgE7iVidZuz7wjeg6DCZ5WgBJuVD1we7c4XWz5pM9g7tnPIVZeD7o
qAo8iUU8YJ2oQqbLfEV9x5cFoZiCPihHpVlsCzCXLcx5Ial7CUXhYYzGX80MwPqgfbLBETTJJlQN
VI64jclp9WOOFd5FJV7KwWHwkkspvRO6FyWi2ZygUEDnBrXQY+AMI+haGJkAlLOTdWB8LHsteBXA
r0KNKmgnbqV4iv+YxAPfTgOuOksy40MHhhNR/Cpsn8KiqBUS71nUvVL93Gdj7fEUntaERX7TZ6s7
3AYxqE9CgD7utvdQa4jgK15rwVlA1jaNSGLLQw5sTD7njqnwTEh7lmuBwOvKI7oe0/ylnj7r/qnA
Ipk0+S5+JMxnZlRv9aTa928VygzcxCn9VDO8GKH/H4X3lC6lQrABKtuZVS9KQbpoG0xhJFA8eG4/
FTaqlYNvtKrZQyMNkYPhxMnIWWbRb+x9VfQPFNq1DUVOSDbym6RKlHSm3lM4opfinjJVUvu4HLv0
ZzOiNftf3G80nnYy4QRe3xwzbhldvtXVSqOYcX3wrGbT+/gb0EpqmhwGXvDX56LqoEyvsPQuzJq3
S2Qtp7CtcZYWyvfdoyaTIwaeqAySfuicjUjzhRY9wbHwH1zYWkzscyNqo5rFuw1YID8Hd2CrH3ea
MW5vitutlp/Emo+zp1h3j/GGHdg8Ui5BnQ8LayQBugpu19ZSN0fQ2Wh0jqz3474crhivmULfBhqV
joSV9KeGxiLrcWOSuAdMDHFIzRsdFAgGLlJwLOyRHDNmTJ0aorDYNfAxG88/GGw7OEvpPJqifJW/
4YfkVv+rdMUDycqLrwAKq5/48VTlmeqMkyloptB0X5xKRUwZ4Mh0zGigGEZgBOIwmobgpq3Pk4LL
y+H+k0zCL/5zOFakJ1k8dd1oicjtRa5FhB7eFZdH7hWRoJPp3Rb9oyXgQMwdz9vXFW0lMoFGyL8j
BcPrPWOA0kXg0YPvO8jpRJQZBwI/Tp8J3KbA7UQ59BGDZe8wDvjVvM6Pgh2SnHZwyY3jd7c+XFVU
ocXeXOssOp7pPzaa954/bYt2urI01+JkqxYLkcCJUbnRx8pTe5N5BFmcpk+HFGFnURJDZgiWwHAW
I/iQhe36/BlHBRL40pYgJi9kxsjvgfc5QrEnTf3VOF7wtpnMovHuJlSaxmmi/C1NXA+xawZqoePS
Yrvo9847Jo1e3cK/Q0N0CYTw4LKNDtjZh+ZodgLtd71b0KTcPA1g60rbNPHtWBVbiQ2vrOUQNvHg
3SGbS9yiy6FfynxQN0kaUzng45ynCX9KIp0LbZy1VkEBgqbZz50z+D6fhAHUBxw6ozQq2IOzDP3N
La4DKyTUUld0id/JRH3WQurzzO84d4LxOaUVRFSAkEuQh/bgohiS1UEXjZz40G+nBoatbCJmowBb
3taiEtM+bx1tK7LTkbvMrg5Hk5w1TEqIuVdF7CAnXHLuK+5L11SdOmOuPSKFVxeagfeAC8mlet8T
EGwzn4eoH6xguKIUhPIc/Sc2w1tktWeW1Gv3tLXr85gn02+zhrcqjwBrX/sl/gP+DAc73i1YvoAA
6MQ5IpxcrfbyfDN6/1aGu5MzpAQjIHzlTcs+RcXp2SSraMUQwWlUI4SzCh2FlYjbG5HWCV7oxaLD
vyMhk2rPDdowh1HGsD85IDWpO/B+wfCQ8oEAcyoiDXnVsTrit5RcKa712bxu0i33lxMqkhCUlSgc
QR5sRtUwtO8re3BybsJzp42UqL0zM+m+CQXfnTM5wvF7TYpB3YXeJT3Hu56AYM1a4s6TnvOjUCyz
qpEyBQdV6CrjLymLwiyEo3mMiYF3Ln6PsfPic4wo+AnotaQybJhjfhBY6b+58dj69z1g5dFig/kx
d0DSc+hEB9u4iY0Czi4izWH6mLvnPEoc5i+p+4kFQlbPEoxVIDY/LjD9/SmQikbv4UPsnWDr2M7C
Hz6yas1R3q9d45IS6GAwydCt4RGEYzHxnZcRx5uF/BJX5MfZXkcmXUSoly6MJn2yNTSFjCJMlwLr
s9Xu4jwhJYH30W9+wJAC0TYJmJHawju3//gn2fy1JFhsWWOx/E91AL9EmZbEmZoDG5Vv8qCLmsaQ
p58yszhi0SNfhg/EsR4vPxXaI6PR3A420yP3TXe8kMEdQCi39zLdKt9PP49PU171hI7a0RFZfKcW
czaCf+IcWP1yBhZf71mBWYSGNkX8woohMK/Rr8zlvWVQxK3qz4nKJ1Wo611K6jkHg9LEOsFli+8I
+QtzYTjLkDKLTvHJTxWQ54MwbeZGF39qPhC1okFoxU7GIb88V41yKl8z68c/NzMSpO3J8xWIqWlq
pIdRs94875Jcv0NkNt8/8CnWbS4MEDlwhTOT9NYAFqp3ynlIsJMVoip6Tt5CoKTOwLZ+SBPrzrc6
3CIkUr/ejvVrbK6aXtynrSkvMpjFlJjMhbt25F3eJWM14ZRwlTRQDKdQkzGyY0ZpKKrKDy86mQlm
04ZgnOss9dvvH16R7qS8h92uk1b1HaOn4lEkJrzezyCyYvKjdoZJkVCWxM2DoARgQyEgDAcBzSQJ
ATiVIABL3R1yUIbBmYAkV8PVJo5jM1hfPlT67FAyuCCLsVwMhlj72tcSLonQEiHMiaZYvVLKskz4
Y8+RsU+QwenM+r030qr/d3lxkG/nePCMd7RAiKYG9FdvHAcHFhNmmxBk02i5YA8lUmcSxkV24PjA
pbMoQDjvCy6XHw3Tk0XNsVaIBbsigCl/0F5XDFIyXfwC+NxZbv/0Fnvc6+9Rz5QkKXIFHVIliYWJ
9k1iGOIG62dRJGZ3eNQy/71rUcSfs+ADUQJ9+yVzgoaaXmItGyrcxGUQk1yamYOzluo/tCa+HluZ
m60ppJw4vHm0fU2QGUiSp6aFQY+SYif59pv+2imiNLMa8ewctnf8caEHaSCAxxK+USpGJdN4O8CB
VvcrGLaM4WKscZOHbvp8g5GmUgIjnMMHzKfTWSExJ9CYN9rBtH+lhRmo0uIbDLPWLSl9U+GSuKzD
Hg814Azmt6CpjyhrkX6Tgp2qhZyASyDyOYL8OBEpBhNwTvTmPDS6uarz8DXdUER0up0MM2KLcjkC
IjLWSGXjcmVZ5R/VjIfWXktizHehLlmhSESfEBJXz+BWI9Szko9FVc7n8s0E5aIoLIOhwKQTLQ5L
i07YLIwI5ZnD3yTqVbKlF3vt8S02RQtTmwRRB+Mi4MhYgH5r2QSyLsmdoqW6gh5gTNQiXX3h/37k
rp7Jmc7d4GahwSFaXzJ9KVPyLe7vdzpYKjWFDJn8GR97d6RJPIhF490kWJV4FyrNnUzWL4cOjVke
80XyyHE6GCaDYIzHnr02JbtwLk+Q1J9LW+pqk3Boum8CR2KEp/9CAuVyB2lNn2O19k3aj0HB+DEF
d32OM5/51EocZ4SAx1lgTvW9s1T7cDBLVDilP+9836o537eyu1rzYCAz75ITLBQROcmHKImuNe6S
NhX13gpayS5tNWhdEzwh/y696zW0/4CBLcOmT41FAzUOTy/ei/cQsGjtbUx7UCC+6OHQxRhP/WUh
c2U0hUsWYxVfW1yqdPT241bPjS9uYiXH9L1O2bSdWUmUlCEyoCKUPMFYWo/QF8dOKR7B5M0QGGJf
anaWb6FWBomKe/Rs+ShLn3n8KvBlsvHm8n7dtSomipx3jgvqUV+y/UrWIEDhmhSxJ49ZsmL9GccT
3NI9u3OjDsuiG8vxyOkwaBZcGzVlT7hwtHNvpzGqdHbEzaQxgV1mAMLFnBWDbVeucTG7Ckeh7PzO
7XfL8UeQGLhGGVOcNi5Exn3Z8fy4ozZHnmzbAA5UkHkxavS6dKCF8g7e743/A+W3NjrcuDxWiizc
iI+7y5GhAhTII9plXWyJuAWPUklzYaGTpnA7n8d1jUCVrpiapdFfKPecgB64ZYGjv59FuDjF6eAO
yYg3pTz/7snC73F+Y4EnMoiW3fjFCW25G+hjHF3Q3h+TFSzGhgAxatsN6M8N4Cw5i45qFkjw/smV
zGh+gxbgZoJ8jMu6Rsv5o8IKyCVao6hayC1IkGnx59Xa4f94tBTNKqhme6YKlIWCWRvlYGCYXP/0
tkdKoMY+KdxneTp6KCKEUYhwLYtBzNXqur8dmxW0RVSXdjtkB5gUATQbwCc4yB2z4FIyutwvjg3u
PA/EaK2sgeged092AT4o6ULxueAd1+GGA2v8v/vBfeDMzqf0aieqRCKj1bgLUPuyS8SqiAUfg9XR
d0gKc1xrpWDWHPP0OIuxPV8CaHPvFYZwIRF+MNsbPvnpKKkE5ujenV29778XKO9mMZi2DoIgJM1B
CLN774UnAX+FWAhXa6HA1Lv7D1UOB2niYedQQZjuWzeJ8ANSsgTG9BHzmSTy7OB7cpFna8cbqrWm
M3CpJU7AQ0t31mW6UpQMcov/MaXvHkV3Z4ClzTxd6iFkW5GIKmN4fE++53NTDp4etiG0jtiM8gUg
A8gXdaEu8KLlMEI9LdLTC2Jwcp2Gi37WMWO3DBEMapJ9crVZdY5g6PkJwvZXhCkh5CWgXdMij4aX
nzQd69xu5vGZYrRnDsJCtMp+LUl5WA67I1pxeqrTktFU3yV1LYXw8o4IX7btmWq70DkTAdyrQ3uY
p6lHOUNewGGCER6vzgS27i44Oed48oJ/A/2+WoKUoy3jCbJgXwwEsNbbmeIgQ4t9YN3Dcmj1aKAE
kH7kbJe2+8z/f+7KcAGfCw0X4VgmI65kzRgNo7J7M7WFlsb8umuInTBIGkBfwmX2AtW2lpXJkW/f
FmgGCpOwxZgeHg9YAT4Wn7ztpzbKRR/i0BysqDPcMK3h85DCOwJY5wzLpmuCXcyCmNYCwXecrHxQ
9A861ozpnYBs1IyLZCjjzZY/woABDw/LcGW+pffQwyWCzKfmESDjituZvUZfgMfF9WLneXqa0wjH
325IZVPwxMDqA78YFVZsOS+pxvp1R6GIadO4kM28nU8JBO+oqSWm7/+UQgtLuvNPgL7aSWdSh/cC
FzrUqASFhLgx1GdowAq8Vhl6lObPQ776AiOicAeGRKQJnXeLySyLZTOfJNYisvVJw/xc42zPjaZG
it0H79a2bY2hI2hbAJW3UBBRaPWbiJg6V/8DH2hZPm2LIyU2LqcLbY8pNvNZiFIqZmX7x9Q6qKDn
DzhxKkip9B7X/zCKh4r6zkAZpEPKGbZl8Qdqa8u6mvh3MlBclQ18si2WUI3ib6gMx81F/EAtgfJe
NqBYi/i4TnRnYkvknxI4+PiSwTeaD8gWj1r35d4f03o7yYp2uuYq+OmB970Js2iQYigNtf8MSJYF
v5FtMoohkMaqvJQwmYqExtTxLiszma8divEoiT9TV1tO7izxxpbphNt/dwTZ1w/1CY/KuJbkha8x
aaL2drEH9CjTn9HI1fB4n3IvtqOjunJQSn+X8H40lukhsIHH3xhYU4PZ6KS3/ew9YlDrxwjYNW7v
FkevdKDdj4i20vs0421c6vMsUzfDKPLCmrw6ZB0Ig/qUUesmoKT4tIODQFKEfbX7Udcxnwxr+xc1
5W9AYQuqlRPxNozyy0ghqxXnukVVEDRc0BlUgrGdpOPxPFM+/9XIi3cziqwYzMmlgsGm9j/tkVBL
j1PcSNDjseQe0qPDj4zvcV4cDuTJ/xcIngBJ5jnxPT56vV9kCfGQ26Df67BjYQejY+vzH9y3MfWj
d72ZU1/bWrDWuzejM96PKs0bNatljvWjrY9BMaVv2Bm93kWd3xkomFFKfhUfdjfX4ma3GX6foO80
EX8I9b1hc2O2YY2xIGLjJtqxC0WmngI9lyRC2lys1M7+m3cmsIufPMMbqy2OvTxHtylbPyCtSjv9
CD9vBZQN50KW/cvvNf8Vu309P+fspWwBi6/TSqSz2m/yP50T0wvPayMn5QaWmhASL9E5s9qkLC1F
5ROjlYHfnCxOG+64cJzhCziyrjv+Z7wP7Svl1KEVMTZSaepjeP7WOXbOJWtBD0KKbjf7a65l4jqe
56SsM+3PosCLwQXAFSEDWu5sTkIu1Ia+3kzpdUggA53NyoZEf3A2G8cRdwksMuzu8ZyweCpGxW5G
N+RokjX0rXrMNWs+6JEqat4dmQ9F7p7I2dWuXC9oIbsE5tw/1IVQKd6vUyokJM7HXsPKF9Bvabw5
Jks+IMp2Xlr9qVx45n0K+wa/swsHMX2rY4lglIELU+ypWXOyWbnN+h9sstV1LDqsL+/nrm7wxb5u
DWRbN6BL1gka93VGoLpGws5vql4JH68eswTGlOVIIqWvGZ+Givns4gF2OPowoY0utQdXKcfrhekV
iil3MUFMJLfclnfEytQfTfe45oUu1qJRAKEHZBuL2kTdANl4AV9Mf2sq+xZaZwmWI/v3Zl3X1Bo8
0qxZy6UCDJY8Fq4UwihOuwGKfC+JbQWB7Q3bHP89O1IgnY1o/El0pyZieseIX1u9wO6sHE7svi/V
kWsnEvZiZAgmudMbfBUg1eRV1AlvmmHkC8OAgTlPImVZxW1+GA3Ur5+TfYPctDe+O/dG/0BFp2sZ
C8k+Muk5+61Hx24zPN/MRZwhOAPOoXHMRvU45YDctimfnFBBbpPsVwa39cCKVPLkrldmw2N8CTNZ
WAhln94EeQ93Hp9IoboBhpAHbJZe53s2MzwbkBtv4bD2+uUtLtaFbqW4EkctYkEZOx04QDt2nRVt
ogrGOZAoYun3r+Kkd9GLNCI2+bbzT6HSa0ziuh9hqY8IUe3e8AnxSfho2Sl9mGid4aPlc+vKt5zP
AM2hsva2/xf4IJ470YPfkZs3BhcXUvu3oAripkC/2/vw9J8DEzoQ3pUS+gQNsuObe/a7T3ZCkF+i
+C0SUx5n10Z7SqAZOHUH8d7+sTd6oP4g16V5y3tcTBJJSEAwpVwmAfKVERgzqtMXEked7Sa1KAnr
zH4k5LITXU6F9shhOGRudsKiTQj3vBrcg5CuN7W47lVADckIiSLfTCo5CaqPdZ6mFp2Y6l/rfRf0
ebJdS2oEpzMIe5VS8RDjdv3S84wsARdyVr02PdpVnQ1Bc6+n+Ac/KV/xvowToGagUxiDyV4sp1Ig
HqYO/WhJG2Vtm6l1r7ZeNlyzOSt9JjoyjF+kYim7y5/gQq/ufesJYIpnlWUR6gi0PZZ87Ltw9abg
7IhL1rlrVf9h41aTLLgrEUnA8ckrV6MnXNkrkv8MYKixy5/U0Z8nVPGSeqq6GeO3wWq/f9NzCkQ0
CE1sdzpleXW66YCEITEVKs8n8IoCRkfTMydYWo42cmcFwYETpN0L82q2gW2bPH+YX3FZut8oHJAc
wkJK3CS+aznUaabZ9OcLBGleQ8ZMfsnS/fdAJO1Qo+dYT/n2cEnJhhTSU1yYC1wepYYy/2z/3Lfp
D9car6N8o1A3bjUKt6qY/XNYR7nPll6XidiihbV9/eCKD/MGkhS7fxCnzFSMckIrJ5c93sxsrbkR
zzYQDTlcT3ptBpQ5BkXOr4urHVihwvfZoUAsN1Cp//iWIUoknTflMiY/xu3Rcffens2ZqonPA6n/
aLRGtbrLFXQDkbKu3d5v0qbWgFR0Dgs5XuNc/eRU5bG2Wmb9GofMjvF++SUfw17NOJEGvGkDqVDu
Nir5IM4BciYEZkNTghEx8HlrwCcgtwvCv5XHpjK7vYA+dZOXprnpZssPVa36TAcEwOTxnsgS456F
qofJD3WLEXiUvkN/mLUdVV6OG5/soiYfcaKfh3hZ8wgnuE/5oINOKw6Ja0VojpeT2dQQv8YgI1x6
jDvAnj8x7veN0CDXBlzX9loiV+PjWMkMHGxzE9ix9mByyWHkXo3CaLCkDzPcYcpyP6qkg2qPNALN
4w9IpRH/MtUJbDb8cKBmUdwZFABEDYih2bnmijOTeBvDLt//6dMCDJlIdLQAIEACU3ismVHhuB5H
D/Mdg/tptislyREW9S8Y5isrdU93Gh06OGqlPuLAI/uBXylLZJLjG3UBjo2gWVe8apcL4eqRHXUK
X36AC1tdRjT/V+DOJtvENZcH+4Q9GKqUrt7exif2/3SwYj5X4RSPFtyUIDEAosLCx/NIGGfiXQpU
ukq19AQ2XHbF8f3fVoVSvcY8EKfhfYQM5ilfKw75H2iKH86oJCxyen9X2IF4wUW5ARb+idzm+jE3
cDWJkvfNQFtrGqOgpTvo8ahJWGRhZyFxiY+oDOWy0Yl+1tmmRsRtRnN8XhJjGsCIrbLeoDL+Yqys
1GQRAqXIBokiRFRiKtaBEfZW8yvSMsnMB81RgUrWOgRa7OoeGKflCd8Tk7xhsrq2QbheOb0dyTOX
G8kUHktUfVi2Jvpe7Crh05jB8Q6fQXg7SrteJD85BtkdufqSfda6HoVeRGNFgPqOQC2fZ3ecXhJZ
XfO0wxtsd+d56NFROmJCEzbB6qysG8xvFOJUeSk5Zo7Zi5yCzkGISfBCoFZqdR7KyYiaFHeM+fTR
FZM89ezArDPJ/2jYZIBJ+ovEAJ/6PDYPmecOwIVvUfvap7cyJtk3OBklNmpXwFyA46Uc5OgoJhZX
TPUhKFm14STCwMgmNUmW6ZFOYNeyBCPrz+zL/oIhzl44Uy2ZbmhQkET3Ob3s3/UvW7Mu1HjPcMYQ
77ul5D5zlQqwG8P46DfianVPhU1mfktHlPSshQdh+f+JX2na7OLR1TicI0XKENTfDti0ZDlo/c3F
UbynXTf0UHkXTBbBCMuYansIdoKCdlGQFYcXWbBDoBv5+S6JP4znkaMaiexdyfL9AsqVvI2ABi+g
vtvOW66GBOke64yfYXNaK4UMn+d4Nbql4aayc6d/RQxrKzVzpTwyaKnIZKhCKwex4PrVuGup0+Ta
jc8EV6becX5StszDy7JEuFFibYKOzE7vccF7AT1BmEadDTnd9MtdKvlgscXGFTZr9fW/q8DZeSi5
3/84LsaOwiNRbZJq8B/TFOwZ2jHThJqXRvRE6Z/VkS7soibw6JkRjeeKwCSct0MnA3KSVbjjjuX6
cVsatdd6eol466GU37C6lskfTkbRd+S2CJuTZZHHwGPl8LApCeCthKXtY1JZGribZZlot/jSomdc
7YrsI7a0BAjTpmxLuRmde6Zt2L2Gv5oS2zjIWUIbHE+Cb/Oqtcvj1x3RERD3e8r+EowlSp2uWwno
Rft90HxAz3LGlIQt2P1ZfphWUZ5YRSzB2BpAu5LxrhmelCp2FX37xZ+EektUX0NtrIeu63aGD3UJ
XB5YjrQy3CEVmL3XCcWtmqqqrtvYgbGh557AU4M0DsYjIVrvqUxVv73T7xE7QO3w0kwCWM3bMaUv
wk/CNH9zZE/z7U7H6OpXGxo/oPnMqkGPciG+3/gmLokaY8p5owBnRyY7B2b+d/c2FhSBq6M29dh/
9UXYnnPLscC0iJZILCX2Q8kZW4EMdze1dVztgvQPuzlAniisMlyKAec0V7UimAz3n25RhL7ug096
Ispw8bnwY2eWghRdKhtlmRfycHzwmeCNrVazG2dllL+0fFnvB91hABYiF8SGhLH26bTdBAO39la3
XMfZ13OswPFBt+My7XiXiWo45/2Pmmz/cDs2jpUGvxkvX9dqLTwAwqgZj+j9to6B+wZhjX9QTN50
usW7iTmSpo4kndhPjoI0M37O+vC2zi2WGdfPexRXRxHwuM+QaX1aPLDn6NgwZQ9SbDZNnLCTz7vc
gTp1YOGV5GPmlss5iZL++qtrWOrubcsty8No35dGW0GvXke6Lj6jeeH4SkzYqK0ZxNtbUHLrQw9u
9Mki38xRZaor9Dki0uU6Wwz9Mr7SOmJroP3zs40Q/IaNMO7ShZsF/4YwclIg9b7D8wKiogS1FxqU
j/hPw43RPVuSOWh0H3Lcm0Y0BCoIHWA9esUqkYKF++AyUdK2r4SD/whFomFm1CGnkW/+K39VWjCY
F0QHuusLWF9zhsVWzQUnhsZDPeArCelmIeuzbJw5E23TcKd4WFz+PpAFon0S8HLsNPZ3jEut8uNV
iVLuVZB24LLOmuEOj+Pnyx7a/UwQFZ3Nd0zmqb3029YWcutlMmqdRBJx9ch2DA1yL7V7IKEALPKH
JZ9k2RnrGBuUGQIddWNNjK0zcUgyXA2JnuRjPEHmLTyihLq1m55UNygUhmYytGf0p6W2U5k6Kx2u
Gpdt5Y+0GY91I1mLrcmTtQzjzprESl9vUyV76O2vCGNAV3s4OB/mkyjkTMRxRUTzsVYOUXJUOxn/
PNDLecwcP6rwTF2GwlVubWdMCxeavf28RhhuqaQydHrzc/6PnOxws4cM4Vz6+OTKNJVWSGK5CECL
seVyYPtgOZIz86dNBI+dz0gQsIGwslsF5PUtWVOdkMDGway4MfLQ1+eQ/7qRqQK4Eqot6hX1ufTH
xy/1QzFHhgeN79CBY0jAPuIaeClWlif/f2KtkEF6+K2AEeQtZO9yv03gEHRquv0bTRsMfGKVScaG
J3oeL94SJyLsjaFfEU/Fu0sH+0zxZx3X2yuByORrKSJL6O5LTIW3aRFCWaaTa+M0bW6H6xqC52o5
vx7I5s35Z3kN9FXXYYqItAxy7HR2XZ1iSfmmGAFhHy43uQ8+oYdykgvoanhfj23HG6JId/rEu0qR
GPmrB79v9DduSF0p6nypL+SWz8R+8MOlYk+eCUbpPeV7iYLSm3gCZ1QRJexaiJEobbjwts2ck3bt
spuuUOjfNuw7umgYjW2/IiucAtSrqBhnj9UUORWWrLtDaLBCbpeiGmSEUvJsZ5YYnF+f+TwFbGv7
ZQGFYL+v4b91rKounzF0VlwP+WcLsA+2FtozzOeRUHP+MQDQ5ZRIJsYa8l2/O+3iuocPc6BY7Q2N
IZ6KSRZxLJLCCKQahruzdL6nR9BoxY/roTfPz+0av5ZD12UOswp8ig8uKWNa8psLU/Neo8cNgCl3
gJiivjcb5jOPQhMdrH9ABiaJ79s0IGUpZZNpmciPyl8eF48QGOUAZJk9RgtEfJkUFaMvHFeSsRmO
u4TS3g0cH0NpfRJoBqvVcgtqXMUMI4gaEjqEIrXJnE5OpjTBWGUrfpHZOgDIKhOZOpH/1yC60IcW
0mdfOwRa6k3eZCnYRUh080XIoAcQTiZmTNUTgNDpaJ9JVa3u3aoKvxAbYT/JjJu7C8Ar8yS22Ide
0jsKBh8cSisTd/W+WOU9N38yF1+LLlmptBYpNtVvGt4Sim5HPPftg1kNbuhZBIS9PSfotwoFj8Gy
p9LAdGVWdGL4DeDvlgAbsOK3Lb8ZMtk37C//FP5sKufpiuiiq1DWKDa2dnFpbVC75l/kgrdZVEQe
GWmA6RZLzoUjHr8lULypHwJi7nOMV0u6RDmtd1Qnch+gcntLIEEdeAdD0GkZG8D2GMjYP4Zxxsld
uFpNmdpfUp8fvdtsKPt5XI2eKJ85jrVNckmpc+yxOUgCxn6iJMRyZs2sd7yzwjaYVUhB7kza7G7m
qa+0uX85Kr5S03nCiF7EOnCFBmsLciUOUtIF1HAr7rjX1oQaUOkeos3v6NrAGWGIVDN67sXtGTu6
3U64Qn0VChC27MmReUhDuu++ino63T/5pVvyLATqwOzNXievW66XTZT1GE1rFMBeFu4nJebxemjw
IPut1jMyDTSBJA1zqVPGzn5HD8JMYnN/DtrsUDsQoqG0ltWwhg7CvSdSWesnmqYvNYO8JnoDFiMJ
spL/OSJjeMRtLYhxmvP8Tgj6Y26djJCRwD2lS5k9EmXPIUf6eC5YYTbaAo1aupr3lsdDYQ7Vv0u6
BimrRmKOdizMEZJICxxpnbzOSKq0j6QNUTs86GSFQkDew6yr+b/5mHYQnGc4w9yu2D7any4ctBcO
JW8usAVuSRhVb7z/mDrVk9G1wFctFsA3scrXwq5SML2QOTF981mVlMUL9NrYlq4quzk+FfXsYZoX
rkj6nDDqAm/zqBDDzlKwo2mol/DkVfospn7LRElfnL7rS1Yeq3Zedbxjh/EusxKrh6X2PlQVui3H
LAX730ATY2ZMEhre5EzzrXM/rZ2hVm4ksWIIcddEXl3oIK6UUfORRgzUq4EO3wcJpqIBwFgv0CEj
z0gp2FlssuZ91yUOEXxdVuZeS5YtBqKtSX6G7sul5LI7EK91tRl2jokLHqJk/wSvjSmvAhnpGPij
MJBS3yDL6c2Z5yD75dY8wBbwkVAUsSXDP8DTFEiLwR2Qlz9Fe8l32hjOGCY7Zwakt3md+AxczHbJ
q3teEahBy59tOAc9edflWgtcPWwhIyZQrpUAE/q4Y4HwxcS0VD7ngwI0pGzqyrVG1395+Q4Mt19v
Sdk/VoZLbxA714pQz0Wh83C0QjqW6OijxkWqchD5Adgw7iOPw6VViA16QhDnZ2HesVVw/jSzWfL0
6hlaBn/Boopfgt4lUHqhQWwSvbFWQuR4OZanvLlEbBZXw7aJ7OwMExdhT5TAADU/32h6aNT/j3k+
p5TojBIT6KD+WTay3VLpoOfrwdUjDORzbNXijDMvYHd/iiRGFVmvLt7rClizWEi5JvPNfRZiu+Ts
GPpsN0PG1zdtY46huYbmguOCwyqLCANrdqJ4KulGaDA0V8W/x1dpFKJuypw18EZQRs5TXAmGNvts
3Ng8Q3W89VT6pFCoGYJ+zlpOpC3Oh81OhcBQWpvDnlvkEoH/ZqPV0bAUv8ny9NYU77l1wpnwapKB
hK9/1fmPtDXvgCXwRxWv4202jpIzEdX5MvW/eaLVBUcogukA8ysR+giQDv2mkdQ29xmyvLQZvkDJ
JJRRSJm9N2F0Rdl7c+sQSg+HVP7qXm8ElI60yvuZTJHZhF1fFgZIpVhuuWyfCEbeDe80Q9Q3Cl6A
Xu9vOdaesgEZmhH74/pFoRK8oJAQ/16A31U1D2bFLOgbvbNgMoqaSxQhlC5OrQnG/1VxHh8DXQYu
CJWyPifldv837dLKeFH7rnj9MiDRUm4p/zqoLn7aU4uzaOMGTUvoZCqEfhJHxgry77xUxmDCbXGa
rZUfzzSnytbXE0N1duSv9/VS0SlSS4A3HNj4Gzj3/ySQjFXt6GzZCfpn3c1jeM2fxSW6aI9e+fni
Y8oWN1/LkkfqXX5k6oLD0rbWT5grn4meBenu7U9ZIQ18/L/LgjyF/fIBhZ+zapptb9xKO7emjl6r
PqSiRfO32tFmknSsm63VsFrhM9g4/ErpjlR19DZToJU9kZBPLnrGl89Famm5iSUPYXgU6mFJBPX0
mmlmVpTpxYcziffTOQBQX1QMSFdNwWoIntIylyo9oJqZrmBAxRAkVST6E9IyLxLLQPULMeObc642
8Zb93Ois7RMcSzSgNfjEL/76664UQUqoqEgt8moFRtQkilBc/ntJJQzdyjd2kCf9/070/9tPpidf
81vKSbGtQ/zm10iElRVXbmBo5Tc8Tr6QZXEr6dm9BJiryePh1APj1KAtnrPIRoFjulCELJISsmUL
PKa+SbV5h+LifgdXzQQaL0LZFPwbirjJS0k/9A7P1JKtJW/a+EoH1zcrh2JRkKcRZbF3qZ4VB6JX
IdEaBuPMnqlu+nJh6eD5vep6f3/7/CSd6CI5rhHCfD3TYPhAkaUbMU+eQNQzIAl5w+HhgPIHgh4P
6z04OpCVvzwm2EAMHjswvtXaI0hpCY+TZ11vmX3g0KuDcRC5dcN8Qo31AyTMt7loFi5JMkWys/zd
eTSHJmfYWkHbHAGQd6zbZGKgmbAcBaYORuVVVwAdZeH06FbCkxJJdBOs+DvZZoNXnPQZq2g8gU+j
3q9mxrlB8U2UjFYKm0YQH0uKwFBsNi9Cc8jNLoMDJF0RRltj7qHqqXmP4UFKDVWWDIdSJM2eQF+B
Z55PdLBTpBiX39GPZrQ8oRm0iTsTVfSrE0CbhmsTBf8aZ1jJPXnbVr109I0QAwxSC2TiPeTAVtgE
0PzUXKBd1ebZiDkSGv7yBPXdkthI+gTpgLprgGNrPxNmFc3dGeiPFRSI67vNS8zbbI4wkY4eiwkq
PkVPl3P7YV51d7sL7mzdgjy7M2czs5W60I1ifakoomXqwHvDFufL+Sj0uicqMRDXgMS1GX6IxC6i
VgB9aRXDM6K+OCmZMPJzkrocuWeZgl7SMcSXI1oBblWowszvD9crsmAlVQgaHTttB7nI/c+Y+dla
qlkN4Gp20wkDbwoqqnWQSYhrqvC2CjqJGgbmkgvzuOOU6jDk4S7+kjuC6UCdy9Vy3u6MsO3moHdm
SGL7PDY1/L0m50seG1NBSgxzvTGBACk6j4BTotuG1uHzdsQIT/NC7dnVpZWZF6+pIwsLK3MFOGH9
shabDL/7f7oWf3tGzoIPeeaxpEKcbchm/lOnBZ4lJ2EQ/eoH8FdUjWLsoH0e9vgAhCs0gMHkMu0Q
9H/YK3bKAGIv2I7Ln13vV8GIfCZggaSYt4DX6uUcf6ObGBmy7CfmCW1/MkNx7PdOySts5BhYuOEA
Z/8VKdkoUKTjvRE/8w2J4eNitit0502TNSAep4xhsfF/sypnSLDPi4aGQpwBCleUva2Qj8wIo2oy
IXNihsJ2oAH7pcxwxxUssZRe+5Z41eTLE0XyAhygH2a8ZOd3yCfUSAm3rErSvAmCOcVKFnANp6tQ
2u16gsOp5SgEpiCYfnpmy+G16tTIqbQWNQT9uGufECWjg3nNm0NMiHaiOzb1hIlBZDv0MpmQs6Gm
ZjiyJ6KUTwp2a/gH1czQDOuI6x72/AHUVkChFVqE17GzRfoX9R9GOaVJiTdojNbNGCKWXpFRoKCe
ItOdyc9igzWHscdXgr0O+0PDgjf4ofavwXwNojtfjUMDOgs1mHa75wDLjW+panyMtIVuEh9od3FH
dSembWsYddcxRRqqb4mlLINNq0RM9dmrE5Ehu2hiEnrymPhcf1x4XH/E4f2O4wlmpiX6h6RcEmyj
AdEt5vg7EAxQB5nKxNW6DWV7NshDWE33LZHTu/dFXQbMcTsvJCIM7QTwvxDOmXW3ghVRZPH0Qrr/
MNYH/Xnb9su1ZdS/EfdM2swPepFTfwjyhAvjm2uU70/HCy85UEAr6m8ZV7YtQUJiwF18V8BR6vbd
sGTnOSM0Nppp+Srvpv35UMP1g+3URo1DDcPLICiwkyE5WZUuu5HQwbUfhegz17PaID0bXTy09hB/
ih7RqvJ1Px24gmAboLPb+6EABCig4S+h5q4txqfWHHucUATi3Oom6CyVjnoXO6O4uB44SamWqxZ9
CJrNIHK2ezXSV5kE8ISfYodcGkCJiNhpuhImXZQy6RbCtE14DLtERYjWrRjwBAsa2Vs/9cYMD6dy
vew4OwP0NgiWKFgendtvKF1UVEJud4T5WsVNj8IndAM8LGGli8YTwCktuVw7eAYqTUV4KAwdsTL3
ZaIoB9OB3Vn0o/c86VXTlLCxMVGNuNu4aQwtl3//FcJNWQCGhyXZDAn2qEII77y7Ct/Hh5BTqXAi
ibTmV9twc6VOU/NVLHFWfxaJdBhkRaI2jChjN8w0ZAPSLxmhCbBq1LJD9zX2zJXP2PpVeZdjJCv6
iWYU2HKnsO7GN5JOPt0gDs1pXCfAmuwgm56htwJV9DuxqH3yo8wVyllFW4R/wr4Ixi0JaHuVlfXL
PpadF4kxlrpaCVMS/tLgAxb3NAdb1zyU4HGWyhXsZQweciA0D09NHzyUqOyPWjNwoaO158W6Dank
b6CylRKkk6Xy29+G1XY/4wROPlQ0xYdxLpNtGcA8BioPHLEV1zlcO8ki4q67iGyklpMzHWQvjynS
es+2WND4mjLTdeCIjAnf1HI/XGe/wAD2dHjfdC2OaDkZhqpf73nMVEoS6xN7VRt73eqTIgmlW20T
1C1WFJGbt+WL3vGYZRjb2s61j4OJj/GOhLJ3uaT2GqOdPm9oc98304acEGWTBdZRukPudmysKCVD
MGTUnmTqRLiV1RvM3uXPtYcybymvjAARN5KgJqeRISpNwy4Y6FPY3pJIclALPC8LfA8UigCSjlMd
WBfS87VNvFuyhst0gl58GfkicLmxZtgG8O+O6y2up65o/rL6YX3RHXIXz+jsp2ndNyrCveiDOtFc
+FeE+1jqhgmVIAwLg2pEdvI7ie+IB6KlCch9l7Vati+jBN0zflZxPtcIj2jYFaTT034sYbeS7S1p
8FCvlsSgkk9mjj6tujSojLLExaF6jMuOUe8dga0plnZhDdQiyvSbsIVVlWk23zYyPNDILu3vbNIW
hVdyGoxDfH6+v3+5Pp+zZJctcbJkanhHnTCo6y7uzcrwS7wyY0GQZOcXn/x5YXxoE9yRrTMsQdGu
DU/sZAQUJEb3Z/dNX+5IuCu6aPw+VLGuV+mlc316bv+iWIcNpz8HQ2iAWaqSJLh1Qnpc4ZFrYmHQ
DdOm8If9Jl8CCfQ6qEQFHwXrOlPsZhG9jeYY2kiUEEaclJe7Yw4595anPaWBywCYgx+VoslfivFB
wNtiBx63kTGE1+rKaWDv6MxwQOuEzec7cQ6YZnCjKEdew4TfLfNsTFfVRJ5v+21hh3sD6agdmDVg
Dcy+NNfvV9uMMJ0VL8S8AGelvZZUKM6lGIb2NbJGKDhnXDwdlhmJG+WRUy2diAWBadbNlkhi56/u
IBoBb4FOV5D/m5yn8z81ugNBE12i+25plOKcX+1rjJqFqS1eBIr0wC0YBdY+XRE32Q58rID5oky8
iQsjWWDl0UdYGRHaLxbv2O1HhidwBbjtH+Dl5IVq1wCdOFYNxOVWN1oPjJCey7ihIDrIjxPbbnBp
HLdeyZsGLaERu6WS0kU/jczQQ1/TsDhqzGmSbNfRq2+I67ivN00j+6rZBScbtnFUFcxUls9rHr2a
/4ByGupRSHlDvwHLg5md8eoUAhstMmkcMxU6F6S+38bFP/gp0cXeKiLy1D6G6Xl4QnbL3zWMWbt6
tXEO8L3XGDWETItLItVmnnCQSel3/RRn9Rj9i20OKuTf/rE57ymoVoRq/MmZ2NAz4dYb+Q6Bfhcz
lqwPB/Lrkx8SUlArnxD//6J8vqwiOFO79cf13+NTh/HYEUVX/VtZULwgwqZH/P10wIDcFCPH8k/A
4OUprM4KiVa7+fI/NKv4jPgPk6vIo6jWiF27XuAG0Qf9EHU7/6WzFY/FUwBkP1pZJ8/ioXk36s8D
ubpC9Px0Blj9T+HfjpOqzbHCp5W7Asqo8F+QaIdvPNZ2JiDgTdqyvENWovcUBBXchzAzPWd/OX9k
HxIr/GaqlMwGlatmMbj/D+u6Z07w71X640M8B/awcciOvmTQV6UxQCa+93LRdosOhY5p1RPUNRDb
LgoEh6ULWSDg3nEYcrWh0VQ/WREQmK2zETHlzZmWFtF5KXa6uqNRYcmoaGts+PVbO/J+sd51uYgM
5PbP7SJDrtnrqYxyIXzqi+8EIbXxnBT7A7xWfMEp53sD0d2TwXq5jmmwfxUSrjcNwL5l1W3eYgC6
Out/tz2lA9D7oAXrJRklwI2tIdb8O2iWczvWHFy5A6LFuyi+dP8u8qhqFhq00u+6QET8nfkoiyRU
Cc7CTNMANghL2WVpLTKGy78kQbRK4Qp1N3eA/uqFFT5VdNYNeuNQtoSh6yr+Fcy7gvUTDYQ0jFKw
wS75nFpPRb4UVWsJ224N8NCjW6rXd+ybD/miu6cqOox+HyNqe6E9gwivDydwl1ZHrZVgx5b5BHoP
361AbSi2UyOwp97Ygx8ZaOgtxJSlry2MEWfcITfv82zzhFHQXROoi6+v+ORLZSwNH0bI6Fo0wVqH
zovqhrdbc3I1B/kxpM281gdBOMqOOr6tgbhpisruBl/37X1/Wxqk+aLHac8x8ROb0ADZV7h4d+FC
wdHl5yoBgHl2204elU9QvpQuivAy4SMKCsMFcFjWZxJBamXWGjMCVSCAqHHIZyUogBjbEqpde+IG
8OO9hU7ClcgweFPZExc/OGFRNzv2FyRDPiKQ1IuZh4QkihjAE2Btz8HK6UDs1Rm+urr8Ddzkb26P
jhCQYwvbTx7RmRSiz2sQ5IWobvT5BGRDc1wTrMcYSkGZ4wieTeetEbhdC0tkGvtxV/+P+bDA9AWI
LJO3KOtm0VCuUogHLJ3rUccspNCVveJbPR6VTw2uQY9V26RmD9qs5tGm1Nh/Rpt6Au9VrGCwGAVt
5uoiwcCVAE65tdJCXKSxWL7wjDdWiwZfLj1PZSjOX/pqY8Zl+ycUTPqN1qU59HsVyipfdxmjQtww
klmyT0IC1jIIPj5A8QzbQ+t+1fKiLFb7uZe0sDerMxjPn+uN5f24z7ZMDV86AttbPh2Y3IGh0brw
BO1Htwl5fd0fS9IPlcxugWDj78CALlLh+wu0QovRP/3L1kICpqR5on0Nq0as5GWFxpwlkljvJXfc
jkBSM5t1x/Sa8cOZASqvueHonNSF3PwKfnyiaPak39v83t+R0iIjK7kKHHR5IiTg9VLHi1ezpC1K
G6RMP/pn/R8FHpemhn0fXuJ1MiPovgxMnNLMSqfp/1cOpe8Uyf7B9p/TnC3oaWRtLdhaozGKAmPq
5ETnisDH/Jey9h/P3idIfl/LdcjXZjavMjHkQ4OPBBGlgPIAUX946+GRwYRg+8lAzCKW+mYKzJqa
5D/sKSE+BSlW4yeIP5DQMl9iB4KmOGmrxE4qx/YFEi2Il2t4SD+12JwYR3o4AUyxXTJ43UgayfqX
7Ry9DtThRiKVRLe4qm6bRWZ5sUBFTJagFvNon7yXNceKVkPLMh2aNt9TwZJZ1S9CGcQGgpYVuez4
dnjysmGo6YABiaW90FwfUU7nsFlkwsINwVlzHlGynv+J1DUWzMc9QJZmZEievpnoLh6ro5rjS4wb
QvrlKIJNS4itMjxWRCDQZ09fLPfMjV1Fi1NEOmX9CGz5kAGYC6UguTLYDV1MuJucx7ikpOXhE4s0
A/ewFP2b3/jpSX3m8W8yJRNbRjy+3U66Ggg/z97y0DWzGgjp/oOgxg9UwT43remFme3GrK1bYuCy
Ks7VkLhUpCWX04KmV0CAMQfumOCyos+6dF8bLm6vZsI9qzO7Ba6RYwO87d/LzhYGAtkuNq1/c/Q5
hvY+QfWyFiRTw5upwfqVQ+E9t5RpKKfSWvNSVZLRQVN/VEcrVynimsvjwTIICGIu4US1nJaqdz66
EeCQ2ozpn4/Ymgpvya/6QZzAdg4Pz1/RNeBfP2+p0rgfGtLu3jTEsYZHumxFcsoTJDKrS8lf0522
BdvndNSSZ2m91m0GTxqGfNuxyfsN9CGHGyKuO0//ZPjEUGIGaR7pjfYydq07cuANZ5D84RBqS27F
YCzbpQ1qjCk2MgbET3xkCaMzoLWcpXCSf4st47qAn3N3EIQl1FvAMzn3ynmTvbWgUmI8uBr24YuX
wOzxz+8yEW/alrQGtdiuL+PuF0fdsDgjTqpBCV4sGDLGY0SgDs2MszPsFtjOsdXCKsb65ZQDxBrd
5Igq+Imd600AFLooK99HAplKrHRG4+s0RT4x0IvWt6AcfzK3HdRuLb9KVRULuOHCUlpMnE7cP4pu
cF1sIyKJ8vPY394uDnEod++pl0qXACPKx4jwdPpTigFEBdcVj5ON4kuuGYyHPeKusLRUiiYNkqQu
e6Yf1qmgAs0vCk0bCPkIE2XUbXvXnnHFnPONyqBF3/GE+Yn8iS4cLfXuta4Fzk5NO5/sXEN6tAjG
AsYuCMHQHuMCeyM5eXVm7tuyteHmE7Ko+8a8oX1TyT4U+9nI1mVwOIAAy53BPrM8YY7+RRwnNAR+
cslMO37Dhk/X8U/sv/9ns0pawVUTzrBS8JSG6Q/gLWjYJPajG7vCof9QrOYrgCVyX7ppRcOwPoC6
Y+z4LQv+Lk/oypewbUs1MTWSFznMRQHp+2t1qmkddTGYW429Z+F1WUEnAv+eBcwogVHj9yhmQ/YB
MFBljkwZPTj10B4EMYYNvLLiSruK7CMrcXS9BBE1P4zrnFLZfdrjTu/SwM8Yz76Tq3HC9Ade83z/
S+gnSewpCBIGYPupwHStBpxzWGMjulKje+QgvxCv+549sUoYMhqwXuuCQXiaLPG/4cYiFnKpg7sn
BxmiFu85Yk+oIyb664/JaK6gSdxbIaof3x+r1skmQhDfL16i7lxSISuJoVnkIyirUjdOD0jjgbox
0wJmTnY+FUm6pV4Q7adocMmn2iD2yxspyX+XWo8+aUPOjlXkIMrV6gk4WtLkR4HElx6giYwZPeN1
ZaRsakBZkCO0DyxTI2dzADkK45ckKqBoRDktOAGNdmDIYyPUtBzYVexT7nQ51B5DHrHg3wfjBdeA
r8qgVc1URnAzz640Jr8TFDoL9iExYyJVBHgerukeDmcqzuFz2466ZYNvmtOGAeXznewpMb2MypPb
ZLsUoJpn8HXbwfMl9PrHJl+ko8DneBB/29p5gI9YwohMq91xQTGEcCdzQcKfrm+gnhIBfCVWQd75
lNI+ECIQq0UAMF2tkWmhOM60pSHOzMmagCgHmToqH0Oy51RQzz2Im7kSCtpukPz7fRZfNej8tkzv
rezpI3PF/q0mnTKfqZJKLApgXGwK2GKxa/8U/oUDdr5PUF4Z7q01E/2KZDk2zqSBC1jhMqHI1WIH
DOulL/JBxvx3FyCi4aA6m5Z9L9sdBqb4pb/hgtBdIpalA+3nTJVWHrhwpfDrRZwaLXwHiqevtwsE
QNKK+DRfWxy7cUy9oVsvlossCH1wr/8pRhNJDWxSZPTGwQ6fBXruDv3Jrs991OnAN/Nu0sMolpVV
MGLIeaD+NwwMBcZ0azHqhk0DOvPidG4GH2/jzLx+Y1lsJk8QjIE8paIJQPKom457FrUmBIYRYm0k
u2QqR42zB9DvWiW/KmJ1qlmgCZTY/vzfjbqZm/pCeJs8bHfVsm4Ahxhk5+lm9XAgEqNxFBgV6uGQ
LMyKNeMGF0N3AeyXzLHpcKpibdeUkLNCi+Pwb3nIqx+ZBMHPVek2+4i2YB33e1IMA29Pqkc7TG8y
H2FDPWJXu/ede7aCfuU9MdHtjZxs8WiQgUw79mN3HcqrdpcnuF5oYxxIfK9rEp+05PpiAGNMjaAp
2vxhhwsN+gYzNDoCAoI6pK8DrTfjrlkqEy3hc6jIDtX/NFE8wOXM+hbGCkB1CDsm+GZCJS0tkgEG
6K90T7ZnSA3wLdwt2wxlENvOCgoLTmHcYUdxwIAaDvtlcPcKj8m3QqAhbbNjBboLcGnDb5GDl6l2
RuHmKBXFSSI6cQtbEpoqfa/7oK0f2TTiULgFf33reLVJ9n6YMBZ42jwOnlpHbD7E6pTsteESlRVj
tDcz/TMDvA/dFYAA+F588pbkGdlttTsFNhh7bwTwg86taChAE+GnVZWA+t9uuTk7PjJGV1kEoFFp
8bu1rfIzXPtoaVA3ULyvQO5ZfF60PV9bF1t+9CxBcfh+nv+0OalFJ1tf39rvUUDnu2xfloUrKziV
WkFLosc1Ap53rOKYJ/R0b3sBDLFzywtaiKO0+XR6bhU7tLkPOfvhwo+Y+NALdPYCk2jK+UojmTzs
57aFijhlf4sNbS8/lmwPWEMPx4cSpbMc3QXuYgf3Yet3wc0WdXVnosq18gp6RqaokKRdAFdFsrqt
Yi+ou+HTbgH9HiJ0CjLTxr7NSsdvESMTjdLcr9lRiVD2qFjQaudSMGaPvtGEdgz87Ip11pmIYFy4
+zYhDjn9eA2+VWOQtNs+WSddyNdKbYJfJb+mocoaayrF4ardCm/c3sEzjR+Cm+hFCt5hBHVs4diG
9ToV7LHE6NMq5P85U39WBUrIetqrRQFohhQWCzzkLJDqj8cT4ZF2wqZHCq3RyFzE4Y+VyL48AQKr
MlIYTTyFrS2oNbomeF1azR6lezrdXEmrY+llDRsdBDOsYORjXyVkBdRqQVQiujvp28zfK1Tch12L
AMzSMQATPQxwwARQ8R02YGvw0cuq8HJ/eCYzG9SbKluql3SJWwV9nqbBscm4Yi8YbXRfnQ4ArqEB
l2GFUAR56c/GdU2eZXqv6DyCBA0od+kX6aegAJbAsAKcWVr2F+KGfM02ekwQatj1yrPdTV98AgwU
4qkeI7ozxF8nN51aP2JJ0tCZP2iMTN1LIhZKJimONdjCTdZn2+KtXD4e2fiwJ0BOP4vp3kdaGj2o
gMnM+TH36Tt/xb7PAc+G/uhrgkOasCDLs4bTih6Eto8GxuP+o7lRWvlVGSeJTMRbfRdEDjJClCH6
2U8azAiLsBb1e4wqgS5t6WuJ8ODlemxWTHRycgQSisH4yjD/k/fPMQQS4Y971/zCQOOBmJKiOOCK
qhTyt3TFHHQDmBa9NJNvbWMSAADhE4uX6i0fFhAnlAg2T+96MTuR5nHRYu5MzWufNiNVefgRLRo4
D46bpb0yM3KCreBGcSOzrov1wvCj8kqAXnCPPoXo+B+VprSsx180cMgLc/cJEgA/e6Sc4BJy0kIr
MJi0D+kuAhEJD1bvhW23MJXBRx6X+xFd6Qc8NksaJ+Hs8eI0C3HjsWL3N9Ewd/L8U7io8oXeSqoe
ibGa3Vp/wxIIGzqHN2A0G8o6nkwLLi9clQ/HNFJkKCWvdlbjl81urhr0o6h4828BEMECKGdwQ3PF
L/v/9kA/UbT2mnY8yr6LPIuXWReVR3xW0vWMA4t4BoSrlBHWzNwlwAleNH+fTDgm8XzGTOGxxRDW
gCJVe5NMKG/xin3+JT1Nhg7RMNztQBC9qXztwF48E+RNR5DxTjlTLitH0masJhPlYuiEcqR+36bG
Qrx4h8NHNopr4Qf65//ekcBkEPJsapJf3JJA4etTj3i4GVL1cNWjmya0EWrOsyWMyphpCGmHigso
YyOWyIZBWaD4vLeBhO86m59GvPvKRj4DNQF8fARR9qgFl0wEnZ5FhHmsMEjP4oyE2JuQ655F8N/z
bgF8yarrL66SXlN1ufB6NhN6quf11LCfx6VTEz6i8ZIZseX0G2Haclco5tbVEE0ON3uMC2FSEkdE
/DjWZ+nvYnyn2AcsOG9e8cij1CrqtpPqC70DlxIR8DVLnyd92AFtQspW5MXT8Jzx2a8QmWZH8klf
oPcgzn57Nik2aabrGEmgaL5lcrKIYVrXQDhZlD5nWO9qAJf0TqxTfvYYiaw5LpHg/dWiqEfLWvAi
bZSwjxqrh0nmuaqmWMQsPqBmCYY3eIRfnxxWEcBFlpTjcd7b3rRv0DvIm0hLCeuCZNU3XvhVLNyR
5i8PVhpw3bXHuMs10nrgIuzYZeRfx5DBuiE8HOKNear6n3Sm6pP9RX/zdbIKcQHOo+JBI/VoU/Sy
6UD08Gu8PzRjtxgdzy7EfK1qOGoBVNtWOGbzoFwhO9l/KFQJJ7WubUULaNo1d48pFIlqL2Qi7UrB
EB/27uxf2B2UvV9If0jfTEX5ggCB5lxptly1YjVCK4V0lIYwP5NrFLJFHM82PSw5ISJN28B1fgZc
ebg30uAEkSus/uLJ2ng4GxANvzSciISAWqRgdKjnD3tI4TpTfANlKmb/LlGMaRenvfnzh580dhDe
gNNWc2093qly623XcYw/SrKmJDCUGTbi5os957YA0IcIvxk79UahNOd0pEaEC+LAa8WS1NPnxk4Q
twDIoHguMcImxAqboeGdXaI7UZvUrfawP/tzF9EqWc+thdYND4nbqFrW+yKj9IJB9IRhz9GTFaYq
8WMB1K/r379Huv3OCIWI0KyzF3wCoOkEdrrOENwpf5FpcuPx2Dy4rPN1s3+iS9SYsxj0uECWw1oA
u5OGLUCZ60Kv3K9JjOJUxBA0euLLShVsTLsL4pfNrFUmVPxZFd/VexScJECds6srXh2VSPl9nqG7
yyKXVKH/B6tZTiCcIHXd8dSOveUhjUlVBmmM96yxviyoSlDAYEm2//qyiEkqAwZH4zjqZNm5/516
IyY9Lg6Lix3I9vHFNxhoSkBzF+a+M984c19j4eDQ01LXJHRpOnaDCAXAVXY+C5KYPUdJtmUQA/vV
p6gnapAUqbECAeZ9bkncBhntP1X2bLqOcGxOneTsQ+ynmuVum+rPNDoEFn+Slp+4UI68+y8wwMHb
WKZmNthktOtPfVlhUiGm1NJHVUGLv/NGEUCMsy2qfFZ4F3mUXQH+ye4S1jT75nh5stIBXZXeWkt+
f6hpL0Xb3y1IqrcaL2Ma+8KDiC237vApCv97BqaW7uVOAkPmRogVjz3tkB8knEIE+Z9rrb0HBgCI
6UWvwQwYTedDv1M+m/h1WVCfU+yRm5K7Glopt9XRIPzM94so4AyUGR6K9sr6XXcWN/Qrf+pIJ/xL
hi6iADq7x/as4o0YCtPJCz36c2Yq7OeVhJnb6mxANnmPVnQPEbwfWN/fTdJ2PtOtl/rHkp/vl+Vs
wyxnMppk2aJJHCe1syj9MHm4+8ZJoVNZSjf9N7BcSqbbMHJ4NcJN3GqT6SELMnyH2bcx5JvwbTBU
AL9ZKvJEHrqY1zFbdvo4VGOzWQ8toOs/J6YiZqA4ok9q1DrYox3aDsTfK373aDV4ApB1+PaBrFDb
6d6GSqyJ1Q2tI95VQJrFlac/NlwV/33/4Fi+a3e85UPP1ImpKPixM7gfkbfvzjMF0KSVFkv9xrQZ
4Xv8vNelMttU+m8I85eNmKBm6Ea/UtbZKJaG3V9vCRQFfTBlno/I6hMwaw4ctMylfgZQLGmPeBBu
dTW3bxYqC44E2zAyn9W/4f724Dn4vrVnIxyxM8UUYz7XRN/A8ee72Gawin5uY9o3hLvNgkhJyOO8
+Qy8yXi5OJIUwjrxBw185trzkXffczvLSuc2EyNksL8+mY/HLbV49WamDjEJT2aoZsJnWeyzIJed
otEXMrkjadp91OqGJo81bfVTVN8gYvGXEkDqLhz1s/0KzPvPwC+lesGFTWL4hd8UarCMD36Oz7NQ
aaYgJlBoGoNRKvQfTBe9mKHWVlAYDpZr6wA9Ks4y7ZyebueGh9xpYuflQoUBvuJLevvDIckh7ILC
SUOUhX+0nyXg17hRfVhgGg/cWwPw1OulJTeOraeICYWTnir0Xbyrro8PNjFcTaMrV6xTJGodouhi
ZpFSFhn7e6YGIY5hmJMTfB2DJYNj5L6qCz85mGpSqcjmLyIOhU84ZmbG2vRqTpXsNj55GvPPEsx/
dDmIAJCmrHCRXfoUmZ7fBqgEoEYaxEfhAEZThFmJSK+YcDdNNBA4maSHCzYDZOymDHnxKslq/iGn
wT8kG2tinQJMNeveRYePZ+t47F7+HUL0iyvoJxozKiLKdSdkiYA9/4MEFI6LRk6UAQOT+VB7LUGW
EXe1eZ1aA8XuWAyU/prgM1TZe/KyJ0X13GdXKcM+3OX2gVzIBXbFnohylh+reKA4H1gZ7/YuicJT
hSRiQsEaeZFoTSJCfWb1xUtWoz8kuGLXNKDmGtv6jZpGcOabdB9I4/pIDfvXMghDtZB33RdLSGYn
Iv13u5Y98LhkNbD9DxiK1ypvwu+oCNnyY77EmTpKZlYNvB67FrgSm3MvbqN4cZKTO/UIVVTsVBTA
AFaZAd/zQcpMdUn7P5AEI6HUnHrA8SiXTiLv2W9jIXCsIa1zOZXL4cfP/h1HOclnn3G6+45c9yue
S5BRoK1kCWr3FeIItxThc9Xr28wIKm/u0A5sKMK2XVFiHO+kHffvBoLBVtUO6AR2ZhsS78EG2Vqx
e99hq53wEzjC1C22E1RW8DtKExkW8hla3oSBA+zdk+7aj5k5X8VeyADbbkFxM9mqvZVsG1vXrste
6EaD6kjgbWw4ReUunnHMuzI3lm6zBQ4hHsUk9IEZ2fabvkPrdsoJHMx8w+JlAY8cQj42JVIkcYxm
R0hIOKN933kLwM8Dc/lMTp4F1I2FWr3zjscvf7Mpk2eYL/GPKis8Ml7/IBikwdeQdBMHkbqcn06E
uS2W92treBl7Y4jU5dR496AKf6ZgXmR3ExW4glcofZTw3srD7D9aNg2TJf4rdaMq7AVuUu+eGyBh
UZ8zWs6rV+Yd1SoxanI6GbaFTszZvCvF0rfPJXS4D+VjveYOPWzYLXfsySx2CxtAfkvBjKkHYzBE
lul5UxHsajHP+sCsKP+T1z+YSFoRXBcUP/uqPf6V8iQ1LXSg4MZg/7+KrQkzbiJdq1uxg5SZYeGz
07hOW4ff1GFtLHyL0suXAIk01KMhGrmpr8CRLgShBD8UJxvJVdP170SIAf7yWc56aX9vFcasogf3
CvJTcM1c2ZsXN8HlcktOi3t8pSE2KcCxnGjoUED8RzcbP63yT0a6LNB1M0C9fGNLGrJiGRt3Az9Y
mGdBkLMpiRvgJ+iqifiFtDfBn1+TKUd/buXqO2ImIGHUPqKMMGfR4Mf2KVP3+h3LH2gUNC94Ls0w
u5JGxw0kZm/rplED7x6SGIbEAFa+bQlrkiccfxp2yvvTi4B9b13KZ6fPkMaV5mIoY7Zf4IstRIz1
rk9+IsJGHiyU6muv9k5zOAO1G8EQ60SmA1KgymMMN+vBwz6opZOaK1I5L7pfi+9LAHVi0bjIwjfV
dnWZnBuyjzFcOQnfZuV9gwQSOqU+PgPYr5MPh85TgpUI7msUdhrpXEYHabkorfECxESxeul45wQG
l7ehNNuYr/wl4kMZJm4I4NT0MkqyrgQPVWQyC7LstHxLt2HNKYnQ+TrNG0x2mtEmlNjKaTiJWzyq
ADxedSawd7x+wMQ9lG/l9FXn40kevH6lc/36N6BPenhSPm/KqFSq2Q9OOyqC9E1sLgc+oF80m8kX
QX3wvrzrf4nU8eo6w/g1GrLcUm/AqzS8B7KvGKW5+1Xq0+A8xiIlKWDHDu/ux7NVKfzeQIQWyZ0z
/oHkdCOVIaH7z9yfG+z4mArEPHDnaU7q0sZbK7mVo/rm6rDEIW0tqzB9fbCyTwqfk5XrtoegiPGW
vQI6OJyfe9fHMqhnRBhm1oTNd25ZxJuKYsRFBhfy9E1RXddMWPkbab5lL9NGpWcmp0KJmMS+L9SE
yIEbN9M6u+F1fiVLRkydFtfzNa7stiaNQEGemUWuMwLtXorB3uicIrVG+hWnS/p3UMbYhyNfn3M2
7T5ohFKArfMsecn9f4rojsEMtPV0aobDnHMyxlG32OjLILAPkjDjEr2XgHRV1NrPQ7wV90Kc7a6D
3yrar7p20MWYIYCVQhjOLkVgHtbJDYthLeSHXFGp9xu/MeALI6QpfylkkRfCP6e7mnLaVZi/hOHF
8NOLdQIWaAnOPCt1vFn1x6VBO9eAbM3R/K0MMz4CRjLpm0U52MCnuL1nveu3K8+lbJQ0P8GQJj0R
rA7itNleF2/vTWmCbuE1TmcS6m7CaYFezF+jKqpNfUrlVTolavDtorMCCeQSd8uSg7eNVzS1m610
L5f6dCT4tbi7ObczzscJ8qCtlsmGD5HixEFcqpfL+IUfPVBLGerR5LUEFeH9ZxVPc69Wz+nXOrzC
uctmER38hEMUDTC3ldugYG/DCoWZOZ6jWalMHMvRq5ugCePpI81Z6kdgYtTNf2T0DriUNnwqeFpD
CkRYRktbrsq6NTVVuPwGJtmxQDn+C/pDtiEVf8ktGRB8kldObQKn+srxXIcjDSb4lVLJjviJxJEi
mnE8ZCBDuk6fBO4JUt9SmNOAwCPl9H79u6kjOVKKhvIUIa2DSgzEPn6ElAvT27Qo8BoIpYjBivO2
svMgD7QmC9HYBH3LhkM/035jE4Gfu6rsNwXWLL/HQxkoqP3FggRkL6FOq4pa0HGWZ55iTkaBqnB9
Xnax86chSukGs8bWQpGLvnaBdQAK2eNEQGiqhEffTXqbQwIZZ8JTpVaagW3j1ZjHBz2AwLfhkBM6
gRsmX4HprdeH///qC+ZyoDc7H1Cu+UMBkO/znx/vV25ybryjJvK1QZK37mSgDLe0+rxdnOTomMvS
X+DRMYbu+fk3OTJBro3ILNscfJGdhBfao4mH8m6oHiIhluJ02qk/rEss94oBEHo67rAOTxm5jDM6
MuTqcVW2D5JjQENlXtE4nNgj7SPYX18ejyxOAb+vbWxqxhLA6C313FvzkWXcT5m+BiXSci0gt2Td
fVWU9lTT0xPCzkUVY3hkoY6/cjAuyCAxClPJD7cN0xzXDBy6OzGh4+7YAwbTt+FN6qLUb90XhVda
QA0zjDb/11qgL43xHYEQU+E1+zG8sIOC3dGFiXyKXwxVqPvWxBabgm4sdYjSpJmRYN1d9PZjHEZm
Ztb0/beKOHBedltLG/3hHj8OHQHSpVfH+vx49aFgTpfOYyFIChZ3rxoOK0KRCqDz/CjkJLW5gHjh
R1KiKf1vIMcRJqY6ee7y6poNF6WZEzdh6ZazdICgL73U8zhwUrdNkKslxUGbaKVjZIH4Kz0me5QL
ut2m/EB1JKl5tfsMCagpW90fcpMOz7nq9wTJK/DaEPC8SrodR53xVzJpRFZh+4Il/YH89fRX5VOt
taY4NHd5I4R0/dtIC96vpZohFNnqznX7XkEswHY1gwJxEyoSW3H006YDMkVTUkhd3UM9WKP1iH5L
I/9fwOh2mDhgAOgD6ec2IlSPaSLneyIdlwVIfHWVGmQS0Ezu4vuPMnPHmkgo//yWkcCBbMKczU/P
ZrQWbXqfd8v7JTRzunKSKmBssslwAXHrH6aBcju4FdU4fiJ7kbX9zT+tJARaSSadUVhTNwe+HmXg
//t9hSr41wS6xe4jMnE6xCTsN9mHB6uwDawnhipIUEjEYBVvm+Ug1A12jMtbX0897+8JW4LSo6UB
mjh5lxRZ7PElfJOweneGlHvoT6N+al9KgaNeNkhGOy1Jt8cI8WhKF20bHEYdLALHpL8dsRWa0O0z
mPJO30qsJENjOebeAXvTkLHeAVrfBsGRzSEupqGP4/oM4K/aRAKzi9flq8JX6ilZptdN3STLwg90
OVajeUYcXJufElFjX2v2MFTn7TYeG9OgXVy5vf0fh7R2ohyuteCBHZXU9Tq1oQxd6B8bfEzdTcBV
km79haOwadKktXaRNpbwZ0WKKhwd2HA1m0lrJfiQrTqbIXmb6Uxe7dVFXU1kov8PWG7VuCYm88uf
VPIAb4b//Kq28g+SPyRBtvaydLxs0clPf80fOXmz9qWyflh4SRp47RabnWlebPwX1b8gfLuhgphZ
CDchoZIfv/InclEQevFe5s4LJEQCPxFu7+YsgKdrgqAMdKDfT6GzEBUOR2UqsOS+44w42OX6dAYS
nXtk+a3nMfflQQyQIr69cZg9XI93OFxIruw29uZYzvNtp/xCRBLprBHlQe+BMTqx8SuWWTQwAxjd
sHPx1UeAUSjSEC0a/v9AyWCRpWpJUe5cDlh7kpnpyjlBukXilMU1MXL/SeaHbDqPipzqZO+VR4Ho
AYZulGKy3kYFk3cD5/TKYMeYZErwn3D0QUn0xvj2+2OUbNTBF595qqVOpAkrbxmnVnw5U75rt+LV
N9yoR+D6aaEpfTiOPKtB362J/cyx0u2sz8aeRAQB1Qa5lOStfUMOjknq9onkWRme9Yhafnai6D71
9s4ZAkFMQogZcRGIFQrWEjdvZ4p7wdfXEkF0COv4SoWc9KkslDmL0n/NgtnB/STyv2c6ru5KjbLI
zfiIX0bCR8OOeDWPCRmV2flbIVhGYh5AotBF03AWpvewV6a7o4dX6jjscCU2rh/M0Uw84WASD/vN
nZNkDjUUEOTXmurcbKhwcgnkO7WTtvZEAUj0QYpeFAxnPPlQgxFq/1YOsqxr7EuE7x/Eo5LYBPTp
TrONgGUbUmQ5TMWPPPBM7iGdXd5erCo8YKVB9dPb90Wwci4XKGtI9BwjSJIhAGllunoUyKIsSI+5
sY8i4YJeLmk6S3zGXIKeptmF4wMiIK6BpjIvMA2Utc/CMwNtsVETlHq1pOVU7f7OjzbABzCqCHob
WFTCjrOCJMkdAQ3rJOo3+8UHqOaUm/KuC1Ycre7fEKLdHI9tr478GvYpTFdc1gGX8xI9pcy3iMVj
sD8g64/XetqxLiHY29QXPQl+E5M5++L562lKN5qj0hB34iAwbNXJfMKQjP2IZqlWQuwDqyaR4fjp
Ds+OvVF2vsDTe9n6+QA26SMKRzbU8yQrnbmmeue7Y56KU4szsr5bDKpDNytjlO1OGVVLRp/SpSD5
/P5StVUVa1DUruL8No8FA+Sm6rUhyU+48Nise+xzS24lMsah7oFFm7CpRCpFmMF7M7vjzifrVh41
qNGIEqNWu+Ih30DFXYAs/ztzWlj7goZs7Px2ZbmJUlx6H1g45El/0aIX45Qte8uyR7xtsCYXVMgv
TU24zNW4pB20/PuIlmGSXwPhB2kgNR5xA2P/bV8GnLJVtWf3bQKsp+IWZKfi/aVx8IBkNV7dawqu
kmK8kqitUeK6Ld5QwYzdVxdB0IxAodvX7kdKIFHBDrYDXg1Kqu4Qjdb7OQbof2+kvnR8ac4KWfiv
8KvNKE69a6a0I6r1fsWY0MXr0+oRxKZTlm+3Hpig51vQyZ7E1ICX8aex9efTftosB4RsEJDB/ifD
FNhOelohwqaWedNXMq0N1yPJCkecCVYKrYx7FPXmQNrTYNZH5z5XMhE2CbQb/u3VY4KFdjnEVd/T
EfisuYtWIU4ldqlXJgouW8UT1B/1ZKya5vuilitmS+pKgT9uz4Jsvm5P/wAMcSRJhE58B09Tlo4u
eoaiDTAk6zw7pdijvoLQXwjfa8vEFjg/dBMiYT7hElDg1b0tRi/B94oLUf7VqOYIYmHYNLuX4FpY
W4bzjADqb2GqUUtAinwcZAynYd/A36wWmGzIX6yiq7vfQSkMW4+Ik1OCDUV16kbwoc/jGktE/kLX
yrGdySSecJK9GHCvN8E2+H4EzNQ8jwQPe60Mx3kDJiks5cEJDyfoc00eseN6QgwNgMNglBgjeVMH
PDT6xpmgcaCh9zptX3VNlxuo4DNhdT4fFG28neH7U9ptyra3SZ0B8PwDLZM2kxQLzfmVYq/GqsJD
IdFmpeoCdpSwKWpN1mkZsd9iHeGgel0ruOjACJNiLtP4M4e+gySXTQS+ThSEXINtujyrg9iS81US
7F2vIFLPa5xPuTxAGE+AAOAd7KgRYTYeIKDyB+vKNO56nexlFO9KY3+iBPRwYmj3vmhd/MR/yEqq
lptabtajpjv3Kxvg95s7fYUqEkvIQkF+mkinsvWMsCQv4MQVJ2RQAuLTGYMx+rWlY/fjiOx4bdTH
gS137dXs6IdN9+6AFN7HAGTPYX7KTIr1GE/pb46d4msU8YeIWgvSxQfdfv/08NPIwuVD8vTaN7QI
ztXiAeVrao5YH27xzJyceIoYF9dh1ORutTTxZUrbSwpMhit6rPWiS0UsxC1eWA97Efq49edyixz4
EmLw0Fg5WMhWRw+TZl+xZCbXLfsELeuJaJ3fBqU/S6ViUXo5HbO6QMtqM0JNN7SUdfCKm8LF+dcj
W1s7K4pdhUblaoUzR7YpkV1eeoCRMLqYfyQlvCf6IulDZLbogUAH7ZrYBYAbVaiTgoDj251tZfZn
L3SZLtqRcq22eqz+Xp3HO+Pu3m8vR1RP5JsqNf35yBR2Jbdv7nmPMgdNODsPvAgzgEDNsuAMRfEg
IGOQHkaawzAQKH+nxQiHGvbHc+Am4SxsE6NzXXrVI2zu9qk+CCtcL0s7UpdVYX83wQ4HuaFPcBqx
M6ogWncsA4XCFoMfOZTP8XQOj72nxwK3IbF5guLayHgjSIM1yZgVWYjnpgjwD7kHXjWFs5uFqR1V
sIuJvuA3gLDdxklYy0rtE2VfcUmjDLBfcnbyWLHBTvED4+RsKsRInjGI3EnMsk8WyUG0v98CKR2W
CDo+yy4xsmY7YGRKVfmWWG697HLcH/2Xwf6zzoF1uags38EH+GOQSAFNTtJI8tPAg9deyzmWywDV
5JXh243i4lImwkYV+spkXj6jzr1dnnw7RYnsYIlejTykwZnZG/OntQA8BhaddyXCczDupFaoQVMT
H0+mRrG+1JI383g5cwZ0rERQQbZLepMhphejUV3agxVH6f23iPIZ86PPfVlf/q7ZXf17hkJDC7ci
bUaDFPM+LHf/N9fqZfckSHofmMKWZVoY85tJnH9uGkADVak8Ob8eYxvOTexGP8Z2T5d4V+ssACZX
cS4rQWF/+IIvk18d3KPZliqc7nUp7J9OlZEFvQn8O+OfpILz7w0R3YsppY83SO0FHeLEYwXldpVo
Y6BCjEMFII2xYjSYO43/UaXp8cxXuRxcWBjN7A7f0TLCN+FEJvh58/2hd/5J6zbqvSC/NwCrL3kz
kY/w+lhHXvN+7TTDC2U/P78rzWh5rCcBQFPDpt15Pi8XWrr24DEQHVz//uTqZi9MoYzo/zOQaoBL
V0baE4ACSmD7fdDsjBlXaSBdS/8bgp9DY54wG9t1dIYbJz98DyJ2ANQ3IR29dbQS3NZF9dyh3i1B
ju56qMg13kMjY6ZUosmxv8CClHKsUfpnUd4aCAwS1g0jNiKZgiyRHg7ODrEmUlUc1/0HE0No87Xk
KYdIjuMOtQl9kBOJAV2JLVnmuYMSYgsuAslWxKIDyJ30J/BacmV9ag+OcHPgFTzzjiwCcC+Pi891
BnBH0JtgGdZaJ+Og1De1xLL51awobRkHc0v4AQN/ZLlR+ynCwSph5IkgdIZa1ct+fcFBriuUVxR0
ZIDYPTUZ91BQn7vSSP4WF7SQCpgZ834AkMibMcHrI4GajIgzKY4LOffJkNHzUbpi7G0ChtxZWBHi
u2l231fa9Y2BtaHQmS//8BHr9Vq1Jrg9erZ6CRSNKjo/2skSvXDa9EY5/mw4ljEGMdE3xuCRnyIc
6RcatdNQggwl0ENp5l8yrSxLuepMWdweLnGKGGzKeHj60OYhajO8ILU3CTsVXd5fJNYBmIIsKwO+
X3kz+WzSWUSkygASMJ6jGwKTnYBSuqD9663n/hrKSPVcdntuhvhma13YXRAxxqzF1HKHo0Sk8dfO
Z5tEhnKVSIavg39d0aL47XB4h7NGFiZ3lxS6kuZoJegEfnmPo2Mtuj/1lk9bW45LaJ29qKRxgWh4
4IGwKgOyBi5+1U5JxSXSNbih4Urx6g75xm8s4JaAyDK7WhJhxDPz+p7eewEtEfutfQNvZuNS3sMc
bARBs7Kx3wxW1oWHRSkZoaC4FicZDwaEqy/q32vE/z2fMXs1UZhPs9Ee8Mldfrh9+bW7AFOif12d
Ah9540zb4bsUFRyGpbtxpxdI8rtwcqjeqiPibY9XLdb8rDeAekoQoP1rdxsvGe9EnwMbXVN/MkXK
JfpDUbwso20CXIKMrUvYaq4jk4bMWOvEixaHD1DEwtbilFdUDVYzNR/XCRmamw19zNGQdh30WIx/
mFWGuo4j4VdSu9XDTp28ZYrRWynmsEm/Rlg4Y4Qrp/EkbI+hnYmxtZeiK+KoUBptbXAHCOz5jnmj
nu4keubR/gh6JoNbTCoIg88YHq7t3HB0EEXZYZiUtx+PcdAPyInVkPOos0KskJjO097fHsiYP8em
Jes5Sx8Qo3nM4xlqMMJN5+pmzJPFHj6U6aM0LFiJBsdVfN9T1whqiIDppCnuRyDuLawV28xhYeqy
s7Q+lQOJYFt1KIpUaL8FocKUQd43jIx0AWxpRbBx2ywjJlzdRD5cpiqX5V80fa1VmXCWmB+TWjXX
ZiGGEsHkAjLpuCO5A12uq5kFHH8eM8reluPFbYL1CeOh6lusN5CB2gCHjS/aOtbWHcgTy1MxKNr1
4QCEFCJfWCxNs2rbckh8fz1jz5KaDsD2he2kQXPjRMCipn/Y10Yjm9Ye+S6e3RpkNPdXeMZLQ44y
7rrTrAgtT3nXM2jcFW66mM2FFYPs9kWf1glUnBSqPr9Ct6HkHwIBRcvd2NF7IBUeeiJYUViEm5i1
lKJ9Yqc9C1ghSzvRYsO9XjuHytt/E1acAurUZFA5d6g3np9x1nRBM/xNsy0DN3VT8qY2HfAtEAvY
+lHYsO8xIfMI5HZqVx6plrRFHmO8tHkszzAfHOxBgwF/PrvE11m7UJVT7vwZ49ekS9JIsXYfgizu
b8GVxv0OXC1gvytcD40dSh2+1q+/oNtos4BTWGFzUumDWyntcvsucW+1ZNmxstExk2rSOKaP4G3F
sytQp6+HOVY5Eux9mDvRwIqsI3Kj9Z6IwGbv1HCTLQRSaIG8Izez+1ADw4e+KYiiKigWck4A4jbi
xYLxjKibhSs9IiY4EmJYBNgmwZZ/7dnyFpIotmS5697e+GQWPP80LAglB8gAEuY1oSUPyATzHIbE
ZZBK/4XT60AFVFOgyLLgd8D3XdaQ1Bm9GEYnHdaCugL6XVc6VJ+xxt7838Mp2QjrzEvF8bwTp8jl
90/KfoE4GPzcWe1RZ8ZwV9V3+9j1VDtt+YYh7L0LkT7JoOs8ujn/YTbtCXVfjLyh4I+HzQeVmU0Y
c2NQSn9ytfaXNDRXH/TZWX07XQ01KG/FRjo8Ee2He0N3AZQsOSrUCQTkfhHDogvOEInyHz45h8hz
uIByxrYq9D12Xgjs5pSQaTHqsZtUlOA1oP4H7v5oj5bI6bFVNKz26MjhwkyraTgUjk3JtX6AiHvT
Ju/qi/h8GKObKUwRi8ZYf9b3zV20UA5D8k1bWOmKG7xBh3I7aLVZJ+yCbtRvam5TGe2+EDKDrcqr
+JMPscGNlJoksAw8VrsVlmXkw1iycJmxr73tgSpjSeP5K/XFWIC4yKkGYtZzjLDzd7Ocr65pkMWr
vGdMvxSEyVhcHku4vflx8+iH8Ov99jlooASKpTEJUmNa/XHwbXArAafkStU19va1Wje5QEDtIQw6
sLgwx22dFraP0Riz4NwbLUEhEqdfXqQbzrq9h2QPlejWpPLImRe0QkP3lQJFxS745c8SRY+kXQcv
5q3OrjsxL3tUp5gCtRMILfnfcgu0gqre0AbSu0pFad/JbHy/Wn+DICa8w+bGcSVvV/vFYDLGa9Dj
Uf/TljbyRsfcDOrVoXy5cc0YxuwCK/1JoMlfMwgBL2uZvJeSTrbVnOQjhAoGPQRj8w8flkk6sgrF
dSKAykTI2mqOO0EgvYPh2L5Uf4aH2PA4EVKl4lWZCY0JSD0eNA9hcl0A+zMtTa66Xk4r7aPeZY1J
75/IpGI8ySIhDBXlBvDLxc3/p3d7lYKx3XGs/jTSU//z9OTyGUMUpBf9/1iV0luBY4fTVlxT6JKl
aB4e8F7+Lo36J0edQvkfIEGrGJfofTvbUNt0XJkejjpEmOHH+EO2CzudLOzhvzYlS7D332ox4w+z
XAsjRMTfagKA0lUz1RwVOnV/c2wWrhJkmO2oUr404WOPBedL9d/f15SoRI3rtz5n5i+L8p4P7R4F
1cGiHV4GEc0RAJ+dsJyjUM4Ql8NOp5VMTi9ymso5X8vpZajj292FKe/g7Z3SU9EvLBhUB6Z6pPHH
EHQ146S3kM9iOHbHfdmsx/JNos9ztRK+SaLkV90/ttmM1xtdUqT3qccV7rFgBWihisaZMu27sx3x
RcFyR/pyZGpwwupyrBV5WBzFwom2fkc0F5kYLZMGa4jwfaF78AA6P0aqmobmdNqaR6dugHFFOxpd
VBINjbU2anGD1zQ/HLIC/JzcmlPcXqhsIqyeKQCX3v0BJpWhQfF0yZ2vPf5Egmji82IOncdC6MgY
1XaMlVuPbyA3CXofAygVR+2V9RKCK3aYOTb/+wQG13MUPTS8H/wPNVFDFm2u4UQ09qvUVZa/ipsW
aMlJEO9eDzbdO345pP6ywgpDb41PjR/zvqWZeuECl9Xd/Xs7w62t7ad3RJvFN0zNoeeSSqCdd0ob
E1x0qYgUTHVevymr9z0Lhy+IU+T9s9U3w2fqntKvonG3MxyLesFVj5YDmcgTgprsRsWEurDJQhWc
HsIVP90knYRAf6tvYQIq8CMVz4pRn3gyVIpUE2d1XFzUHhBFId6QlaX/JxSJexrmNoHFKEpLdjrW
2gCiqCdBk34E8Yt+2jSmkkqjIg8Qj66ZXik/3wRFQg291LHBZwbD3kdz2L5XQxo3w6FD5s8myCSD
eNrZxv1OFQZB4yyYCKC+f7KrbK2rzGVIzTzMwQJTLjNOlr2hqWVyOyCSN30hWBQdOsaJWbY/QMZz
4EAglSUJs7r8qBlVyc/jkLy9YDX88XKF4ECKorEea/VN2N3b2PYz7hkvZTUUoJJ0aUYqLP0Un6Pa
MMbZa+rbt5JYtTL/rI3HlbDhKnSwwf+IegEnw0aSp2rtsSin/QkYgcWy/HAkQpKLnSmVWgDc06hm
nqPqvDTNPGVD2df1mU5PATXsUbXDhTAX6tEcoRmx/rzbFaLtNyH4UZ1CrJDsK6kYQQLNx4kNVx0L
kvBA5rjHTI+Nr4StgyT4VqOR46Nf18YjJckkBylwpt20cEj/oATme+bnFdPqb+zPWAb/+4IwTsKW
rmy+joMZT+EsJarAklLd/E1ixwOy1JFL47JsRi9wLY6cTy2bJrCQSLES5cCbendrpQPoPhB6kwNN
+HelpoaG5ZIhvLlvBFAKG5dRKIApQXLIaeWQgal5QXjoXNwGhj4HAEhJe1FUPcISoLQdckeEtPvX
Ta7Ce2mv8n7w+bf1Ae9UU1xZY+xoyJJa7z1iEobg0bHw8tttyABQKaXdcDJh8jKFv2Em2ey4c62p
ocvuPTWb9dAz6CMiSpM/8/pNtHHZeifKERPg+IAbxFbxrRDupcwGG8x4RZHYBRp4DgQmlEVsQXCM
Tt3o0PGnQ8JbsnTRB4td7k/Q3KCsV0pnbZtLRT1AXOWxNiKhrUEAEUdeZaPCOoZACuz2xHAvL4N7
1SFVh0YT+0JT9lR9mUJgl2ImsyjyVOLKYY4kiiuNAXomRFP0Rnm+PJ7EF9WPxT90kyJRp1+jGJCS
Hdiivygkr9s51rWKSpKiLYMRRMo1BRhjqtvRHHwtPskGTBgRFsNvGbqoHf/K2KPyJ9H6Y8Gw6k/0
M7WUU3qqUOfQ8+v5XTFRrthAf+uZ4zoHZkBTX2V9aqboyWF35WIQvBuHFs3s/jRH8JaMExhQDCll
SEv3PBufEUZVVJqdkubdmOqJN3HBe3ekSYemjev+lI/7FO7Yi4Ew3TD3ZLYE5+Ufluvag0UsNyq7
f6skYGoJfpRxzxSYybUhwbgqnQ3j3+qodgl85i5xdsEw3xBpP1nok/AEhPZ3M8WxqWnBPj55s20G
p5FMmw4AJBH2gJ/Sr0EG1dCQgttL5IGgcSYNqKLou+Qb8d8A0GVghfBrdNiji8YdxSFE93q0cryQ
oUGttBFeLNoDCNsmB3UPZ0CFJoNE+PkIKK1cm616qTORH9DziF0VuI0V5bJi3Zbqab5lhsmBI519
LijboNwm9QLD3XWA0OMiwhFJsazSkbP99+r8dIdCZvYeVc75EMGWaXVU1w5GPnHfFmb7eP0Y66Bv
RVuF/5fFQdfIF7daW66Ggs4inBNsTYWrqRpnmvjv17GsZ03krDCKUsX0O73UkEe9BL9FzMkEiGSu
vJ1DOtcaSeOJkHtD5P9YUsxrIholoula94hDZWr/Vy6UISb8pwUQuDrWAhNmRRMsltcOvnnZOGJG
IMmBThQmCyZtCs8qLlkhcZm6KpVOI9bZ5aHQf+XhN4x6YeIc+9veeO9THHHSIHh3e/9GShGl2ggQ
WgHdPu63F/vV/noPpMgxy7N31ZzNDo7q33rcIqlfZggiebdtlkzWk4u9FvmGV6q7fVaZfmoslzAg
/t5nCF8FGwKu8jkOCw4o295dDJ3Lkr7Oz9D35FLJHp2DQd7hOb80Tk/Nj0rbd2wkvWakbsStWbeQ
0BIZ3hIlQ7daEfKjl0xeWW0TP5IUaCDWsdQ1qVlVuZ1jIzNQ7eLFtpJpCyO+a9uLtZ2bIXp0yQs7
UTQMrnc5YqP0Q9i0OpdTpafXycuCwUH6xYeI/u3RHBwS6UoB0bGAXQcZBoMSTUug03/JDZgZgUh7
YkVJQskCeQW5/GhRqxntRlHqvgdB5pLsjWveqe86VSqkBZ3EYz/5WASb1u73oOExsRrhKONjjdgm
L2688MqmQ3jR2KVKy8P5qQd3ixX6m4jwMCSFqcNFrNBiV6tDruO9klc2gLKxFyeuwKmCF0llpv9q
JHLXBb+CDu3YCUGtqe6Oip8B8kqFOf17lIQ8Klynkg4Lk5cERfoN38cQ/h2+9Lru/jPkLeybCp8C
8yJIVqpl1sKBFCHxe+crs+tYRrV4CFMtbnmhMnxF3dRM2wIMTdL/RjKUF3rWg2MUhojTRzaKYtGq
KsBl+Lw9UWcsNXwacnpPD67GTRwHpikm+P45cVK0OW+QaLqnk3TaZfce0i9xXBbPyzFxMKhUljRf
KoQpUhUwfOiN4wBxsJPm5GRsJkG1uHmHzRRfu5Qf/eaFOI5eCm3wHbpq3L6tNdFpYBbh9yM3nvyk
a86U/3TyR3z2wE0jgj8Xv5lb+IMPkVQxyUe2HvykQ7T/0khTeiWdc0NiV2ohVTWBtGMG10eAwRbK
Ug/sl1eLz/d05ZOUshgXgXgDo1dPYpYgCgzd89M8vVKW7+0q2o86W1wTbVDlQCMXleKRsL7s8ErW
5ZRDtfcN2JIOMDTneAhup0l6XEBXJq53D/K+jhlj8lc+rszSjhgHcU1t8/IQ2DGv4rVVryXvNIBS
wLVH5xI5Q2hes2JoRQF6RsLUMUl1C1nWpCw3ffyppW0HSHLjLfY/0nVUznkdafZi25J57go3FxIn
9dslqTuGsPDn8UHWcSmHNq02Vy2KGgMCT73g0bdZDmfspVCEbncrA3jGAr5aSVXgK2zOeeF84ytR
DzDjWxuggd9UeFU3OVz54uj+7g+cs9SYcQHx9xNo8U5xPb3mgHeAey6m7SsXuKzDLfFTiFXYKkQB
Q3+jRagAqOmAlix5FUgWV/9C5edLCUOCL2pCK4+1lR1uO0qDXPhG+c2k/od1spefMqGc2sOu0ZKw
qp+2PlweBvb1oUPoZjVA9grP9DhDm+kMzeQcPPCpXsvBegnq1hFPNdhGo8N8GwBW0F6NSB+XQn6a
R9OjLgfj2C5FxRWkXXymUnp+JzrMzCeejEm4sM1epaftziRRTEbnSoi4LDx6GonTq+ccdbrm3HiS
IC0ScM65B+usckRe+z2z9FShAoc8YxOyd9Y1C0NkXlZue4d6+UX7h55VNcHywF8K8T5fvDY9HBIO
jx0wRhJ9NO3OZCBHcMCYAHzf2WMfTYVnlsUBy6KLqSn0jFYB2jamkRZnY7lCukwkQQPBQnBFQmnk
KXLBOClWOuQDPmmBactJu2mX5ITRhK1TXE0YJeRxDwKwZ9THSP0GsnH8MgbGEfolNt7w5sRcBIuf
xcvgYyxfvbkmFoiRPVtDDRhYiRWOBzqQSSob3TyYEnR8bH50tJFt7w5BxDncIiOWyvox1CAJBAK9
KkkKsRdzFv9P4TJy5u22F3Po9QXfsWhrWNQvijkitWOAmeVo60v6juvAXwT2g7ifwsL42gdE2Lh6
0uFzvFtzIabf0/b0iVp9ByKUgjwln/yst50UpdHZYp2rmtS+uCjZL7JyhMBD2EmklYVW9ofB26cZ
lip69XvD2bSmt28qWjcpkHHyk0v0T9OvjvLpMrWHPH2tY5qBuiix5DOpvOfOplNyU8DPXu2fJzR4
nFOEAq3aQB+ls32hbT+MVmIqGQskS3J9NV3zkaHMo92+ghisQAj4b4mNgmIGz7VgmNYvo0xDpGRa
8WhAkL3BC5qu7N2QpIIxhjs4Hk1Fi4g4n1Uf7DNfNNM4+as2n6NIGKrk2bS0rlhSWhJ45QWjuWrj
J3329IzFeZdsa1WkHD2JFOpINtqWBDfQtBmaDFvtyaWxo3Ao3ns3J8I/36HsBGmfCfy+ozrd8wIB
3EPC5EqFPdobav1B02v8ZJ9uufxLAtuwfWLfsB5w5V5i35sAprhApLPCESfNwIsEBbaasILztlQN
1xK27gZhXbhH9lu0BzLRdfWK82ph68yp9N7joZSFC4pkKCtOAVBBv/g2DGsKu9zcC5NiGeiu4ntl
DM2gieWBS7zcvq9dBxyadWkdgRwHOfDcAAQagfmd2aGxVITNAfKfEM0NGdzheVniSuutKZMHE/VB
oznWAE1aOwY+O2tKMIwXJAZdje7bBtkOCrqYKS144RmKrK5j/XF7YXaweB7N2pHDovWQWQW2FuQz
bMLGBrl46VCOFc8u9RtwPi28BlevdMJkd/HpuoQ0YlvKu2Ig+EoA+je5mSG7BSGLlWRDOaPNxYHq
PsZYintTLq9jDu61nwxWedTrhEsSqp4KiUp6p3Tn2xhn952tFIkkr9wXgCkgBgDQ7yVySuH+6Em5
JIxs1LDLlNW7je7DxzCANj+w1ejedvntU4LZaWxU/sDjbNfQdSAaODzydkft3KdeoNrds9yBrvCO
Ol988SIw3LoOiZDgZG665ryz6Wp4/aotSnBxISiz+go0BIBRjdcArJDdQbK/Y2sqdRh5KYGh0je+
FOgAAWbGGaCFLuzZ36sjqj/nJVdW2P7B+Eks9HHmkDisDzkIX1ExbvPgJAsccQhlvltVMiFNEO0B
JvUNxogl+VzYGK6OrGsPrfpB6C0ZBwNznj2WyXA89PZoWC9qffuec6iAMm3eBNO4f3sIbuW0turm
IArt6kgidena3pI4zUxk2MbNKW599kvj1k6waDr/33JDHkmwVso+iky99+a7pSSNc5bhMewl4z+a
n4CAvZFhzqJ2cKiVjZ1BxgfLRPDxK8FZCfphz9vErXzia8d8bZ2pAHnZqLv9LChlSdZUDud+rpkw
3l5gNSoi0KafQGqMBnqPKBvKjC/MxhR50/tpZkOYKuhAMJedUVzVDmXqlccr6GDXhLlrzHQ33Prf
VbVkFuoy5DGcPKfKaBU0650Tamx3m8XPVEChtRqRPGcWTCR+oX6TVpCQFoHYrCGmTdDI67/aCreZ
tQat96aDIhjs1nxJIftuvuDp7SE4L/zinSmzlGM68R7GWOfEVBR8Bfqq+cDuDBr2cQDHFKOViAW0
QCbvoJyFAQ11MGR28taemHYwke8N4YJV6VqSH2tzcmL0OL+T21dgP9YKuQPmT9z2lAJ1Nd6afd2c
4fHIQbh8GvpLfW2DZCo4esFi91kXra3ZirQPvOTbOu/PPn2CxmL5l+Fv7UQS9HFME+VG07ysARlJ
vWNGwpDdc3Sh2l2ltVegT76cdzslrv670+Ga4uw3qtqjzVtMXuAVK4l3PPgBzRLmFJd3saDHCHat
mEtPWeV7+nuM9NDplBQh2UY0qJB89wEimpKKdder+RQXLA4I/DyivwYiR0iFFqumTnnQ5AaLzZFj
CcZX/nqJjEFKWInZZ7lB9WkP1IXG93ZKCUeK7cZ+eToaTBYtrvAOItR+ZcTZOiSfTrmsuTW2FJe7
ArHUFRh3SYVewq1rGK5VQm/UyENnQOGsZo7w8wYenWYnGNqNkVYuMEN0bpn3qPfjMiDLLOIPQsRw
bt+jEOu1T0xBtPIOffxhtI4MXmZhEeaUU+Vi7ISICJODfAlt+gnetm3lVtLEW9pcT5KgLFe8JQRH
yC9Nd/BtwhTjxDarKZgiIUEdN7BCAEm9843VpQEO2UyaSsVmLxB9ODWawugnjcEEEzGKMC6ePZbS
/+7wAwt6uuVc+VurhShoe+Zgb84GWLyTKYgyk+mtl6v9qmPTPXEk7JCNz0zl8kVHwkYbUYJrf+Ax
E2TqzDahySKZp5A8yv5hGjiwjR4HIQtn9YXD3A/xnAlRw9BkfvFAV5MjXfVZZ5kXioDDYLdAEBf1
jpa9X3g5/cZPJ1RLGG3dqmTtCX2pzhKxNu0SPwMxIKJWmQgUq5gsCwYPo1/Z8jXuLp6KQDdF0335
2UoIYsQgOPSxX9frNEG7y3rV/Q8lziu4GT/NCji9+SNnwy7erEFtlzc4ow3xK+kYdpn+c2v+Mtg2
wUgqVzqBhEHaK5gsft1GGzVvN7mZJR7CLGAr9+Iq1L389PgRL8Q/sCP4opJcebqmFBIlZMsGPOH0
bgM6caBUGlWCXaB5EX5i1nkP3/C5qH+KlcLvPnv2Z1YdjNhemw/fVMoY+bXKLlTz+UWSqPAA1Kwg
5vZZCLMueC7V+p1R3HEVv+FYe4CDBxEhjv4gee83T3pZVZOvbBl07NGTJE+bL0HhBWiDDh8OWR4O
MsPvvXevJvV6Wn5ZvkcY+TVS3AIBLiGq1M84xb/Io7hvhN+/cZObUq9Jh789uel5WGnaEbynGuFB
wOoFQRoMwiSiGiV23o+GqyVRZLIhkNIA6K4r0wURbTo8OjESdm52g0C7kGVjTQhag79EseP+T12z
f1dbmhC0EJ/bMgLFPnTT8OzpILEh39aoPREIQXL9LGGVPSpIDF8CXajyHa9hkdMPTmrZWow5JeQh
1jXbeu5pLAUYX1JmoNq6WW7i6KwLBePFd7xrJ8EkyGxw6TpVGRFaBbLEahVAHDQJYC6OAdFhKoxP
4W1paQi6Mcl5dcm11XrXmXQa+JW0JW/49hsC7/yHG/Kb2L+wqbWUW6Zti/OuO3hMxaeCnFiO2bXR
2uR1ns9ij1ZRlexuEeADjx2DWx/uM1logRrhOT5d0tEf191+KAprUNxntd+fyMwOFiL43kmsqqaG
rChki3waTbhB1fbF4z/VdYvg6ZtmDLf7QuSrBSqTaor8NTF1aXM+vvTPVUEt59WT7y57GWpAU91G
+s6H/ym2F01Q1THGBUexs0zTy+edQGoHpEMxDWrzTnIheE3honUckxLME1NH/9/mJ692aDwEmlYq
lYJWeRarUOLwlQ3UUal/5kLChqu58t4lhs9tO+mLpKJy7IAOFcx9nUznFqoZkpwfoHbaetld0cPK
2P9xZMtED4B40iLYB0eczpTDTA5fVG0LFKvyRSo0JW5vqM/UaXLemC4RzCa5H1eFzTcN30eanqgK
RlEKPVyTYWQPtaP+YSxjuqiItC2PJgIt6rkR9SKdLfGHMxLsO80k2MxXTT1qI2UO0y2NOqEAQjml
plG9PSuEwkSfVUxv3W7gY238v4vGi30fs2QCyO7kHoCu3GCcKXzSImvONH4zVzb39+eQkknvrhmC
2VVshaIR/WBo1a3eUD6yiCZLDDNW8g/aURf0yoS8zSqB/Qw+FLK9Wl9ti7kQL61OWtMg36Fp+F9f
o1nWbR77C8e7BxNwvwg7YHXOXSYnukDMT/A2/Q9Bg6kZP+Nypy1msIJa5MFXz0v3AXBVMk7savC5
m9bh0zCc8s05UTvjRI06OEsMGJuNk+sV/ziToitJSIHvnIQklggMKS4N/q9rbYwsWWD5jQw/1AVF
9xgFCj3JGg/aFYFEdI/DFjMHoRxSfr1+2QFCsC8GE6EnEJXJlwjJQtKFRjc4rEMsYbZlOiMaWRbS
Yrf4TjFwxn5UJBwKmBjj6J3SlfbWxhteUY3jAVDnYDMbboWyEjBGnrT3f08VqEZRthBXCCSMgtOy
a8LC0V3Y4bXHPFXLYqJZDP/vLvRS0q1aioTYQqDT3ghxXih8o4WOLSQ7Mkyu6vOIRONT3qhy0E/U
KbZVZPrwAOIMfJmH+0k0x9Q3flEZTqswPbpTObSDKLrGVp8NfKd0Uzn7tQdaPzByPm8Ygc4eEANQ
sFfrC+5T1R+LdZ2dV+EpQFGIjyH5eHHLEQ3jghZrncmXvNY9g+840EMwq55aLUNeVYLrEdCk4OZ4
RI5415aOETNiHeZPOp2Me87z9ohMEHJFYdjwV6I6IljP88swnk7cqXAWbk94QXHw2v+JWxi3aSjD
YTlTaybVJZ6LvkdBM6qHmsSfoBEL3pPtG7LJDHcHlyCOf3cpa401iey7MbUGd/wfYIWyNrLkCnRX
D2bWk0ax9FBNZr2qng7gVDFolz7WWv98y8FI/KCo4mTxzlhVO04RtEOcZMubGiFYIb6F21LjsfPG
8SqfOPpQPxMirzVyTk74ySVbNzQjyedge370OKb9yNqHr/tCYU3ABkRDPvvSNGTcy9jM7SLZ0UTg
iXHlV4lKhiUHYjZ3u7zkyiyq/e1syhImUzSp2ycIvphAm3G2dvYKFQrunUUDcn9/cCsjIJ3LboSp
Q0o5gGNXmuUm8rVycc0YvxaDA5QQzFhlOVbMgjsj3WhD9ztDv3y12KifFVA8HDoxEXfvFIBQQtM8
4bRk3fq3LQNmoTOwuXIUXKng4VGtkvorW4fBAFyI4X54/roQE3AC01EBBSHwNjUN9vsXKeGn0E2d
x8WMRROG4E1WMmLuJsRCMj3mgoJvJjpr0BZVFQKLMG5uf8t1IVgyesHJxh6H31Ipmwn8J4Uz2FXG
i/JVOMU7uSKP5tihDlFc3JSxeC7lMj7xTrsgf9BdfsnH3cwlHRt8nms0QsJjgSSwHsaKfeM0GVHL
Vean1PKjh2CHE8/ditzeYyh4QTX6B0fr+hZZ8NBa2K5U3zEYmehp7HZlW95O8M/We/me4cZ4XQZm
Y+4qixHusnFkOoxtXF4bzSDDm+cLmPZ1eODb836ts4iTwAU3KIomLlHS5e+jROZTYIPr0QhehHQ4
GMcKsXKwZ22nrHK+EevitX2YQOF9pBDt2YasAIeOeNcStFEBZVHZwXdiHDbsgps7nwEZHfX0f9im
sANQlXResZMn6kcCSzVeG8FQtBDK5x4srbXPdPMGwJlokDtMnDr5I6hDDaT/r+lnnT6Wc/6Z+JS7
en9y2JN+CgCBI5dhFyL989obA8EhQsErF03UqlOQOrWQJioRnagrW+L4BGRbYi9ywrrWtlVIuG8h
zjE5spm5U5V0UD9dgC4uQBKGOJigOoMV8h0IiUl+xsoaNR5HlM1VzNfAyDMpmW8z/pcBwsIr5NKu
qIyrYluGaJOjftgZ/a+AlAUDB1pKnkPeRVoYOinq7HoCjPMuX66FyzAV7xkWzp+H9nuOgK/tyjuR
QJ3KPf8UPNIAB773g8BoIf/L4J8cGeH1pMzbNKqPZWyVT9eaosj1jTqV5JDXa2UeHyg734Iwjmis
wo+EA6eiYCoNF80Bfz4BloptBjHUqQftFra+xWkDaNjzXKfM/kli8PCA+o91QsaGnwk20bFKKGcm
N1DSrTa2KNfAASFjWeLUUPYG7UsgoYL/kP9UyFmV++JspclOEygRwAnGLQgfs0jJPf6/28kCNcRK
wBN36mOL+Lv70k3ID1QJiqd7W/8MJ4bhki12TQ5kFk4MZBabjvWkMJM2AVTCz1XvWWkdyEjulADN
oG4sw/4bdn+OkeZUD5Hm1DfW/SmHOhRKn0APCW/7tP0N2FxAhxqfD1xw77z3ns0rMfHgX+IaRUzR
qqQC1RaabcK+HfIgoiCKQzko4h6NHG36xUI8WK9PuuN+MMb76DwvalcV3hbPfHhAwE7H/IoXWrH3
/QdQsqP2gRVq85riirWZiOy+J3ta2Zjqip3vu63wNaepy4cisigTBTpWh+CzOXw21i3QXPfE5mDL
HGBKyS7o+bdMYK1oORRcESNB3GX84lHGywFnT1MqRVMdwm8vQGda4ixN9DJCpGUZrpaLk+Kw3wR8
d4bErWOEVcku6MdtzlZfleUmBmQLPFad+sAbliFwn5OAyd2impkTfKvj8U3rvLc2A6PGJA05tvQ9
4UOyp2xjijHn+zWj0fipGHkURDwJgpVRCS2mL0dXzm9rU8jY1+P4HyfUtG0udKCQ4yO5ZbX/JGLE
6q3HVmjhShW6hkQKCbu+xzDfEOkUWRNgNnwLKsNd4t6Kk83ORADtnv11ZS91BFgDX6GsvBTYpzHm
sr08nWgZxEa8GU+SQoMpmKYAJrmhNU9sKYP93cyMgZ0i3ALEEHZiCRyBXkfiQDBFWd8CrSWgkXUW
CVwIAi0g+FR2zO1NtlSveFBenF9lD5Bb5Q+Ac6SsaFtsxTA9M+bu3PP58fediqLXWib5bcrlMPtk
36yuU8Miyk8Rv3RRmb85NftBzvQ5uuM5Cd5oVmzD8uPWmhzyvpFmkgyufEhcahj/+di02lXJMxYp
WlIG+puaIco9oini7x+/pj+Ck+CC+rTrFNa4x0FKqZ0+PaTMa2twbxhoSIvhhniZAUDn9RhMMYwK
9G/Y4z9Epl2346k33Cbk1NsPZpexWTpkehXVUfG25xpTuEooetM5YR/y2sZ+O1G4sQjmoBXnNX3a
41CSxz8aTVw4cG6431Qo4R/iCpnWk+l5jqdxpMTEFMbn+KAdxSyQd0W9/7kDvs3v3FcqCKDME1bY
K93RMktwaCrgPUbWYSNNUj3G97Sfi+/VgEtcIdeNQ6PvMSyQ9cFXfWa2LnPITVMAK2sGLm6Spb3c
g/fBAsbXZqevj67kO184Z8RialqSt/n68E9ohVDW3CFUt41v1nm9RfBQ+QiXacDFvSGgf7ZxUKnB
jA60VqNQOnJF7ZUe2kriU27Djvprj8ISQUZQ2bAHPCpxt6Hs9feeyyLeT+P65yKF9HCnEh1zC5gB
4pXZCICGJLiptQBVu9UaCPtlZPEvpDKiEOkaE/LAxhOcXDiOnQ2L0FxktzwatLz8HFIqeklyLlFW
aVcBgkvkicoMbCL/uJDbvCMy+3uGQLYgVHZ4P+K7+LkN4sr0VUu1kltA8aQMzHDGxB0NJ5uhsPRf
b3n2GMVtVwoOQetAlSqVWbkCL4rTPHlD1Xp7mhat26hnd83gCQHfI3Tspl+1IXAg7lrIIi9HpY3w
fcRFyAZjAV3vJug4nBBPRes6fxUNkPzYQze0uihOjzz1gtRRhVe9ejFhYci4IxR1VYB9bTOvtieF
b6tKDXY8ZSE07kRGBTAdNlUJ9LvIYGwMZEN+jjL+t2mPgJ0ifyG8oR1RDm+lqXtyKHd/k7OS9uW3
NwQ4W2JrB93+YMgBjfLM9qPxj4w0awwdZKBmDqUQQydCIO0a/VWTHSQLmgJHHUhSOQo9fdpwpdMa
LpZdClDxoobcfX+T/C18FqMzPcm+67PvAHb0QgjNyJiPjVva1/F3dzSRYAbV4F10XiecTflAkdeL
AgqE9B+xsWxJOBeun0hFKeMeqLHbNinKdaP2lGSCqDC+9DAMM0aoUjN7oZLgyoBu5FsQiGyT1Wlj
lAob6Skn9mRCYxgmxrQCe4H2bwSTSlvSUVi8HFUbcsgh6dABs0i8KKBZkFkPBYd8TxORElBktwKZ
tGYWuCjweqMqJH/JInpRlPWtTtSn3fvfo4EUhyoV3EpMBoewg4HbEYKLvqwYr9UhQ4/mgCFLXQlf
cA00btsE0lPhGbrAmfpnY1O1inqi1FedW0GX0z0CxdwM2wADXuCAvkmuRbsgtHa+VobDVHKnNsqs
LkUIgdDS/X0PR+FxGusZYukLF84Zyp3Tw195SuH+3MrAJUnnBq7XZfkhuA6XkcI0IYMclBJmIXN8
Io7sA6rWayk7vi8mgf6NKEnCJ9l4t6U488jum+sjua61CArSMqv9xAtgq8T5DHKOqBS/Lp3j4old
6BZsJEzJuZQ2Bmah4gpfZWSQbpRoavOn/jao+DgbadbDld2tWXne3ch0VknWjjTCEWwHhGAd86RE
Wt1+zReq5tgLU7uhgNxEPOiaKlr03nb2G+rrt3cCUNV0J3BtsX+f9FTOZG2QfYDJZyVvUx6mo9ow
n8hK+KlkzBC+aKYPPerRtUwzNfHfSHPturx1tDj9B+XlIkuTTvV8jnf4S60Oy9+HIBPK8GWa7FEc
34m7j92KWgefXCeQLwUDsyXQFQtqwJfnkJFZdmaBzQjP2cH0vOLa1U+aRzUsmeZeI8L1HXBqIAuc
rVwXQLLFPpXzohGri1+6bO/JTkxdKstHWBsf0s6Dhs4o3ZSSM0DY8L3CRcmZwJNmG4RkNYUk1fXA
jEDxotvJBl7aaTgTfoXAr89XkJ/D8Ni0+aq28mqKvzhs1J5v64YrDNVAZCnROX1iIPY5Ru0gCDSm
79laUMN4iDgri2QboY1CErCPPCvtelUlQZYI3r7xv5AZHh6les752IbM2jfjjI9PHctfE7mrdEK4
7OqfVyYszcJBNozkqY8VzcNTWwjkNs6sSS0TV82ra9pHUA7hypwco8009Z85XMzODjz7XK6hTQDX
FXVLpN29py7S62gs+bZ32Y1yavZ3rUQGY9phobtPnk4YUROhHFWRRPzwoZW9+/Own+7EtIo05ngM
JHkAXxn4jcNxFUfPAEPn4VRKJIL2F+kRUmjGiFvhbu1D5fwEmeUHTmm8rQCok5ZeQUfTJH10gIX0
3TGv3uKLohTF2caWDuxQ2ea7dzUMppJzYfX60J4r4yTNnxzBQrzt8hhLTE2W+4kqpZLyDS2y1+yS
TstK86jCbYr79oksg8M2TSyf+4OacWDPz1tZuDm+5cvJJvlwuNotfqNYj/aDdDMyJKlNwSuLwVHA
dWVzo6y80bYBD4Og9zuhmxCuO8G67lBQqSXV1tdbJ3JNVxEYCVwgnRR27U4n7tMv080VD7oRYW83
ZDKl3oRL7hsO52r/6tZBqFSGMVcSjIIFPQc1JasSgl4jAvmDN2cbKv86isgRi6k9a0LMmbTXhrnR
eUadfG+xk1g1drZPeDwZ3MD73kdldUKBpElUZUU6c9/fm2c/hfzWmA2uRZwTqsICQfXVHST2Dh6e
+yKlurL7s8g16yCpOXVJM4p+IsIFbqQ3afXDF7TjA9fCvfNI4iNXQN2yxW2oQRNnX87Zb6Ihu1cx
flkChgOnCct+hWbbirJETImBLU15c77AqFBNHrq6mAS3okNhK7J+nr1jQhpfrCo2HzUMAmHfTx5J
O76nm2y249XfTw0dgCkVSOs42D7bz91WZhCRi+mtfD8c8iFsmed3kOpzERxQSavrv/5CEZIgK/Pm
gUSDPQAI6HZzIgFPgwFAfdnIEAauTdGqcqibKsQc8pO7I0dZL6o28qvLaQkhBa0TkJ0BjvsPCkH8
+TQv3BLYeqOHouh6j7ZxMS6RQdIb6VjWMs/+901w233XUbNoP2xtbQr9Cj7BFGuhUtd3kTgRWwTK
uj30Uro+CfL+U5vmrs3SS1mmOnXupx8XYoJMfQudLjmDib0FeGVqznyNjRwt3E8Zt9DischJa8Fg
upGVWLDN9NBAFFs8HXX3NsGvBS2RYnvz5NmELYUb5YvTCTWilZkiJyssyOoSaW3ziy3x2aX95R2m
pqQJonGdoNUq6s9o0c3RpCalkSOIyMNhWzA7+7H1coDl3u0pBcZLJHQv1mpNIOkHwrX58SgOhrtk
2vRkrGRDwvCb7ReA6/4UWP/FU6+mx1svcKy9pn7GXie0wIrGl0Q92joLRJaCtK/EUGcT93t8tBSz
HNTr3TTmlbbmFRQJVCNSGOHCodJ+v78PrXoJS8iQTlhHbJr04PzJe1o9+ycK+Hfz5JNYZFqCf7PC
P+DSLnS3VMypMItQFx+nWEjgdxH3e1WWcEIh65Y9A3/TsG//WwE5kp3o9dLFMZSwGX1ZV7T2mxDv
SU+maoLZX9g9pXcEKAfmTvYylGXng4tHwo7wr6kVF1dL4soS0Rw3yGPHQJT/4FKQNE2jTpKSKLfb
8hf/fLovlAqRTFDDmXwwyzy/3hU20gNF5SaOoVq5xbTWUzffvcItRhbXZ+Md9JQMNY6uPctHNhnp
U6P8fQD4gBNl68mg/GUTOm7TbeNzoyWTvSxqxOiZpIgWrbEcuvjhMfcISS7VPb0LyvVaskNYRMRF
K8RF++ayhsan4cZIZXCzLj6z4HvdL1iotGcRddys0JxO5gtE9NVX65VwmuwKGi/GECIwOpwkKER7
mNFlKKO2rVLkp2BxKfG3G0vds91/eQF95fcP15+UqUv4441d2LvZajnS3bO7F6LoWGoXs+f82Yt/
k9Dj9hUCpp6Nlc6C6mO1qYTM2SK4KljOJh4MHpOSU79IUJKcDmq/xTdjIyyJXp3bbiJ15U4cVrMJ
6isAqYxKlXwtpIX4pMpMc+b2qh50INcNQsxEqLtVQ/HbjAW6Pfl1q96vw6mMw3rDdgqkkfdvOpwK
8lSUhUSVlMgbuijb51rguqrb4TzSX3PWyqJbwSrl6OovG/riIF6ux+rcc1UTgfKzeGMSwVWgksps
uSuSBowADDo8gRxeMd5xs76s/KJR+w2AlNG2v9c40l8wnlPbFPHsAaw9q9MCbHzDsEIL0GaPcbxD
IsyPSfY3DIOQwJYUhH76thJwNYVDaxzgtoY5Lur5nSBjaIKk2CEePNLBftnVQqYG2hUdWjzG2f6D
sjb6gDHt1HqYIX+Q1prvqZGd1v3y+Gqr1R7ZcATDpA2ktMmRPTpVy2rnhJdfQJmHZUG9DqSdPgbl
hoQCAYQxgXPg+LP66gHZJbItmLgq6uk7Qj+4JfB4DHMjy3Kr5MfK8rWvRGQ5SCnq1URO+AdM6mK0
a4faube0qpiU+dx+JIxVej1iBwnyJMi5dJSflBvkKGHoI8hRGeqpQqCKiGeYtcOe9JLwOFsjxay/
RXWpjWBDqYlklvL9uKxQgRf4NWhNdwZVSwvi2rlfQsamcqEfyr8QvaTgJ66o1wEhiiZ6YsL3/69H
4SefFRTth5zKcdrSBrtuDUM7saioeoH1hYDgKIckcibR2cVek7jg94lWoiZ/Zj8MWgBwPGKJi1in
A8zXOie2aTuPj3mYr++HHItoPDiurgvBb6s9h6SSWaxkD9K0U/8GXjfcVN35cEAImr3Ui2SklJ2p
gfAfHh9tsnGvN37Rl8x+TMipE86KHLgjDzmFu6/+3IlInhBssw0uq2wT1bcHvoepD33wpCThSn41
M7Ns/yZ7bOIrPfApTTIN13W4TxRLG59ZCJRXrqMX1A5Ewzzzuodbys22MexuvhMeirf5fEK/K6Qg
f9aaEhayVeUuoiXs7qz8ZRJl9BICK/1CL2zLNN0F9oPC1o6PfBLirgE6J+770J0f7xrEdZ0TDFQ9
VSGCXDdDToIRMf7aUNwXdta1+NOD3mvTIS/zk1CPEFlvcIn98ktOQg2vin+lFUTz3AIugXwT8il/
/EXgFdMzy3c8snTI5zyj+xSb0ELzUdscwUiw2gGyeNdmY9kEn6S+rexWh9114SEkYqUORV4ODj94
9sjCo3W3yo49sjaWRppNBNNnq+WzDunU97FDa8OHosveed9iNohQQko412fBVhHN7d0SePSYgghh
W8A6uqGxdiveAkHrARJz+zT6JalvhOR77Rc1D9eMdJe7EqPTxPGAQyTsayMRiA970z79WlmVQqka
0/EdZUWZnhFwz1i2nDx4SIjhDMlaxiKdR0OOrqSnW6KueP0g7s2y7Jzhza1Py6/8Lc7K6ExOz0Bq
zUJH1Mm4JVnLsXqz7Xmi70ATlaD08HGO9MVurHa447sXwxbnltqqeWrhFsfmpqx7sXzKJ+rUbSMR
gvFsbLlv8uFpqKv3rBFrqtOCNoxG61hsSuO7LPs+lpIkCPCSUQ3dUjGoN6T/VqGp47gAXz43Ij4A
z1A5KNeZHiRNfRO1SBrxack26fJQF/JwDBu1HqQ5AeHihYFc43KBRw6I5ZksVHtgD4F+Tz4a0bqZ
GVKg2FJ+wgndmyxThysdEGvB12no9KnqzgEM0b+6skLms4f9zjAv7/OrSmG9QUTAQkRZNBnPvBxw
MTYRutLC8JIedhSv64ZYBbnO0+2digPr4eUZFiZi4eqeLxYaVslZvT5INLOrfhtmnjw49JTdqrAW
+zlmb52TFa+I1z3Blcc6mS+HkYgrIeHzGA2ilc6lmeLbRnoSeFgtw4biuBmm+s6R7TQqPn9CnYJD
XaxINYP205vfnDR+NIF0mcuKGfiXdaAp45yXjCrlSAmtXqAwwDv6CvbiJ+h/81ZtBJbQrQXtR5s8
kY6bAp+lLE8W4F+MVAV4fBFGhqV+Bkog4Iv9lDoSulTOsqq8zS0Q8qWzGrl4xEzY4QXcRzA5RHsU
PaKpqLkhmDOQKHD2URoz2BSddP2dr8K37pnH3JeAHgchRQwho5HFM4bl/4jEqQqOzuq1iNgNe5Oa
7Q4SF0gOAPxx7Ef6Gugzy1bZJMzGrBH6PqbhqPYqbXErBUGwHAAZUD2kvuqnzzFOSjmzWBv54xT6
TCCRTgoiWotRF0rgFbWlMeM7KBZdasyIctt1Z5ZLk95H0lxFuldjnWCvjcPavg7lqwBvIlEz0hQa
C2I0ARJHLQFF+iVJMjBRQfIw8pTjbM9kyBEhgGsH0dPgLJK3ol4qWEjqbY2gKeuHnNVxEINUHWbm
GcDphdRUILja1Ed2LtHeIe1ODDpKod2Eexi0aZIdVcTBiOjU+P1McY0xMga+/loLjGnYVX/3sNnN
GU7i+/q6i8VdmVo/DW4kL3yiJT18HRDb8AOAdShw1+vzg+rAKnu/Xw8t+gCPpptzjBUbghBRxulP
1YnnGXsBGBsKU/SvMgs/fj3XzehYXyhRfgxxzbn2zaWXy4+UoRrWUDsH25VU1PrWNX4/m6Lyc/4G
3WE/a7WoRH/p2nmt2E+ePj0jLPGWUW8xyTTcUQ4wxa8cSkFsOCLl6Wn0+aG62CYEWxTHHHNOWVpy
fUgtcFDqAyV6GoRs/pj7t/GgvuDnJ+qniDg+VeQNU13lvmQTxPSnMD0GkvrD9+8ttE0n7xqPYUpq
zA8QYNjR/83GA9oMRBB6wZB11XNzHlkgVtYeMg0TlvlSbkH0vwpd42qSvQY9R9dFbCDp08Hz6P4T
93+8oc3EODCD+tlOubBi/uL5bvLVkavGuIZs+MiwHZyK3zOpHEW+VrkHTm7iOcOBikbwK7W5mlnq
Zc/gWjMYHuY6giJq/q87aqV50Gg3DXNvIs0PyI6c0UAAvTXSYYsnm6NlZeyTuhdDKkU5HuiCjyRY
XcQ2CmpHXPOOSn4JNcOBzxbNN+X/a47ub0SD2SCbjq8BBv7ED15T1201jeqwMhu9gjxCIbbPQJCk
04xrHH6k4y/7POb+cidVtUvr7HbjDvdCvP28jTTii6XHAouy4uCp25MUzMThqDTsea5AhW4cpqKZ
nfs0o5Yg0QL5Ou9CycoArurLBKeYpUcgV8zqC59uOnHBLusQkyUPYyv2JLBdU6I+4QT3FvvymQDA
dPbGmPsedlbOg/KaoRVD5LLqkewHl4Z4D2Pvc8bezvZmkF55MQMPY7H3j+H9d3/I133nYtcOGgQI
/2KBfjpOhZikS6yRVzQuBKp86uMULdfWfpzgJxbPsZ5fPoqNVIHanyV5mLG1w0EokvYID2IoSxoz
R4TEh1/ABRFApiZeoHLb1sht6I+L8g2qcWZ98iKS6mNt40jW2WNMwhYzTY2z7D6TRYKgmXgXYc13
xamXH2gtiYxSg4CW5qfxbF5a+hal3b0IvuBI6RFscPPFbx73+NDUfOPCaMJFS2yHBDWtODfGRsjI
4YN6RjoJxebakX1XHRYduxIBhXE+KiPuuqTDw20lGnIA87PW/NBk7l6O1a67ddrglsfWYDtaKWt5
0KWQXuWQirt668e7Iw+nQ7Jdhbap8m6V1YYWc9WTc8j553I5abhFIdxb8f3x97dowMIxTojIQ5Cj
v/1QueySIzu/XR5+6C4ZXaMcivY58efk4KoYzIgo9w2I9pFAtdNDmt+QfAmG2YNPM8cO+rpVnOKU
TkMPTbb6LlSSYGM460V8rj5hgGbs71m2+/sEom7MWNOTFKmPlS5bfPQnXRi3MOS+mmXyv5zi5D6X
AjAEUJhIZSvhSFguTtYAIuJCPi4SN0WCdoFnPEvGS9JRzXzZLbonhDRtXrqPM0L5ctmQZYwxAiDI
s+cKBVjdNIdm2D/V47gl3eAMfaE2cKVE7sjh4QPwb3aEd5yYBUOfXZb//uzWGTzd/ibv1ymhGgKH
WTyySCuJ+cKWkv8PMHlUdERQlwlAArcKtXUTTAxuB1bUQATRSXMHo2LG6XGeII9RmhPswKRFJFjX
tL+/0ak4kB55JAZDeQPIN5DkxFYEE4wRUR+nrIPtLWmMUPUyYF51JmroJlsVDt6t7MuNiKk2FJng
CApfgZbiN2xfFHIFywoCeNewGKQZ+dUIQw0eP2L+Z6njyYT2Wje9oNMlG7GBnZIIwLeB04BcfkLh
lydI9ZBEffWlQojvTw4Xq+QDIS65EQT7ioCylqyY8B3UEPKVdukRns+4FsNgQm+6EwEtJ5QeGURE
BSaVQ/9DyObZAxRrFoGF6IIdIFVKHsZhj2568BtlzeYNYxeoJVKgW7jYuET4RqUau0vT4G+vgCuL
Mo3V/dZhlAAmCSb1syqoF2qL3f6rYygbIK/n1doEcVmvcuxGIzyWk4K84XnkM7cQXRKMnj0SEmi/
93vioKniotDkd8W52Bi/8OG5+dayJpjGIfB/BWD7H/tvgJ0IXkPbemhhcIgAqwss/P85DSiFc1Ng
2qUXucqeJ63EsErMm/Etx6Q/x1l7GuufSjRzNm6uFIQMljMhs6q3H9HuiO2YG+UiE/3qtbGGBpRn
CekOLJzBteD0gkiRuUJorNgAzvemFphCSMPaWTPu4FaKCyQNphcMIFjBYcHXILIoIBErukAi9amJ
UnEMeSYSmBGW18D7deXgKZwW0Yv6DZS1uboQE3UVqGiGNlBiD14AsINNaWbuYj//y9F52WRLoU7f
HLW1Nwy3F6kFtHW1T+T7nMQabuU/gWuhuVkqMtRZPfwxBOacPx8RvGk8+Aboq6+Ih/3yJOr6LleX
s/ncoW/DurWrlCSt5SEHYWfpTSp1WbkWlp++YxYun1cr+i2ZroLHgtg6XapjKLQlmZ3biEmu7NCo
UgznGdj0ayIxjIB6vt0QkMNrWe53ft1R97qQHuyQMMRYs+Zm3vdbpPV0d/IoDAOIbDQvWWVqtO+z
3kE6bK3uNfT+cXUG2nG9TSIVRcee4z7Xdb+9MEUMZsuRkLFV6Wi7K3Lm00pQDZSugwsmnrex+zVP
GV/L9Hbj6tlY7WWxq14ovLTOTN2SYNja5tutbixJhRefivkSY2DuE9izzj2eOQkAyElWUNt9+L6P
sOGFdjq7N7Y4RbSV9TUidUKGyHzzAna4HmQ8+/VnT26WkpV2mLrNDSdW/CMThDYzffC6mPIHV11v
5rICRZJqEcHgSY/8PD8Gwh1AAnQv5GEbv5Z4i0R/T+BVehDzP7ny2iS/5sA9psDrDLNW+V5TwvEQ
PXfw2pPtYSzzwpBYem/7LpPWa0kvQb3/hs02vrXtAh1hwliOyAW0G0f8uC8yZ/T4vgc5+w9ZxjQS
cjVOCANtJJJZgUXO4RXh/IoR3UsKB7lDtIGrYdSjn1ilzAOc2QCJr88rSBf/Jj5zJZHwgeUAtt6J
FQ1fCMiVMH+vzxQLy4xZ5b+DXd8d4pLvQXrCiuAQE+y+tlDYvhnLxqpGJXKFNH0WRQy5KJSemH35
LE9DeBw75OLUQJT4EX/9PrT9+M0bFV/T671Ot7sHb/HykbFiiqBqGo1psKKbeoirviBg/3BHLwVl
+EpUfzxGQf42lin8k8cyn7MkEROGKzLqfw0X8uPtZSFRiAivF7Hfg4V2zOEJz8/qbmBqZtZaCE8j
TUtkmJJSXL6j2kMuGbdp+J14BzL8Lj8YSqCBeKf6mdKBar/oj1w/Zzv4T7NdrWrrEk/qKoFvV7yz
5Wyk1kIwTdpXvNpTzF6A7i6T50ckeWJAOQf1Gx4vvluJM0Ci6mOYV3Cg9sR02i2/IiE89vAUHGDD
7DK4zKpUi2UFQX1Gq+GHnM4u3f6q6+RbMzlNVJzfd9NSbjO0ekq5d3356UXLoH9/qcpnb/gvQ5Dm
p3O3ovjaTcrnHCDqd8QwcieuWsmUNbskuCfqPz7zll6PFoDGMYQa4es9PFvMKhwTe0hkuAx4VGm3
rmUxZJ0HeDuNgJjrHwOon1cxUUwcJ1q7H+p47VHGC057gwhELsGyRYQhBcyFzDKFbukHnpmHja4X
dtunPyWJh+/BkHpPTXgKMF/gKF9fsm+Tp/m4IqrhJC5kqeq4YIGNP1YVpVscIZ7P+rCt4DxflQon
OacLN4gxqqQhexz0wmOOV0rtJT6gMEGMSjka9swoAcUhOR8rpRKVqn3M8Gz52YQvJeKl0yeTuyPZ
AffEz5KSQo+WDLhuywqm9PAnoccVKbx3kRvTXb0Zx0SffgSm7ZkCR1j3CVWInKEfHC914XB5jXcd
v8bncgHe6MnhbXtLBGjpsOcsFWYEqE/nbSOWQXFApVpjBgyGu2FcWp3sSohQwu3M9DWhGC5hoXI2
6s1Z71ss7oSx3nyecHb1mGCzN98BdQy3UV1Ikv7NHupsxn6kaaJzmkYY+x5AEs9PmJ5p6dcgc8/p
QMBPQ//BCE8uiUBwzS2Kk2yaayEwu9oq9F29XPwEaGeaHRfiUMiO/d3A/J7GaeJ1zySzPlDhw2zB
nReZ2C7ftYMk3bePrNKPIde1tGtyKuZ9m98qu8WXdRPExw2m7Zp0eRqxfNr5iJCX4gIenwsvobF0
/T61Virs6jkYzFd1pNFaoYB0JQ3ysqv134kDiwa/cgpkIGo8bl++I17ca3CJsEpG04aksQOmKMH+
5/4ov2dWdwQi9Qn/myC14OAWGvb/jFPCxFpNRsl70XPLEVZ8XHjM/+U2PbuKMrS9fXRvPFz1wFXB
1q94B+HdEvF4mjyokAlkTz+wJFKwxf253GxLl269bybJtnl8xTcxG50BWu/9p623RLqMs1pO7mYy
re4YU2ZOiK2PwCIp6NGNyrSlxrCLGNz2bOawjMQqoqce8/ddvit8IzE2KSal7wt7h+BVmcY0QYCW
F4rbmV+kUEtZeevSrq4Vv20DXkJSECmvQf4kE2aQoL98Xq2HdaFU4vl9/JNyfzbf6l+EOVgUasN9
zDOTher8p0j7hCCqupww33lbVX1dgO71PTxWgcS0ezeia5Xxy/K9BFgyaj0WbtWxh47DKh26DxPF
UbgNy8vmbDEe2BHPspfw/aHAqh9wc/Ikusdw9rYRDuepTubvTDkKKb62Mweb1Ve3yi6+dhjAdBKO
QX2I8u3y9Y0pUHThOK2ruGgvVKgVG4//QzIhV0SBgagAc58nm+bohJRXz80Y4HSHvCAFS5Wa8Eay
fABluo83yzPSP6TeTPm1E4m9fLE9ARbmilY3s49L/xNzr4tPuXGIX1T09X7mkfP7tr6hSd0K/mKk
w2cYBgpJhIkWi15fdkwPp7CGuYAjUJiM+gZb07Wv1iKTnDZGJFdQ0FfChgHxIenrW7CNPc6YiHGy
CR7DlKrEPkoffjp76Ory+DfuUSW4SB9Z4CITAxZF68xVSJMoXEjQUYxHHjKUcuuKBKCGP94YpQz1
KXTo08UU1hf8mUNqDz3wFesPb2qnHxSCCLIipUjMso/hTDsrq60pOPLDmGCRpcZCb8ia7cIi+swg
A9+oMOPtCg99/jc6AYFMDyH/bZWZckeV/ERztqD+XHl9LR1oAG/egANbIYiBxQK9tU52byKAl/Bx
X490lxexsh7zSqd4fr0CNpNv+C6wjQ9ov2q7vyo6FDNJuqIZyobJtukCpYVsUvM2VWwY+R829AVQ
FbdhKPjKDudhnn0p5woBJwCUYWCylCLVvSi8uJyYCWtPvvghwcJE+x6cT8AiF5koYRyD+/Yk4xQG
bgxxDlIQqsMPt1rVBVSTlt1NhqIgU24EqaM7xEPcHAIi+mPfmjjxmb2gwXaY94i64N+aEWZlZz5C
08d9JirgtLqKmzKo0of9Xeo8IEDhRganSR1J7wdxXsKz4xp7LnSKV2glIpaPMFgZQANL+T0TYTL2
tHKSeDbUly5rRZYulRA6qHrJXha1lwI8Y9SIOPCol4q7HtLeAKoeEMdyUyJWiCp9L5oGj0IyAaaW
cVXKCxmOCx8CPdwtiYGKcNeGTepWUctPU6p27vC6h/SdFSDwgjVC72eFD7EXfqdtU4Irjldwvo/3
kp9A8nWsk3MgNhgNWX+PKFYuAkIkCnt3uA43IICqSpESx5+YT6/80s0zcEZQrYvD/F/Pefk1le+C
SEGTpMmaYY6wDqcWp86sDGcvYYHdibZ+8lp4JJJp/ajHkbBMUckkzcotouYfQoIAg2mhN0zFg1Lc
ZfmTTUJ4IqqkRfb+FGtXFUHUhbDd7YDmOQqVb6sNKnhnL9kWzIFLGA/d23Ybqg4hCIiNlMRjwQNO
8N0bJG9yAkgGZz2Vdx7CkRuP9FAVdpbCGSit7bNcR+jdsJcunlGgVBAHDe9BmI0gtnaBSH1Gvkue
5mTZNQfY9jpagNkTxF7gZrugEZzm/pyBJg8WEXsw9Q4bkm/uftNd/rrfWRnlQvcke5hmYoRWrck5
5fxVlQBnp/GT5iLCZQByiP/2ap97xqacm5ie2qc6PbnUitjhFCcMa4D5TfCWjGqRV49t28LNgXMb
LZNkmouJUo71bTtIhqc6ZC/kw/JWVJGiOv0SWy0MaQXFhnfQeQi+4eQJQ/UadK1VGTHgAxk08mxB
oBPt6XDF9pln3iQr8b8lUG388Rs8gn6lCQuK2ypyZs+EFHPVxcgisLfUBYSY05qylUsOFaYIK/Az
Jpd+ZuHlhGRNCeaOn0e3ZEU7NlbkUKKeGL4rGBS2FUA14wFe1jar5FpgB35vajNZ1RL93WlHrK9y
n/OJoToUV0A3mxbVAIwWadodrB5Ja5nXmx/ODcfPOkpeu+NN4MPRKvuk4PUiRp5jrypcxQ6Lb0A1
DEeaKnUfwv54OO7pT2RL79q+znth43BZC4j49KHMRf3qnWL+peWNHt0odOZxY1Ya3yvvjUbD85Zf
kN/+95/QLvnh6xgzXsBhwM4lKHCtOS16TKyp7SSTmRoTw1BZJVQ004h9LgC21IeJuWPmHsUhT/WJ
hUNRgK6fNrkDLPT2ZveSfYYYtp66i8cCVq/b5NMljHEdIRs41ItcrRsLhY9NdbAESjVM38kFMQSC
md9uyvpw5WSzdZ+/t2YTbPmIzSBr/95g7Bs8QoheaPj1HdqGlikvESTXJyXa8llt1TKTFVrYR4pH
Y7qo9tMiNrMJpLgQe8gK5Bwp7uPIbINBm7uwCPnCYvDcRFdnAGch2vHF0S9zHYD9R0gKvYAzSL2w
tWM13W/ZEm+FU3PYDlZ50xTakZTyoFTYqB6NtMc2YXZf7wVbhPUpvEsAMVCJQWlGMJGjX11xYkwB
/dL0VFlYcL0cZtYZIemOgwAb428HH7qxSPcwk0ynRky6Xkgq6lKwfMAAYnVDeqfxPWwane/CngOM
eMwCvheR5NusvtmBFAMqRVNlbQR6Q2uw6qdj6DIusHj6+kbeoUx7ov+2/14n2WCjbikqpO+523Lo
5N3X67cY6dN87rlawW7PvZmkuQ7TuPtIMOfw7WRNrzh+lL2qzuMun7BlEc9p83fxqGLfSQNpQmgj
e3pm99j5avcGI5roAht2W0kBxcqBi0Xcg1zJ/1gZ1/BIaNCAi3sxZjN3Pf/X/RQG9TaKQx+xJgWh
pKi60ovwqKeNF/0PX/OIbkiAjkAWztMk2ZEHX1nc4czt3wfDcE8SG0hZSOgGxDBssEYFGetku7O+
3HZFiFlis3+CrP5xwYuuHU0Rf5BoV2hHGraI9LsQatgn7B9UksfgiS1/G7C72bbb2J0UQXWCTL6D
HjZQPO5/0Andg4frOycNmI7QfBUARlEuq3PlurtMMJW32Ouo6xyolOmhQ8IdLljJh6wCk77LQr0H
qQNEu0CNn6wUuEywJ4GwCIdjizlChvu/OXj3u+NI53q0KyyBrQyTv3qi0dCT6Dvp2O9OXBfYIh5D
aPON/QPT4eLk3bLw5+jz9sbWTAXldGdgv1BbngEjoz936IIxBC13am4vbSXJHwfGUxbKrftJQ4MS
9feSOFp5WVQCbQNuEqJiugreKqWUYPMQfvTtLanEYgCjUFvTLMgeCOLEQ+PTDUNrFfe4JclFcUbi
ipT5HR5PGZ16ENAeYbmLtopU56p4owXV+pIwjsVOi/B+C+ZgGTV4zriDZftZpP4Lu53yOPCIrKKo
cb283cNLSho3xiPRGi9/84O4y2F4IltVuXlobkk7ydBWWXX8XDVU9V2rzWLQoaOrlissTL1kMOQT
VNHx9kV8/cXZDu64nOxvBcWbSO2c3k4aev/Md52ODGVSOmxQJy67/734EqNmsB+VrK2MrskIpwvI
YI8O0BWKSQLzlc7Cb+ZGbrb6rTbY4RYb52m8Vhd0FPTpxn4TH5+IZdT5yWfNSsCpoLGllEE08jNa
K9Nvt2edoMQsRF5yX2a19fXnfyXiup41+QObVAmNrppUWA64W9BKyg8/WjMqrvOgenx9BqByVIU0
g7O4cphcOON15o8kZ7hGI8KdgjnsEO1dTBmqVdqN4plyaCuAiklK/1O3mOjNi9go2e+SYC1NtzmB
VMSa+B8B6TkrO/zPDy8v5hJjMfAjRvNsfwEYsVjk5Ewa4A4qEq8IKyuzxPuT0IWB+qxTGVxET1iV
6hpzsUjMNqygm7uZ1BUkufOlqNXGl1StUDGkOGHB0zDCpSDZcbtPM8xOJa8OLT8zH8XejpJ/OBx5
WR307s3gpJeihvbkVtFeTTDOAlhePsyY9ieMN4NBq3O7LwyAzS+zWtMDcenzkPzLJL3Flthi6CBD
AEqbwKjs2YgsEcgXeUSQ7OS7rxg7NvdtL5OjMz7eh2dBjPgVoI5NG/+BZoNz1bccBg2hfWwmXMkp
fL4KXsuH5PLDZaBEiogL54wVZsrMlDLs843VJ+Gpr9XdFjDddawIDPUiWZeJ0mZx9zBgWxr5jgiy
kep0p7Wd9BCJfBrhy4VRA1P7UTBblFBewmnyCg3/rnWTL5v5LGhT5XFYtzNdQFnJhUJYpliEKg0W
QNP2lg6aLuA934st44rvmShdqXD6WQPzIbNdDuc0kgQos6YAW1uKHKtSHUGnGh3OU+JW52Wmsu29
G3hdP4rNSLqnRFk/jOn7GdkrIEcrkmNFcbQ7/248alU6gZPvYz1fedBi9AUqT8AurVwAT/9wPGEQ
lSQTG1cl7cFie467csdSqZiqZCMk6dpSpT8CV8z2AtOch7Y7pNC1xJkJ7yVDjfIgJDebayV1+euH
09wUrHlnA5kkcap4kvlMSPtdPydNVWZn5uxSd3ekDcpRcAgEpIdQcQvIkNl6JfE+AdeP2hr9MQ7V
pIulwNmffplRdmDQ96kbo0kdYGEZueqR4iiOkQqoSVFHt/aFpMtPiwyzWGThyN2Af2OvURnxNK05
kQiiJV8HhHsJnUcegmLuW5kS2z4dQzlIRpdENzAn18r945g/z23H/IjXO2v0lhqYTJ12D3P66Izr
ujjqNu/M9H7iFo9A7rfN3dgd7kWic+WZFgtiYBgfeaYieyvZ437A2dEQ/d+lhaE1jgu3Vgd4O2Mp
U77PgyoGbmuWn4rF5C01CCeGLV8LmEcpUWdrO71DdFzR/B3bUwgNggoVq1TRVAFDMSaD7tYvTAVi
0jNJ3/gjZDYWBqYiIdyWDBRO9J2u69+IHswQJo7mlR7Brrp2CFY9TX10QMthMhAy/gRsogoBeVQ2
Zzu1DUhs0ssD97eZdIK3dad25dlZwkxeTL0sYfXBrQgo85bunsO+dKfUAV7idHtcAbehwcfbnHdT
3cpwIF5HbHk9LmORC6T0InX9ynMwoYoMbXvAWllawbPIGiW2yz+8d3myZQLV5tkM0BCnqIncp/GW
zz7HNfQTNqWKlGeKawBfDQfbZ2lyTIJ/3ql8R/SKPkG3BS/B7v+Co0YfDkoII5Cbf+gKM2G4+1hg
dOfEt7CtOOHnuZkVIkewGx5vi03IE5D7OD8BQU+rhupTzo9g2TfVQoPYH8JHBS+9FOVk+spCDez2
sB++CKNztO3VM0/f7fRqZcKzeHMmM645cL4Sq4tay1p2Ppbk1z/Bq6t7HWSUPFqgACitCaslqVtb
+mzOXVmQcZSncAqCho2zaWUVTRehghlw24h48ShYB/R/J4bGIDq8iU2kl7DGKLbkkaH+inbKhjCR
7YE8ZWfOcZWkzt3pUbXPdDwvhy+sV3jbfcnLwQ4surQ2nrNAS682Ct/UmYGF2GulTTfHDSdFOBUR
q3Lj6bILdWjBsVNbhba+MSVW5Ya5d+7slt9vOBHnez9hKeYsvO3OrfIjtpxkWwT5zXX1E9YZ2m0P
Ki84J2g/b5zV+n7So6YI148ANynpJh3e9HYaSKAF+D7jLsUOAOParQPVlI/5asBpzEGjgrfaawte
rq0FxvpucxwNOg3TqnIpZymZCx2U5BYYyjivk1VhiPmF3Avj+ZKEp/j8jZrILmtqo/FXIyg7DhlD
DsGZZyqs3oe8ha3duw82cspNWOIgGVFu+v1vWF07h6RLou1afoql72zwhLpJN99vsqPqj8sXWTTI
TkOsvdZz4ww8/hUPMe1GcBQ8Im797gEiUb5glLvr0N1h/NLRDpCXg2wzcKdOV3iR25o5bdm6H4kG
7JtG+TVZwoa7cotaW3e1BRjP/L8qOyeJJS51kZ1+HCgp+kytOA4xZMoB3mLY7leVNWC/Qp8g9Sm7
lUzJdXHoEBc80q90iUMNYX137C8w2Yk8qAr/0J2ZH9CbVtXWBABXnK/yzVYNv7kqNFralklSA4Jq
l4LSHjW8WLoke9XxfgSdVlMDBfhsH6EuTwDb23L6LfywL/pJ6QNn2/ZfiS8326ZwZbpVAxoreLef
TSEiV8OhU2Xnvj2gEhd/SzCS4RshYYwhcoWsNypdn+M1ajmjRlAD0NBO+ghZegChH3OllAAuq9py
rH7K2Ps1rGlM9MNUEkzqFyhNo+5wkAFVqsuBpzZobSuPJWOvUgSx+TB1jY+8MxqCNva1MKIjQKQ7
z6/QToUz84qyNWnmRJnEmi8ZxVY+qJPAtxP9MOscT7lUX4gxgYH3AZi40WTGem56qpslAB03APVm
2kTCWpIyGGGl4Ii367wPb1IPSytppg9usENwxLJVR0gHXTETBQvCWi7R/oyUL4OrpY40heU8E6Zc
Zq/L3XHXILyxEaU8q/VxPObF72lUAwt9+rFEVJhwPznepSu7KOAWCOQ1QuWcSklmRfhd8UOHGLdH
ZvpcSZeT75fb+FaEqAdWL39N9qir7KvFscJhFVY0fz+B0xQhCBCB/VKDvbQPWS7DEVCuIokUt7sg
hIu9B4xSuNtmUjYU7fyNU+GsFQtKhah2nm/UCUR28/JRJUL9UM4shMAldB5jVlQqH/BXk0dW/d/g
jpd+k/CUZu8tqlbx7N7hhiie5+sHWHCNoOZno2e+B7720k0bKgj47+OPBWbRUyVNldCoJPP583wP
Yr2oZP523eBNj9FYQANhPqS6n0KngOm5zlWCb8dO0J5WxKYinsyd85UfQGqH+3hJwVt5AEeMyx2v
Y1452qhL7UnwO++X7F/ozPK1BvSk4vha0S66aux7ENYb9HT/9NrZJ+Yzp7ftQxnLgkgTW2/8XY2k
zWeBWCzHSe/Na0nZ0Y03NvpH5XDqBVRhcDID4Doa6GfTwF46MHGv5H0TMwBgEfM4vXFBu7vPolxd
QyKv048M3u1BAS/dyqrHjv+cwg05+TR4knYIMNEegOSFBvW8ykzZXPXCqM1c/UmAR4wy3oYhKDDt
J44teNm54MskXXiW6yjH0Dme6E9yBeSuF7BPDys8QPFPUcuFavvPLTZyCpej/C+DJC4roeg1Q3+L
17xchJSLmhKwV1fEiyNxMJbEKBb9Qi0B9+q6komoNxMGwEX6Bx1qqh8VMYUuXZoEqchpgHwU3jOe
e2K47BFeRda99yXP2+PVOB9zEIvEB7vpyZZcgMzdgQFAI0gQPph5KeUv4vaObenXAheT5SmxEobq
SdHzfxhyWVGrDeKSChIPtBJ4gbGeFp+ErJM5zImiSt5TKmf1A/sYa4bJbNBSVVf9CkyAVusJ/HWA
ihpbOhHraATLFPH3FAhITgIwwfm9VW37DJqgW2AMv8EiFTroGVo69yWHz6jvOVooPdT5y4/N4Vcz
VnVsfwFr7PZ4S459dZcQuKvmKz+8lKKmSebIZFlur0gwtgjpY7eCBOrjIsccUdhPF/lznnGKsLOV
3mxxvkyTnohsg5xUn3MyEp6VaLPXPwu2uqnuCzbbyqsHuIvegs+ovfo4MCx7r6FAWFerVFdbDols
7gkpImfXBhpwUIPs4tsLoynUctD0lomaAjd+moHqB+OEjQzl+ka6DjGB0wo7mLJxRwEgsdaiMJWq
aypuUfBYQFsG9S7ph3EPmRmOubol35NKtznFodn4ix6UerxPhnSZclo9L3ylMgtyzks6+Ag37x3G
wUHxev7/24MedWY/jdCBcYswsKgBf6uORkc08pURZRuyVsYp6S+ASuRlISwYp/nzLCH8d0Qhv1DQ
y1+xw/uzxzhOEWqtsNqMxci9phl9FBYfEXbHjBwMncYyaS1dLKmCT3x/Xiyq+4BVuJzrYt6JII66
yHYnb/+66asbMq53FEFGWHjtzb16mStZcvz+yH0Cz30GwU20Ak3jGVqmZYdlNBF5qKUwYXHQgzgB
SbEfmdgS76VteUcidOPTiNEGjHocgIyc07C2PX7ku9I7zpQSVLZHd/VOX2s4JXEf//AbhgVyG/ba
0/+Cc5UzghkEG1so/Y1AKtaLFucyCAPxNlMe+seDMVNLLlMBkyZYG7r7T5Oar57Gbjk+HIDcM5vw
ORp95zpaT0xQdGAGhs+yV60SMYrk6fK1T4X/lMkWrXIxo23RSoG+EGHnzURTp6AP6xYFr+LiNBTK
zcR034wSPZYFMVVhIVl2C5st5OMlCsCLIZVw2ny/P70u24BJUf2YQoL3ldNSxuWJ9L4XsQC6Af1c
JHkEQssmZBqBgApBN33YWCXg824v7IP8pymlJig2GrUQKBOiBNyvQennR9Ual3MLzRVawaNq/Dj3
xB/CHpimlyE7ANlj2Tff9Fx4js8pXD7qmKyEcUJCBO53Md1R5UANSCeRUHZElzmDubO//6v7yqe0
C9jfFBIGJ1l5MVbBuhOvw7Bh4j8dOPi49lX3PXoUMgMk/piE9i4LLefpSfwaqjUywK94UtNBPFP8
ZOM51Yy1lEn824jgs9p4E0qlCW3HSefCq0PPYoFK8VDWzSujhyOiJxxamxgFTAXg9jugF2pYYHGG
qpK4ClttQxPiyb7Uzk47S7muubzI5X9b6YxIJDl57HbsoTdvf31+nKuh1IUoc9V5T7Eis0oqtzy/
ai4wBqc9U4sQUTNHx078ojUcGuoqcemfrqC+pvCetBLIQbiKWHjNk1DRmDFs0ruprg4kGgsJ79Gc
fobOSvGBNSxY1lL20WMgI6MyGpSZ5gTjviznZbQuPgIyaqj98kmlzhEZQnfY7OJwiLKfygMpMwJ0
VGTwTQVWEyW7mXsyQSJw/pTbwHIMtEl1QYqMTqbVIVKn6hIroQYEARNY9TG67a46774TfZnC9tND
lNU+y3iTCEXH1rLK3SQ2Bwi0ipypJOMry3Mqc8j+74YgdkB6sxlY69J6FrVl7JFBOu04yHs6gERg
jGd2aB6WyYbehT5GjxxUpZIvcEVgxRPO3P1JSvn2je9qfyhKyVnbRKZZhRza8uzNYvFGSJQmlGZ1
RMhH+r6POPGm6EwHHhTIOxoY0DJhYL0wrHohGUGjt4DYMuWNCt3dcZlywzYtleWQu534e5BJrCx8
9i2LfvYT9bftD5wglfBU592fT0JSQe8hDKntqo0N1k3sX1pIdN1LHnSz9vb12uyQ/TW7/XOVGaes
5IpJx8ZbWnJfYdAz3RdCcSlODg90A74dbnp+hpLm/s7QdnDh9oYLbn/k5mEbEZDqssLeexTe04B0
NGF2aGNSA+pg3MPPecUYnVPVqvZ/V/zcuqahf+sBfuKre+6brkm/sz8u+SdqGHsjrm7LMi7KWWIE
fnmqauW3uC4T4fJI085aPhQDtbrnyoCUhSMwLKEG9KUyJnxmc2PA6IjXKJMVWGUUtoG+KWe4lZWS
HbB1HSgtiMlCbH4WUmBzJIpun5A5rG1is4Rs1A9l1Zg33v7pr2aWEpU7VyivSlXYD18NwwEKI1Il
xnlc48Ffleyq0XVmO4eEgQRnPoiBV3Om4RaRbWCEEa1eVBhsSBchN2d7OHO2Lg1euLvJuhrdxqFU
IwOsZ7jLPMoyYba6f/5ZsgwM4KZc41la07hPv3CEO3h5I/zFVMVa0J46MjvVRxhlqDZ6ZPTVM0UI
Cciaj2RKqh+knz2UCehCoSD35EMn0UkoTDHDR8MruCuh6G2OkAv2IPQpPClM/BjjFU9tVNjh4lxm
2weJ2YbLpFe5utYI+zXNPm9VQ0KqLG0IiG4W8myZV5oY2bxWBpL2vGD1v2zSTLWSDVYvUWWl3m1I
1FDVdACeGJpTd8pMDjdjkwwrp6/gDTECCHUC+Ukifcl+soWrIFs4qLa841DIu5+aWXKn00Dv4y6+
VvByUojLQ8yxllqWUGM0RuyCGy7RpU9PHla4aTFVruNi6T7OIfyYeOqzfHBZv8BiNK5plbXsd0w4
hCMT6HkYzrY0Uep+SwjjFHXFnMQ3c7bbBVYdMGGZ3JhFGymvSjpcEtoKJnlWoEv+eetBOey2KlKj
0AsbO4BaFvF8mj4SaRy+EZLJ5RprJHji2sUdzbahvpJI37bt33H/NJmkM1DmI3XzasGJhQydaS8P
qCImBgSydN4xaftZwYL1Akx1e3F6J59ceV4el28AgQre5eO12PlHKJ0pN+hfowR0YrqNyMdfrSkV
blZpokGeV8U4itVCzbXs39zynCGjyIPIcMb6fWyCV0Hrg+Rewou6Z/AV5us1NKJJjWtNabzW9/ce
Z6Df4hAmycsk7UePfj9V6YjJsY+7KzRr+2nfN/IwWBqdiFWA+tVAmhjd8sJs6CQIzYVE95k7vs3p
hpw5FZZgrca5vj0aVp2tdFOnHhhbNQwwoYH0diFrIiUOQNrKWAQX9/pzsTaUrGkme4PRXyR1ZXqS
tLF0UMMvUp0ulfPka8QvWbmrX3ATM8BYrp8sS6nGViVYOt8MejJ1xLQHlIlQs9Akjda5bSEAqUYp
8AnA7wbsxsnpv7D0w72l6rvN/+zfKcFrp1TGnHbYsorUS9RMdCCtKQSkBAvunRlchyLnvs74brmP
j77fjOhOYKNGwxmhjKetC6u6qXLGea+dvQ1R7+afP4wVjZPvWOei0oW+ghiiwhzXZyQEbBa/YGpm
CvHNrnLDakeIHch5ccxzVCbM7HMBfPeUT18rT+apuBDXcq2+dAhhwMLmzqKdr0VIHQia6tkHqcDU
UYLLb2gVp/Q0YoLuEDuGQNWQ5ISFaxln+5QFx5HZ56DIef6NMh7KXR8ZJBFbRUnvzvfHl/1FahB9
MeHJyxbuCxObXF23QsLlnCknIb/gEFeHx+2u6w6ySpoUwTtmqc6NnzLY4Axfd9sVF2c0TUNWPnnE
ooOpd3v0QGVOZHwh6ZjESeJicKoKitsrLutPYKEWU/Au6DIsRUkcQN2eZtCvlOC2ysUl6fwz1619
cLFSbr+6LQOokFA1U2zomcNJ+DXnycw4QKxAaW96fkHwYrChydX8Z1BppyqfeK3xvUfJprxHPAVE
buK+SN2HMgnl1t7sRU9oC3pCOtzY9bKU6cb9VogUTjZVjONrvAsQu6j130Ru5XJEBdr+fojhKKPy
4Tn7hOHAqQ7Kt6mZ3mAQSsRmEp50xX+hEaigjBFT37qOvsV7XKhZyBW3CO8/vWQryBt9M95qgyDd
sdggm2YR4owvgw3symi3ZZpkh/Df+e7S0NkNxn+sJVydTNameXq2tOyu90re5io3JIyBFB5RtcEN
VNPri0h3Pl22WAZIIgbVtY0MVdZnEt9BJHDEwR3+zUbZtQv/RvNBwUZhHJLnkALn+FYkMNDd/gr5
3ZAtB5phl+6sS3SrhJ5f9+5VaTq/0ctIYzTSlz8Wy/I+aTSDj7zbR473FTnzohM5DNIiQEQXbBNt
PqA9z6PzFibumh5Ljg8wD7Af7QmHV4EOXCPK6rZUuHnZknc1CjnqE375unPM1NtOOjgI1Qct2wM1
zXCqf+O/JINyZ6LaOt1qJ4pjc7+uFtS4DX1GG/o4mjYrqVIiybnY84dZ4IFMXY/STPE05b30zCiv
Z60PthwnyOUDdpS8VNUQithSf2G7SU0Cf+UXuPVkdYf+v1IIt2ApnsJsGFI6PQmJl5RID2BC44Q6
DUlf9flfdtLrg7vIZlXaBqqdSKTBJ0EGkgNDehEymcwABqog+n7gMT8pZOlssGc/mL7dVUSfj8IG
xBV4Jtmdxc36wgM1wblhsAonm6WNj1mNMRZ5FCIPWad5oxFNHRdHj522VDAp2GFmwLztMoxC5iJQ
T3Sp+IETlah19/3tVgv4bP5GMTXX/Y9S3zzNoOO2MOu7ZwnlR1uZSLAGbCUxT6BZ7WKJq+LsRQNa
mKK2HVFHssqrh+e5N2BWAGtMRoIfVS4skS4scKRVpeXVrVSP7/bXwlzcuUIMFDSevIeIeg+tOE3d
MulyLdNCcQYzqTaTR3tEjgEESnuxyK+kWtGT1sxrRBlFVzOcA7bDt1ZhPz49hOv4EFN6Cvcdj7ou
jiQf0LPKTqlo1zABVe5GkDBnyf1NBK9EgBR1L2UHRbSvWEUN+ZgRdPywXICMP6yVBgAV0SHfZZWb
8g1o63SvzDGNGK7z/8Pj3WHp4tTfc3wpXz6Xra5hxx2qefqhgOPCcaP0iwbpyu5/D5EYWokHTXx8
nyi3781Xyi7eHOd9lwsVmWhNGKFKcgaVbNpgCitiYF0KHEyA71QYCdVw0JzK4FRLl2FVpr8QYlem
vldZZw3taSy1RsqOkLfwA4sQLJch0kmn+bhXTXa6BE/G6dqFEApkLOqHFEea//dtTHeJGhqJDaGj
keGew/dMwwSIWDHqXo2/gSa0G4iXM+XbUJLBsRutjbPPNY40EH4VI2CMd07c3z2n+QoXMYbjBM8L
BnHIub1IJjNl4QWqGyXpS1BCZxcUyyotVnTWCecdwmydOmatt0sGXiycGH9KUhmKVjTvMu2RrjaO
V6BgP+FMFsVR0975ZIyuwaXo3CnPc5o2i7GtLpTvFq6q/WPPlorZ42iiwKy5UMVoTfFAxUU+KN0J
2jP6SHQp7tQFCdwmkeWKORQp7Iepfo66Fv9bvxTln6p4O8gaJUmaLa7OFIF6ztL/ImsNRQ4bBvEx
Kq6u/iCaoSjd2Fvt6XnQXLXzahGmfgn1XwT+gaqe4dW8gKA9qDnmJY9hEYv1Xz3evmi3Egm5eMe5
UPq2Kk3VN6hRlQ7ezyIxO1RDIjfzmIQZ4cTLU2jlAH1jfrWVlcniUIOkTb4jwFBwlfo/MjwbD+Jj
DUZwqcxnxLOANsu0rbjvJnyIyQcr7cRC1YRu7F/mH+y8PBUMIsAW+kqitZXjnoX7LzxmLygLyY9I
RMaZNvCBJipR9hdry4rV33TeVeUtj0jKftz4FR6fk+IDuXeTpwF5L9RFB7jf2egdOFye7UUaFQ2q
1bXsR6W7oYw5BU3eNnsMs1fZ5GeaM5R7A6hGjTOBhFfB7Pdnj7kXFfqI5twzWU1TmFWEpwL8qK30
WUEFPuoySeSHhV4axwfHeQG7A6IHWj1E8Jyavl6/DPL0wxAkgqwAb35A1DUnTVMgfh9DvsBIN133
b678oLjzwFWZ3SyOarJ/+HJW9wkEUJ7Nl2p5DMp4RU2v4bs65IRmVXccJ95J/27QXMXMjVyExE1l
ZDI6YRRR/RH+CHAHpiozR5E2uLViZr/zanZHSkow2TLQCKeBk9jUdWyARJLQcIox/8b766LSU0ht
aQLwyGmRalGgjo7Z+H/tOhdmDa0X1he/BpDIJVKWZwWblGNxoVMVjDeUuQCYnk6dSpgBi8wZ8YAU
T7GwWpXm2lIruNvQQJiwtjlprHXuNWmUyJmQIhKxYIoZIWfTF9/dOSR1ykyHjRk4xNvWo4U/UVyW
V6cLb57KjZbSySEgUer++0VietyoCtiRXrK7ck7lOIhKBU0lYwQ4VVKySMeSQFoWjycmO4ha6FJy
Ey0jYhc0xXr9zxpxcxOf7zcaCXFJ/8DSCreh08MbFoeYeQA07Guy/PBSg0U1H3dhtBAs9jv2HLZY
GdRDqYwtsqeUAxyF1sIl/JMvRB3azzjcAO+swJmWA2RSjzlIygNWqDZcaVgg1Pm4OzNVllXhhxbX
2sv8r/MMwjUWHjpg+tbX8GK1RSa6C+5EmZnh/e/5q0HJJk5M0WwTBuYpyweD+HaqQXxvZcNSW9ES
MAcTJ0E6ZqcCRebrbQGY8JP5XTE25meFfl8VafyLeXiw3lnS32S0JnFuZJUI2kGnW6wSmUtleAY1
n20AILWhw6Pc6keKBBUjsCbx3dtRpOxYADwaere7DVIPbzdiGtBD8UGE4mbm/fWSs4IhOeU+o6bX
75sQq7KJoSQoLz1BOgQpFYwGkqnohyW+6szsKV52GhV+s3qm7WLRma3LmddjsUcNZXzz1VQnhycy
f+HwbbKGEyFbwF1xbanXOodLrR69pM6mASMjscbBAoDCWeS4mwl/LyYliwbrA0HANoDEEc2wcCzx
s+wrGwum4GGa5Tuy+iIfjiaSm1KWohM12AJS6+1DMlBsSqyaZD6Oxlo/w2H6lR89D+Nz6oK2w4kq
x6j+LMHZRHfZyYL7LkGN3IwBpIcZuX8F8uu7T7xVe+Q7jgGqC/MIcUE+mI1TyrYgRquiAfndiUpR
Z9w8iCcSTpFMo7ivTi++LSd27+wtOMN5tWYuigbcJeVplRe0DLQBE9rrrV8t1xl7y58JmxaMd8i9
X8jPZXykdzaalXnh4Fgo7s0eQuU3UeCCjnk5ZvZGo4O/5AoLX1OuNFh0HqumjXFyMMwGD3GpaV1c
xaSsIn/A5zlnaWkUD6I71+z6ml9mY4uISeOIV4qU43XQabThWkP8u4zxWEYqOst6iYFfyakD0SzZ
1M6desktLSe4Znx64tIjVwLYFYSfI7X3SAD4n2hVS4PcIqiDuaASkG56t8Gip0flr8xo+DqUFNuc
KhCNr+HQFGiFE/fFPenRTR2Mj82JJ4V6oOX1TIosbtSrqpJFzWc/gpKMvZt4BlI5r2jUhSFvKuLQ
RhGbGnebi44en4ahL1u+ClQ7OMnlh6BZgk0yXlrY+5I1pcjYHXLqwtt6o9NbqIGyerfq6UuY8De+
jlcGWzXfC4Xl0l2s7QgJg8lOJSsygYT0og3FOE1gehKfXwEEvSYbv0/4Fwyuf+NXPXEvCHv9QXTs
PJuNDX3xCiYI6AE+uB9i+GiMRNoY2Xb9o2NjMpPXCesDdRC/aWAZqwzit81eX6aV6dC+sSOMLJO2
uAUSGKWGXsK1guRQmcawWD6ZLNqbpfq4Qp5mLZgBWkWi/4omUDMhVtkijDU2xTqGdyyGFJgPkgpK
hIiA2jDRXkE6ItOqTM9/5AKMAYNnxqjW0k05lnuslqETpALMOTKPm8DgpkPh4o6taRwL3N0equYW
BQOnoSVVgKSxhwyKoeVIzVuis1l2IAI1TR+anzJ2i1dvU5EN2AoMq4gut3FlJ6d1VUNCyg6OfNsW
1xAzwSeGATOTpBwurKh5YJPUXMMUvrOciAlYQUW8gr6DbMoLx1tZ3uVTsnnXuUvzo4ku8L2a3SJe
rbSLH9n4KawMGiLKoprZsQAqKb5Yx9nZYt+l+B0gpI4FLi+SNs8gkC5+zbxnXFbbkLp94DPRUyKQ
QYdF/Ql7sm/6Uz9PbTxxvwJ816NTLfHdDXT8klGYIrge6OPihkP0pZC/Hoi4WY8FCEkrysyHk7JW
56LDgWJ5zsFWeHoMT+cr4YUYdUK3RGam/1YXfqYqk2lZhdqg+r9KauWM94e5zhgnCUDzlOap7BiO
sQpNUteThoXgyn/a8Mg6/hNXtOEY+EqufR/0EEMHAqL8CSYwqrk6kqBJgqPuZoaDjbz6IDI6j4Pu
J8QxTKezqkk+ugLeqrfBaV2nBsi6JJGmlmlOLckglvmp4SyUhwit6Y9DU1dMhioIJpb5P78JrLTX
Rfaa1xfF2nRVqlp49+/8sV90bdf58rB+NBBH1vYSuSO0nC7J2MJ+2RH9tCP3VfFl0v/96cYOkOeH
Ft8fo7UWfhfW4Zgiv+YvO2LvCCLOvN2hQYco3/qReKJWGnPCWUiXybYhDeA4Wwu1jCFFwhAx4h6x
56Y3u/1XwjA5TxXqBXdu1mgyPyWm7QsbRLGGdAfd1lPcMywUBYh4g4OluwNEPGGZn0fifkT78fyf
FB3PqGeR2Rcx5JKy9iooS/7J4EdyW7YsMR7lkzhmJrgvWi+4TIVzofaF9QqRABIDQqfbAwhan2cc
DKyJc5Wpuq2cWO+OOJDW9+4TxoLKrBPS50c6WZV38JZAoBDz6yPXPvupOb3V6RJ20Okp36nXCzZ6
OfqIVvULOkPKJsUKx48lryqt+4H+vAV6SkDokW6UIVycZ26EqgkFYaM+jhRSsNp75/dFHGTjVuq6
+gVVfdY75ohscx4kqKT7RPTdaTamCsAGz6jQmUVTTd6mqCmdTyA/SXjj6lZfu7J1vQVZL4Ria9vM
9M3B/o0wluEKOIog/4i01OFu7byrKgWgB/uTn5fltinN7ee84drvLp1BvWqZ4bLnfZdypyIqEjFW
sp/aZeQaGLN3Gn/ftobkiIIrr2vly00ZicHkTXmG34BnsH5aCCtuv9dKM2jKHP1nGR2/TY/cNzsj
0VYg6/RhwRieHH2mmHIYZhWPzT3qpOyl3g5oaEsumWqAUnWLjMN4nIoT20wkKwpgQvQfI/++n1VL
U+7jMmGDmudabkmF2xbHC3lrDIYVUOzXovU8mh4T1V3YQYiiwsf+NMsZJ0qd/OZ6Bab9KD79Uv7q
gg8cn8ywk6XyGOoBaK1CiIOt0nKnabPJtgMk/LQe2h07zsVosGfjeNoejERD3hGQ+gfacX//DKl/
JPRflLoFrEtQmFj6E0e5NqAuYcKonLxC8mkBDmVwAMxnomP2U0gXkmO47zJdiKidZGGppIayeXpY
G3dJP5xMbYug1OyHtEybKyUykXsKl5YJNgBl/RowvMfKAKyIRVEtSST/LnmsAvFosdzEJ7wa0aul
vbKAGohlgILVr/ceRQ+WyNlyVIYBUUgJ7eGLcqGI9JSx1vYbtH5jEUAVfnDg17mB2disNKtM5cpK
oEtYs+MMMVO/CuLIRG010hd4f4gbnkXWFYxfP3EUl5pzaggqCIey9shVKZYlyvzeCdB4vVlEnTqK
ToY68zrKl5cPl6Jq17Rawlig10azaZ06325e78kHD6/V12g/w95E0s90fRkHL+LRjhOTiMikL0V5
9laeNBBuntDHsJu4v2JweqH3be+m0qb9vjBtPG5nCuigTCODQow324adGTH22m3HJ0wVLk6AImAU
CIAHrn705SjrXkprwk+wk4GLHPe25gNiHDN3abQ3BjnBbnmxDB8KUKdkfd2TqArYaXflYdeCEUUk
cukRBxVtrdYQDPSymOCga1W4nO0xWQVy2raiMwHWvkhYN9zV6KYfS3/ca1euR3rLjnaI0+g0pFEg
q1g8FTszMWfURrDz2lO8tqIxwTzS+hdaHMtmx2Y1ySCKwF9Fe4yiidYJSYY59qwr5oSa/nz9/v6o
I5yMMvMeaYUe0a5H4uHM+Atip6FqBUYrtJXtHGSZveTK3ay8p7U2ngE5oKO3xh5c0G2e+tSiTRz8
pqKbtdhMrtPIxzEPJMUChhi5scMe8eQoZSddWh6AZAoJNA4hlZHLAuLO2ysZyb0oSBkkM5W/4ubU
zKQ/hmZuEg9VEc2NiTtiO7Ji23MXn6zX2YEX4QTL+jp9QOBkZCibIIDD4sz+DHp8R1+K2JqjRqD3
dXSEMkLVqi/serKEiOIQaP6fGSvyKdOHeiUHl4xb8csPkgxq85hlxm/SV92eLVXuAkSluQnqRU1O
1dDQs+afunIk+fFx231PD+jqd+5WJTF+Ayy+bHMytHMxEqm4jN/DIGHHfrVJNPQrYPjPBbQsTEkX
K8lPofUxchJqRAsoe1ckPhlcGLIbMBzE+uOfFI22lfRFF4n9jbZmABM476Yo6ZHOkjRGKNfYD/sr
EedHBv52uhjIzJmeqFIMf24vMxFZPtqgNA1Zw398O+fCZ7BVlBpRwNXTL8knduTq1MiFau5zbciK
zcHz76EUfYWGaKjXLY0sdOSnS+5k+b7LpRMdW+BoPoP6ydUX8kB/IT3Fpx5ascLZZbzB2MVaPXZ/
W/+bAzi220q9+rAXrGP0xdvZE6Ou5D4uKSeLSXb9A0/+7ORj6AM/J/IVm4zsOiywT/xXA1Uc6/iI
es4nS0DLsimIAQykTbgFQ8SMFLoWqIRMBSqatQkSmYtWCLRUESxAgQq3CyafBt10tGh0z2ViHgsg
np+QSQEilnBTPDJNnIybVUPIQIDomjkujpeoXkx445vPWgACPXz//AcGXYBiIszzpJlcg6sLps9A
LXdNGQeDnOhQfjcJmbmS/ynapFoDRt1rHcckimgM3rKtyxtruQZs1A025vuJYriv2e4zYEivb95L
scAZUUSNVh4gPobVZtr/3jkfDvODqJ1mSujq+78OcnpOSG+wtYBSt6q5V6+rPNNg5M6KGH+2TXqt
ms0bP2yTC3BM0USESzvkMk+vna9MlNhuiljxFfOgAFmFbOnPheI4kdKWbkB1TOOjnDrbpatZSuMC
/P1q96JJvHbGvZR2Tx4Ns5OTQkWXgfLz3duWGgZkBaTarsbbnILPyFdCUO4PLnetFAK0rgikovK/
+vgH4MgbVTN83RWMxZCLkBySRrE6vFxJLJpqPj5AN1kWuVRgw+mon5/59wM9XWR5W8j7Otk1T0SI
nN2Kp6LsyVWIiBWgCbur/QK+n/ibM9+dsxwu4uE23jZgkhq2iaoEOdgRJ+a5/CJ6LuZ78PTK9oku
GSl/ETmHQxLkiZDd8ka/usrW9PpF
`protect end_protected
