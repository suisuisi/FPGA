`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SFpyA3WDAkH/h6gENMNzEC70V+GWX/AuJRjC9uuhJRzuSJx7LjCfMePfd14YnV5eJpUmzZ71W3kb
9tnOI6KXTg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FappTG7uNGFdZRwaHkH1xaFvi8BC2aKkPLd6PQ4xkTkeceiv05HkyC3+B1zcjatywH/Tgp5My5jL
RzYpXDHCiS+WLEnVqDpcElLtP6A/XLl3ajXqKvZhmMUVZsEI6d4wI3wE8drV6caY5dK99YnGiCxy
c/wD5JKxsx7IEFSu4qs=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LRNAkwpKrud10Lp0Eq/NqP5B49JnJU8WkULh5UDIksixm1tOfz3iui+8sx8gHS1R0x2iJMsSndD1
7xzPuxZn4a1eVkZa4n4EghKA1iQCL4jIUagjOF/A226osIvTkxPBVZ56YpbMiMwMMgRLER5z0xet
LPBfedO96PfexivUiLv1asz99hmC5fi5UUap1VwJdrnsIHsC0bEW3N+9FFvOSldno8glOl5txGSe
hOwrv3syYadhoBtySSxq9fjTH5UTCT6nikZqZkVb5yhHF7eaz/U8CnmNnm4+vrB5n+GG7KIVkI6G
7PqaCstXyxVZ0I0FOvUz/cqAZvJcffVN4NdFGA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1B6Vk0Eso+5EvY7kmrlz1476LggIIsaO8lHvFGJ+HKHly0lYN/LsIll2vy/lYtCwxTSlrDsJgNk
NtsXioC5DfcQQ4kEDu1f339J7HYisXvM7Lhemt1gBNgHhAmdUioIYx0fpzcnzuhwqs4zH51jdAXH
PU3S8K0B/J5Gty8ttFjVJwRIoxIqhWdYqBDiUuGzr/SoWf0A03jx+7IJtD5tY/voAJ5g3LhC8YQt
AWy8nfe7i7XNQN6Y3WxajBwMrXsrAH821hCM6aadbQ0v9Rva24HNcIHmfKUDspzFekOzU9yGfpW0
fWulISNFKBsu0+/BoJRhSZ+oJMcibfGGrXXNCQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ufS+qjgKdn2oE3oh7EcYzivo13DkHjOXZdvg+7gUZzbjFQGb+M3QU6lNcH0LrOEXll22KbI2ohfG
TzYR0mnCNIzsPfjq3uw6taFIWJM74+oLYtSXEeuY6ANmuCGlqaVPg2smc7PFDAPdH082wsWirRmd
5thR9q4u83J5L0asBhDI9ZTgri+q5MwrlbJ05yQiFPUliJgl6amNWt26C09sTCAwIMPW69iBKeeW
4vt5DSJ6XyglFS9MDI6DvF+Cy8vysZSNzc8P7lm9H64JZqo1p7yTgGY0TjifISAPXC1fHwrwfQXY
BsZz6suWdJqjyzpfb60JVTQ+/k5D70Xj1MXLQA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TI2B3m1FrAeKaU6k30ykyHfDnWZXVLw3GYVFmPwE7PU79Tu2R5dzZ8wRPsdfoPSTye6ipaIAsPtr
CwCMHFOrInoC4tES+00nqn8BAlNtkgIns4JutCAsylfO0tbo1jdQM1s3ZfLRmzO8TErqp7qh34cJ
cDScSpPoqwYzQG0FgIs=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pRy8ixMxliZyP9cGiEmLhkLpE8BPUs0NUJLS9EUfKEgqPIYh3TC0iGkIkNMUl3FvP77e0IxaktFA
/jqS+a9b+rZb/lQQUSJMP1pPdZyeKNO5EYTlJkeq4M/QPt/jHeYrB9fa/fTRWFaLSO4suMctHSMB
vZbG6s1wo4stlPecixWiLDS8vMBqt9xY7MLA6d9rFSok/TUkwwve+vf4FZtQpUFEhypIh+/V1Yj2
bwgtk5lfZpX3tS8eSCYcpYqNluL129jpVqEYjJIDkcuxvvuRJPiKMpRwiViOhJULCVRU7pAOu9+4
kiLxod5VBhsHJGbgGwc1XTZvGawHjedADbu7Tg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 124208)
`protect data_block
hA10iBF+ZRkqz9Fi3dOjxIpURLw12xqxgAtfe4my1asJH2ow9FYSvBGw2LD2L1bH4Ih3s5lRleLo
lqPuvD2LcWvhBX9LtKTv2GERHH90Q8dQJPq2g3WwFBDsp9IJMpVirpFA/CMTZnIWZ3hnw3Ckf8v1
9mKO6Apbz3XZRA5tzTlWX6K40qw0+UKXXLti5FITwKfg7GfJfPp+sqJ+kGQCS4rOb8ymySiDsxH7
7g5DKiiS4G3GGTDvAPU6Uh6Xd5hid9AixlXhMI5ld5l1OdpgitoqNb2n9dE75S+j2/qKTKfxsQ/e
F7zwHMqkjwZh6ZYPaXo/4pLPSjGEJYizDio0Pye5E9uLVABmzKI8uSBRsaWL+P7lmeNIq/5BZHYm
QiAGAWxcAQs/V5q4KqyVA1qT7WTw1yYyri/WIPArobYpbYfdD4kwVkrcmUK8fmYS9lJKhxAtnFSB
Ysi9Ko6RWWA71CFA/Xz1iTV5V9J32XOKzCOfA23ZO4vlJYbNjcjutH/KE8sZfFVBQ72SoTDsNEmj
jXQygX2d5Pqy+UwD5+ZxxXEK01I7kc+ISDtenqqxAQyBk6xfZDOabFMleYsAYGpBpuMovepZVa/c
XeCtvi8OkppxZJjAr1Vx+APqbZDvKK0ygkZTL3wQ6dEpWbYn2FqmXC84LJYk3hi1WQnPYUTvXKez
57qB6FC+aypaVmogdQiinO92GNPflSfT/68eMnEKv/2p2mSF0c7ipE5k+L7ewmnEWgsspQjDCFlY
ux9yjvnIcCWtO17CdKAJ+ORXOM/GiwLbKoMf5uulnbkkfsEd0RyYkbFbdqW6zL38yBios3Ro8lYQ
/JJW1PEWDwVc2HK5KjMHXRhSqgbOpDb2hc3LkXPGIeNcVUNSy9MjDwMZdkdV5I7ig9EwV49xG+3P
qH9Kjm2fh4DwaWNy8LFPNrYlufQkwf+T03C/LsTSA5lvpIE4JXvbelfJJvEmZSGClWIWkHTFFWpq
2emV9ioSMJT4UPWUSGVa/pBunGD28BKKZwWJNFXHj13zWIAgXQyREC3Ube5uD/NY4l2Q05oHmqvO
6j/fR9/JQAZ4vn1CXDRyzejmEVCOpv7BajrIF0VaQme0S8/zTovPeyHxaW2IgWhP5TCqpGhyMTfv
Z7ce4s3OVyEO4nlnIEhQo/3d9sEQlIKTo3wwnm+pwJ9ZUSKDOTcs0pVlr42BS4GAaBgKFa3hUlTp
pbzeUyHsS/MEXYedFHu+ZytrTrT4JiM9vTQ9HigWHVfg79oFI7J7pvQ4lOHVh3aZhlsXSS01AFbp
Bd293+OK2rgK2+kRNXdFKiNLDR8LR47pw3wf29C0hU1zy2iBcr+PCdVE0UJwdlP1K7C5mWn40pe2
xBlGTRezpEXHNsJgoGMVOfM6myEv+h4ihS6lrkoRmF243TW97BcDf4ThNq05oQe5CWuC/M0Momuf
ggaKhgPS4l5cf58Ggfwht2btmR78l7GaZPMiMlOPvPfzLp7/6SynY1NBxvC9RNqceDcqGo9rvEjN
6T+++8V9EmM2iH+61EictvGWH0Nd94G76Tao7iUygWqt5K+0aYCL4UxnPmoVb1oHX7Gg3/5OjJ2Q
KAIumlZtVIOCuiOKY2tNctb+HM07IeREB3TSZ0CB4nnZeDrPxAAxck//xrNaM3tg00/MPzGk/7ig
DOgjmeTdMEI1CGtgekyQfWty+qXBpvByLwpiXjAdJXs6c79BW3h8J/hkf9fShk7ubBD3NgrA0uqU
ghnB2Z0B5rvkt75bAvCmcKHCrOFy+KZB1trwIZEUTTusmVWY7k6zmC/gLcyCpxaS2JK6a9LnHXpb
Wfm7vxIKcirtfX/H16skyBp8lr/UWR3M96LF++nL0AQVogOAsZL1Hzyq92q1obU7DiTsH/CkTQac
KWvk4NPmieWvcMv+h7jIUGxOefPwFhSjWjtVrc2lfSU9JykZwomH0X/BnlOCUxQlElapX6wWbTPI
Zlbjcifg+JDQiTL4ic2mXJ3qWvp1OWhjDZSBXdqEXb1nw3BxtKb+n8r0WTQ6wF9OMYCKdfwkK080
jb3IQcCtrLUoClm1fvZ16DwrZfcwi8g0sc2b6VLKu4VbmravWg6DuvX9pEneY2Zxd5vEmuVu1EYm
IAIg3kFLXPHr0oRmaaxH1B/zUoda/JhcDcfrB17TcuKdLP6HQHqou2cdqPjT8RlMPay13Gzb2KiR
4wrr3V1xF5ur6+OuyJL3qhCsFJTyixl5TGaciPSZ4RB9FfkeicUN3df+tXXSeOc4dpXw6IvvWxUY
aIo/MIK8M/N9Ha3zqxBTXN/KF3RNf5w5++24mnzeHxNLcpZUOYuximC9pSxY1thsamJ2vR9+k8Ex
pbWxAR9jKcAEyWIrHe0V9xw/uaZWKIKNOzqcT3mkmnIZC+Zf6FR/CJ1NeyqckjN/ceXD2Z0v+/1H
PRXlVIANIc1Ey4g/DFTgn2q6BisWzGkbr/Sn5QreaY1adroxXsbDBZBmDnvShKIaR3WFIqBs9Isb
BKKwpxCc1KVKrAuVxXnfrtfFVbLQa4yGQJxUra4iBG0d/fyaALFQ95xDoDrFC6ME/ZZkGJVL4wF1
fLpikEIFrzYnCyq9i5l+E+D1edh3LHUpLe4E1R7/tumiq9SISXal2Mk4j85M2EYNqnLWCCZEmXVr
loY5CkW9hjYbM3lSyxRGEzc4+liBYPGfnvkceznFwjW0y9wDthDL0gy4mkjam0oH00HBLsjcVb5r
pzrzjqeSbtZNT5cGnn/QSqeecsvBot9YbCihIZiwsbvSupaY3HFMJ4husNzhzJNA5Mf/ZU+Uc4ys
CARIFOURgO+V3L1rN7goHSpKGwEvGiV2FL9xtKIeok7IBSmAB8/LA0FWSUPqJGiILr3OCtvJ/Zt9
STk6vW6CcZzX5NWEqHGEyHpmkI7MpS/29aBQRu8iVsNlEZdTln4a0YmGQra8vcdTfJS8NigA/KHl
8y8yDm8boOn7X6tM+tl51zRIDXRpTRIYMGvI9xX+W6nksBOJIMXJZ2DKi1eSuYIezPALONRA1nGw
BmH+EwZIct1RR3w6QQEhtLjvpAMyXpBx/S33CKmX9hEf4T56bEPMgpOlfUnT1mEGs1CmSRUb5QNr
UwYBea3Tj7zQfpB7y50+zJjETd8AzjhqK6W1KGnrlUQDqpP0di8YGV9lJqQJjIY+YnTZgz921TRN
J8DFAtr+HzHtZ12Qg3uIJOHwUL2FYsDYMQR4scWVnfa4oi3dGioyPIsPsjvKtrpSRrkXEz8tL7cj
Or+bgmgGOH3Nr4KUgW6Y4x8wf8K5aluSMgdMQkKOQsPMUln/JFVmTt8xxIKY0Uj9+5o3uNsqiO01
hPGiGSRu8A50mj9WB7q1hHsIbNsSi8B1A5TQotyugaKuhp+LPzTXPKbR3kcl3j7W6vlBW0R0DkI1
ItGzQx2GIoj+1DBePkBrNk9hSobNgxlgtywkfrW69+P3ZpP0zfoMcbb+KdSOiYi2QfT6H+nxl3sr
QWVshCmOuHvoqB7b1+FDPOfCR4ly7b2soz5T2M52tlVh4Qq3E5owaePEFhLau18fdTWzI/n07kA/
tb9lxEu80tEElQYkVow4N2jAlj3697GKZZM2j5W8D9s197dv74FDKozefbvx11f4tvBiFa+KivRS
yX66XPHsZVXmWYtxaBuBA1M9u7/gjYgTv4/LbtXdiflrhszNXzDdk2Vu3juUBMQYT9XJrh0/WIos
/ORKeNPvRgZXIhUv2O4ePktxGU+AuFQ39qZUKMXxzn3T0TccNU3AKv6vwZ0mRUVrPOm4NndsqMlX
HeID6GPOnl9joAezUxQT/LsN28T/8kOqDYyQhsJaPsDSfrdWX3i/iPxg6nPzcHmr/RplinhnmboD
HObLyJPGGWPPd1R1CmtcmL8rfqox3wt8y/z+Ps3jFBPFt3QiqJY4AlawE09D16vL3gT/lEFmrVpR
OMrwsE9R/0Iw3c3FRIhpo2wtkd9cYdW/m38/5VoQcjZtc1uUjUeqxL3u3IxzTipHxNt63x0axBkd
R7oMTOze5ONmleZV1Ee4yFgEuzIoKu5iVBiBO7MthKg8ooDNSLZvBcr5k2RtytXDMpwQoHFcID9R
sVd0zeowItK731w8SrLkU2VQRMeNcW14fKeWtkOBr5Bi7hYxSo+iRtZ4P3TbH0vZfVS0QhWPywO3
VNhFVHLcYl8ws78Db9RJJcbJpHrRWk3Ejxfqbf1DWseASx8qhvwNonpfRW3e1qjgseLx0NKlcqf1
8t+ISEOyZNGXPhKFlrSeu6xVnJiFqLll8433rEdRuRXII7wUWpVIRaLNLpx+Yzhdx2GFRARGYugn
Mc4g4o+KjmcaQu3TYZ+cHSjqtXsYF+/0v2vtoAe2qDR9Y0Or5j01yQ3Z6fVO0pZ26X8zK37FUbK1
+CvgqyWFW4PQE2Jxf9ESgZdCC+c2WeipZgH1EIXJGqJkvvQQQnpFrPyJqO6GkyMaFXF7FbxslTHu
CAdeKCTo091zn2XE8+ZF1hoH5p+FDZ+rOmtwyz2WufJEJALmo41SrtzR+95ynpymvMJ6bM1eLvjj
eXq0/rG+lnPN/o6lyFWLRh916i9eZIfb+DlUzyBAnidyawFlumisgxG6ScjtAXM9JWFVHqKveM54
XBIcVPnT1B8qfOzZgp06fqhgIixE8Q2bvdtsMNdmXY4UYwwJ8L3PrB8h7ISCBOaZO2VmQ1l6nwy4
fdY6oB9dpCeLFQ9GCi5uV8u5anyz5SlDaFZFfuvVOhEM45DaDf6RidZ3jlJbc8+liFHAI9OqTucY
coa7OlBL6hYCSL2wl3IOyN6tlxkKv2ArJUgO2av0cW4yy0T/feUddEcLjIu0W8O18Km75wCzP7SU
42/ll+ZoECZc0GEXWLNgwTB4GQjYNw97l48TTY9+1CwY+OOBeFM+nEn55iB7YnLyZ5Nziftyq93g
zyxdbiQL9L2rCXS1bLd7PIEvo3s90AEfbxu+jMkLvzUP7o2/DA7H01XBhnmHhCFNVqxvR67LcmxK
yErg2Zd5/MLEQ0qlGXJ8EyxdfeqyW/WLmB22LnviJtywd3PsnI2frH4yrGiNThzQ+/47lmRnAXye
cLU8koI8l+6aLPt5P+M0Q7b7sSyl3Je6mUx0+kDxw3AM0Z0q3NzWddYt8qR29rfEiUB2SSegeaao
yXvn/h4CiogAAPo7YHAzwpalrFMO/Wzlt8Tc8sBeLCIqwn14xxnhg0IsRuPOk6sZkV/aKXk9J2wz
cpRZCxeQ1eo/c5YxPaGk6tHv0l4SpeG/Ym2W8ppU4OmaqpBHfOvTJEhqSPNUPR78+bMFhKuEN0T6
VV5rDLf/2HA2p60c9cGQhUxfjYoxxzgiwz1p33jnd/DjdscEa4FuOTd+A13ZhvSBjJ+r/VuJWfgR
izlnXwpU9RJTjw+LbYIPEYnVrmmxUwVB29nDVMXZgqrahsWCnvUZr9WrLemXl/qS8trFrOFWh9VD
VoU8ZvtoxYzyWWnPwY2TOr7AZ1VQOmBTmL2riS9nU5w2SOHkR8pT6FrJ6nQheHTJMfxKCLPgGdyD
8I+sDRPG9vQyKcuhJ+w/oBSt8sNPIxzIGHVrAyFG1DLTKJVAnyK2yKKG+F0R5aDfCkSX30xzy1ry
CtpvMos3GKyfmtNCTVYKNv89mmBdrHCIpIZGodJB5NbmwFY8yLq8XDBM4luIWk/LK1k/90T3tK95
tTazG2MmBjnvCWOvrQgYUi3TwusW4LevLaN5kKPp0U+iMaSTVzFzpGyPr8UyhMIlEzAoT300mpGB
Yck03DVi0/JL5RK5VifJQn5MKFPtDPz/Gtf4I9KzOC1aemcl+boZJOghvb21YpB/71554P/i0CMU
cXT0Vb9U6/lRAneZv7jBw2eTtl+3Ff/kQzxjtkyM6w3nXHPyxdYnl0L45tyBpNKs3WVq02nAjwES
tjqSnwfID3NGfrc8ZOev4q25rfvigPfdsHhUzTwaghz2v9CIJLpv7WRpdt/pXlBEuWqFCl50PvYS
XyPtwq8OMJGzaJzEil5ojp0P6c3tLpZZPXE8jiwfmmTOZffV24ABcXV3fngnEXKnbmq3MSlvgZbQ
oj3hsUQOZsAQi6IdU18a+7m7B5FnbTXe+ENy+h0YdKcqU2UanfXps7o+wyZnO3uXHn4/DwWKgqFN
3KIB0T6oVpfuwPd5Ff9dxH1OB+zh2A6UGtR9OKjB2vMuWX3JNbS2ifcp2xyRtLu6oknRzmy2JKbi
UFQojUXbwCuUVDVPNwuLRcpmj1eiZYk2DtaqhVR8MN7QpeRwxPBIExo98ncO5HZPrLUee4wbbziP
2C7u2UQtcMSOhmhmz1soc9ZnMWh62fsKuanxpeJ/wIhleE4THvuKW7WjVur20wRfR1LG47oIgbuO
NoQ1hgCn2EvgbeSA9idgOKS3pZ1SpD9YrAYV0c+M59te7JDH3D8gvx8WXQkdRIuXVxiQ5LoY4TZy
e603Bf40ZYnCCJTO0IrkfwtRjkvD8y56OLqNeuSc8gFv7hBxKKT+i7ywmr82NcVuqmSuEq417n6a
X8TDJEd8zzyrfq5TQeSLeim2KDJ2Kv3UXJkKdVJBmnu8yyvezNr1ylYdEkbVxS9hywxz/TQi39X7
H4fR/beSbfvGQKuixIp8q2tceIEzYhKpcjzpuYf7eohnM+/RZNzwW8xPwMXorwxyLPkoDYTt3UuS
cGG7hyZTEj4FvgQp7WfeTr5uoPd4ZHiUqqebo5Fvxnv65GVDlko4mqf9p26AMjdDCOrx6MCwjHcf
fT8nFC18TounzJco6aVP/gRhsJ+a7s/RpPT9RfTT2PKJAwKKHm+/bAkPCsOwpY4bTQyf831Rq1LA
12kOuXGrkFPm+zmibbgVlI41TMSlsfbYvfeLhYYtUwtObguU534zVePq2AafZ5PK2mFqEwlKkRG2
6jZ3Ob4HJhSJy7KYe6ZboWUtewBEmauxSXVuW1sKHd8nTrhBwHSwv1s+nw+/TCX4HNO4WDvsdoc9
kdxGZ7C8Gg4l+hI1x0qZ4CXxUzzQbyDFTjFf3M/3LAKY5RZjp7IBZySLaEfwEggQ23NtGzG/6t5b
nlyF7Yszugoa9C7AJ9v3eEQX7QE+Wc0ybgnm6njRY34XBxonmPKWS8BFctXt02NsV1jDVZGWUPkm
pdAjmSd6leObckno+1f+uCOETg9OD4QpWvQdfAFPTf4MTrfepTngaL91vd8TemFz1/62ptGmVblV
ve+WjTQuXnPaJG3IYZ6oB85taDh4Y69eaaoqmJgNl7bCN2MS+6tFLxbjLSEnQbHRHSmGw7uCMhRu
NXPi0NqLdUzKb2LKtB8hqXHaAMDCZGM8RM63W7S+43RclR29AamAXGE5ad8ORi+qcqdYIWMfNHBb
aEH22Kx4fLXojKYeyWtfX58WUl1o6/AFVaBsSCkEl/57xe6FGO4eX6inSchefvfbFei3gCxSTt8C
fo1Hb/5S3T36mIW8XCU2cWuH/tgwlf3Qxn9G28grJfnDkXj0Ax0287NpmMsQndY8STADPkT84MD7
pgsx4Z/RwMFPw7Y/86LNePM+27WwHU7P0BEcGFrkp1eInaPrY2zN7ysLq8WoB5hkIuOBiLtEOIwZ
lJRNVA+x7ko1Chy9ISXJn9y06/qNqIhITf0sK0MhO8c4ryotmXMEFlibmWi/lzJqrWLBV8Wep70S
2ole4VgupqIcJoixPptmvdx6VrO0q5vyyGl/dWCXO0cWLFzvCCn59wfMQQX1LhsfZ7OjJLXtkNZx
rDYqyrKLiWG7USFaAmXb6mHAelg3Th0MBr27fD7ZUTzvjEzo8kOxpDeX8XUjqMWoY2gMgZeqakQN
fgRO9elbExOwFcoerfvES5mwsNPkdAV+382woijQ8goLUH8tTReRQ1wUc/qUrgdiII7bBxdEXTtR
DDPfMNz2c7Ub6H2WEKztjcU1Vnl0TMTI+vsfNvIglhgf4CyYIC3n9U5s5CoUTyMBrczbdDpGFa1u
Lp04ctN1ShkNFH7+1OmlFnuLFSbBX6Go6n88GG+hofmpC9QsbzTWR7cSTdDCnQ7jg4Mu46jE22r5
lAu/YEtnKYWvFD05JtDgBa7QglyHCHeBjfmqmJ0BwHpdD+1WilwG3flAIV4sX+ic5WjprBIF2bbG
0F7VRjMY3rlYUsvKK/hY/JdTOL11O75Y4KL/1he21WXSNOYb/jmQIrnmV/4xMB1ZkzsqThAQIUP2
3/n7A316oqMhXMhb+xj00w2iyhl0c30x9949nbDSn1+jL0zhZpT+Hdbfc2WSkYzreobJMX/2oQHn
y9FcBIwoLVdkhFSoWH3pKRun5S5s2QNM+8lVyX2+1vAsBc0T0oRU4NF66Lz+Unny+P7++0Y/gOyX
X1FL2y6POYvRIRuCDIAwlSrvt9BuPIiZ7hlD5cg7ID9F34vR/CFRXryLsr0XchwJgtYJK4KC0u5e
r7+HTsWvS81cLZefVxholU1izzdqAcRTDNu16gxo8VP+JWe2bEAPECdLpvsrHm9Zeuh29LfvyCNH
xl/XsUdY6nb0Pj+RxBVG63XctZ78ZGsDzhs3AiojYycNpzUFVHcX5k3yLtmR6ckBogo65+Nkl2Az
OmTVY2Cyo7dEDSrGQEQj66889GbF4NQD2uAZv2Lt/emxIcmSiSEKjdhznQv4tfiP0spLhv5zNQNj
s34VqBqzyQ1eyijsjjV1jnkf0rlluqEXDC4zm1eXziFc4ObqWUUY1e8yRASHjMqjGn9BGl7CQI7O
nqBV/0MrqEOAlEzzX2XeiJsesew1TpaWyHoIjk47V0YthzDkUWU1fFhjKyyW59SIoGH0voWlNWLr
+fC4lHagJ6TFgVlXrPZ+v/wI4R/VKF37fkB0qRvPPtnCq4MnUPErQj6pk2Nsnl3EvRroe5YDHAQt
5lwyQl9FZbdCmCvEx0KZsmCtnNcRNc12fEbp2KPZdG16elt8m5wZ+/EImegQdeIboDJgS9y+2aiP
VBHcbV+qWxKU5zH203trHXyqFzrO20w16JeGKqnIPdltzmK2RxtSLDEyGKz2zpJL6RBSKeKAWvL6
jtMhj8PC9II7H9snq9CSkOYV8tHQlOQb5ZuFtl9Dyrz6SOlwiyTgJ10XCE69mk6oCpSuBgfpW6lx
Do41ZrFavOXWm9WeXu2n2v0I0OW9o+YRfUwQIUQ659b5pvQMhLjDz1vc+iNGLQzlKJaT56JEtSV8
g+MlD8/CmFBLHBvw9WG6/GsWV+pKm9Uz+bIN2wPXf//Vc3k5PXULLvx3U079WmF54CwOaolzK9HX
6VJmTsRFyiClG+uNhKxiLKpY+EcbqIMYh4N9+ywYJb2zUEPe+lbztrPmei5tl8unUeJx+oW2hHsS
qxgUozmcYZ7sVW3Bh/9qtNKGEq3pOFwl5t7QhlHymWznfw/p5JaUxRPG9SDNWNlKFxrCqI0eUrd7
33dgq9DCTnYKI7Oo7R/1D+nPBN6PuSs2hZgvH0wvnS16HRXMnCXCgUSjQSAB4SogCuwWSMvwkaz3
YEK1GJJ0lWdDax6N9eHcSR0PCFMjIvhpXdwb4f5jamIOFHSQVxwvDAKMbrpV9HHPY8Q2q9LfmIkj
kab/4mgygH0qKorO/IobQ9F3qd/l4USmTJRpTNPLdL6u1m0STYdj7WPmM6G/bnQr5tEJ8EMPkQa9
2pBLDzQv8/7SPAx1SBWMHx4ybs2OHMFKNaeeM6vU8t4hhrX8usGrExtfdkxpB8zMG6iU4AIwDfg8
68bahFrv5lBb9NRC0tLaqlYocaL2xqFuhtxqNHYXGLDm5wXrWAQ/PVPOn+aYGkllKAAltFyEBWty
N0S3sYg7XpqP+fUT+9icDPCdTOMtovQDcKjINiolCVa2aW29OsQWF7dI2wODbTGXV8hiYB3qxn8t
GqPLHUjFqiW5oSysWKEvT+kulxZf9tIXcXD9r2pdkoHDnOkWaf3MuNtlTnsSMUAbGPdyGonWubwn
19ZV17H0zPxMaSp30vUon6I+6SVs0ECbAGs2SAWu8ALbNdMePOwbOsxqj6wPzz6jPgOx/Stb92xG
bee7fwguvhfdQHeOcvC5L+Y5zCWR9OzcLk5+Tm1hu/+MElq63M/IXR/3usAljxZ5OJMF5WC8VZ/g
Mv3Tae/w+66OwIBoPz970sVsFBDDbtf3ac0oQNhJ3X4Gd1nplY/kbFYCRo44H3CeNB1EfSXtSzeS
w9B5RALcfofgaHs1GccpcOoVpBsFp6o7mAIC9J5nG7eJDJgy5hpD3oM5WkkcJ6KWTfVQX3mmsG8J
1D+GLrhSh2SFMUMlQxs6XoZEbPFaauqxSbGk/Wn/6aEAVDbM50hl5wxy2GMLB8ltSriGzlP/tcke
EYIZi0czxhnpc3MRCB26FXUSmN+9gVznPleapZknpM8DiWDKfXaRuSybzgBceBl54yAKimYtFVqt
96MoY5lPHq9DyUjYWVVijnhxobZzO3axAh9KuNxFibDfCC0CQ+epsPGTheLHYcIj44f0AUVmouHE
QIimRUe4KRSJC9A4XEGgS3NyYPzgpaSr0FJYL8PBr3kXb7ogW2LjUzTUnsQM8+Bn1nZP53J5Hl4F
UPhOzANVnP/xSgb5bOtbjmh5psemeiZRkYlVfxXU4fTMgqksS4YV5mV0s7iXdH7XxYZpByF1X4Fu
h8wXlHmZijSZDEpdAAjFcW58ZDFl1dvQGzW87hOZchHIvPIasnUQ4SWpVp8cnYqAZyJTVRo7YDyX
nAS2CtJgLNJeNx1B2xKrFfYhkQcaInpsJ6G8DGuYHVY0enasqQ0Y/cT2Mdu+CPSm2QY99GDCiYgV
J56cBXkPfjPmORlvXcVf20VbiSWqDqiA7aLRYiOp9fQkX0XXyy1/92NPX3DRZYExrcuIuFZZdnyh
2u1PecHDnRmcnCuZ1yYSGdELoV3eC8b3qCBjFVGu6kX4qj8zLzVXMel83nguccKCLaA+ULqr6BT+
1H8WLicKHOEwSHFwv/rUjU1rnpdimunwKSkx0HfdSA/aDIBZDvtEs/LoLwW03PPSUj+KlHY00eaG
xYBGTTK6mpZJgoThlMEkeP/w8D4lc7nofWo7ImQ0EtQfLs6fYgguF6T5/LnQjMvhP+bOu1OBKttQ
cpWsHQjgoHLOzFZSmq+fUNpSDR/MDURiu1pQoZZFHHJC9fEwaKdb6Wi9P1VgjQYSjyu/hCzEIQgx
V4SoPik5ldu4vKZBh+QeVVGUFRMB3ZKwgFbbijPDMi43LePr2q+Ft6lJUllgrA5yg63Fk293DqmT
rI9sA0O9s5kI+OYg7tZOjkAxHt2oPzWupvuJMSsmzRZjJeS9081eXFt/6M1uwOBs4YwtTqPsDyfz
DFT1gIdfrIBbUhqC/ZbdCSDbMM/5ARPCDRIxrfNqsqwWNl3rFrsOmO9+KzWmhuxehe0LaKCS21JV
LWgqx+Rn0LIfzNZcTl0m0YcYBZo9jk/s9lntcWBpSX+wsbPv0wIUctiKTXENUZJjNr8VaYVofmPq
9KT4u4JR3S5M3CWMWYN/2NA/1Fte+jHGK4PCkEi/hdT9UvRIUdDZxJz3Zt7lniOI0kqQ9ulScVq8
KHB9WU5bapOOJyZUHGEgS5Zr7Nvi3bPT3sfvZXI8wXsF1tq2I+DJnQnYQp/lO1a+PqG38WWoSQZI
ZTi8mb3q3EEpnMrEz/wDFBf0es+NZy6/0823ck/QIxrGGRhu2U1bn1lU3b7kECB4x0tTjvjNMB4C
UUnCopyJ/b+lCx7zWoSwjVUVhyT0T0s/L0JbxR2A9Dj1Lks0kzbrX2pYP6TGcl02w9abVIG9QzfY
4zibl/yg0CiKBpf4SHhr2SU1udrCIj0nXu8D6HoFO636q9RmQiKqLOlM6eKhklC+QNfSyjHhILFR
TQ5z+Wf0vkRL9/PGY8zgT+Vj1DfBZRpUgJfdpHtgbeRy5Ihi+xR9tRfXphMYIHPUZkh+cJcluTnD
/FN50AkIf8XNiWIZcCCWmtdwYJ16uFRAS++Kg5bBuatVuD2+fhMxho9BEqNsCFYA++xEiyQmh9X8
T6FECzs/8WzswmUN5Bx/YtqC2Q5UCLRGKlLLO6Y6G782Xb/onUNo7PDZZf+S1pNHJIU3brHzakyD
sSLB14OtUM1XCPKtZ8Ee3LoBUzmdHxOHvpBfElahUnz0smH9LadazMLd36CGOBDjnrIwa9tG2YAA
YKldRVSvG0tlEfC2fHdqJoDGTMC4IHEgRFYXfOJE5/QaVWFjYrws+G0/3lzXju8GrBOgvFFVBQ9R
oHhuel0IMU94shL8td1e2JUdcIna/BEaj1wFnzjrJWfyw7IisWdRIWf29QgJQcPqlgNh2BwV6Yxw
PiMcfhktQJhZpd09ntrtZ24MhqoaHAnkiPDu4tmzmjcIznFp50vjRYJagNBiv7HjPCdCNJxIaw5W
4yxqc8+qU0/YYHTa5yqg12h67P2xgulVretCTGZDPqqVuWu/dMJ/mnjcVHlq6YzeYKZ0rUkqp2pb
QILy6pKjlhG5O7VpKDq5A06qLI1j9fAmPbRYrwN4LYkkpyVIZCwPjJRL6bpWFpgk+mNrP75jOc6q
hJ6nQw+YRjiT9dTDde++VgjrV70MnP24TK7uKxddgpNPNnxvW3v3aRImd66lqwUOBjRB3yuiHkV/
cKeeBFDkYiumKwkUbet57TVfpt6JuepmBiCvnmLE0JhQgQC0t9AG7ZC9VOHV0Me6moIlmJWIwdtc
SZLiGuCyVoMzEntJff6qQnQL+Mq03lA5sVpkqd/l7l9HA+7dmNLqrI4dCvFqVv5xp2X+FM0r2kpN
BrgBYimSA9l7HqHJOze1ieIRXTMdLz1eWxwohQBB8vqW8X2J9R9k5I6jhc4Q7/GaNYttciioBvHa
maezNASlkXj33CkD9H7JsfT5GZR+sav2ykjNXDEYbZl5JLi2xD9nRn1jyBJKSp8UCld0O+KX2Rxb
RWOci5oqPD1Ndbjk0i1BOtBSe4CWIe5fVKaS8iIYuE2wwPoLS2BYiAvgrr/ydD1lh1QrtvEA8Hlz
5eM7PVz81wiTfOxD5tVWttv3f+2IC91DP/cKq3wIcKtXNDTlZosUlvvzCCQhuTSiDvEI5mUsmsFk
du/88Rlykxz6rMdc1zsmWZVQvJG1KjXzHHqTf0JXFv/u4RLCCpGCFaM317RFkB/twmgiIMq9gmgL
8kQhKQ/U98E68JPJJDPQr7NVnlDAdrUZnO+zzAgLHxkFX+s7u1b6eQG/2Q71d2oDWafG7qESjwsC
9d6BwtKVMTCLuLJeo0GmjCWY4deu9afFNnvB/kjipX96+dotEQZEzKaICsk+iaQuVbxNrQwAY6tZ
mnMJuWVBa7irJOxrCiSYCTDls/G3vd5kq82ofnhvOU8v39hx+KddaZeGvQJuAjGQSYo9I97IX3ZF
CuA+7emWy3sAWErOTAKYgxHwZHie7cVfHMwGj66+806f+buP7uVqIuSK0BV7ZQsGXB4TZIaLoP7n
rxkUIYVPBaFq9uUgTydmQbXkd47ytY77SPKak6MheXF27aEf4E9rfx7SHuEhC/YFBXjeEqua/dDq
dcdYBqCfTfLPQ3fE25qIQYc59zDDjZz6cQkg2CJ7L71SIb9zWWVJ3PGyIw5V+xAeMmT+vngKGIb5
mb1/kpEUFBFpeCKG2t7Gt/tyMcJn0mGvmsn6KqiBbsW8isrkVdKMITwHt8CPgmTNmNHKqnMo/Raa
KZEjcH7Z/x7MJFsMrvetd4bSafSjTNne4jPhyav3DYOeWTONJn4Y5bV6yQd5WVY2T7vUb1iS/ota
pCn5m51MGBP7iTbIcRZMGUuXSDBGERl0Emw+zuwLQOFsAZl43YcsC7/Bq9xfpMrkGd9oV7x5Vbl7
z/bsRgNI8//7k5ET8XUwMSQjJiKVEeGM9SAKGsj9VWIpuJU/b2f8AQCrPCMG7LPDKB3fPvr7kiy5
DXIzR/cXxrx2q6WtPsgkaIkc9XplgTg7UNRmiKi4LAEVgos0UbtnhGf3+OKMnEUOCQj+ftS+e7HY
4kX9Lj9rRT8BFSi5teLPcmjr447jl4Fob/CJlevnH+LjNT3TQM3qj2D+JG03VaQChMXftU0zG4jM
h0GkoiEqXhRx+4HZa5f2Y+B0hIUL7uU3nRiPzNhAExUQKfxl5H1vGeUx4EsLWFrsDxZdWTWmNqsW
6gqHWlzBDJvg6588jZnZnhRt1P2r4kXJDz38ZwdZ4LbSL/watmOAIatq4aw/ARcNa2wtESuZMeDz
ItXNSl0tF8g87CuuDelxtq1waQVj0kjasX2Qx/Z7BOfoHxS8XKQlk8ZpOCGCSMpAlZkA112DvU1N
8vWnWJx2YU/KLzdlblb2s47bHP0sJS3wF6xKZ5cTe5Yqqr5hPmpSPO8KUp+8+vFw1TEUYyGJaIKY
ZI06cINe7Xd5tgHF8vPvefmf5uz7HbzQ3vBbdLu0V4f2TP0kaxzaT960/U9u/hQiY+foLUUuioeu
NbBvFDTfHRLVkH4OMkDNwoNp6L47AB9tXpxJJCGpRpSnTHgw8HBq/nfs5n8BKtWHLEsViQsU2OiT
tVM13GeJaMjsofMkZH4lCcvGZOmmYBPI9O9aHBbQ0aNtu9jhbCDOKwZDzzX8BfpYLTA6rNUUhVM2
yqIegtitco+z0gTxj/WzqSUo8Ch+q9GjAnPzEs4B3HDnMgY4ghp7655irf0R3rEkpmXWHxDzkWyp
jSMF1dvvTbC5UuoW93rrJbGrU8TXypgj9neGijzQBuPmcGSXmehCQe8gA/UFPY8kCb1RvgAQ9vs4
IGLdG89XHR85H0vZPsW2p/U66SQYLREpTPvlSHefQChiwLS9J41p58AZ9qpTmQ35mruh9gzF15PO
wydewfFF/xt9pWUSqNMLwiFbgvth9pEh2NTjUV8B1CB1UPzzTtvE6E2+MYWxF+kHiXCYI79MWZ9k
xolzANW7miN+LDQlaocrBdX08OfjGzat/VwFBw2HzzR56/g/VkfutgyCHdp+EekJfGjnmf1VowIQ
bcsRv/prOrZpBQIq5vNt1Al5slGpXqxu1djekitUoD4lKqrgT+5g8J9bMzCd5l3zM1EpvAgTg6hg
QWq///E9+A45FVBuD+DXWv3mZeWGMnrOKpTALH0tz6HFNhwEh88uiwtzfYIfPZ8clbYCpl9BhAmI
KRLwv7N5SmUBK5dWCRoOfqyfJOaiDYOJLuC6REKKZmq3oWL+tVFE4hca9k1tVI+krnlB8H6mgYb1
ZSBBjueEMnqSALUxwY9/HvwF1IOitOw5v3Ei/ca6r3Iwn3zxfQKTGaDAuz64u+AIcgH3o6mqE9iw
B7X0GmLnM9yTIZPOFGc68n4Km+GWTdn+hmTmcohB8mxe+TyGrmYyucQvaJZg0EcQT9+jF5TwnThg
4X5+DgTvvX8wWYT+yFpO1C2FWJw9JSocNVUYTCEpeniLenoHqH1KGKuENRVVtUCyD2L1Dqmi3+4v
0n6AcWXuhn+MKED1+SL13Fo0cNAeh7cwcuYOo9YKVHPLl8FyXBqv8ZwbzftJjhpdh6klfTpZUIu6
cBUueG1RzvreLdZRS+KZ68QiLKu+EqpE9xxo+Io7uV7+tVKZNfDEx5Uz1wSbadfYdMZEgUH8oAmA
pljMWo9BsrzejHKN9xeEhjXAxMgDvUJAH6egRshGcRcRaw2ctBpoLEapVe0bOq7z8odQOlzfSLfO
Wlj1BuSBJxl5NxUhEL8rokrFUIJmhVLzbbQWr8Si6SU4AhdBQLPJ8VVGnERckW2E3d7v91HwSIZj
dYfjEhGW2vZ5sp4gZJOgzh8q1mWXaz/YAImJToies+tkSX2JfzrfHmWCg0NS7SHgZktzAjdk6BRp
KuOa6DWzxcvykzbTcggNAtXAIOiJL3RV7Lk9u4HuL0SeG1pQuRkXDHWApXlV28RD1THPiM/8X/j2
sIz89qrEqbS6TmhUX6sBYlGJSAenSfmFE6GNNp8fkX/Z/y+Hh0reZYkQFUBtCrSCFFnJm/jQN1Vg
ZF6EmsVNzXQlg6hLTZcb5Xs3RUH27ejnPbfh5B+byoQQIcIqFO4lIWIXtSUVIqmc3VwkoNRlprmM
OIabDTRaZ6KiFEOhfAc6a75jd0x5KvLHoarlN4ajP2NIkXuXLF/ybVBb2YwvqlTIVEzCraeExvU/
miS5vO0HKtZ7yqE+7GMp4Bt8MDPs0U+QT1B/+4GI9r59dmeW9Fosciv5NxpX7jIuJGxFMR9r2Dmv
Q0HY1Qr63Lz34ihdDuOwc59PSy12wBMfcDh2qh6q9yzyGOfeaj60lP53bpeK2XHmqMKwL60ST6uP
jW+9D1JPciTregCLy0bzoNVQ72FGI4QG4BTflmmIoCGJAcz6gATSLK7ZhEjbAyGRThnCCfQ2cC+p
mlyYwo44UxErYz+lYjMNIa24txVaCKhsGbhLMI6fdPYKeiESGsvkRJPQPpylausQ+x6AUREY530B
IzOOeDtVKARDTjL6jOny6RTkOtwaw0bs6wz3i9opWtk8a9vv/QMYVd0oHfmMVAG+5c7kvI+n2yUe
uHB7VNUiMxc5lPu4YTNneeZZMtVfXJDzmOsRcL9tJRArL316v24/eN06KQqwtEWbArWCW/WO5q6y
9FMr2hxrNN9vBYjy3KD5/els8/Q/vDzEsuLm0bRZtAkQpXnsEdj1rIbTKstqs2r3KFBVA/xsPjSI
faGa21dJP2lEsFTWvIvX/NIbQJyAnOWZeCZHY/jWQAgtehxgc7et+/f2ZOdwETpHIzLh/OL+LxYp
vYX8nRR2QpsGqD9kX71DWfIqtxrdsGjR5QFcYboUgbe+P3emX9WdAtzMHQqM7sM15PxDfigBk64j
sj7He6UHY3QU6atwojO4z1Zy1ZaAwUPUbHUp8cte/S3gf3qgQ1W36oYKJ/lOkDMWXpogdaaK+oPP
QaudWpjNDfiiIOwXSrYVzBznh2gikxCpkTjTnOygSoyGW3r162JqSzHcY0U6rZwePbP1Gb9wAamn
s8OyodXiCDhszdMRGcdhAR8Gvd+MDWWolbZDNSlzBJ3dND9hFCLj0NuIgLVI4mQLI1EU9/bDv0nj
vc5Dtp3KozbXHggPnVaSXKAyR4cqY/fCn9QjoMTl9rH+hSaWTKElCpgduSaK90X+aZqZqWeKnxXt
AgJ5dztccn6tx2phZaImdN8k0dC2Xe+l3Oy8+8kZLizoxgE7VecjFEEtAbRd+CJVKsOBme+zZir0
TS4uv4VdRSjdBEvdtER/ebkR59AdNohSwy+5wXdDWcjldDqBOJAk3PYheym4qOaIiWhVUeO81wL8
wvlhN+8NDBljZrvyXz8ULlcVI0GCx4IGdDykJMFTBs355HymQEFojDZsQ/VFjjD1O9pkIeUXuQ62
j6bDNHo1a1LyCS+RlTZxKELN9IhDAaoMRKoBDhrOEjGPUbvX9QMTysP8xNAFKEbYe1/FNFzEoM/H
1ai4KvWCC5Z8jae9naEwEJTsYfqXVNcO1/LILGUHq96l8TyTMlEt/1uDMimfVk/5CcCuQ8r+AKJZ
8dgy0hEJ3rtMs9K15NhAebSMWhrnHC3Kel66O9wehtCx8OzfdNjGL6fMaM/EblO1SldOdLinBhk9
O+nyOTZP8sajaUuIZOUE9HrseVk8dRaJwtxsdb649fjBOzpSPp9hr4DJgyNhWBKJENcGnRSLq8if
1aLiOxWvwQmoN+JngPxQdPPEiHdpXKqDFo1O7kpuwKtNHsFXwHIEVpSFpUnunTOV8aO358fkm5Sg
iGWYVKRvb6YNzGxVkYIRYTAqtDGAvthk1ywYnIElRHpXBVuVo4lcBCqeW7iMcR09zGsf8SM/DeTV
p0Z4eL1sVTc4znLNhHoWiD5/wCmI/TL8jBwBkgH7IDJuzkbwNMfi6tSpAT25U0a7PQY/4Q/Wr1QB
J2AnsVNpNy/qrgGkxmjE+hgW3aVmMFkSaIH+NvlqppQS00P4IEgi+9gZ2lE84VaPloLPWwfR/0tp
q89mF9zOWVfX7a8vDoNmpNd5870aW4NEvq9qSZgPBRU21hJvLd2Pdb40TjYjSCiUcAH/ZiOxTj5a
GAr870ZgL6vrfvWGq1TPaWEg8bgCyDcKFWlauHwCDNAeF6xsccuQSvQSoDlPLnSTBD1Poo2XDHd/
A3KElZdZq3kYhAFcxPuJNFQy+GyH6Ntm0wdORdxMI0XejOuk5X3DraUj8kkfTsvTneXA7KQyEZBU
MKk3irFldYvaJ0seSo1c4Fw6tcqRe5w7GjzFCfwIPFRcYyw5cuemI1g1dO50S243LFWDQee1pWa/
5N+EHThjIaqVy8snoB+D2HIQKXJebZRFlEwBZYz7d1YWvv1r1JOEDQLMzlVAJyKACFk8IUfKhou1
07WKsPB70xb1fFkWktQU6HZrAm6MNQ4YFBANxPaj7AQpq14tAXT2NMesTCnr9ZiputU1LlXfkMAj
/GvwedsF+W7rk6OCpczL3GRB2gStkRvmTb+BCDL1ya19bGLH0kiWq5XAvmx0OXgjlgIGJ49Djjz4
N81j9vypxXBH8iw2A0PWctgMH+CAN9Z0sGDFIRN/dd4cDlU/jiBCG/FBhQFxX/6R5LPNc10KsHKm
w5ZRuEYWXSsdG3Jta5wZUw7xwczhltvaOsP8PXkysgstSmppOAqMisFJqmE6yExbWq4ARzSimDdO
zajISXXX9ltQrvLQtohvtgzCGnhDhEJZ6TMszvCMe8FbknolKzp3JdWcIopGJnv4/7GZiJjj0kFc
BiyJsP+5nTDPOORNL4MUTxvlHDDNyFTMagxrqQvnDMKhQL4g0WTdr9Q1DoG2in37y/qxXzTPrb0u
lY/gVI9VjLyqEsa6ltM526boO04J01+egAprlq1lt2WtdLbWyDcDx95Kh+irtvQx4I21mvXKSDPR
dMRc4sIb74/b48saI35DbxJOSdPi8WjQp9NYSpwh6y5yYFetZhiAnr41+6VCRPRlXj3xjvTspiQ+
g9BohwwCtwJeejQHZwmCvPgA9XYTgVkkcPEi8QJlU9tU0eX6Hctjqdb6siIR+vlllm6IXceHMCQg
xWxhj8baJSIGLBLWbXebDtugzaaGzpaWeJbNtEwL9iPIGUMEP4BUnan8O5z3P+SVQ13l3IT7NT+Z
zpPXhpWodX6Cxnb9WheHUlq7Tcqci4+qW4AL+lgK2GYMquH+wmTnSwbeffoEC5ar0lVPpqK5mBT/
eJ/8TCyyhxQanAU3Ib9gTLFpcFqKTj4Hqw8N+QhP0Pt8exb5hW18QXrmlWy4DwfkSFQ0ByvEWNPg
VUxkACvE1jdAbFmd674GbmRlo22VQl3qyz0zlN6FEf58vl/agYZnARCGr2nkyt9qvn77P4OZVMwL
EYsFyxaGPv4ZHUIAdGm5PLVWVaKUwX198v5JC8GVlictM3ri7I+ZhGm5d0t0kj//OiQpW0TidrGZ
wtnNg7SwkHHlq6T8Uzpx9k2zWL4rP7x1hetSDz6BQsJ0iMD+b+QehzmrAjoYC/qxJ3SuhCcLo9Gg
VoBoFBtpT2DOx5/IaLMrX3FCWi40W9zijm9euAyK1gj1wmkPdCrJicQZ1OmUNXVl+T6VISEYd/+7
Ld9ABbt98x0EZw3mw7dDWsoS2KMSBjqSrD8euKXFh93t97+kp6X4i7B7C1hfCVh6ONFFEVz73fN6
r224DRJxVajO2yDrh3/6Q6g2IaXZszhmhsYm91JVKsceYKqYd0vxBEyGE2W4YP6B8W3N3o/EIYJW
0DHQhZMu9uMmBunifbrANcOxrLI5J1E/OdyLhALDwKVT3KftthV2rB1dtM4t2AwGrIKMGOJepMg5
BKko8Iimc44+N30fxyq9ZgJ10rMw0PJ2uLPqePU42oCkGWXtK1rEn11jNJywzlDsu2Uy0goYU5aI
onzExkL/8xM3NegvZNJ+wk14xpp8apcN9nFllEKRy4wGXiJl1faKzn3xGNSputyVV/GzVGGuHGPP
QVwbLRbDTvyxjK6T9lDXYJUGVTrCpFL5nLiqpdx6rmQeSNsTU61Rn4RvwP+3e4TdBDKgP7POUrpP
diumZSD/wwiNw/m2KRYEHbnI/xYeIT5cppT8RIg0nh8HEXZEg0z03qX9QwLh4FcxJQwSJ5uBvKwh
IRJRtaUiRmvDiy5tumx6Kj+IyJgX8CxE4Ui+bkL/usA3zQQ/LiY1QIqXaTVEoPp4ge2UgbzsBY1l
IsC344iXJDYlzsDTVO7YW6/RFdIOB0zgNNRngT5x/q1QO6ZjD7AWof9aVFcbMOVXF4uvp0J5i1A6
MZSBhj4vA+DSmUL8MAYh7gC2zhI+Z3Q9Rf38iGPohcLcCTTyOE6fdBjR1ll6eFfP41Qnct8wTSWa
+0A5+YBpbtY3GKKZqz4bij8IT1vKsiM2BAan7xjtsz6RgEdAyfhQA0HWrNtVEYmKmOe6y6OOxxZL
/te7w/x48cbNK1Ph6941v6D6FlZ9tdKS1Dw40j/C5hqUKaKrJk5rGHtwEjdGBKSUtLMY04hKZcWf
WvCtrvaIHki1QSgDTwolpqV2IwZwS91RKU5IOAhvXHlR8GAnt3SNHsFNylxLoIutPDyDaVgwiI/Z
vCTIq9LBnRbY65259OKTzpvpCfdfJ87wyrn08ywqpZ7T5/Pgm+AUcaqvwfJTg3AgTnMfJH7jSgC+
7dXUd4tKxjSUK5eJ8N6yBwvOyIU6Kzd3QUE95oewq2UwPd0f3fadKaEHfcUGOxlCgTpd614shqYn
MRBEO8/vm8Iyqj65SSrhnJasQl2GPT266HCyQV5RKoHil48EoplC/mu6285rLRt08PbjzO6LCm3Z
Ose8YLORo24jkzRWMRcABKFFVk7q3kRHxkAfXnfLFE/XiEtH/R5i0p+7jJHln1E3PCuL+B+QImCV
YNOVRukHbJiDdudshCU6wsJrOu17G7TP7UZ5j/M6SjWQ4SPAoswadfWMYKHHQj/lr4M6x75CW99W
lEygSzJ0sW/EkBhbF/9VDSo65Qgg+IXIDkzkNYha9gnc4li+kSz7ogbKDSSmihNl5YrrW7qnsu6v
b30onxt9GkDtdaA3fEDxVXj/lmi8I6039oPEZf2VdP0wd4exp5kPEzBAV5O7ZaR41fAnSLu4oEDt
bHRZP+kqeHK17OFhFUYMtiaUfwqRk3HqHDoseekAhupZZUOPUBlY16Y5nCe6miQ/UbVAS85vfDVs
CEi+cgU8zKT+3Oyi2YVXhZ5ei1hxp1gE/8BpGWudCQxbaZp9ljjOIFuzG13OKMlYPF7zAQ/jLzCO
SdIsaQOJwr/YPKYHpNJ3bvMo2NPRnKmeYEfPNpsd2d9m2lMGZskAN1aIuPUbUdxmp2dzyxxqGGgr
oLzfNj2bXV29ZaNHZVzbz2BOejrKRRxQdWekNargQsVXEPwG8lD7W1zq4wJxi98Ihlq5+djXZBfI
+RBw91zeZbD4o2ikbMLUGPTh8vPUX4Qej3+oFOkyA8x2L/FeTwaVfN4HJjl7lzI2LdF0dcG0AcpY
InnmBxk/dlO5drdMFU081A/RxyrTh/ximj20NuyrKyFqzqedwz1WYcFqZo9D4A3XWqpL+VTI0UBN
eC1bJ2FUn6t6WAI2gMDH84OdGN+ttmieQDfiFcPN9xqujwkGjeuIyzlkfwuWzgZ6rbihFeyEbUXP
4LVutXj1B1FKLFDdyT6adlFbZYOtTCvfPcfer/hYCdSBO3Ovu1PUEMAYQATOerLS12K+svDkM2vb
p1KXY10c9N0SoUf9pQUMnzgsuGtefCr4Y9vZhsPCqUzfT8SL50OylWsugO5vxQA5hWeJoecxxWqg
wZQi90o8fEwi0GG5Sps6TNrJYJD42Vc6o2tVveXKiSyQcYesC1X8pVwaQCZBlruFpXh38MiSGEPz
e8GHsAMZHxpG+6ONz6i3GNkoXwmMw3GFT6BLKC6gdDP/UMECTTdQEqmFGLhIa3ngUdM0skZY4cxh
01KUej2JCWPwxYyyjMlRIg2npAa6ZkEqv5kMlwlntkNrwNH2zqstGUjQdeDZqflzcPx3s8r/whFT
cEv2eiQrFqvICTtVlKfa9bkS8MSCXsR0QeZI7a4Rg3qkMUKqKN0TCeeg8wI5QymBrn+BsBLvo1+k
wsbwX1Nrik7lGx9XapfDFC4LDppgfxT/Tp8NiGcY37q+ru/Eqyc4XBIqixOT+zHAU52s9dF2Vuwi
hw+cfSDcII9Ndd6/wYxcxO8FRpXzNXmAZNhj2n4qyinH7iaD9sVgE8mZJMb6kjZIDpPWI9S9jIeG
9t1+SkJDiOxq8qhKoRRGmvxbN/7zjjY4f1ZMWBdFjgyHVZu3W5aV3Dg90axy+AlQTIf9BMZGYk69
PmR+iW5BADRs7h8js9k9K/qvlOA3MGRgUhoybAPWi0CMdkPHszYycacDOeaS/wnYAimTVlN0sVpo
XvbHGrqGAZfNuC8Ocq4D8I6Z8/viP/Y2R/OKJIpTZ6OgOnKnCsJpXraUGLGozrUpW2CESiB0fO3C
6sWfjzN1wIwW5sj6PzXN2l6ja22Hwlp3tBfowyE0w02ma6AXe2W+ldNZkrKPQC6IclKybVUbmGqQ
42afdq94iYmRtoVMf2lCtknPdopmWLzRhlC3eULAlK1rXKARGn4ApIoh9pP3d46oRl7KJUjRvnYi
BSeOoGpyDzSC91dS2VwwMitu37qVyyFSsqwyiW9LgTAFj2TBgMk0UwZvq1zc335GA2AM4DEu5GRz
HrRbB6mv3tmOUMHNcFttkLus4L3ZT9cvhjJ9DVMrpuy1rYi4N8wN4e7YPdSLZFlqgj6d2gA93JcE
Yd0xqjFF2F7ohiPxHY+z0Ds3lUPSx5Sb9XH+mLdwKTAkL29Mt5MNo/bS6Wl8qPK5tsrwDfo1XaC9
Mk19TurkfR3pIdm1z4dAYo+hGBDLVQCPj9UE9bSPJVL6FpucIaJtkc/0Lne/DrWzo02rwiCoZ0Nu
InPhmIuU8EyjzJORgJgNxOcFyFxiObmvZHbBZLqk1Z1D2ziCbCloWHQnrbHRyseYpsw/JID4ezbr
yDs0AJKBuDZx4E6sUfMIgfxyvyHugZ8fmrMtjlfs/tqJ5gKuZTsI2VquMdIyjBqtHPtwSVITbS9i
k/zL6f02O2+LKtwzcSlzLVULntQ+h8PQWcx6EZhTmDFkZ18Kmxoc6lbSm1vo6B65dYnxuXnlz0FK
+6LPgoyszi/fqxcEe+WR6uo88EoqbRJbNNVZagr8y/sl11hatddWgvQ8LeGHEVnG2AM0td5Nq3rz
5n5UBcrVC0d8RYWOAwhjS698luj0O25PRxV6JZboX2dCLILxq2h38NWeITOv/wFYBSKwAgZ9Alrl
5gdfXZ2vO6084/rEkUG32OC5uhGqZJhcEZ6w8I8HOO+u88Yo1NlKcSkH1mkcn1DS6sCw8569abb+
3h2UfKiflP4cJC0SRsoMjgP06uuKGA0AAsFx5iqIMct3TMS3w6qs4QDY7wFE3ZtIDuxdBoLn4ZGO
yOsi1F5sS9LAqI6LlF1+bjI7OTvvKoyR8bZWLTlZnZdcx//MqTwQl4jU1b385qK0CjSIg4cyEN1i
Mf8DO4dinLeAKxp6k+bZIJZY/9Umivx2/5WUI6r/R+ieMJlFFFnVAOTWPBnHNThbtfpeo1rmsLOX
cdV2qbt6+5Pw20o4vdnv5mZB8gBG+rz33roRm1pRQW407DzhtdaUO+HIUNWfysGxe9LoOdCuzFE5
Ex1CUMwJpjzMLG5RmhuPIMosYMxDK3zKAX2XoCdSd8YOUr1F8maswcJ/9xBdQIYLz53MxBo4R4SC
G1N2I0Oa7U4tQkgHFFpg2wO/o8u+VmynFc7iPTZxEqeCM7Ngh62GS8IoFIMwMuWct0KjEptGnnAm
I9Z4fTDETUWQ2ReJNax/tgyYCXMxvJBYEAJ8BFJjP/DT28wzB7XnCH1m860Qmms78n2Bui1WZ1Vm
1PgcQkRq8F3Mi3DRhi4fbzr9big+OAt08Seh3MzeuIRZuq1flmGVaPyi4YTeg7JCYnA0707e4HhW
s0YN/mm8OzytV0hjM8byb7uH31GvlRkwqdTVMcyXxU0mpu1WDIq6hxUwyzg3vo9pwD5LzeqnJngb
5y3TTB9qze2q3JhkHR6XU2NNxIwN4VP+nx0qCj2sLCi4qIJf3vHVRoaa5CRis/dd4Hq3bkJVLoUQ
debDOpmnsY28ynrXvzfIjiZw3rY+A7/tJ/zsc2AeBWlk+cRFP9YLlM8QaM7NipZKzfWaJK0FbYZ5
YCDnT5ikRefg5NEf7rn1Rj3nUPri4DknquZvyPSoGdDdg2Wv5l3g5J3GUKbgoqplE3w7fPEGnS8I
HGmmG68RB8wo2o+LGvP7t7JEB7VOF+CKBGLOflr9BMkN22J9VQBzIzyUE6wHTT0to5ouNrpOrpXF
k4rZsQDmVczruNdvPU2d8tSEki+SM7YMwOdIlRSbeCsexvW5Q83VqPvdYqaImutzf0oRZv+z3ANJ
sHNXRUEldnlC/LvG56qoCSXHdZSr32uJJM+ebHwfE+jDWjBNM2qj2bd9cc3+gxR6SmDzx07lTYm3
rHbk75G1mNCCjUSj/vkf0A8ypz9OUsWntBdfBdhWRrWNmxSRVQdIQQrxSQPwiToKW/66BT7b9YTx
qviitoPgzNQBQTzRvdzFU8R9fM1hWX4V7g8LzDpb2RGpTZ40B9IzdDkUjQTUATSBzwh/jhAk2tnT
bdZRg5K3U/95KyI/OuJ32QQKalGOsKG7yBL4Ne18qgIItDNtPOKNj/vyXsEVsNtOn944Ij3bl4qX
VKUuNn3NrHsPccTuxONCuoROpJ6wxudMJB2eBnUD4ys3kbjJ1uk66hUsooSy4lIAlXsJmN7yzkaD
Oe7x1m5WZt/WRnJ+GTaxBBw8l4aGpDnBHit4o1RtZnzNr2D5yMhmmhiF+VaGv4SgtaTUgaUXy4Hr
MUYUL+btB4VzeOGrrJmqykCU7yKkWlFosRFetSj9KXj3D8TtgvVMQJKZTLvFHiI+F7NUTPoqI7+y
fc32EtU9WfkSMzOBrzAOZvg6Oqu5wV3oKRJRqrAIaxgPEBKTZz6lvyvjODWFyBm8fJQWyYbBUb/5
5prc1keXwYnab4olOOnphQVBKFRrTJj1R+YzeIJ+3WNiX4Mmw1Q8IGRpPnQQyTjY1RSGdE49e/LS
184Bm21eJbcMn+emq/J9NDqk6o6ZKgaxBdXe60pcTt2v6An5e0QNGseNCW4FjIMuvwgJejFxY+9G
CwzaAkPkO5jiBsemcQo3CYf5L3RZ8K+PAq4/mdMikIBHZJ1nUHwCXWSmwSNalC0HGlB35ysAEv4j
GbPGL3LaFByyj3mA73GMOzvjSB86CvWsLDz7tiKaoopW2VKq0FIs/hGp8jDAt1wXZ924WofiAcKR
nv+/9RdVYAD5BLVX0nbLTCA+QVAF8u09x1JTCBp6Gbjxp8mIT9sjzntYOSIQQD1kqKDuk6DI9Tck
aLjFMlcachqOVx9ZEki7B9+evbkaJz9o+eR9YRfExoAmfI0AWSxCrOAs8rJbrYpIhyOqxxg1t/nh
P0HbbUtrCUXgNjnkHPiRXI3OOJE0e3Fbc/cRb/4R8100hPEwOFm37ghUoGz5yhniTn3lA1Nz/lhG
eumwCZyyIYm/v9ePgccjN9yOmSKUh29sTB0S71WtIMcCPwSMts2j+hQ99hZ+Ku11HS/Ztz7EEHZh
B0nZEyEkUnaZB9YYLu4KjsNVWwTOKrB/+Y/TrTigR0mZtxA5DiKxX4QtGKPfPFF7KYEkRj0F2fgm
+OWe0RxwxR82o7Sc/r5lKR9a9/kGIm8uCNu+zMGXSRSHRniFwLp3+UeNTz4AjzhtEehef+lHggoS
iEV9YjedHbEZN1uLcSa4Mpy8fbkQaqk22f8BAL7Jm6m5PA9DYnxLYs7UyBijGw8CrLgCXflS7a8j
QDREc97SGQXuRxx9LYh23EaJ+LMMUP8eUe4lV/OO27I7psxUYqAxzFaJvivz5dHRrGvfOF8kKId7
fJ4xXdnXy5/PCb8SmA4Oh+l6NsTGmSEBAkiP1NteogppDsqudSdxdV5tKqvWipCvJSFmYXDn4sTi
h2r0B0vc0bk8afNOhO8/Si5xu5ldl98Te1haDapmbE2bVfUU9o9q04EEo4ACO448q7IxxNIiW9QU
y/3UNvEOe6kvAduY543g7eln15vsm4ybCCaxAEDax9vetIla04lv6lyOYdBhaPRoReQYarFlWDmi
IZB5rfbrLRKLnH2axC4SK66bS3KAR0KPzDszeM9mvv/jzxHNmH4RvaDj912pm/KLgpU6DbDH1sYI
6YTA6E0luP3DKzuukAT/IABpsPN9pRx6uK8fQOipxCaa5NP2NwzygfOJ2ermob7m2F6w70iDYx1y
RJmAwWGy24JTASzOI8q0USmMix2qnS+zpaztDx9dow57mhAFveA908hfzzN7WZom8V2vRRBAUV8y
z0dMoem7/Sw6sYA90MCFJESSo9ff0mpLaU8ZUUpxbuxkkwErDce9eUW44yh6E8l7nscH1A6qBkuC
T7oCufggvIiuy47q4DRerYqD2XCgw5S0IGqNmC6LUzJXHJd+wLXgtMxByB2jvBb2evwZL9fvzG4J
tn1ZrgD5maVsDVeUgnU5ougepe59nHc/gJZ20AW51VTpSu2MRQL/2KCjZBQ1ab3QUzpjX9pXMre8
0RT1kQA7XN9vw3ZIm3r7sYMxMLyuH0Fujcca7PriuETtq+6/qpggsTYffEguwPLRicDaXDzObXeg
4rcqp6n4tk2orhWi6Ha24iJBBfIyeHG9Xnu7h+YMy9PGqTcy9Mybd0tDtCUfZQKHaUmbms7L5ZPe
GeeiVwYrzDz8NeDDBpN4lfqwLwrP79Nzt4+nkGoCGrTGSOFHNHffN89lOU9QodOAkb2S7e7lOb19
Yd18v5RQrw5ecQnJSPwS4DWC2Pz6+S4zCTn5eG2vRzf/UXYMzgAiAo5JgJlI1EY/s/e3UGfQU3Gu
cmsZ4HhDQKDLP+LnrjtRrQvBvkbdZh4cWEbOKxAhsUcxoK2CnZitWtix/qBElGeYbVEV7n/ymWar
7guPJA4RJgBrbpB8EXG3lAWfjjQWEIG+FIlXmPxT8rMVbZQ8YFrch+Z0IJRkZRWIMQarJPjbCXM2
FrsU5o83FapaOpovQkM5f7z3mcPZeK7RvqYg3eM4iSeoxOMTIf27gSn8/CKlZFnUOY3zAK91wHHg
YEReAcvjX8bSNb0CaTraeMfTzUHg7FaBpocebMhYoUyjkkIEQWRmAiFyN9YZv2sF1MjlKLrz9h6g
BfL6Ss6/zFBv/0BYW22b+4wWQ3Vx3zXiLQ4u7UTb+QnpNP7g2LY0HWLwSyCiSmH36p50REJ76cpx
TcwhZojZpScnukTD25txq25PiQpfpwiXrd6hh7Z8TM+Fa9Is6CMj/C4yEt6R6xQn24kCHqwxQXyq
QE1oWa07ZbPxTomZuPbmjMiV5AdyfR79aUQYPhcFPIpHeyh+T4nh/EAfyhocggRxyCMI51H9KC1H
+bTY1NMR14TmHMCWSVOhwp+Ou4wVjNKKFhS2PdBuZ/4CIlzij9JFmMdyNkQ9EIMxjl7sFUt9By5W
0bHd094juHfNEN7JVESiFhkIFzMsq12myFfQSjc6j4xOv681TG5Gca5B59cLdXREVhIfXRIr3rQN
UNiA8YdGvzlLyeIsdgxCArFYR2KDenh3hICQUYDsvl8Ag/H0a74B686yUcc7wR/3U2ylIXv8TqyW
+shNIui4rojhHWVZApwdBXsRbxD/pmGZOpz6AH3dLp+DTuc0sb5KZfrvVo84PwUIfNZGsTBUquny
2BEBeNlkzblzJhQTHoqC0TIfpy41Jq0r4xXwCav/7wkJoNgpuHWZ4VC8XSVoiSfCf983skzn9qLe
BOjOS4lgaapSYoDc2KgCnzuvHBfEQoXhqvSABfkunmdMmb1mr9I9XJA1zWnTZwIbxqNwd1bcc9aH
bfnGekYWKaAGoz6iYepsjeR9jWhkHK6XVGTKN6UWoptp0SJTvoHzrsecP4JdMFgtwGAk2Of+LHyE
1aOUIWABENRXbgM2zdTr2pnvQ3vQRD91zmOrZHqLDoLz/3GgXeETHDA7CGpJmvtenwF8R/Ow+DzZ
Tn4AFqkqXxRo7jThZjGZwZx6K0LwsLtSdF5C9ukPecnOafwNwPLE/kMEDBkvQD8kDmgtn5JoC9ex
YWEiwyhDT5ONtKmfv3ncg7iZwQGIRxLZPoPZ8vBhzmcNhQsiuByzT/Ufe21afWtgT37qX+xcRo/f
3b4B9MuuVHuqo7vLWtAU4vnTrV8Y0KBqh0BKCpWvcA7ZTibaMOZvUOHiHH/RV65sBmh/6nRDHLuD
0GSOiKibYn9KRGKd0sXyoQX0rvr3HXRTqtsmEse+HDo1bB2gsZRTgUsDp54YothCQKR6ibbUL1M8
DXwsTS+KjURWNExrk6FAdOSbLWkq48fWIwyU9ls4YjMfE1w2FbYs+S/v0mqae5QaD1RYaEbeW3UL
1oCRk6YgpnIAyjcEkuBFRKYcUXj7KrlNrqeT5/R57wwAVOOuwBA7EzVN2RjX5Mkjk46VPn8qENuT
LmQwxUWwG0toIS/Lz5h2/STY+AIi8SgcPMzYs0D+eOtwPCHiNkZ24lD8znL2xYzvaVvzwmP9pScm
cLPtuuS3CT7TqR8P59x4qxjFfECkTVa0YTbL6ocSzRwUsV0uf9SszSmvd5GoYUQfOeiD+PVcz0pm
IoZkNC0XIzfzo9LIjhJOKlYL7oFYELjc5+fl7duqvFdg4z7bwe+x64BJWx48I2Pa8q51Mx+SrfOE
SPYcHqdaV9LDlIgbYAKhYc83tmkhJ+yRZiKiAO0DXVYv2A17YW3ypJzBpkiUbr7o7KJb6eZjbYea
pnAz0P9AejnnmKjshTyTRB4xoO3+s8O0oG7MsSmz8W3Hx5G0Qi5pF7E9mSfFDudcKS0Kfi1Di2WU
NFcqju7glky4MWyz9X2Oh/y6xhgSqyD5FqEMCOQRHdKOw8whU5cqzzOdFU998rd7ju9YKrzMGhhE
fxXFlISxvaGz4onL/MkovbZ17e9nL6/jvftfWJJsyZmAwt0rlMUp88MqlW0TdSgoPFQrFHm5sf7M
2y9Kgm7c3lKmARqQlKbWSWE2PHjqWm9+FbFLSJ11+LrxrtMGYqZ+/zOxREkNq+GeI5XgPBFIdDx6
ymfQSB6SOKT+3LRrEnOMZ3U2erAprse3+My49a3VqO2l6HkFFWZQYaNwiPhY2QOMq9NIyvLQsmcE
meyZoVYKyeL6p6vqYbh48hIOeqTHlWaVjdTAuQxHBXj+dTtjPUJCowNkJbFjRrKNUGcxOwnKxYd/
WRTV72WUejZi4SEzmvkJk11bVxydroI0BgmAuXlrj6QtMcbs6YYLesXULaswy9qW4WTHebM0uW3S
t82chVy5mOE8ZV+GHFgWGzCIX+2zR1axRdr0rd4EiE/XA/GdeTe03gdLGGcV3b8XjtEfEdBQ/l03
9sq8R6XIIGWexGcRgzAudno49haUbZic55gIopcreGvdE3Wr148JXEE5iLjSQz5CCZMskvO3Kd2X
9MOqlLCjr/2EpxvJAUMZBgrTg0r+9l8eFlOglx9jtRGHWdfIRD3lHJKam4eIXBRpfbnUNoxKGu4z
RQ2FRlxZuLk7wBNOoTycI/4n6pOvUwcZVqeXZVo/zArD1TZ0HSsmmYH64SCA81sFBYyggp+YAR7b
Z/Mr8JJIsod/z3LcvW2m8gC3qiqlfEUZE8ieIgt3J7KKn655N4mpLckXBPigc37DGI9o3S3ZpzB5
ykr53sK3/XPueFzk4zyrKMUI08/icJvagnXP3545ndd4P9yJNeYX8X7NERgUdb4SYDIyBRm7BgSz
CDY2yN6mOe74MfG/g+OkEh3WKLxwIfWUDG5LQVgTVebsL+d1t9s27kibXw8ub0Z1kBjmTDhRDfYr
dpThe6QuUsaCSOrQF5piuI+yQjnk6wsShYck8Ayyh4EUwEJNKjVuaFH381DGoppT0My1QJ64Pz9o
ba6OmWujyu3MkZ0wFgQHiliVhD4Z3YXArl8VvXbtI9fL+tw9+QNB0CzTeU5erC4jig2b5RGuKHvP
HFk2OxB2+skoYs2pMhxhSyuoqHbq8KpbS+8l7gD7qFmAvz6/Cty2GjMrV88N+T2kLWkPnDvUbaAC
heZFxdUbjdxnZSdvvUVHfuLFJl345tueKPGq8iVmoHMC4gminCjQObdtGvxxMBmAgPLM5NDHTgTI
7PY+si9QnZdAT/SbwyHoVQ7FhJkHHAFfZ/q0WbhSNwGH97xC/g9vqFPJk2F6o1vNLrkBEvUKdzEc
Mwz1HXrL6dzyemjYh/x2diD9SoGL7RsaDpu4422s0JNYtXmMjJnVD0HXQGBcgcfdq6AXIY/9IJif
ytmkzLnwOC4xyaqMTCYudZtTv92sNQCgaFUdk4iLIlms+7/cEJ/U+2VhSMlCeCE3kN3+hxJmaxzl
J7L7y/OBrDgs1T8D6M3EsVeEjo8sl9ERT1lgyqNYzb63fO42jGk45Q+SpfbwUiiB3i5rSq7WYPFi
7cBPZCfKftZNc6FgSdtpcpA89QjwmIsCsBIyN1YLdnCqlkvUTj4rJb7NSKDOLbLg9afMLgrMWFSU
mdWP5Y6hGq14XmYluX/gicUmVfCOz2H3kOcU3caXh5rl8xw75jg1V1UIXwUQiVEe7joSuUOFtEWP
at6JRnAlnxLbbGYxqL5FmnaGa8Q+Zy/AkdthD4NKUUxhUTipcN0YZroagzHfMQIBVzqpNuCyjGso
tW05B8OxnOpwAzj7PM6R5w31cYwTJMxDl8D8B00RZ0K/LPWwRRWhUUyKf0oX8dKl9k6MtJ8sA8JW
B3ZCT2N1elsFyWsqPVBjqSnNcyDCTR2HTL8oBMoE+tGU+utejDK16oBxRpvkOE8HfI4DejakqcC0
z/p0QIY5JAoM7IUGZSPLOHBEHhc5UMknF0bPMGUZ6f6xy0bWWy8gv24A8P3qKwwIluzaMDfMCIMl
4sJSvTYKDMzdGgiYR/vY/3UFSRY/1d5tdFq/YPG/uUuwoVLn25FOy7euXFsm9trZb8mu7mK/XecD
lkNjTvkLwfjJZ9vBh/f13fAH7v5PrtM67Y80boRB+iXxf/tGuKcX7JVaR7vRxHTjYCXuNPZ+EMl+
a6l1xlajuJyXoMhWnFB6gYmtZy5FttuyiJtyKNPnn8q/mOmpJxr/bOn9A01PyjIG1U/6CkS2PJqP
1/jfKmPVGCyLXGdqWJ9S1/3VXt5avVb3o0wx/hfesHayKAR7pH9FSRtO4h6CAfWibvRLXY9S8XMa
P98sWFrkXJdMe0U0YovRueq1DUTOclDMdztgZNEHFtkb+kzZ+J//jz7Us+8aXZGTQFcu6nb1hx5z
x6ftcCOaS2LoumRBAA7v4ja2mlHZokYrNG9M4Ga1XSozRInA+Hil6ThhYOONrObH59H7IX0hoGwG
WY8XqjtnXnt8oZ/XCqdIkCPB9QiSBZ3/JHjHoJLRhl2+ryYMfLMti30074yIm5J/RSXzrr1eHT0p
B9Hsl3jLRaoewdIpPZZYvtkCppVCtPgPRIhvRkcwgh9ysr6QUN//9V6lDoilTGd5B5qE1rGGAlKu
AdRa5Bcp/jaagWLBQuZJxYSLgBj2G/5KKHEVtCTy6jzGsAm0cg5e3s24SKdi6VE2XqqOgKNdfN5d
BJ+zQt3lwdo+BuLxXiMAAOPzkvpMCaivG4feuD0nmW6LznEiArYMY5oAy5ogxzqbkTIfDwgW6xQX
8quAY0GEEY6kwXFeibyyVkegFK7nKNQj6b71adt6YFuIuaILNRBDAbMb1/IhQr+dTZTaf0s9qQcX
uvQhs6dUVz8vFtbzCobrUMxfxZ7MXCaiion6nUtoysFu4Fp1NgaBCSXaZfsNmav7TGW4CO3aGJnP
t558uKe10h+Pf1U0QAN1owi2R1rY5tsQIjAPsK8phhiStBSquI/JANaRzPjX5F2ZsPRli3Zdlep5
IcT1NRqO7icCW1BitdJtLmYui62wyBXW/asDPneE+CfFx0/pxAKEsi1KKd7hcS//mL4bcDYjb4Jv
TtvAwJzy7wQuPOeQn0xMa/9fonv3cpj0dv4dYNlrFuQimbb1QonbM5mEuqhIOtfahvdODHhMhBy5
20rlpfHmO7gOyX+tslwokQGMpIn8LAnNh/hLCc4+UPfZrFxWjoi5OCyHzbsFHNga2e/uyq5+/JNN
Jfl1f6rZjHIhZ0VB2nU7vmAvPplwD+xSFuORbLwfrCN9Ps401Pk5RKvCKfVThnTsMbB/WEsjZjVb
Hvst3WAj5i2pux8Qxc8pW2S8lp8gGAWepzVsu+KDjVT1EF66ofpKbumhzEEPQRKxa4sTx4HwGpkz
BK+uV5Unq4ehbukJTV+mtzGC3TEWxCdKNGiAqzp+uG3Nm5Z+18xMq4cSbTEbzQnG5xkmWUO79dmz
8C5ODEKo0e8k421tOFXMaYpGIQYZx640cXfIsAlcBBqaJHutu4C9JzpPeffL11x+xhdXg1SbKYrK
sMxccS/++G2Ybt+7sidbsdBNeuCKVUqZ1L/n66RqHyeosejfzkE39l6dwKTBTFvmX2R/kRxzMBaW
ejBJxdT9Xik1rJktvjP11OEznIWKcMwkyXmV6agBnW2F0A6EgEiH9xp9np2ZceLZgxXiUrzyhBfk
VPbaATTLXGJC0pu874dihQdhHRveaOxmUhXxR1uQ0ESOyrNvhVKyPT2XNhpSFHvFws3tWJkkRUXt
qFhzFA00WlWNfaCMRIQl1KmxqTlredBuijoY9lNJ4SsZHvzHpuIRqM7Ozw0eWoeOsJ9rOklWp2CQ
wfTZFVGIeGfJTcRIs9lB4C3QHF03WfGIPHTaVL64yWe78V/Y/+2NrSYuhIrUbOI1wMlrmGDyHYt6
PT43wdgzgftf4aLK1Cu5nrfDz/wNPupWUDai202ZspcR0t3oub4UzhJl+CdWVOsWQ+jyOz8LuWwy
HSSsAcRvCooYpduvbvV7lPCCnrw1iALDkfyYrJRhaGiAIkI6mQhuxI0iITv+zKu+yhBXHy5oNipu
z3l4A1qNruV4pslH57AaYb2bU+46TvhDgpS8UA/3Rv6MMkTXhiIpc3bkPxjbd3z+mP3b7HVltTry
TZMSGTtR0nTT5pIPZJOlvvHUzIRgBK7vbsCTqRe8fds2lZtTdIsFH0Z/iYiE5PMJjeDhOtMKCqhP
Eb80vzMETIzYQMbHIK/6e8m51UXzk1hRuph/uY2g3wo6TQXtX32wLlmM80oYSEbe+4Xewbfbl+73
4I7Sb4XTsG78gUL4SJVit4siSnsWxXh/mgYCy/yJPwLpvIiWz9BpQCsjI3v8qVQY846fMQrqXHKI
nCM1CftUwp7rI011x/8i9uMunjyXmEaHQMRNpgdCKR6O44G2HT2J9Y6ze9eg7igMPLPGN09TJGoc
Ohr8KkQ09dBUrog7xXE5V4rYxEmB5pLmO1QFSwQDkkN9rq9KKYMFSppyKkU2EJ/PIjQ0oxKOPm4H
HJ4uSIi0LVOp/4ngeiPSFTYDa4FoiQzTuu/DpsjwkmMLTprx67QeaZ4855CDbZsQK9JeEPLC4rXx
LyY6hkefqL5Zp5KuWfyv4y8l0CtUByHkQGrEZAmeqdl1VZriCC22o33QohrqkHcurRyx2k5wFLBb
9JOv/69Vpn/KlUM7hFVS8zuhzcX7phnNngQYA10vnIZQPBzn8lgdCXlBXDckRQf/TX0CNb5faCqY
rpPwIk644OYABrcDxuAcDlLKiMYPfGd4syIXfYY8Tz7PCcCvenj4Wjfy0/kZLrNvstZbTcaxFXDe
CFL9VY3D1MHjNEuIO7o3KtvbRHhvBIBj8KahxwaLt8UWsdkSEKj5LGpZkb5R6avGapEOgV1hVE/u
akJrGHiUtdF0N5SMI3RwqpY2aZEGpTmY4jERH0X6d+tPm3HnceCJ03x94WzC6wqAbtkm9xQPEgOF
rIW5dnv5Wds0aVyBx5igOdjksIX+9/9JgYy461kqEpG0IHxC8jnDonDDEE9ye6UPXkBrC0dBmZL6
X6Gl0z2XtPSt2X1I6FKdeeQG42zwWI27U3IN8oelwWPV1CEOdHkdMKB6zmgp4NsHUJcAopYYHr53
p7r+5BqOeOfQ64SivmnbepsYBIVzFDgYtmhDW8yZZgg4qNHJAuHGP28rRNDuhwinjk6owpCVvQRr
PKlwTOsskgyOvlZpXUdFW1yxDRbBDk605CtzJrqTezWth4N4k/aFlTDoqclvLaaPrFuVq0uEhOl9
BmcDgbT+pDCOhGz/bG9i4Uwt8J6VZ2Z7bzrtcdlMvJd8TrFgjEKoP+uqTWIECID7+zm6MmvcofZw
pQJtx7yFWC8qpkIJ7PUBuL//ml77OUMnfkvfROkxPG09W3NAa1kFEZNoPAG0EHcQ4bTertcvYw35
WZwlZCJFrAxHm5NAANT3PEz8P7IZtY3w+8En7Z9tPuToPp0W3GSooeboEdTkLTPx2gxo6XkymZHH
mYhHRyfhkABqiW0ZPZK3nQk7nvyH3nsgMxUoXaB0Xat5n4XYaEXXb/WKw6KyAULQeP15J3SWofUo
u7+Yy7B1DwL9YnbtEewF5b8rLQsEMTLhICipwSj60d+aqeMDol5qjPWoCLqS8sRp4Hu47Iy8wVws
SzWRvPE+wOtWRWcZzXtpl/uCP1vm95W7YUmEFI2YIExcq5uOD5b/Ws3GMKhqLZNxcIikljgnlF3N
gw30mYn6ahC4nt/icspU4OXWukBIhXwNRJI9IoIjXceu1odqtffxSGK+7ik/aNMVLCnw/biMWmMx
phdgfpuzkE7YOgYOmwI6G0miJExTRKpmXfSQGGKelBTzPUh8eBipEMcSmvDKyVTbxx+sZygvAhmm
m71mT17qygmv1MpGLH7ESmYhpAArJOz6R2JnShbpuDeiOGp9v8Rv/iD5n4wy17Fs1IZBI2SbVW02
3rubT4Kej/dCRc/hW2wmciPbrhmquAfj2EE7/CpToD3jFZ8r25+FQngvnpIEW39eO8Hpi2KrN/f8
Ryq/KPBDrixx/JWMiUafINcpsR7jIMobLCVrNFrQ6KHZSiOpFXY0yriCwPms1wBppzPqlhHaSk6W
Nx8kOFWOI4Hub1OcLvY12d9rXIROpS8FBfueKi65Aa9laikFgtteNvYGZZIqvf5Ru52PuzLjlxGU
s7tQCgoH3IqnANy2cNWoOaahBGcnoT8F0DC8w73JeU+AxrGc8qwxMj2vFO1icPXSQH2QWmmYaDoU
50kKiMCK+BACAIsn/uxs06QafE/PdL/yjHR69T2fr9e4HzFEh3pVMZ0T0nbKMz4C6WVob+T8SSnx
RS6xAyaAcWaCTQ3J2SB7Q/Lw1wxQnT+Q8+cKNnD8I7jSGOqa7lw1Sq1WsrewAqeMvWKUcf3nR+Fp
d0/u2AgKd/GouxsndP4DxPq93fKJ6+GyAfGGP+iFyahKAWuzQQEQUbNyQYuXPq0/lQZunXLBkXxa
V4pc9LysdaSB3nV+wSODiZATVDLx/8lIzAY7XJU1mQp3OTvdcCouzEdMmMioGb0VYSxMsPrpYLsW
j5m/S7/6tR+gPaI7c03vrh7xQvlZFOEhTodUuyb4FxjZyJQ5AzFxww/j12C6DHDtLJamWj6aP4KQ
cw5CK3f/MLIFPp3l9dfl25XIQa6o3TJ8FHdyVKJ/R1IX3eQojMAUbgid6lI3/URJGdXg9IDNsOyk
/F/TrmvCd0oJ91gBGGFdRaokHcRbGFjDRrnEFsa7Y1Ls5a1mV3rTfgxdiX5fuAaNKj/qmGa0QW23
R1d0wFG4mqB30NVLx84gk25YgJiu4qzW2rz4F/cJxVkuq0KM/F5RzEMEHOehtVR2mhA9U3SUFqFs
OOfCK+pwWS8r9yReDrHv3+JVh5PYf6OGxS4JKfOhzImII79J2La9deOd8eYBwHvosj6LALF7ur5Q
42HYrHaUg185zVGprlnhBmBUaikhBpWDEFguyC1bfDCXmm4Az5s4ggC/EpmW+wzT9nVsKaszKP7H
vq6SGaVvPOd3vZSIYxnvorvL1C7c08mztJ2RZSm510VLQ3nnu9GnqoOMTiYrYttTEkmikU9mYYYi
d0NkogL85RM8LGqhSUDqgD98Lj9vBXoTFg/GCcasM5NRfFO65xlQElojdkmc/IZmGJg3ByjYLvTx
MEAKvsaLE6lyrIdzd0fI+8wBWL5omZwA627/NhSZKhfV0AUIqpeAaP3E2qqTJ9LxUggzHG0iuLfL
oy26uAsb9FcZTGR4A1/Mb77dzwcilNLP6PJOVD/aBmFv+rnIfCuPB0mBjhEWlxwiJn2zwNnyEO2z
fjh84haPn/ysiu0FnfWDfsGIuCAOtOm66z3gWaZR9IB1uEyFqTEujIW9cFDqHxE+Yy/M1pm1z04J
GenTD8R6Kq0droByJZkiuwrKlAyVkZjS7Zn5+a5hvDPghI0JQIuaLR9OQd/qTkTZKHVjSUGP/Zih
YMLQmYjYpmvDmq3e+umEvyP1l9n9eeReJeCz+5g5yzKggPLP1TOeWr3cLC9Rs0OsYo3ybbPeND3l
A0y+ao7jwlSPlXnp2KdVJ38vdrqHkYhLq+tkWyBwTyvzjYI9xomeWih/unupZ5fGClJwbykGhYMj
W/nOJmxDXclggOyr08R7zQChBYUo3M1sa9ybpTrs4AWxm3cpk/oR9hiSi0dg7MkWGRQa57XUi4c1
kfDthLmA0SsoAcQxZLCdLJLbbTNizBrV0grfmsL1St/8StCVSG0qxq8vx1hj6Wh9QtfxbzTZ5iOR
JeJ5sz59oIO6TV/eES9JGpuFS3+IqbLO9M19BrhH9dWEM8uXVZWPohC2d4zerOVm4wnVe5m8SIdU
IpMeL/OY2iy9O90pVrp4dJcCe0JA3nLdJI2xzbRK+aAc7uQSA7LIP4+GSNeO3JBfiliExTt9yoU5
IOHoJmF5eKUOEvWo2L8gZsAfCJw4pGoOYipm82Vdzi7U5wKZh5D/VlAUBtNg3we0YTTg0hO5Je1w
MJL/e/tbPtXgoRrR8I1IvAVU6P6nj4vIRBtLRrp25ZDymANoAFpQf9i6JOV8T3+Zebr6/XCV/PpX
VhXNniMdsDRpzSm+osWON8wROZJ0LtEpLQ46KOctUWXPPM+2hX0DZjleeHPHJmeYU9ep2prY842l
qPHe8p40sX+5dxP1hoonEAQbCd6iygeW50BolxeMvc0aQKuAiey4jghII5pJHybOD74YoNAKNEnE
f7S0wKfTZl0+oAlZzOVGdXQ4Ok24NboXSYR5nujXcNbQtZBoxWAGv8PCGomqrXJCpHupU6/JWsH2
FiwjHRUzDJeZcaG0PhvyUBlnmJqbqezrlZ16xnLJCR5zr4KTkY3vrd5jFGzy/NGZb/uizqs56Q0A
oDuxnN+XUCS2rqu4HE1FA4DfGZg+ddet08elRYnlgukIA4+rMYrfGqNog7/oVoHe79RsqrE4KF2R
lAPSwo9ORcXls5cNXorlQ2cxkOcmUurTEvG8BRCiavs0NIcwKzw4R2CBlB0ZJhDVErxt+8Bqvyhg
Biqgqb9RInE49HpDWvxX1td/8v/cyPbjwZXYordK+n3stTRiViMz5yQRLAmZH8zxJeqHFF6Ea57M
7Uy/opxmQjth/81txLmV2zaae+HN9HtFOtp0ePcDSglytvpgubf102vyTgpOoZiV6A4F+a6R5jx7
zMssuTGja0kdeV9UOqWXc4HGGGjR71Ox+5Ix4Rz11eJyMHFA6U3Tccr2T9p2MR5D7USUeVE7yuUD
nB2pV+fcd7OPFya6KKtihxNq40HbV5Dqv5GODafwlxRjAlG9wyNMxA1hnMvn2VydsLThYTqdct0h
zzQxLaaTJL4l7tnlo+gl7w6AAdPAmricrvtgAL0rorT2yGkJ6ZzqKRdnF2Md3gwiOY42vEpkA8Vr
960BdP9IPdQTxpb6NUAperBV/qmS4Wz0rx/msF5Opwhp7mrwa30XM0JnCU4bJOVSUdZJBg0YPC74
gvHewYsWb2c/SOqr2MJ6FjTJ8V3sFc3uygrXDqY1W8/wDtBGVNm1CIbs/xc4wQJ1H7ZSvrhCj+Sl
b1j22gaW6bZx7mghdA0EjLLJ/lu63WzeR7Lb4BB3zvYVMtCuRswDJ5MTjj0j0nenzp4niwr+28AW
4P2SzgJ8FpYnfw0vEN/hhXwbcDo/l+gqvSV2rK9Aub63wgpzMNbtxu4RA6iASDmE45jwNARg8dvQ
3SJGlz1/QFG4CqzCKe3HgF4dfSfk+bLG6GUNHsCxlctKA5GT9wni+mvtj8G+qKFsSlpKr3GddUDs
FJWBBkVL51mHNsVvzI/cpfsk2SlfARpUNOvqGeqvKKtWqRcsRzXr8meLmATwiG3QApnZvRUlYUaj
twGMbZgTnG8wko17WBdu98G7jHWA276KTvcb+Tw+Eid1RBiBgfG8ImFTDqf5wpaPaEe9kV/NEQJB
cZ+1kC6J18DCmwS+fbZzVMhdKVOxD94BhDmIgwxDl2AjmoOqdIO9zkjmqAXX1SMykyISMwc0LJrT
CChMe+qgYQ/0ShN49KkzATcsUSdH3QXSAmLLtyU0BN4dqf/XQD/RQnwpNFt9kSpn8RgkscIVP6ss
ohy8JTEY8pdH5woT7VzXmi06lrXyQE/kV7q80mcRRBDGJGwSEMZlWUqySJE3C3Rz3T3cJ0hIm/dV
4KwgR2xvvJLrYUv5KWyzy9pjZrfvsDSl2PlP2HZlkd+la3QnvrH4VxW/cl6iR92twQfh5nWTMNEp
Axxl/iew1z4i72b+KKetjqlXD/BHl0wcNtbcLX6hBUxrZgHeIp8XI2r6Rt1O8KtDuVJ+ci2+t43W
IOHtMwiH55qqWsc7Axd5NK27peEEGNR1Pft/xxhP3+/2xYUJE1jS0o8cJDRYFXQRU6x1H6RrLk5p
Nhkps2D2d7r9n0Tf1D95OKlFDHd+XaKZOvknqSSKPAPAmaa5gTD0JVUCfLf3bG+p4vigbNV3dI5/
aoV1V/rOyXVKlXYpHs8zJ1OUTGJnJFYT/T+ynFxUp6qMU5mq6dVg5uYTeB0Yu+oTRIz+vxA226oC
ckFIPYmcw4lYkEpovM2RPILTwTpTo4HNG6De91nH9KfZhioj+eWk3vmKi/1WVJkaUFd30Hgok8Qz
BhfSiYV3sEMQbklNMspIwqt4ul/ChuzCduD1Uo6IniiLjg+TPsvM/Mvqyl2Q1B/kxUqkRoqR1SgX
ucXuktsgt+JodiOOP6FFWS9P07m9PZ3FM1gMSZJiDlZDi4mfjjzEcdQKKpABM19TWF6uyQbES9N/
MlS0jtQRvjPYz7gpSpDualnPIOiWBQbn2YWEkhXs6kho1ls5kuneT/qYjIre1ueDB5L8oBnH7Ua5
XPWeovqDb2XCU/mWZ9JnjWEk61uQzf+/cEU5OSkL85L3DWXZAG3z2izF4p87iZ+0HvSnujmkd2Qy
xFIQGLr1xYFXAfcPq0Wh1jAjw+z0y6TRUOqWbd+xfl8L0090ks860qSDenmWbLBhPTeAefo3Ejkm
sevx6F5JIM0tEgj2pWP0szm/+K/uT09y6EorBvWs8/rPjGGB40OQYD8MPJcj/bU20jdUAwyffk7p
uVQ0UmoXbwq8cvpM8gmiUVlqv4i2D+/PD2JH6EC72kB0U9IGVnriF7osSu8buPaEnHP3kgP5V7Gl
dX2jNmPi5TKVkuFA4Z/k26RNqatCLAs8SB5XIkoFgAm9Ku4RRWKGxTWH9WBXLSQUINzEF/6lCtYZ
wlTVVpLwG/OkbFRZd+WjGo+24xolcWU7m9BBEzIh/6wu9TJfdPcfdzT/rp2ZzhDKSw7/cfwkXHiG
cmnYO9Fynq3DJv7f5gcgO+uY5Jewg+iQLFeNCao98/5Deq3BX3Ta16Io6IJeCL+Ukg6570VQ4FGm
UJ8yKUZoaG0J5s5EOz8uMqpFjPZMssALirL/9GGz3BAatNORgQaBLkS5ZobX9mUh3uS2jng8iIes
Fu+aZJwhz0BV67yFrEe8F3RSvwoFvwNNlw6jgkm68PHwQ4Bas04dhBfcrmEaXuKZ3BPuq327Dyhs
BtAVDDjmBpUh8f6MJKVpTc2MyPAwZAPpcP2siEWbdEJwESqLZKBPVm/eaRFXt6aTByYCDPtoxuPa
bEEqptlhP/u+DKbTZ9ewqk8Jjxra4OIaNTUDMcCyjS7j+E7jf1Bje82vC7lc4EveU2UZLt4QEizC
ennHQ4MrLTK2i5KiCj7KicwfdKdg29FzwzIvTCIvdCfW/hk1lNQPNckoEXxJProfDCtXAkKlH7WB
2EXDE8XBLNEUxjDgW8o+uRoWFlzMxnLLJ5WZiPOY42dxiNQMKbzdSc5yqSEmCuU2327LhU15IrHU
8ApVhCP/fFrLeNIc/4Y5rW9rkt7wNFIVssfKKxVI21kPXggsWhAFVJ58CwzTS8TNLPCEWs+rvwEv
xagPrjNbt0XrqfOz1Pws2JhmghXVKNNSWWRqrDLxQNANnFMwwbHWgNeh5HmmVn68bvu57wLIZK5T
hFh4B+b9CTMUUdJYDBVUlScyLuDGraisuIRbUhYGdSEl8d+WP5JpPk85LNG7Xu8WQwzCIoPzegCi
F2mT8Qfc3ehJbIDulcpgxODKrEh4BHmo3kcuFv1mjc7iSBFvG0v1mlLUPFTuHzP9xJ/imSOSx1mQ
JMLZnz8SaiJM1CJ4mVml0BJlSJCZaq1T6jdk/dn2EcHRxgcrPMjtdKimWgo+Bru377NtZNI4XDpP
uiKG758QPV16vXeqSxgLYQHrtkdeVyJ0YrDa1lhI54IU8qvB5LjCdJrEVLVDSOjnT98e0y+a6TAf
2wKQoN3TBORi9CrZRKbMrs45U03uhvvGe3bW95WX2axbMOQLsWG+YUKzSmX1fiq5Y7J9CiHh0OdU
ZjZhPOcHUX1et14SyGYK1yMh4dnVHRYH98MOtSB0bCjnGrFD9bsU69RHCbV6f4+F/uD0LP/C9pH0
K2ZEouWGzim9EAuKLqVkFQF2thBVFwHoDcjNlVL9klaEZtlVez/IdY9NApJdd4iEu7J/Fo5OFhHh
Zwj9AHFKTj56YY6D8oOhQz4lXctLep96WDHP3ZMbjsW/xD5pJWUftcHTKrHP3bYJh7lOPsG3Vf+N
J1LPp6xaXBOi0/8ckMJKSMDGDIuPJyKl7oKPPRXGG2A/f2VXQsUCNCH6VtDS8zg1ZlbYmAP8wEb1
yvBWmkNrtU/raxoWRrilhge+F0unzZYEdNupvUHpUesBQTkIcxtPkmAn+37idVF82JCuZUp9UDcL
PuB662SNUfCNMT2xFTcff/w5y0dj7HvK26aDJrEelUoA+QHD32H5bY2Gq+vLC4q9XzilJDQVkuwz
SmQcQoUK89ksHVHRzGRUw75scy2r1tWmIVPXhH3G/nV8vAfUSGhMSaLeQZV4lr62q4QJUbEut+K1
a9F419WTbTCu8gBCyF8BAMHj4kv8T0suXOox2Csngiw+3SYx8XxFQG4zPbGNGKa7fJbwQCQPji+n
qJeY0H165TGvMnQ8acLiNdcR3c1embe0gakpO5F/00Xd3FhYTA9QNb8ntnXnmpi7QYyHiq7J96sn
AMpChhOTkyhl6SfaMPq/wuHeolUYWhSIidOZDP+/26Z+Nl+QsL0RciuoCO+DIiMbx5pws+a/FIYJ
iIiLgNYTeFq36EZBQECTX/v9ZeuR4TVb7l+eW9oUogjWb6K3AxoVOGjgdwB3RLGkBGuT8VZQ3QQr
FlWYQRnpXKpMQ3oLtGFoW/y0poxAqZWy2xRM4J/KFZ0i4onGqt+q9MVUQXAvvz3Fkd8d/icZxzk4
v/1GChq0pVU4uDQW25kknWsVHsWxSWn3UULqpDCxcAt9Dx9W51SZTIiscxWo8rpHPbAteIRIJNtK
xKyFMNm9+rZE4aPTKhnobrIZh3r6Os/XXWkZ8Zab+2z66WCaGThBplGLI4pVRGT2a3BKYSiIf4pC
w6Jv1pyZxbpciDm5WGKOVq0dVVZVQRtqMnIhV44Oip+DqMx3zCaEMmqUiPPA/8Cmb1Z3ejP/6Pty
Kr13TMpmISoAyrrn0yXrbKrHIfnb8MiH8mPc2q5Vg/6HWf4g01vQ1wUgGnpmlmMzCHJGorf9fdAq
/YIeSzsmOtOGrEG30gNW6ijPYCClL/bmMArD+1N80iEHVK8BJo46RDLE50MLqBMmst+KFwn2XjXc
e5CqC0xndwQEYkY07EzraFh3iJvtNT4oEizUyOQBmjFQBxzj+Tt8WdoX6VYAllmahL0JDNHa9LVH
03c75Q4CownH4caHFABLQaSciOzZHdmGBP7PPLvsIIU+jilfpM9TLekAWb5dnCZzSqB2w1cLYveV
ESKZTGckbRsGFqNNiITRn57vAzEXKEJf6yLfntYnTbNwoJCjh6FNu3JWp0iJ1huUD92HDvmNBehs
FwQovfOmewSvulEWX5Hkfw6fOVapghLWgqSHtqdOYuh90ytZ6QutQiRRUW0Jsntl+aPpu3ij4LWu
Af4v9AKd9ahiZLfAc9TJJaS1zML1qTS4LHLNDuCkEhfO5tIWCWGzai0RyMDirM589nNQVhJahkwr
JiCrE3Et2Nomg9+l3n3BNfbu21gNEWyDyqDULnZPLh9aH60As2yopnhvBAUKi+TARfKfYM3C5f9W
RQ346kEg5gIJzkmSYz0l5FN1FlMWvjA72Zrp6sPfKqIIH4cGn1i2t4VCGiHp4GnQRWwhL3us6/WX
1dEJ8BNjmcNZbzwgmRxf/M7I3iwWt1M61Dj0IMV7uXzR8Sn3kcCcnsTb8TUNNxHE0dxgQZLVNt1S
cbqEASI6QMnT47blpaRMnjnnida3fbTVAC16Dey9bV49NwKrnZT91SSA3Qf2bKm6YGr1pzsH4Ujz
IT1xY3L/PxnJ7p213qLvfglVTrKDnkoohhANZj232OleeTdVIRrPu1pqgmRiroaeFuKzwKKjzr3J
v4NdVbpkPVl3kQB++UfHntr0rv49nx7GzgdHyEjpvChde3opeHmEXXYErlrVx5XJZdOYW/Rp8nKh
iljtCISxKe/Sijho8vX3xcMzrcIIDHhkKcSDk0k/0qGSSoFG7B/GRX49dJnPEqA56ykG5bgmoeBc
fGt7wCAksNYt+ruJGj7ZkBwPwSp0IFwvoCZLQwZSxPddrluAn8l1WTPmHQGqcgOaqw+aH+rupHD8
4eYsZKnpSrDKZZB9VvXd6weZM/Rn3WQd0jRXFrC0C1rMLhM+1KB/2KRFMW7yxIjeeNJ54MJTB+Nk
BIjEsOi4am7ZJ4Yyzd+r2m4mNoYyGG4R0oZ48PfZaWHZ06k4MTa+RMRkt5NNdGwUvvMIkPWCKZg2
ID1TL1U0fINXhTPqSEOHoj2ZJUlaJIPBuKOIYhl736IC3p9NBaR2YnLHDzU0gyl57WVlXZSTQSaG
HRrfv6oYeW9HJjUoNvKgoPDMqNn4ZR1XBRT2bbKl0TwDvFAEK3hCMJDnCksg9Gk6EiQyZ4LMH5JK
uTC0QvnQ1Qv5F6iHwKwuMXbnPbQcDJwSEd1U56O55uM65U/8dgQ6o9pX7idgkvFtGNc8eWNGuFzl
6JEx3mtS9Z2ks8ZrIW2SCwJrezissL9zxezfbVuvmMGKYtVJDgF1Irf+Zt/DvdvzEciFfHXTF5Ft
DO/juPxOG/TTNk69+1Ep3Byuvtn3wC73Twq9afnUaHNctyFvWfQJcgCiJjuCTk8VjZSFnGWsWNte
3KutAEa1tg/FyTk2nRLkAVAVcyficDMXo/W6+yP4k4LsD1BhtlZ0qHrZzxKEje9W+F+yJy8jhFrt
c0PoITVRHY/d1PjAyXKHu5Iv23E/emi7d/5Eq4/Mj6Pz8EqtJJ46UtE8AV0LEwwhQBWS+A1m1WQI
7s7qUEMYjt2gaDQfDh1Ymbwxu2LgJTmfrjymV3kbLWRdXTko89MCp/9rXNfFipS98nhoth3TSCpk
xD7q40MP7r/ncl+4FgCRDfdirWpuxhjmkL0sb0GZawBb/216/SfascugaN9nXKGUJTQ17isYoA4G
ZmGSVsKr7sRDmqmJq+A5v8aDrYDGojq2I9xOGxh3mqxPUd/+2jyUfXD63FsnhVX993UAkle4Yf3R
QlYsqqK/uD69xy3jAz8QhAvjyX0PvpRL+wVY24Ifj1qObgpjoGVKckxXzBxVX1V+uX2rBijW1gtd
tpJNUXeWIAjYoyyLdhF7rjCvwdMOyg+WtSJ3F64BWzPGKbARDwL19f61Vnh0wfWpU6s8bNeC6Y6l
BbP9bwfaGmhgEVdCEQGMWc5v28US/uWqz5EX9vHgRJLITVBggI/2ZqKWQtVdr7Wn7ENuBEbH7ghH
LPW1aYg85L42uYcWjuGcsI8O1fjBtOwChSn6Y+6+KvzHd4ARYvmAOmcpriHckEaztV8GfroNHDY5
oohqYYXqjKb7fvS0v+hSz9a68q8u7P+8QZDlxOswNH8R3RbDBTr+L2u0mFG3RneBcpLmJ4yibfey
yeqNY+OgzwyAe6kaUoYzxQ99pUyAL9tmqc8JVfIJ9y53bjIiYXB7yFJaslz6XSyO53zQ6Mp2MlLl
BXstyJq9cnj8cHdToXACYYVIJGIsg8Tukvle3Vg4/oetcI6Gz51d21j/1wmjZ1GB1I5byKbADyyJ
TJpQhbUZJlN7PwqeCzO6KmbXVZVuQhOf0gAtcvHp6EkeljuiGoNLFyCBVcaw3mU3mgEfeAbx+cXf
Jp8mbfAwy6kTVhYBWkSczOXlgRDzYTpoXPXlV64jWH9jLR0pwWdGkSOeS/DIra/fOD3xyequ839i
UyyrjjNQJ1fQ91efYOjva785hPjad4N0DFDE4Y+J25vSRVd/wG4srI/rVqZCeMD5JdAnh2H2mp20
fUY59BVwW85RAuVvl9JbMcEVOZzEw0xt3lS9VfpcS7fURAdQWbIeSoIWrctW0CsTT8ItCmx742hl
pPCMOgfAZvakQprJSYnz49XIW7XYKT3tJ14R5jz7L4e2aL29tcEdYCAjWga70BZieljxvDXDmxOH
FOKv6EN3EE1Razw39LhtXgA5nEVqUYDx5aYGVq+TBh4JS9JVKdK1GX7IwX67qDQYEF4VGs6VklTO
R4uBAuq552juDwbcorQ/lMU/p89w+GNqmg+4YjTTmtI7PpHvq4GmAJzflH9ekTGfxquMy2K/gKLE
ikn6q+FTRDApLMD4SIhLEpNak6YgnpBKnopLQ7yyIHbbvGJsLtHHSBVswC5Ky5vPELiA8+V7Jv/r
s3nFcb34i5MLwbFiu59DbSvxkhC5XpNQ/mQBzgBYggmNjK6yRGfeRl3rgyD4H8HP/zv3R5ogc44H
7jACz52G2r9HEuX1lJlq5qpv+ZOLdJX9LWDP4sqNdKdKNLbGRHNsOBkYh0O593FBGXf8ePdTq93O
VbFE5XIKrNbDkuHIpxFSxmtVbT7Hkl1rLqkkERU5u2OU3vjKoViYtP2B9r031UCrZX6Xha+VpA1W
PglUH4SlzK1qSuOkExZUtEt1y7hRxeiSbM7KMSkmNdof/hHymG2zAccxX1mqQCzgj6ZltpQG5NUj
1fztlBobFjD1PEpXY/DGmcawiucaieZxZm7quTEQSnmeTTJ/GFApG9APM9WMyOsuavDsqxMkoidZ
d9POItUWF7Xa39eEK42cj8TzMuHy+RBAQkouIcgM8RYCVqlztH0cpUOyyCIc5SDZuwIB4dI2nufM
rZABIDrdOiK6IRGQcu17LouzgbelAhK+9L5nkZm9HFEQDMFzUy5puhO/xUsKj2RGVKjhZd4FhTpM
Gw5GAnuKShOYqqJweq+yF6vv4+SpDpLwiAIOjaXHQMBX6w3/TuX4rt7v5pvbnQLX2W8kSJ/yJU9B
DpUEcFoITqeeDbjuazZPVzCenE3cf0DD1Fc8DMbcvVHr8N+Qug3MIZBdYc+OkM1bEJDMHJyjQhNi
fTN8rpatpoHr7Auss5k+PdbJjftNhDVMoNaqc38ES3H/TlfjWrhbxEjzin+F+jhF3+YnspVFWEZf
d4Y12pRWxOqiJAjSrwbzGrusVgLPXm1JF6l3hVNpBYIJtt4Bdfz2oMKe0kYZZ3IkVtuD3W2et0BV
pePbJlPMSvZSGSKU5Q4coS0NCzmLXf91Nrvq0KZ5YlSyPwc52i4UQh4vTK6dty1xhAHeIN2QpwTA
aKNwy6THPvIxHXe0lw4Qlp36A38gRTxX8mlA8jFqJpSOS2VXqPUvD+phFHGJus3cKDy3wW3ecrDP
AmvtrCeyl9WrnMoujny5D7YJq5VSW5rlBTr/tQfv5RKLaNpSAy/xqLaiStR8EBRhT7wDqQBKNd0x
mR3l+7gWuRG1Sh2RFUfxGREvoz5qeoHuxxPbkQCzT1E+JMvNz14kjDkbp7c1zZ9Nod8HhtSP4llE
D9iH8VdMy78fk1o/M+2rf8v6QVErsZet1mKHLRPCc2HEcAm4Y6QEDsqb7zVgPhziYfGGZU7Uj/1e
XO/0x46e5GEDzlTja+ZJkHhFAt2xLKgpnXfV21Leq2EW8btYKRU0jsg1M68vFmaRNqKkUFeVE5XZ
Cid0js/a5/KX55HfGpqd/BomlG6esD8z+wveYVwGyTRVbgqlrWYTAcPogzG08jqrlCpVPR3w2bX2
iuJnE5SEfgwqaHyVWKHnMaCYy7mTApiuyFiHkPrmcY69/4StN2vDPN3ewqtndIUztbLavL1351nJ
NPesJOuNCrKl4m9YkBMwP1Z07SD+Pkhv8flNC/tzUm2Otc6S2uc1njBMR7bD4oHkc7l6O98kHb+1
iuUWL6nUCEdS4e0Lkj+ndxDLZh7pn7LCy8RjUUdcWOajgrUwgeqjtTp7ZmJhREbispx+Tr/xam6x
Bkpne1YEnlL+uBBZ8aNiLBG7NPxyKHy5DDJ+du9VwpTEF1ZiIU4Cwvr3ycN5rOAx9/o9zdLeIYrT
Ny93XSbpjaooLqzZHfXJ9NYoj6iySb3wt2wcMgDez3Cec5HscctwTTA+xZRj8wyT1gmyoH6jJ1Bq
Yyn8Iv9EB3cuWLDAzJM9iZQUDVq5iOu41aETvVQ65aiJvUjzVD2oD7FbAaaKTb18NPyvNwxz8DQI
ldLr9Tagxt3WGSCFGPEYt9uryjW35zFM/hJvPsQalco+PR/UdxZfAlJuGKdAdsniydhF0mYGdjeS
EBxD8U0yJ2vJpoGwyVsGlHIDry9zcOBMfbcAZ1+yx0WIS63JUqogzSeYX0mPicnogYvp/keVYYLF
vHEjnYLkwP/SpeRG1vPb5Zw09nvP5E/NtSf7F+xRAxyW/C651JmqbtONa8Tb1nJVlJh71GY51IG2
4OFO12KU8Fd77N4vwB2TbNr+tN2bzSzusMdLWP6L3wMT8NwGEWzDqAGfkBWDPqlAzeo4YPpVU7Tf
ysCPU5yrYhO/dPyML1mHyWF07hUXN9DBUfRYc8cN6QcLGKqpmWTG+gxmjrY+1+YibWyb1rAcSBeg
Sfa8Wj6LlULc25Bs91IbM9b4dUUqmvE2BpPzQAYroyTtdiN1fcysjA0nP2tVn357fH5SszxY+JDP
QVLU5jxXUHi3PGeqByEWwhqPLECQVqPiszamUB8ZRAqXeiPAeXABDNaMqKzZQIHuHcyRhL+YC2HT
ecV+0VpfRoLcToxJQV7TfR6XZlyO+1Hphmf+2g95Oj/Fcwnh5pjkYswRwc+K/k2fEbExBslwB7i3
EK0X5hHUBwMfogUK8zEYbjBNimVFfC4Rjp+10ex6QcNuVEB7p4He1/1kWZLmoxwJd5sqihQad4+g
Fn0Z1oDW3cqAx5DmDgvvNPQMQxmBe3EwbQ4FesNOu6jFSZuAOTzhVyDjnEJB0A9EmHO+TkkjmO+U
1NwhATJiBKhqT9RfVehBY+FZ6eWY10vrBA+m0AjvqO4Bz0K6Xqs0Pp20l8Hhopg7K5XUz0lLTLN0
AQTZpZ2ZmWewKsSDta4ZYMaolmu7wdDGu9248bFhTQ/A0eJkzhjGeKmDA2R24wL+XGkNIY/RFaDV
9/T0doBOvtcGq+J794hf/Xkz7fyX6nBptz9cu7aZM+adg8rPl/NS0v4c4MeALH5plFoOmZSdP/Ks
I9AQsKFMaDHIgRsc9Fimhj60bcsD/Hq4spz01eLBel6n2k2h5elPeSo6HzWAclHpBr2iQORrVTtg
PzN0890qQp+nfbGvH1I/w44mhFZdWa4L4aBFGZT1szQGg5lUle1yirN2aBPxIRVBf0z6LfCiBbtQ
1NZGut+8t3lzdXZe5kRX/wZlmOBwP+c5u+XRyGErBZYwaow+UCOwmTRqxxwf8b+OWADtlZgLEJTo
tSak6ezDqXupXrj82PGp+np0yTFtc1xmuUwcjE1olCwqGTczoHoA4TGVwQUoE/8QmYK2vuqzwEGl
rNDaAAz1vduCwvECOV5hSoLGkk/3q+Ox5eTtueomeshZ9F5dH+ai/SSavuu9nhFnZ0SI0SDGqo3H
hk+q1AZPEdOuRZ0y8TeyiFuCUv/TCjEzaWUHaW1R4muCy/oUMnUSEEYZ+Is8IMAMBiF+tOfFXxW0
PWKk8chYZmzjdt9B0BWz0RQsIUBy3wxxd2thOp1qrEmJQwboGGbSpKpSPpZtx8mhxzPFeUqH8ZHK
YKnh8j1zXQh9h8+WWKieJJS2P689VnwhDjpkfe7ktYcyq32bfXo41qO8jnwk+LS4qSyZPn1m4Wp/
W1Rkev6LwixP3beJPGgrIL3I9mrU2aN9tjR1iJxxfPxrg7GFYIuZhTnTsp6yB5E5uAwm7/kqYSdB
NwzTbIKAg8/ct8YM1fj0aR41fhqHEa07FEEahJcx6JPmHX+s7Q6I2F/qypRtOmVY6QxURE80NNQm
um0HR4mO+KK3Q293nSHLRUogEToiB29lL6Sz3Ftw5fGK9vUfpRqdsATb2IZDVXh2NR/XlyboAQYK
1kjr1YaMND2Ph9yn1M0RY7XLrA/phLQVcObPH5WDZHcSROVvpHdD2YcDTEJmlOMR+9IuA70NPWmo
YJEfQApOR0ENEhxuMKGO5oK/D50rT5JlzeDYE7hXqWkJxsYKbJg6uIsON+ENTaBTxFB9sx51uiv4
inhZBH27J2xQsiXqZx2gAenyHVqlzA/WuO2gU47+v/P6mTur33THb0GtadcbyXd3vc0QHaHDZLWg
wMYpuo8d/n8kE/k/sE8a8k6bhM0zLLdF37D+kuBAC4N977DmzRsF9zpOQ6FCSiPOzr77PVU+EjgT
bh3Yagq0mn0UubtyTFBwGX/v6LYGlebSa1OZtmxqH+6c1lbpWtq30d2vrPNXQPCoPTpMCPVdPrwx
kCJv0tin0M3vUqI+r1pltJ1YLE0q55dnR1/3/WvezDL80Xy3QKGdFtT7QiqNWg3Sfrt55h7I52tK
37SX4oc9gG6SNWMHItz7GY3DBFntcss6brEZqpJ0LUAUJspjgYmUpIdlurEk5f9ewOsA1dkXnofG
hRFmnz98t28XFQRc6QFZsBMFxY9GzSSeERmnJ8SnHFYt7WwI5jXiWbh1HfNDhFKko2UIdd4ECoeO
mk1w9nUdVPt1o6FQYQGM9E6xzytmlh1xOD6VbhwDYKPUgpRIRQ5mMwi8Wj4ltm6yN60gMmIakuOe
zgUiyUxo2jfPTd1sMacX2nxY5JhvzsXatUX9BG4MLhdu2orNUL/NONXhhBVt8R6+6u+7D9fGQkPh
Gbl7MyL2NxJeimp9KZjENQRU4R7aH/Kgr8EZfyAkNICoQRRWie7o740STHIXlBU68NC2w7QoN4ol
NnILE3P8vk1EwTeRqRqI9veAe+8vijhH9KQytEr9osMCTe/hbxWGAfuqHtmeAodksU6LpgCQyKOg
EYMYv31QB9JyhP5F4Io3dAFdMG8aulNwssv//zY74urHBKY3T7ErGQIfZYtocfgBueChIrQtQOfm
P5v6cS1EVuMG9m4LGJOczlnwTpNU9vmF6G223x4caJ9nGrh1BEGl51+kOSMR0+kCuolRPeI28cV2
Gt+zl0Cc3dtg4S/gQTNKyONXlDyTu5UE1QGc6nntV7dBJdhSokuY1+rZExhldlT48G2E9gVk1JvY
xg6e1vHZVZldB6HYz+KNOwpeqQ9FCqvIlmhbkJhd2zewL1Y5HjMxkhgMif49ZMnx2OvcUq5nhY4V
JKeIMVspfAUs+MtIh+UXm8yUz7ycrd/1eHMITxtciF38NyFH/qApWXDa2KUFR2IE5ZbCKQoH5ByO
KcGglwXNT5OXdzWv+Aua3/BuYwscKlkGgdyYN/hx0Qv+k0PL5kHzexFdPulqgG62Nfg7ro/gAzrX
j7FZaTqDiwLSusaFKtKRVbrYmI/xyuqwDpaEytK0vyIoMLoMKGi0jEn0ctCQxSFg+O9x/b46fCaE
o2k3MgBtxFgreS9+JSN6Hwz03xqyN3YPHPhWv6azL/4vxM0PQKm+cCMyuKDgdcpBBvOba5HHF5h2
C6XfIfpR7KQd2yI4+hQ21oh3h46p1DTN3kYe9GMvF93Dl1xVh90haOn1uU007WX8ktqo13FqpMlj
H5Q1SRlumxtt0RGF+2b8tYAQom+7d09yGNyY8K1kDQgx5cdbJkfsh7UP6LUfF7JY9Ocm6DWbZgrG
5MUviXBQvbFu7+RIdEue6HJhCxRFjU1Rzz62G99FPWHgTGCtEsP+tI/T0I5XGFMdqYoOSL5Bmhk1
PtpqMIxuecztqY7FJbh8eZxlDh7hbyChLOCO9S6k5eATrbXBns4hzOgfz4ZBWuBa+cTtEa7qQjJm
7AAS5TR2/104PnogBJxERlYKQC5mGreQ3goXhJcNQALDzEBR4auSHpxscxCvQzRx1I7tIKpYT7gD
VkNpKKOPUlyanrK1B2xWpojdT6xUARb6Ba+jqBgKzqPi/3BY4q/A8T6ccXyC1En9zYJrbw2Z/u7P
9pM87XRHTLVy7XUTax3U1gRW3URVfOynNrslOMpBcMDBkn1ShMoJStUExpv4M5KYxWwMJZHHXMPg
MgmdwAE9e6wpwJhgkySyfwKfLFikMjF775HZYHfXJW2iKm5NJwJW6SttVU0hip23bMDIiASXaMAH
vkqf3Tm2C5pmZ9bByCfwXdytZBv0fjGCXwcSXDo7pcDetF0x6KwuJKRW2j7bEsM0CdoyE2wgJe1y
q2KO7I9LBQZBvyPoje6yfN2W9UXaekIIAO1XiyBqU7OE0OAAeLErjzOVtZrSZu6OfY2/qFh1+MoO
rCNfl/Y9y7fPmlBpb9L2LDAlpFa64y6QpWT/lAcwKerk2S5wqjX8AKBqlgD7Ngn3Rs3bGAekPT9W
yTiW/QXuVJj3g7ZYsGVr0tQIA+i1EQTGDrl/XavlASL0g5RSuZjgYt2mbBC3k3Vyie81oTkFy70q
hqHNQwNgfbCs3lmo+zf1TWHmZq4MkiB9tPMGLb1RIX8LERgE0Jdb9gkPr9ajTrBmr1fiwm8EvKrA
ByYaizdlG4jkjyd/ZfT/T0vNyZ+sb2VyUSD2/pi5QydcaN/3HjIlIxOfLfqCK09F1LTqOQursnBx
FN9JDEWjIPu/5MMxoEo8XjUbszahc9gnkGPA1AqGLw3A54dyKY1wmm9zK29YkMsvOC3X8oX/1CFd
a4SkyRP0exgg+pHIBrYI3URI59fNc55qIRL33VqBcZcdY6atgDVdz6wAymQEzb4Cz5/7VRbtWcjZ
NeutnnE3xbFuVDoDFI21uVVNzNQcn7OjYTGgJbEwsHXOZuyTbgqMXeOzLQDxRRp7kP8UplSWgkUK
rnt2nCfvprcsQyPKqgeMbz+toGq92CgfLrKnrQoP7rwPAy1+A2l2lpCnd4+Gfxi7uowgHpM7uclq
CFIvlGxbgMcBJpLPycTLisT60IIUAF7RizIxiPL7fyGk7/lsLJuofhZlRjZ4BPPiwjuPQB6Bh4K1
+u1B5oAdfZcKq4bmCprjfyO1FD3yy/BVwbduyTajBFJK5XOXgqwv1bk57X3LuoLqQz/r5YET0O2T
5YZnF1Sng7e5LS+aJP/idfA1p0sgAHGb1ia7E5r58LobqqwB3OTNByrIbu0IcAoDMZ3pacBzCU98
OZEWgHef2o4efm61pw+N139DQH5LzZLZl+igFykJgTx+gMvTOvAiGlrC7yycuCFOyg8Pqa++8bSW
I8q+SgRfL/J3sMtkrr78c1/O1QlF3Zmt2/WeAWB+TrJIHRErLbl7/1N9oWYaEOTlEvNu7y/NmQS9
tX3tBTLKAfDuFLViwG/+XllYlLzq9vldbS4+ZYVero9lcaGa2ywxhNey+VeVOoJmytyFmsfMC6No
rUCpNteu8wMK+ZBj5DNuR+jDEFOi2INdxVt+pZ2aq94s916n0rG41zcv0hhl9P1GKiflWoLXl/qO
ZM0S1w+RIu6DVCR0xMmu4OKac4yCQnZLo7VLTN/NOODVu1xZA81ccDd/mkyOyTNNJsSsWhjBT6ew
Gksz9XNhEXplyuS+XIdAyIftWOgwu4tsVnA87uUY2sAullsBpyR7pHKC/0ZxplZH3WHa3Jwe6seR
kKHFkh/2tB5VyU8lk2bhvl32V4n7ch7XH93G8rUIYCIB9QltSHmzyHCi21NAqDGO6VVFkk8TRWon
T3rocCl9Mldx8c1N/0AYAybEtTOmfaH0Avf9lBYGLikNZ/mM9pc22+9XkkpBs7WsBWxDL/lx2Rbl
jY2LDo2QY2Z0i39SlLiJQMYqe4AVeHl7wdBZi30a/PFsyTeoWWG5AvhqGBJRuRXA7PuYVQ7JYA6y
D4haYh4guo3FVOz2fVjynvdW8sj8VVw43UJce0jt/lFlxN2wJwI1x8C1Z60JwOMKsHYNKrbQt/pC
a/6O6w99Qt03kXHiVb6gAy/1Fhhyuk4ST0K7n+Y3DnQwt0q1VSEXiAXDuuWHuJkppFB31Il5evUL
Pd01KeB5xk9Xtnz3gl3jspvP2b021SqfOa34u82ZtVCjbXO1Yn7bYDcm58ZTeC1AyiGHXM8sc8nG
8RgjAUOz28DHR4ab7EbXtV9LxwL9L6lhUpZ6FBHpxRnbGeJ3DgJF/IvNDI9ax/yQdq5EaG0WiKv6
JcxhZb9gLC5CrxOem38VhDbslCm6m5rbLrE7Lk88cSwIezI17J+pVGY0TG7ScJbI7ME2m5JbXy2w
jpVLCZ+uQ/nm86BSVNVFGnypXE0vTXqX8v3BzLVjIBzI6tHfB8yangwSuN78vz8mhGJIISpJleC5
9uo+ooE5a2QOqXOvZgN1NtETmmfy3W70T9+Ult4NhT32koBerDbCxQDYG4jtLRcj6dwxukru6K6k
AyNQdgeXobC9dTjY11FWgQp5bq2NIja3Cho+L7+Kg7zb2nNirMQa2rURZF0i94FtKiisykuwz5we
fcgzEjkU+a+yWWsNrMDNRPj4SdXX5jcE16uPdHdNN8ZOHL8gglSpdcPNLfT4Qo/fyxJZ5+LFucOi
ftcATLIqMc3MztzMz7QbVjQ51LIrNKN4LJU5/d6cZcOL0Wfwru+jk+RHeIot6KM3Q5DUCwtOEuJ3
zZorODb+pwOgSdPUl6Ij6CsiMHYLdsKJxnxXWjwTgb3t2sG+q80iB/dZ6mbVqPZ7xhQtq33yF9Vl
PCtrVevA1Qv7zsoPe169aShlYq7DhPXWZW3c/nWftQFaUOHPj3LSJ1TxVaePumSKHK/SrD+X5Dtm
Pn4Dt3KTKbsEXRSsLuuzMIvYoUONOzZVFwXPoTVIRUv4wkwTd7QcZURHwl7Pi8kG0W0EcNdUpU5e
vXv/1dk0cm/kEc1TVP3NZn+kDVPKAwWNvdm2qgIIKGY2uZgnSlc4yTKZHOIUUCGHgQaL6wlDqSmk
BXqWuVCRBkJUJbXRV86azzujTj8JkrqwhrIF78+O/rbr9evVO4sAGeJzzILlR+jqYvWFIt29leyK
IdDLybyT7+s3BVoemxhLbAc22eEp5icOySJMxM7CTm+MFQznsGNryhrmR71BVf68adc+spwANNPT
0t/ZQf1MryyCvayT5g/bFmV/N7avWlVLXf9wYpIMKMaKcgCeYP51g9hTRUdynhmPYKOl6kpNdoLs
rvZ/rYI/or4St+J7pjrbgBM6XAXAKJkq6yOXXSEEksdOcQLYAPRKCExDJCVwIvKgdjIadPVxjdXP
bU0f4crkACxO2Rh4ORHtzHnlx0js1+zqycFxuFa6BxWL//ER2HUQIFaQ9usbtmJW7WppzmXQnp5D
sZ5TNuvZDIxbctamCIBi695Ua3iWiWvQm8NKau/KWIkRObgNDJi60WK8V+kUZf62uF3JXTRnIi04
48qaZI5kQFDec3SQeAWFVe5UcrZxUlw9QWJ9aQSjgUPSn6N3GH9XtrE+HQELQKfrwo2UYZJWGWej
KegsOromq9pPvh8iN8E6yjxlH3YcKyKB1dpWlfKDpHQGIIXsSLCpM+Hr8WyiwD4Ijp9nfZiZjor9
lfgJErVJ6n5dyIQDZaI5zknfysDqJadM4Sdl2FE9OcEXX5VD2uy3CpxD26cMAnbhNUPHz3Fo0VyC
sJ413QDg6xKO4PJofI/1hKOVbKIVn7riccB2fZbAE/BcP6pQgVliA0A9+AblxtfC4P+XyhjBaop/
IrwOZPSr4WEIgYLW3IVQdQ3TxHgOTMOpyH+0791RE153ziNbPqp//jKjraq5IL1oLcCRnFmw2jtP
5PFjar/KHJPlIuF74P0xJuU6fCl28Id7IBVhN1VKZ9sjOzv/vO9ajRzmowHhuNI+ZsVubjSVtV48
KTz4fSW/mqgLfQdZjknD6mIW8GLhatzGr1aiP+UBaIgadxhyvt2QR5NBxLQ9hhyukiUYlRc8IliM
UYNQ+pyirpmu/sCKI2T0UsmZlGlHalDtpHbUni8NOGdK8a0dDz3PnjQr53cdnjpbAdJu4gzksw2v
DlIzSqeAfy4RGy5582ziHI1RNYsf3ZVa4o4f3vr20B1WOA/pcuRtL15riIRppGn8eenunuauJ2mO
qRFAqarO0USv3R+V5S7hjuHxg62IbuRWoGdU62mB3K0eWbkcmuFcr14tC6fnPa44H32yfV3xGrTB
r3XfqGS/9opTl74UfYwIrQH0OTfq0i8hUZYMiUPeawDPJtSKdAQd9w2E8pAqeNFFTSwc7GPEWsak
5M+Re2UTx7RND89TtJJXUUU91Ar4litEyOiEX730dQnnD80R89Rvb6PNdetpxmc+Y1XzKiwQyzF5
n65yCATFuZFmanpKnDBGOsXqLBh4rd88KJIRMirS2XNYzclFb73TBrnlcQ9b4r2zkX/Cg3u7HqVY
kbQnDa7PvILomluqiEAmWIk7tW/Y50qk6vrPhU7Shg4xgf+KR+8IGBWzk4x0xyN+DJ3tOSq/BTp4
8A3GgOV175eeNbo1AjODVYjmJP7Lp+IJoVhTjJnuk9KRtDRZWhlWLty0/Bm9FSRHQ4UKnHOyrIYR
JDYCWQYy2lKutrn/a0C/ySuF4/GGSfZonDcgXjwkfez/O/66G6ShWJlEcb7j7mVGIGienlFtpTi2
Ihy+Vvjx7iXxI5U0Z5Det/toBCQVFMHUkEbzoL+WlLvMlK+xSuQGCZ0x3vsWma/vyDfyYl2Ok+rE
SwIoslwq3kNX4kJAJX3L8TeyG+y/9+hh8/x3hipvkT9uEEJjt7Q62u8YECjQ2YzUCTYX9UALIpcm
1jlkCKruChRjAV3aEEK8dgsSECIUP8CDAbFTPmLIByQ/XEYCEB+Q72CroiVtQryaSgAhbtzsU1kR
7r7wl32rLYVIx1RsiJpWBXIoDcRG0XiaQbgLc6a7BdoHjMkVfv4sJGKz0BJGBzYy6G+DRPDD1Jyq
dBtIQQvPC1mEH+jkS0l7zutqH5yThykS5+UpWZU2Xn2hW5ITsAFxBIYQxnmtW8puaQrEbrlrYrbx
kX+OSm3RxyYH9G1A3YvbMw+ol8hXhwa4UOOE7uryNZERVg0I4m6vo0TgfhrtWDmQZHmiHQMdywun
WqApUu1T7OqTMBrXV73LvMKY9PEYtPZDmy0I6LaSgXsjAoAUeF07tHOIQPK6Cbla65ak1cAKqi6w
skyVpSkLe5n1gZvEcO3trtL4QCq7HssFv7UkPBBuWd/CEs6X0+hlRG1oVwLhUnESeIx8w8MkIQLE
SJdbet1CzCd/vW4XLBmT3zzaZrVW9oU/SxRkk42NAUZLoay9uUmGtkCOah1mnLzBPmckATeWFlEx
5UWTudy9E2IoV8nKXhu7BDVPDzyVumoI3dx7TecDwYZlrzs6eNKFpz3m11VtoqEdBOuTkWnf5dQS
SSN9VffLeCfvdX4HDKoO7r+JRpY94QfJXyGvE1mgYnepFM+3tG/pxHTmJs6o32dke4xevojAn75m
MXJe1cMf3/E6CsU3i0Le/8mcrQnyjIioFl2I+PC6ymwYSgIQ+00HrJyvzXTpfUgNffeU+GdxN0GT
/nAl9KQ+KBdIsPXNMYDacvs2MZ6d/d0THhD0TfZfeaqfmtljPoBWmv1VTAnyAmiLFJXSDa06gj27
mXzK9Ealnc+goRIkBgPJ0wkZzkxoUZlhHAmMoou07s6tjpMOeXk2ipgD0T3seQR9kzfuG76Vzx0W
XdpRAf39HZlF2+HbwD8DJbjO8v8DmFDmC6uO0fXul5b9QcrVL3SeBXF8+uWisu6/vktYz1zobsO3
/rcOP+bNH6FyT/b3TBYLIfszVWERttLlx0fxSivR4mVh+pAhY2vu5Nadg/N5wO0P3fhH1VYrta26
frP6tv6VCfOSbvz3+DY4hZtOM/qrXy5S1TcAMdgUBgHWCaFBHCpho9GjgeD1DDHcR/ImzYp8wqor
QLjv88pSNafNPJSanMQtBvYqWkv2jq7ip2nxeSMeHr82Xr9OHhzkkAP0EGJOBL2CbgQpwMKCzXzD
7vJIT27/IMO6TdwiJH5yrj7Ic6SCSm0x6OVmiEcTWw1/k48NaFeSqlp7POxppsU8npKaNKNMPmDE
IElwebL/19k5u9rEWcP1dQD/FALAoKlVAhRqux5lxk6/AP1so/GpbFX8EnD9ml8Gs9bHnyW5XM7r
gSCGE21a3RKsigKgjYpQaTvgQgT7lzosOFAurveKy7NnIK6ja2rMPtZVgN73P+pN9twQ9lpOvw1X
zh+YUodnbMUl2jT6bsKWRlmMs2DYqy9y6fsDYKlifBpaGIWkqE5J+33Wpwgr/gNwevSllRSfrvuy
TqT3EUbICsTLbw6XEPcX7lwOLyn7EclLvnFOjHNV3Y9F6ZgYuZ0YG9kt/YoMq0D+T48/wOmC9K+u
ufCddj+bJlsYXRetkVBzK3/VgAra2yH27mda8XrMaDi828hauCG5OCQ1AhkPAv78c00VI8sWqn45
K5ui2ZrvmmNYJQlwY1QQmsPLvN3QrUj6anto2Aga5UjJuBBA+bSG6jh1kRJy2RhNAHLKfHVbXlWS
t/fO1Y9uee1T4RdyZJWIUeiibEjLmzErdenxCJ8b3Lcx6royOtrpCmhTTKvZLaK4Bo0gy6ZJ4QvL
IeAm+Osu6RTiIfnxJJF0A6Jvr0WIZuPcIxNbLRWOGKpiDJCUzW/2ylNmpfPgKoxTYtq7cXDjhfXI
2Rf9Yr2nRZ57rAf+jG1gVK3Jff6rotIZQhrMkC1fxpdDLD2pr5mntQqrFUsBnE5ZfyLTUPpCjLX9
+/cnxe1wCuZ+MjrJopW1K3lhzB3sVJ8fq647x65NnmIZ4iEZ/ZWEBeYMfmloy3g4DT5BaeefSy7R
Rcec424Bf/Ir6rnaOcde6zoPLKF++j75MMx7RD0FzLWkk3EGFzV4ldGfmGireZbG5Narltleq57W
+YN1oJjegFO7j1QnfQgGL+rQDe8XYKKvSRT8CgZe5GOB/KoNS0jf9P4M1m7wlmzm82eB7Z40p9ac
H+jfQpjBFDRDxeXovX9Mba/O+XONctWJea2hi2NJbkrv4bFunSlN9ITyUD5Gdv8otIGlu62Kamlm
HiODpYV4G51B1RX3UMGwp/nS+f2UXIDbFhue8OQm6roPGLP1+TBqwJl0nRZekuLo2e1kCNKBpp8x
xthbU48Q26prFo4qpKcmpdMtxbii4eAtHWKXq/sX7o/+TsnPuWpCroFOcsF9BZRZk0uCGFlumFlg
TnOZtiu0uUqcYxtEivm6i69+imxnL7d1k+PxtQcg1nvBsmUpeZ+tPLqlxtyI2d4KuI4U05yYo3uQ
p54gOeHd6ROToG6ELUJlDxFHDIHLAwqZLt43d7cUSMP2hmcXLv4Qr1RW9cgAhDtEeTub4SCR/iCY
F55PyZ7FTIzrqNFTnijMuQkleM25uARafoX0NFtvsTRdMKd5ulfif1H706s+m0DwZ9nYKz/C9zV/
HTEteU5awD9bNSH/We05iUf9v1GeGxVmmYFZj+DfzZxwZDTtlqo1AobpxqTOOPR9cBGWz6sFsHVK
FZlFb6Laq29J+CMq7NVlFWeuCGskX6XabOq7WsiZqzHmClpn9xO4ia1wlgG4mYw1qP1pfh/QpQv0
2YqUJzE7kyedZJE/11U+Gy0PIsIkHH2rNug/2FOqH5NFY4EoQZ2uUPvLLS3uwZZe3/EiMHXzA/VM
7LkETMQ1nCpOO5lihjXSeMfWmoGG05HNg09yr/gP9lJFb3f0PhwqSzrppgZjadi8hrBT4HH82BTS
KiNfKAsUi/rWeydrUCQDFujNTiRIAkgYK0HeQR4B7pVdOIb3IBHz7O8wUgMpQ4gnb9wWVgo/i/+p
TIEEvuhGdOXM3g4HvPHYE8B2/Q2ttCHoF1FMVqw6mT738C9FQ4pvvPnlh9zyVxwmbzdIkBE90s9v
MzyqejrdOxfhMBv7z7ssqPxJHWDN1747JmEd22dePMjdPIOox5yX+3/EP0CXQlH1hAIrIJviDJC6
B5fPCA//38RrE4R9Abnkyte2PAMVe+MfxPA+iOjX2A0W1nJQ1WRp8EdJHvueyBdflZLhtFImQot4
YxWNk7JvdoLWlxAhu0T6fMCyap8EKYVFZWTIfFn0w7INxuvSbAdhSN2b5YfndnDE3C/tal2/gfXP
0zSQdcwMnVORRvUoMroaqQTyxecA+VZILTY4LeuH3Ba4LfImA9TJqhGMsXvaNTYO4ZJ2eJIF2Xzn
0kMrHTFBeKs3hQyPDhGsOjBzQR+ViuSO0q+7FJ4TKXEBs1Vbp2kJYG/HFHdkj4Nba0zlVePYWI/W
OQoSk7UzkKrs/XS0Ui62wS0KlH+QLqRxA61LANL4he9S6wQ1pFc1E9QAkjZZ6JLWx5NP7DHepgaQ
H+HpugQMsLNpzFJRma5W3Cm7KftvbkWwNZbNvhRmdmBxrEjjpQbMlpwr9RNM7V/9kRXcbuSIhzEz
t2I0e7IMN4CA7eymOa908GjTbTQrPngalojtsbepZd48Ldd3lcfhL0LBHz7MIAqaQlxJ0183lzQy
iIcDP7HUXDGpDLGECVbx/CkYfs7t/SV77MUTktx1gwenIU6ku2FNRf9sgw7+r55Rsh356P3htjzi
dX6rTzpPdxoOlRoEIKQJPyKZgAwNrzGUfVrMAVl2oQznlfsjMVlhWuJ0Xw4gpOYnmKCm+15+V32i
fh/FXgzCFIO4C8KyEbD7MXg7Vva5ripymWfuvr+CpceVMoa6BhbaGCLlkyZxef0mYfvDpaTUWNyq
2QVBI7rtfunkDqtvDFZTNIr+maD3vVPd6IvSW598JYw0oGicqwA1W/WqbBy4gC4elTx2ZH4FY84z
xtHlDoFdwLNrtZcDKikRxQI+c8XlZ8qF5PUjx7BAcz39H5R0u6+lK/7OmqqjmyoqX1LG7kgXobkl
J/7h4e5mx6yVvafx/r01MZm/tnK1ClGWy53X9OGjXY/nO5z1F6XAZ7UV43VhBuHCWqlOBAAgRBSJ
3PRdimFWMl2CWyl8CSt5BRedSnxfhAz0M0WlReJBMZgCLQbiQxOzOfc3BwIsRU3Y7q96LLKgMlTP
w3uNTN9uwbNChbLwPw1UCWOs0C9thUYBhK7pRSesQ5Iwrylk2NptqMcPKITVyhZDSmb5uegVa0a1
Bb2YftWXLtBxEbAg4M9eCM48jvd7/5NV+3aNdwj5rfSRVM6uCikYYvKF/WD2EFgoCDrS/hB/jgh3
QZ7R42Tn9BSu8CHtPp7Z0CFmjwQm4rNoe1ateXQTHBubj3GMyJ/j+38QEo/gCmiRHQndvjKyEqri
fkt/Q2P23zssYpE2jlMheD/W579S9UPlwsEGmb5UEv7++uZCzSt1or8HAYAUve+rGaAzaXRaQClR
TTe3K73uAc1OnFi36lT2teA/Hd9Daw+mpwwjnq1eIvsIYPY2j8rtORwrxhFjztmH4mqHzgIM8F2t
DV2m4t35QY1TZm2KtC3qqqGXzdwQGn3ZVjhWPmOR1xmTydIBPnCgTwjzr0WOcUhCOv8OYFby+1Y7
TqRsgKWkQMCN01xbnpP2ZTJKAHJoCOPIqdMfddhx80CeeIjO/K1SJFiCIYV2U96IW/ufDGYiQksk
k4ALPc/AjgT2d+7UYRNnFN68momsDdoBREbP2k0D1cvCjlfe/BVkvwGo///cP3ytJJlo/sDaVHPt
G6CVjS0p91KqmnlU3rplqZ91Y0gngSSDwcaapBT6FaQ3spgThwaOW7731h1xLUXVlv4uQOaqZQkt
BWpwLzmXXBV9yWEjs8DdAuHAnj95G/doLy6gra1KvarXSUmNAapMfKcgs91G0n4q/4kqsxJ4rCyH
AcDS5NzvdVVitG4xS3CQWAn2eT1EUc/LAjOeiiTZG0REnyuHU5YvI0jSoQReKtdp81GzmGdX6qA/
oB5T8bMBvWKcNOU8I1WFpK+Gb2fmkF/1GpGs3Mzje/dcTz6EltW9QyI4ZsA7AhrK9wm9M+sIBrj6
dDxlAYCtKI3FhdzJAIEfAPo3Ztqj1f2ZX+KoUpOaS/yYMc8eySQDILLOLV/HhVLeHd4+gBBPRjdU
GdUScl4saiWlZnqLhvx2pFFIL9dY4KqcQDzSmrE1mo1qTuHHluZNgDNWhxDgbIB9I8ysGBX39+yW
HY7M1bbfirTGZavNQiY2BXRPVWf/PPC/z6JhmRzp3pCFWe1PhkRUFe/VNIXiyXHOa3AfNDNreYxY
szdMyckIG1Wv0HzqBbNZWT2hkGOqUAlbVwjIAa+a6dOQGryPB8MwtNhY1LQivHNeSiDYxzZ1BJgB
Q3mwHY2LngBAeA7/REh0vjgIB5nVsiyiNZVVYtPp0ZoT2qy5B4y4m0mOOFBtqLJ2Ojq85QTIHCsx
m5bvOM39vBePm1eWkrfIeFM728E3E7Ue4C6LZSH6QuCp7w0OyPEWjNtHQ/c4egDxrl15C3JMdVMe
1C51vttve0ScIJNuBKPBWh1JeR6eC32uo0nipdlPwlpZibRnN09O4UXgUxPrxmJbK6Z2QVxa4l3d
eHtE46LlTGo8viexYVBS96sL5fPVttChY8umU2L49Cc5/bDFnsjKQ8p+45SV8JSYWWUfmowUsROz
tIdQ4diAWEUoXo49btNLGfYzWb/EHA22ToBsn5VMthHnkU2YdBVoEzsbExnnB2J6OttFMGukyNfa
KjtBdal7BYt9fir/HXw1wQuZKZTXiA2zxKbjXyF+mSennNVVyIM4y43S5ZDsJDFwQfNgHjJPi4pO
cJ8WLzqw8xdayaYCTcoSE4W4+xgK78kpIKZsrgzidAxZrbZCAE6irxj3bfXB2B0Y+6Rc/iVuRcqk
vNnqaQchb36Er8PCCQLDR0qKS30/llVc8v3yymd5MtIajMPCptK0SxL+HIHwQq7REzmbjDsbOJ0K
U/oNMkceJDZ9IO/TU5xr6pURuHa9puupRkrZMC07GnB0M98U9ihcFq3pojkUdw3ASfJSq68+SUGp
N7pwY7OO1HmTQ7QZklvDYFlXB0QvQNJUhWeUQW04YF4bMY6CAf+XE1GlP2Ko5mqcDmvfWByVsZPN
j1Ayp26qdJcX0G85SlaIr64rS6UYhljq9y4o18Tofk4krSEd3GwloM18eP1aMGjX/60sdOx0lJ7A
I5MmfnzvwJ1E02+S2fL2ZR8CRnzxNe/4i0s9rV8gMF3UX41m3PWywYzOGy0Fmy7r1ggyiztYO0p8
LY6kNy3uIEOIuQ3rG1YSeeGbNC++bXNxMHsIIi70DxNKorrkwB5sQcATGFlBi0Iwupb4Lq4XCzfL
0YFsUK4aGAbLMGmgkWylYpmJ8RrqbLJhW+CoyiDFeU97JLlWdSJDj5vFh7EN1XpIJR5WH4o22PeR
uHddsFIkAklf+RyFnZeejM4junG8XM6rxG9pUMY42JllXtuYWnsoKWoetJx4yeMDN9wjpxLTXylV
WfE3DcyKXNomnBxKTNC0XfpzHwsBqyrUVtBTpXOHp4vop66HXj3Dtqgk+0OQbr/oj41sYgyJ2cJ+
1cZMPj9UkbtOkeDfNZNH5eQ98sPCJzMvXa7qbBYsQLz0ze8Jn9BQzs3v6igPZPzNO+hF8f5y2YRH
ytnPIJfAfm+IQys0n1C3mjZfdtWzBT+FTCA9M6vcCWbUIfphVQ6AD4ClbX9y5Tjcrero6eZaTc/u
MvybRaPahaK5o1zoE2d15WcZOBIwLr+/cLlNj5PChugB4dATSHy2BksSdFrH0fmCPibvs7R5zjgS
84oPu6apW/PSWlK5IcM/h7zMXykX8RpmJabAIBLriqrU0GtiZkywxxZ+Ncj1Qpyeu2yWb8QpANub
Ew0Woxs35K2PiBaEbOQzMuH/6JCoh1lxLBiDMUmM2HL6ScxAljSEZIywt6V9V90/8sTg9tYtidNy
SwFPpp6Jw4/F+pOUOkav9S1j+14QQi5lCnrcbAK5UNwRs6VaUJyBqvhDBXAHIawatikeIWx89ktt
IL1ETLP8iWcRkC/Br/RyNDxsmiXC0LfzK1eRNa769YMrxR1e+rVDbfl7S3E5kJfKHL7mnY9svQm6
ZDtIsz3O8BBsbhhW7DARmCVD7z8RPbh9/rtSkjGmYy8PFDpZO4E2QP0fmxzstz1njk5pDSlDjhm8
14H2yZw879+Ec/2TAq0YWGBI7k+bZ1sevuOgWJMn5/BT0h0qBcVXfHZHyi9YIiWYWHJP1xpa40i0
SaabGoCCasMoym4WGB1npdbcyYhYGduwnshQAp+ldi97U3SBp4yUZgNDkHiewLIqh3dZ7+7jyARM
Y0lyKomLI6SXXlxkTm+wTNWfm+Xne1+ef2bcEnjNAlgWznWS6Ed+LIzrZGChf2mUpHhNmNckP0e5
RhRqM/EZIzdj7vAEBS/zBviC0kCWitnm1g5m1gA1CA+kjRV45c36hSUeJn+4nyOCsUCy6UJ8WrJi
IutsUf9KYn9XMN9RBnkHlRotmRPhgKnId7zIcU6a+tEpUVGG+0YTMN0VSxM3w+Y2gU+PEcdXSf1K
PZhz6h1NBmBNvfTiOIUKR7wvwHse5mqUBIV6/OBYZV6nI+kyFD/DbL1gCiygUk/6PXkuNFDFg68m
VeY8aiIAE1rY20m913wyr5YBVCIb/US96halgC87iirQ2Va5OayCoD5On7hFWuhHQJHQTprg7co5
5sjOc8d4PQW5asYIfmmayjaEuHuOnCMrhC9BZ4lDVOXqHQmqkwiv3uHx0PBA+1o1nu+NL+u3GT5E
krHNIzlaYhpw/zAe8ev8/zoooVMxe/4+LjngorZKeaiK0uf7sh8YNY9wYuveMgrOB+vZ5ZPQn4Si
KR8VeY7PeL6Ulb1Sqt1XXICdx9FXE3aiRv1KnDrRUTp2JB/zUZq5spQqEQgqfIRx6F0ZxwDf2nIl
fM3w+IceyLJICXyRhtcf3l/QiLZySvELEh+eRixqgAduM/o+sSS5zhkc/aEez+FbvEX5HhjUXAQb
HMIzyyU5YEw5RiNCScDkoWY8+4QCVWJhy34gwxl9Fn7J06v54qI+k91GXtXC8Clc1ilwrdFGa7oM
iXoceEfXzkfqsd+rR5WjY/7jGlElKsuXlUpZUeF2lCIEivfQxs7bYznL1IxG2fbWMun5yonr7JfQ
Iikm4fIttkRzhHaXTK7Aw1oZK7qCu7ijdmmenezXOV4vweJ3Ej012hJcx6lLKBPK4Uxm0Ks2bndz
7SZ+z9OV/k3Rq+eyK7yQ6k4XAiQzEbJfvNICt0hoEF5W0HT4HnMI9FUzbPo+RhxcvQlhqvfUjYtw
3DGTkdLzi2JT3MRyxOeGQj5WjAVeRRGZr2pWiZJdeCzuAZdyKiw7YYahnadQif2hN8jfbWf1Pgpz
acLkyo2if7cx7STxZR7mlDJzJN4UnLsaqcY/INZ9h4Fjj+PbwzwIrotjNs2OqN7SIo3jruwf0J0k
K5K17dMJ/mCjxhWt2rnr2HqLNU+094OudDh6EHWK7a7piKjRwmwFLC+p1qqPen8Xoos4LSBTV03p
W8tqjvlgd8MtJnXF/SrSMXw5vcLzNLwJNH7AR159yKWGd6L0Kc96zWEoMT3J5tPOWrO+pioqTT1H
7kkKpm/6sEFGlqHXOMnYWA3BggShY2Ly1UIHyEVK0utIiuubNOAoH0ZsfVYNM5SZwnJbRByKKkf/
rlwfGIV5iRh4haNnncpgN8GxGJb4u96FwHKjmp1SlJ4mTP/QJyDb2TMUWk3InvSxfQWlXn03OkO2
jhYUCVV9ksQLj1aBB93jDuEdUocauCW1xOp6LgELWRICLwJzrpBfiNhq5qlMERTFRXZoJ9QJALR1
EGsLNhp0Pc7B0nPufCEqeS1Vbse5WZoNdlAyYa6DkUafd0uxq6W5Q6+dsnqRmzFQCHcylGH9r9ev
ggVZOx0JPG94roqKSEFzXHFX0Ln7IO0lTZunNJx+n9HaXBDQgg6TPpwiZjb/aT9LIB3tz+TmNNIt
msZDIVjmh0pryEc4a4VEG0SsDeFBuCN5/wHBxzK6DGUwcUykcNgFdRrmOM8+XGz/kzcRt6oMASSi
FAHEp6HT2BR1QOgtBDZPwkr1aFDTrMG079YE7e8wgHBCuFd1vfCbHfJHnLQ20WcnohLnpj1eKNpQ
BsrA4kB7Mwr4zCb14PWeut85k7v50WDFplEYp9zTaSCzAuTLJ3ZUCab6WULKngkIRmgRhanuHVVz
HYIsJVXHGFgyRowtenEgcbbDR7w+e48D/Jc2JNSbjUKeZpbjsVlFtPqJOb4WRMiYzoD57bRQZDxI
wj/QMuC0Zko6pAjsVuj9L+2k95vmnfFiVPxzPxWrVK0ZjdHhiwVOpZLiRMz7Ur0pbDa+7pYACa55
rchys4zfV/EekNu3ohkixL2OvQpym10f3zdJS6DvOacm2h1G7GaPGgmBrudvr5y/RTcI00gz4o7z
P7bCRsw2j94BDU8WiU8IxLyh4EgpxspZOBckuVP2llE16aWV0QVvBg8x/cs5lTnx5pQA1xpEsyC2
ozFnncNoUPQGiVzKxw3ntn0gOU+BtGW1IbAHqvnr0DZH2VTu5lsrZJXIurGtOsbZ23IcI7XPtv2C
lGAMCYNtwCsnk6rYmesVmGYkA3IK3i6BNHodqFVejufIva9sbXX9JNzJsYVTgiqfWvtKtGiLtRTu
R25TbpE+MGEUInhEq98ctu1u80wNyYMPS0a1UwjoclVr5YFlwTTmurQDHh/nL0uaBsSJZOvMsz6V
ri1i0TyDk3xi4Df3U1SszV3W4Opwdd+jEoC9dSNwXLyL9T9Xr4abWXWcDFz5h3Fx4VNTvayu3ei1
QDG42c1fqWhcpTbYPaxXOUhIC3QkhvoARUelFQC2RayfhgkjNRZqSNyLWXUpr8f7TiUmvfCtzuca
OzR/IzlqyqpHp824ZyjSUqBfCAenasqHSApY+rnVqECJt0pVeWCN8Asp/sRjewXGfb/ftCMR8n1d
bEaQ6cc0CrG1WGA9qRu+9S1ERdwdO6RhHVIuB3jDRHOW/Uo7fVU1pnrXTp7AE+KXu/DTOu/UV7Pp
8veO4jXg3/Bn+WITnJh2lN4L2m016Kc4HOK9vwvu+rspVwXooQtiIoMMjT8demkCsY6NgZ6BBO25
iCR8czkDU6EpQwD4SouKgresDqT0xaa4T1Er655qlUkbg50VHygs88t5yevbJ8p4j++Bo7iuelHe
et43vEI79n69A7SDAJysjJNN8pMBG9YmFeCIQgBKrP9gHxsXJPd1bsYU5J6JreTy0+9lDK9+JXpZ
cvayc8EL7iikevvHfbxOjy7mLz/GbVPjn6nP2BH+3UVSDxY/CnGkZ5J9guj5udiEnRHJMt/IBK36
2g6kPMq27r26kQxcO4r3ziPS/E0r+fgNYdbYMQPMTB4xcCymDIdeDiFveUu2mXzl418o+jDhLW64
YFRLM/NXkA9c9HEyZuTqhUWSGKn7rNa7ov8iAAXZeyfzLdsShdFbYBSeXLdAdQpXPEaLKAWOm7K0
BWJNrXnosXsA0CSfFjx1Hah7Ve4i1xq4AaXI6Q/Z8FypMx+k8nwtpnOnBqr/gH0pm3twaMU77bD8
7J+tXazqNt77zP8+d9pJKmGx1nrnZbdNidJeOrcc7Q820eo7WDtP1cEV+FET4M8zuFhTlw0JHGGC
x1Y8//Fy0uBY7yokHtryGSY1+pTuKol3TpJn1oiIZ5e1YGtfBZWkF8Pa+up+Fk5QATCAVr2b4ccF
0cHapzGIxv2MzvTizgxOUToKKmFj64Q4HFs5fFzMO2b2Z38wEblZuPBsYpDE9Bln4MtfV7y8SD6l
GUn1q1dVkLK7JnKWSHmKCJDsI9+xggks+n0QynYdyPPhYxlufn5zCALkYpDjK5SK/RmKy4107IQN
yMiIxx+Axdc98Uxxg5lHuzt//I1oxufdIFkEHZ1tQiX4LnpNjV6kMd2vY2Z3zpTAKr1zqqZeyMA2
dtytD6iCgT9gL+LSZCF2tvLNVUOb9eBqDAdFi7esOaMvtjJoSGgs7bWA6LIclGuZnui1PqUcMGOq
Ll4tdh6PAAaVDGIGutv5tSB2FG4EdyHEPstbqUX4UNvoQ4uxkvmRSLKw+cXXV7T+8+z9ObqOwBN+
dhBlVBQJVj4CcT4bJ42CPd6kpoMuDIbsk8CArFtaLrARHTKT+nnO7Al8uM3fHDsUeQt9rHtSGm/V
qGXMWMa/g/l9irzsjJAT3MRHOnSGSE+7uKBcUAL6DBWCKybjQdOD5xL/TOA2594ocvqpEo4tt10g
KwZPH7zvsY719oZC/ACurPAIyzQ1uAb8FBXhICAQ3uA7UFIm4KyCJa2/lSsUA+39xhT1d7fhTXl5
aNIJrTZNRYJbLPsw3VnpMU2jDzdTVQZ+MV42RKeDsNVu1jYoFLJqjNOOtL1pvy4NdRFam1UMZdvU
mjDIPL5ZNcQwpo+YGEfCS3ECfRBldAzjL+c3mDuf3nWhljC3UjmSZFkO9NpfHlVJrjAQr7IboKga
/QgUBE2Ctf6JXL0tFhOz9s6bnJSz8i6Ij5gd9lhQMNarGI5B54Yia/B8Y8Nh6c0azM5LpGjqmPlE
uuhGxohEMinZ37pQjMNd1I/dUX3XGFb1IoIVI4vnk/psF92Rc+/jDCZGqO229GZRohsne2Esdbmm
9/chVc70y7pAnwdQKkS6bCNhyb5+1ckbpVtY4660504n3k5ivmAFRXQm1Tf2Jof2yYGjLKaGlZlq
oIUE9nwQgebsSIOrEMMP2/F6aJ4vqUueZJwGaf4AoDQIWE0CLCJB/vboY4yrs5a9D9VtkfkScy+c
K7RJ8M3HWZReSR23dzMN3KTnWKWm/GyaibPnUPOgEYoINyAXMYh4LPfqymaLEn0wf40Pyyz6JVM8
YYG2siu2bIu5Ts2d/crDboTrHqKfkCMZVUdZdpyPecsKGNwCVz4zI0bj3J3qILzi3U0PVEXq4TGU
MEfOUSGt7DE3krV7qUtduf21vnTdt/4cdnpk4A9qwPC1yiZ/k4DmEgTm/OceLP+V3OVt7IAcnK9e
pE37NmOE6vS2AMI5i6D63Dpoh9iEDbDw/ymMQCZGX4qweruJAdiM1HpxiFYioTfFiQT85PrUPRs0
8SvXZlrdWEUQncLLgIIIhDN5TeKE7mHTV/WStL9mfdUGf7W/OavPVVjUhYEysxPlgMatQHRVJ9/h
QD+GfeKSU7gKZN9JIJN8SZSmXJOCZWT6fC3AV4YhRYCa2vcJiD+rJEiJHu2ZOmcV69YSgXW+ASMO
1m0jTwTMnBph1XWZqublz7gaVCXOBQwKK9sZK/674Qmu4Vdhs8vhu0BikMWo4Y8ITafqrGEveB0K
0KAPP/hYhgoCUxnic3DlJGgtYBR0/I/5xLV4QIB3PllOJZYLBseHvoFGPYx70ZJbkUFDQ/nG2KaN
Z2SAuwOiUpAnmKB9KzC42WuqZGoT6BqzGCIWbiDfyFWU/CpxAAyAoDkZoL2aIe9pVHOSi165nUQ6
V6XGPBSziMhZRWeoA2HAv2FMgMXfE65eiD3UHBbfJ7wLdWl/mom81kA6hE/Y9tlQnZB2cka+5wCX
QGMOu1RyBiwDixuabUf7IS58uobearDPbTRyyOESf1A0mauXk6JRWfSrGFw1lYsvlr15z5anOoUO
Is5WiKmC+JGkBEab7IUWseSbcA6JSI8Sp3MdvoL+TRH5CHafNatAfZX4A8xtxFQBbYcnxxP8yGjn
+9p4YhOOUuW+m2w4T6vNnecKtqoIi5fZi/cteNih0PiJpf9E8WnI4kM15nGzFfAkvxbqWhLdMKxl
EQiN1Tq6RbUHSXZwjs47JsnacSbfonlIQ3fmDND9Y9MFSWDgTqxL+WmTuRBBmMcOgjRymN98P2wS
m8P3g4wPWTafXy+3T6x3RXwKSstDX/+bACETooXOF0hzJQQNJJUSFjQTVw0xejTSsr8ygDsSAco9
udR5jYM4YRAyVHVe2X2EFTmxupf/v+0tJt98MZFZaHz2Uwxs592+ieHZwYPhm+aDyXxZ26JJO8LU
qiZUZ8SLOnpgz6SwlXL6Af0OsX1ItOhaWhNDL/mSg8qTEu3Ns3+YvDyyVsG9d1s8JuJKMfd1NqsS
dKN5VLAOKwAVvCFZG7ADZzdvku5DJAe7lytXAbwtTdC9SVXyk8bVhLsCf6kIJXL6S4agiWjbTtrC
2L5FmRNyPJFI52TX9hI9KFP+g8BxYaT8nt1ofOyrdgBqGBD6VTqQEed3qjSpPbBb3641DkZbGmdD
VQ0ihIPS1hdvF+WmQjWvwvIb1rh8fVKv9sly2VfxNoCc+u90Kpo9eWg83tvzgY0gEg3Rqq5r4HHN
xdaAkM+0OASJE8heLOz5pcMgoLb+qzhTAxEql+GhCuxkKJfr0Q4VU7fCbX/JBJLua2+Oyi57Ebcr
InJcvh7NI5UkTH8tlhql7JlX6mOtgTNBhsGAQ0E0h+s4ocPga+YfCzLU6sIE45qhioOpr21WNkUq
4mrmnphRrutnB5tIPIdh4KdIuiB/4ddCeUhhrKsKDcgK90SsADwGI0EdMLWnTdZA93OSEIGSDbS4
8xbjmncbhTwVB58pkc7q9QJ7XzivN/9g/QnDhXGr7zDzYJSAfHx1C/lLfBCfSeYy7dlL8twdvzBx
Qz97GtFU6Pnuwe1x3vx8tr+EsGmCt856Gd3FraelQ/0Hvi5DO8ILQOtXgKOVrxivY9/50SkpX1aE
aVrqEFNCwI4v9f1zEonSys86W6yu4ju72Pu+hmmpfw2PfV4eF8RWZbavHKLhitM9KbamCBTKyxhN
eFaEteM0zazVbEdZgiEofMPi9w2pdMlyHbOrTHks+rZfHPtnvFF+5MnXExYSycmIsYiJHR+60ano
KhQsavKfwS6p5Ea+ne5t2uictBldUJOSyjjH9KANpYSyRlEhLAbVtYItprYekhss0lC5T0TCP3zx
MgSx9Mnh7NsRTJmWK3FMP+bX07HgDCTo8NMu09umLQ/M54h+IwD/fc0cI95tszT5Mn7bw2vdKhKD
AG9PEc7TIhnghsI5MQC/Nj217/GB8s4XY17ug6qDaUigpxTlNwTY9GXdiLg4qyUU+Q1D9fesUood
q7Wa1TFQtQTT26oIzAbnDF2LvzBI1LR9mUYBm/hbVMGN8cxtVtqy/3YLY46PlyKBuW6RzWyOAlKZ
3Z0VNKPrwR36KmIgTL2qQlKTi84W1pGiPcT+xMOycj/CFW+KaSTwp2AwRAycLLzqnks913DwsQgT
7SybglddLDMFitqcwXzR0GxXq5PFNQxOQ9mJyrz1/DWORuiuIjqhZL1e9DEx6fgsZ/zEhpnYnD05
w0hBoU+vxEXciEtptEqDrR2ODeqclyK0dQq8D8VPITty0pbQcvTQX5N6vBuE/JBico8P1CSQ34bk
eN+drPWA2qTJy8OnypVLUm6T/bmmgWcBRVkBZpSJDSbQeizq1UkNa5NtKDyHKuWkSiK6DKWGVfc7
hrIzWzj39cGWCbec5dyLvh0iizI4ucfZIuhTyb1kOZceJYJWJKUzPr/inYe5W55RPr1bPlWp+CWq
qt/qY/laGaCnLIxNPQYAseHWca2g+LiTdK+QOm2cHJw0Yv5CcX3htLmSoK45b6vEY/SGBs2aUjdA
YcqbA8Rv9K0rgk+MwN0ApeFz+zZjgrh8VSxAh7m36ULQa9gtXPPrlGa8SUzg1ItqiavW504DRrLy
XakSPKPvE11Ui30xHvV4+CSaRTC18YrPCbnBFV81xgouJnYYu8/VYt6yAK57PqB27zhju5Kt3ZGZ
8AOHMV3BY1rPOMu9COj60L8IVv5xZe1JHk2iy6NlbHtAOfAiLXy08u2QmxgiA5OFV+XyXoh/h8DY
q4X708uVKX1ZWQckhb3bMi9xzsP+lS0sHeypAGr6UJjBoOnkZSJsnt5fYV0NrGmTa3nSyi54/Jsy
2uvIqJ9xfCMSuBANYIxYK5q9hUsr3MBJOC4C1uWj2pOtEEEciL8EQhUXZ6o9CAbD+ynauexLZkJS
dEjxhh9e0DL0DOnjVqrHkfjIl35U/MGn61EKkvcFpHVsWRqy6E5n6gnMKSvpZVCN0bR8crPLohbm
CkpzBH7u65/A1/p9syfZHXpy3BfL6vll5YPXylWSBYJtdnEjil3KHn/H57Ys56kBpxc5McSG4uAb
2jSlItWvZCSpKS4+GWpqbaKFZG3AOfhAGh09AaVjv+K1WdA8gKlinU/WApI5VpTe7axfaVpwLT1I
jfQdXdRtE9Hhfs1ixsXbU5y2HNkCOXtrZUVykYmDXu7bFRWkVq92cLZsQjKOzQyfzLkTW8RAP7CQ
xA5+VIdXC+CkFYVpyjdQ2CL6DYJDwH6Gdu/M4GiYcyLmkF//e6x37upVv2NmQnlfTb5DHaqWBT2L
YCFoAzcQ+KGZg8Vb63iL5TxRFgmcF5yf/UKaHV/BZ2WMvxkyn+7pSnvlrCg4jpYwx2071XLk8Oqm
rMu4cK8sGiy4V/rRJTbGPWwuHRIBSTxzOpdVMHResz85B1BWFW7rcKCZUX4Ah1a1dYdoHS7hCW9c
c9CGuBe20DyLdl3jCCC77EZHMloQ/59vZmStOBiFZKEIQHa2thorLUvoFPwQPbWoC+DhTvGjb8BM
QIs00qzPfO8/O9BR5ev4Xe33vkVQO1dt+zKG5F8aRH5mUFCYj2bkroSVVA38NqfSxRJPK3CcZyZ7
aom0CUksa27t0IkP346M8oAlV1mcRYNmL1t3Q97s1tmXIXiPvoNnz/MO3GraLoqNBt6lAF83w1ZS
RduJUeq93w8I6gaRkNd7OB5kztYqrefC5TwRbdScVl3jAjW0hhq98uTXaatFKKUvtWQxaF+dNS8C
n+lmc8cM5Dz3/XeluWftZEm/+rXyLh1DavJDdu0Z1GaNO1GFYxTo0CT6ICX38Qfrs52kO8g/lUyY
Wu94AjeN5H54xe7uN212nxkerBAPsAYiuNoCGt0nIHWSnKNQSPyw2eV4WHZcF8jpDpv1mksYSB+J
RoT1VBWSQqjVRWt+7RCdyzfX19H+G7Uhm1fbKTH1vOABwoplppDZgnwhACcSNtRMI46BuJNvc1Hc
OcXVvdW7O1LkpXO9APTonbFzlr67FLbPd78E3KlbLwAjBaEkFnRGrsVu8dUkEhHzbVonSwbzifur
buQ0iTJ1ChnsKiQNXion78OeLuCBzg3jWTwO43DxZuD39fjSzYn5bZAb1PCiIvGtWiyMSUFajx+A
peyHyFZr3tVuoG5+Eebsq6iv4P8dvwwn6zYLDPZamcvVR4RzKo9E/zUtkXFYnN77S/2eW+HBwTeI
n3mEWxxBoGwl2tkqw4Yk8z9wPlSMfvJ00ch54KzUVA5ndKQexiHKVlFEFqU+6fcvJ7NHibcltPmH
W/1nXbniOTge0VMnsfKytQ29du9/XDRugRb356KKq94qT3vf3jDBC/JtRSXFHOL+MTXkrqIZPvzN
/20nqc0zW/ZLJTXwU3BZdZSRc6hewKZ3O0m0Avqi+XkkRcAAyc/GLMvUGBF5izmRT2NSVUsg96De
rdLKZzPj/5g+8SgQdQUBbf+ISEWHva33pm5xBVhZ0MRJxyZ5zhYJwhCET4gh3YZde5FqP0ALnTaQ
pimeAaRZmbv+5/XcRPK1QyCm8vFlXk0hUxTBJOvhQda7InDacfeL1dXlIdik52C8CRMRh1NYFXnY
6Zz3hoMBsqoXl1QSbANUTdy+idaciFcvGF2ALTpXLDrnlp9dyMIjwF8SMQLIqvlclOZCwISwMJMA
urbL50+XDeUR7xLLpqIyj6YLqXcVP58sFbFCpz930llO3Tx/C59NyfbCbAbJfQqp/+eLFpapHgfZ
fiZ5iCs+ahBCslriJGD+Sub/mEdmbOlOLmCoj9jN3nyc80e2qZBtQQk+3CoOB7L7AaSnlPSGvd3u
XrL3QwYa/LkxVHOXSQ4awmL6czKaSwdV0t4vDGBFPl0FRKXoPliKPv5o02t3U4Wl2qPe3aq65QvB
c6DHldBMi30RBa2zfg3GLOPuJScFYX44EqlYXPlVArCevQphHcAMKBrjqgovSq0FdiEfyq+gSwi9
Zaqnbny2LPkv641Lco2FVn9d+NwpXYdcCjFofpqLGM/gRg3+ROLztrsmM1QS3JvFm/12uJkhVsGY
zXXmYt4VhnTrYP+2iryBBqQ47dQZ70rSaINoOjlMKToX5iHHaLAyd17Ou2bEIkx3ntXrYlO+2CW4
LwNyjy+Ryl8DafBpSbqs5MmS+LS8GnZvNShckmV2svlHE2acWJchGfdpaRrW8qhHJfL/EqMOEG85
UEqbld5/xc2V5Lm7ESnH0RwKy96vw7+QdbCshrIKHNaOBl3gXMmWC8RQSwau93/N+hM29TUuGPq8
guXHv/RfVuoQHt1DxrBPeZuBfP+mum6POHfGhaS3qP4hcJOMTPaBSFcD8Xa/DZIVeZGbwcGgEWZh
ipbrY/AGNGcQ4P2HostB06PD99d2YUFHnYTIh2Jnpr5SvmbL35k0HnVrFJK2lGdy4qCH1dr97091
c37+aMgHoELId5kbR7L4IN4Fs7aqr1gcWQwhKJ2YGjY8CRWLS7S8EB/oT22B7W024lbXlFuro2tj
0jDVmAkD1UBTec9We96Qxo6tcwArGRKMow4FJ1doQ7NYnu1ZLDyRc0+VGDUQk9qv0yy+dT/T9cSI
khoIZ0zaqYpm2M54Q3Fv4CJMVfmvqEfzmb4WaoRKHTsEpQymI7nJ7jpyiMinWf7dQfSeDv5WZpDR
/7+ruteGckIo+VqrbtDApmuo/h9udIL+RGrs+ZcUdJ/qouOaibWZG0oFyy8VCuDXD1phcfnBVd6s
OpQROLzT64Esu6t8dxSDHeciUVUxvhClBoKafdz41Bjs6hOUdjjfkE1Ocmjagz4LF9pP489hl+wJ
SAJ4p+urOLXU2EYlAvY5rHq2NEhQZojN9zFNl55evl4na0bhdqwWyEAIK0MZq3Y3QISr7GS+F8rA
QP4ViyS8UJNtNannoEqSiBEESGet82AoViEjLafzfdYSyBMPIRUMIi1kqt367ZWjZKmAcccQFIU8
zLo6KM+se6TzXcqPutXqL3+WFxT/CPzurUyrd3TBW024MWq74BQ/eBKiUF6Wp+BwRIeRaRFun/nN
oBRENecTSXycbhzebgDghv4sCqor1iJwroUNtm5FqQ5zZfb/wXkAx+96/SnlepSUnZXOE0XMEHzB
bhnGVLUUjP8XzjHZlzYqEWFt212/z9lxGwg1D4uozTYy+MzSJtIisy0JvZScAfKI+rzGOry3Q7id
fkcvFAnA+3IemXfhKFL97VIq37K48/d5jw35WUz7pt1Pf4iIS+HQRIBNiIauoSvagFZEjQXfEdjf
0Fj6J0d4mcadnBpBEI1zhp9f/AiGB1FfRnDQteZA/RXoTAcGbGhJWLoxVK6aM35FefMirbkftvpK
97waB0+dSsSOoO5tLLfU3Lz5G+rtnr4bwVczMeqXnBgu9fIse2Buo6rH5gH5z4zLYQdvD/22cOA7
fxZsJon78I7Aav2AW0kLclCMk9sxuQVM6EKEb0K+ufUDEeKnFLNl4ic7adr3n2BcJmlKiJfgq/ZN
/viPW2crdGTd23y82dX8tQssfSbIYoI4TtttTx6orYlBM8q+jNjCaur55yrLEAMrX1R10OsSazzo
M5dOFSn4y0BmzIpAB3QuLyRy90vwUAc8PKSs3Z22yRUR4Tk2cFf+0yeK2w9GjOQYJTwA/HXpz+aT
+tJXGFBcEwPd5isjZXR9IZQROYXb71biU8ixF+XXyIHABdpYBTVnW5KN1yO/FfyPuxLYRS+pmdYV
sxO3jj5d0Wj1AIfGG0tRjYbs3fK+hzkYxNiIY4T7FW7bTaV6NfGizkYeJvvrVoA/D5Qt1HWLWaVA
kXzdJrmSVak01GCeNYl9yEUoLTNfOW9f60FXVDADcJ6iQmq5yYMiE36xXxWw4VsyRVAN+zYUrP1P
JhLzJnrFdyQY370FVcZco+6Z9ic/i/IXa9Fv4fD+QM8PF6jwB3vc+zk8yVJWED7CKLDsCPA7pJUQ
wtoq4kV8FruCAs4DnNn1agpGe4a3/NiTp1WLBg5iPh0rLg6JRme9E8i8de84ME8SThqPDT9AoFdU
ll4Zs/uMJbpQKCjHeQmCDER8LzSpufHUDSqWGOeV4nrscBieXOHGOx33GHJTkHzFU4UWlvGCDGF5
XG3DniJrwTE2wLQmSvaSnqpNjkMDZJNsHOyySrM3pQ/WO6DT9piFrfTBv0n/WyTmt/xS49nOte/e
NykV7xg/bgt2he3EgA0q1TYCh2gbd3exeW0c0djz5PGS3wHfpk9hKRHrmx8g6PY8lyBbe6Bkn3Tg
Rqf3KPgixBn1rP9Z89ib/5fFhKI4D6ZyppVtPsDBSA0SjQaE1xKs2RrTgpZ4bSeLN2eR5r979SSI
DDcqDk9zIlANz2xzNvb1K7zCDFaEd5ivKo3BTDPZgfqE92ZTkQO1WjL98/efsRv2HeiHELyt005G
8GN1fl5O+f12mTag5Q5dPOVswDICqZrxwqWleNEZ5NoExc/0t9PNJrUklaaJkKxWviErmPh/EylT
gPLAKtqygQUYpQAXootgM8sUU2OMTtc6U4DW0jwyCRqjLevT9sOR6BHLTVD6Mglpu8R9wEQAPOZO
cTL7NWtpIzHUO60++NwZPrRtuWGjldLL3IbbFVbECJnMnXNFa850hLEhHovJhGPY0Amtzeh56hyS
nGLnxBeQd7xqCZJCgT0tD5GONjt2DQRuF+c8gSPwV1kv5qHipmRviDOoSbTqlLCmHfJIjPc5mkdg
TPNnsuShuHVgsxge1x2Sx8ti+fSmRWgBL8by9P06geRrARdfoZFRDy/VeVA0Rhjb7T0aqBE+QPxq
VAO+PzXycnVHvoor0taJQllxeQmxVcLBgf/H+UBO+JKdcdMFz7g35Y8Z/fevZVoesmR0WlgYa/YY
fOkQY6yOAUSDIEhNp/OwSd4nQCi/pGFsFjo1LUOLGQe+K4GpkmXiQHhAcrMomEq2YmrfPplZXjMI
pEbdnd3rEedBoVQxy2G1nuMzOG/UlMnJ1v+9YB62EN/bIw98YU1Y8UyvircvyQz0KdtFo7RewxmG
l+j8b4wju0jSXM8mmZ7X0ghXvxAm+wadODmbKCYZQC6zW2YJ0LQHBLtqiP39R90Zgyh0cxbJrgnt
DV78oIQTaN1q9raP0voitzF5H9Lkdjur9wxvPF+9DfPlL2NeusocFc7MK/subphYz3CqZAyoQxCj
biegUlfHQCo2K6RANcwyl53FrsagpY6ORegB7ZUvquZLTT809CbiRQEKe1bD54ByCLLo1lze8S/X
nhWXt6fkafvhe3E0SbPmOo8RAbwZLR/lf/snrAq0NrULsJDfBK+GUV1Zdr6Cq2iqWn18n6m/gFlR
18F6SMTBu1biEtZ9vWq7WkFwzxS7ZpIbeWjMiuL1gpNq8MrGq1WaUjFmlJwt2E8dvVr/UzIQrsrM
jW9VUHYRKuD4VDNJWl94OsZBiVyiuGoSU0+4jVuux3EL9kMY8v3ZGwspQu7vB6KaHtqriRw8+7US
zIAVwjbFzTUZssSssQq49m6LQS30IkAyHDYpQVWGAaYLyUEgOC/OKy//M7aWNkCJZWjM0b6giWnf
3+YC8MBXSQdw7lR75Renr+YjS4D4lozaDqZfuqR3HlrV8wFv9+VImqtm/Tzvc9bwgH6jDJvVweD5
C+dvaug4buAeUmXjkm5aRMAc5Lsx1ryHDaAD4osKd2+hPlqGTFKxcIorUt6hXtcGBdVxSp4FrEuE
Lh6jzlqSPWOfqHcfEbG+/xr3DlL/3MBQBwR/nqCkeea9zujmrXTQQVKb6YHApucGOnukgsBT6qbu
ih/n99I7zMhKAiRTM9/IV6mN6ociPYTPuETRRQCE3RKve+MkdO1jdDgyqLaTnbRwAKKCySVyP++Y
X2ggU9/TVdftU/E2IXCDVp/wmJRWMNRUFVuzvANsyJbrcs0E+0szxB82lNY1LpSk/FDWnfMtNk6Y
xwDp4LwXSFMqO3X2ED0GYatSuVTabdBZPyg4TPpYC7mPPzzVgG8yZMwT6pcDHqLvAqFcZiI6dvVX
JRx34/JUURUarSb9uawbBORclwwbOrt1KC3XXS5lMgy7W9Vad8a9nUZBKpRGT47Yg719Nt/8uCLt
48IBwWdHRJ1zFolVFY1Bd9adsDzcBjoVy5QSwzjPVBXvgU1JdfAA9Mq+aoFCZUBku4ek5m90tUJH
oXoqcqaU0SK4n9vak6u8xnLDgjIMCkP016KrU8NdfOpXw9lD/jcRdaqe7TwvXYKm9C0SGbRsOSca
uB5fZkhWT7Rm8RMtA7lcIHhTY3NS8OLDy16mn0k0wU/r/LWnvKvMEr84XTwo7I1UXIFImiNlvUDv
za4NM7yFVWZ6+KOE9Lgm+KSL8Z6kkgIFlmG2YPgzqOwyOli2vk8PJ2NktsQtiIajhIGiFvJJkwaI
YaSHC3PVBbn8JOCPkB0DAOnoDYuKUWw9x/pXGznbf2EfxjOLLEiMgBzTkKfuFErK/Y3/4BMArSEj
bayV9k28/VQS5VrYoQQ53Cno2MrxFHlu+WyIybG7ASOSNPzy6DsTEKqikmQz2MgDoAjmuz0QqOZq
JMHLgquqHrZ2t/buYlQ0OZxKOOISYpHVUjA1HCW2JYMkAi7u2XLtC+utrNpBKBTsR9ZPtk7+ky0E
Px8f7LWEHc6UjtqyAh091aiDLmu7sIw9zuFYlyzrdqxpXhEVvA/Y9OzBwKi0qIqJyJ1PtxrbOVtW
hSICIqVoXgq7VQW6cX6C3eOFc53zFHSW7pI2c3sLflHfSY640WSX9oJgfgI2DoulraCEpsgcyXSw
FeLYrvR7YbvCzOMo2O6Ps6c1oT78qIaDFj0yJdlnascis/wUmp1/qQjkDS5a9ritYC3a5ov89dPY
mIj2t0Mk8qq36m0/bf7BItPUMJbbOQ5qvLVKB7HfU0v6VzMp0jOHlKvE4Q2yss7lmHqrj+3FTO4B
6LKmg/I8ECYq575mPWxtBSl9CLnHpPxUEdWt4zKqAMMeIr8ZqcAmiRYEJMiz+ft0ItoChsmmVujk
tzWI1BPvXeEbCrUwFZLRUhDQtxEZfrFAPwUTt7db9Ha/cyeTkZJDgQfDI/mCuiJ67CO1yZV2FUlF
ZfN7/GbWNSzwkfOsmGX6BUXamI/BL4Q8W5m3C7QTY77n0g23OWL5MX5yxXJ9ylp+yvH2MiRO958v
GkzJv856X3JjdZNVVqWaK9RP9/LuAi1Aeerp0tWKaZEeNMu//NtZScoCIW1TQ8Xlmken9A/YxRTr
8AB3ZoJYJpuibUGu0lYAIOR1AVF37adNtCM7zhtPEI/D1FZ91NKMulvwnNLyczmrWYhg2Bk1qwmA
qK4Zy7JtA41GBTwMALgo0xg+iOtUv4pt+RYXke59dWYXV/UuOEh8d2k1rEu6MxvDndFto0A0RbF8
ISGbffZmxnzpDTG+LKDu+WFX4IYJqNtyCKwQCUisQJ3fe1VUW/RlS7wXbpf+Sgaa4PQpsvsEuHUI
MBcvaQ44xC43HhhYvulBzNbkutyxkdPtHT6Ka+nbY5kBlEd99VfCgqsGzIoXfMOx48GJ94tXMtMj
KJC8K8WEz7qeWtnGxQ6ctlHdbhi3ydMl7MreC6c0UQXKxbmPwiGgpcU0Th+/GoINpPeVCsYDeRpi
TS42rMGOdSwVbeCeyLdSxSw3SWs7CQIcn53Uo5sxSu2hy8eRarI9EzZAn7K3v4TDKlX5xHTtqlE0
ZK+NWiChKfK0KNlzwDhYhkrhvQ6IGiAJKDNcJ13eWMFwOM/kAOnHwA9FI5edWlavwbDaCh5vCQIM
9pgHC4BARJIfiIOI4K/dpOoGZyBLGW8jTPAPpIrfeKxbjCduRa4QiPxrbIE+p0XD0sBZZCCHRRmr
Em29TL5i12fzofteOBXhQuALSZV7t0iAzGFbYyFTlOTQSM/NY/iDfSIobabRwGUhyu7b+WS+JIPL
boEZcT+5a2G/s28SNR2PI8ZPCsdz9f8fJ27r4H7oP6rJ+pFbVCQ2mcmfrifAmMDwi88IaXXtBx+5
raHTAPeldywUKeyOqDaepM7P04wZ2mfZ/rQCbAcV+z9etBA0uq5h4GvXY4oPOe8jhYTw65QDxJ/C
HFrv2J0hHbP8gBP+bM9osMrFIl0RRi6qKaCszB5aCQYOy1viwE6Th7jCdj54taxSRtyl7DB0rT1R
EX5aDkaKqaN1a6vCTfWUmd8u8Fx5oG2NnAGyr9lHUF/Qq7BHLC9ULclnfh+RjqBIJk8XBe3qDqdz
2zemezhmwCgxX2u2W5lxp3oaVUZETsACkC3OPFve5hj9BfGppSSQ6MKSdTT0vHaN+O+PdkJMdIzB
HKjTsgZZONpOUEvLKIDT3Du9B3YwDGn5861WqyLP9XgvZieSWY2NFR0YT1N2yVQpIyWvBCluO+J2
gdQFqqh3r2UREe8lGNebGrPKSjb0zpyke3wLAk4aAqUAZqvTm635Ijgf2i0ggS30PAiOkgx5axDM
o3WbfVoY/6r6HsxRaqR7zp/XxMWu3k419Pw+DEGUcOXj317EKz8VikuhmXTqQvik9T6RKXYTWvNF
G51pkJS/WIex55Dvbz0SLaG+EnihXo/T61j85n/ZdzFwsaWPBb4m95sCyBAhq5Lf5k5V3IxSgTsU
lQXIg+oV8IX8DNdlhBKqY8z+A8QHaFVTVlHTbZe839qX4GIRca5ag/RbMpEbeJAjaOhhezQbuPv5
kqT4V20m/DiI2jLQSYg2HAUzNqMLY395mJalsCZ+fZrE5g0e8QmocV4V5pelasEpucQ5giE56o6T
9lbknOiSz7XCF7sLiNFQR8LTnAT9idkNkIc1yonaa8sImrqShhqauAWRXtNt9DgLbm+sf7RbEG5L
9RsDwRgXQbdiEzW0hlg5c3Bo7vcNpjGsuCT7CHlBei2iuIUFnICWCQr3b2TK2UXR4G+0fbni55RP
qxhN03FTjqyS1RLxefr/LzHfjo1AQjieyt+v4SoHItXz9YJ3L1D3xLvrYQiSUCXvZw8vdyocUeSg
b0kPoF0aMkRA8BWI961u/fu0XQ5FZYeg/gr2AgWViNSqqFJGTAUjR8p/cI9M/Ppvca/huUcvl/cS
/fcbo5jHlaCeNJoIdELZUVM/QLgCn6utj+x9NzXveQlbWYNBxe/uDVIhb8Lijkq46Kou6mRzeOn3
Tt1zNxdA+XPPrzAg86lPYKlnbE9VJt3A4wtB86gJtfv+4Xx2WQkY8Jnm3gec06PIkd4+Ugspn8qR
WFCLmgo80qWlV2rz+Y6sy89kTcDI1Vh+euKnhEt9G8kQ05TY+y5dMf3CZaZj+u3df8pEyFnaw0DN
b25RkNKff7NWK3noP74RxHzZkgTZ7T1AUbYPdfDBjtaUlhg+8S3BAQ4qooK6MO9Q/7iACTxCosmo
zCQk0TraR7ZJNNT68dzviGcj01a6uehwocCVueEFzf0cfOhR/jCWPkPJTu6Ao8U9wIdVA/IxuExk
qrK9V1/Y6vosE1Hd3NcshXFpD30aRDlO39+C9QNluZaMBp05uoiS4zxvGQKVRbp0p+4bxpqGyB0G
t5yinRuuS2xdxlHpEwq4mX9ugd5Qy5JDJntXHdWjgdl36FR+wGHsjU4QVdHlvIKzCZ7hst6N+ziA
kUPjqouD1Bse4lRbTGZpxJJhO2xf5gGNtiaHLHCIfogXwYopvI0KlNhdLvspOPDouB1U+9HYbUZC
wRCQCCLGhFQRV1f71GHXmJl1cOLRqhGhDncXzxzF7vXTXXio2wFuY5ao8iH2KNnf4LemPD1qX5wk
n/HoI7GS4cg2rG1TzJZSGtwRjBAw4iITwMOwHsl3SKiI/bN9IFKmptkj22f/eSNdNwBNyikVe34Z
bpKufOMdjLhYrGMDSbjkNmJeAOM+Z61pZRmVjWr8EtvJGt+vKIacvNP0+Nft4CMS/ydbSk1U0dNf
QiEDhPtgeKobDIrlF03a6MbtcDp22BQR+GvG/39BRRmvjO5ybYAQGceo9Tw9jpebU7dDBTmwr5LS
71/fOkWUuO8MjhDT+e2fAy3utn1+5uKce451wQq1j3/6Swx4vo6iRysERFLWFyGzhoTek4Xi7Msg
5fyqq9WeLygcjAoPGAnf/RvW2UuzvuxmmqsNhZIo34Lu6QtrKRiyr9pNgA1bYVv1yqY1u+4OkPLy
lnpqvltebz3VmWaEeYydDQxKIyxUE/k8WTlYu6R+ywUJZiNGjCUTm8zeS5DqP/NhKmNmxri3TO06
4nxlPZ3AhbP0PnjN3sMRh3nkEPFxlH8iVuWSWJXg085q6s0KxFXP3P+Wbi5ZVzzrjznkghPz3VkR
CE5kqN+y13z2nIuY1TaAd91wcRa1cclqFqHMcyFlilnBuvUYlgAYZMeVx9Swvs7QD2x/T66p6hoX
6nWV04VZ/CiH0xGfSljNsiMh890nxGOvLnEIyR0jr+vlsYreIJOp73tR2/pzeMIGsbQXBS6dB53F
DTRrsuC3swTN3qu58WyuST3+dFIjjt5WdTEgkwSZA2fomEA26S93QrFmZae5qomNtFUhOsose7/I
a6cVp4R58Qs+03BxWH+XwQokhn2lCFXMyAYQK9XXK25tZgJZcBYEnQEwLNeOnx8QVhY7a0y51qkW
JLLFOwrSJwtBldAlLqOZ42SjJISkYGUnIL+TH0lf00gmUrnTsNy0jvwWE5IX90igy7WV12tVVAmx
tfMtToND0wENDyqO5m8yS1FRp6Jp1CnGYI+RvH3YYQ9r9gc1qeof2arjvdw0rDLwuAI9NGazVQBP
OyyB+6cY7ZJ4HnknbN1nqtaJ4w0BXFlOB7ql7eUKh6W36rezkVng0l+LwozxArXE9dJ4pHeS0f2r
AFz9dZ5i0L+QXCglLeNuH5WofXJ7EdoP0bAczvN/BWcEHelUfewB+/TCsv3NzhrcqD+sMSa9OaKa
gqW8/AG4Ne14jNc6l37ByrXQi+DRgP8P9QhZgVbW+rpoymaYkxHsRGyUhJbhpQyOUzd2mR/Z0lNU
QuWDJ9J9Bk/bY9IC/psvq4DSEXGOBK+2T+JU/S5K2tzjyd5F5LDMfFgFuz20VheUTcMwRW6+3tpE
cRS2F0NUcr8neeyOrUaoLLrJqjGUUaOeWE3oTGAx2w7rLJE0l1LTAqm7sPh4P1RG/YH6X4fvFHbu
7r4mdAVg39BVeRQkTq7BWwiAUlT5qGKtSWosaPk/rNKUW3yi+jZRB9GQCgAg8YqeTa4/6RJ2HW4f
j8ossPQSQq2taAZoRP2+Dbs0dogo099Y5CPBDjS5rQIG3PREd5XyBdToBJYThJWfC4BqOsJxIwLY
F0hbdAI29UodJebOhl/Dk/bZTJk95nHIWQ3difYYjvfjbK/9LF+E3fQ2K3F8xLUcU4m3xT3agPLR
5HNKxInBfmyeZ4NHYElrITGZx3zXlKQbY9TPJyDuDj8YPTw9yLwY1cDPMpjxvrpwisyBfVh+APo0
f44VViV8NthPk+nsxA+UVjteKXmQtW5HOjrYuygDXSZ3+/nXYwh76kvIR6RNMHpmxP9FxBUgXfLf
ieWY42sFLcsezxUPG/NqUYnS4EAGK37w6pFuyG1oYclES6gAlUVdMuMyUkeY6khK7A3U/0GFq4Xr
oYZ0RdiCTNu8SZ7B81tBKK/guJfcpQLpz5N5BeFagLz8tpKJ97ijo46W4vMk/o1EA6spo6F7ToMb
KUXJTkOWMVWxqCUYSzpUYZ8rKlQvaetFKb6qgee0sPJOw7mHAqP76jQ7OjhjnpLC8a9ACFmkw+MG
exmB+jrbzzptBfrFk6iFHER5PqbxQTakYu2oNFpNsnxIG4josvPhf97qhTt3F/rYTPk+rajlVrkH
WD7eycudhsnZu7+3QVWnjNfJF1QcXJg9suj+KWxpTyhJ4OccNjrgNdyLqGqY/+n6QrhaMLz7Af74
2iEOfmJgxIJwzPdeZTols43xQFCe0V7tUyFWt3siT54Pxx4eUp2zZ9qFgiQVPC8QvZLi48UPpjxv
+d7hWpLCtafYuBEq4WMaObD08A3pq4dYZ06WE25/f/FmYrBQNUYww+qwJmfG82YjlEjnj8UXmHEb
VBQ5FvzVsPnJJmgxxax6aiHFBS1YYeIfkzhzgAhSMAB70HMA/kMWNzB/6azIJMzWFB1Ry9iQEL7W
RPJ4VgFXzbwpDIubiyab6uI4WjWpnQk5HKG4hpgDTtRNV5uqlgjOjTjneBu53DGBHODHNwrUh9IE
8cxfmgcsAyJiRuXFI1IMGUmH39sQpM9CmTDZzMyX7uJea11c0y4GS6xgdvitY2DBIB6Xn7TUPSF7
ZB/LrxrO25Mqd9eYsB3DUqOJzROxd8/a9QgwUYRKH/DaSvhoAd0kf1kpVEH8K9p05C3BE3fne0rI
GDVQVkIklTz7NyOFI4tXo9KLSjXHyXR5ouqK8x5mU0FZuKa6SXuUIPoK71Mxh0E8R9UoXw/gTZTh
WVkt+J5MS0roJbuaVMHB4V0prserggKSxcqOjLWsDSPKmVT7q6LUpRSaCrtvc1ZiYCzxKHx4bK5z
CeTudiPdcnBudY6uJn+CO096kOVyndCOAGvItxlr43QXeKdeguI7r9us9Rjb5GEAhtYkPPMeub4y
GUqUuNbUYmLk+iC+ClNGwtHpt2nY2YlPMUzr4UsA0SzqIGLVYO9R3FpajUE2/lfK5QeVADVenI3M
LAS0TZ56CJCM562M1kQCMjjAjm1RIVzE7zEXjC8QV3mYfiBq9RaCGpylI+MVS5hO0JnYbbWrHBa6
3/cAO/QTTW75BdAslfTfxhq76PmsNDPza7f6X+6nLUY9o2pEhql5w8Ebg1CFoPRtbx2ocnx1r617
8zdtXDS3U2RUFTJqdcYnUA198BeD9BhtgBA5v0D8pgyCK1ONZgDzUJc+M70Ny+6Rn9HmLIDsJdAR
bn7uTwDRvH3fwEpM72NFtwl3rztWEOk34Da9CPGZMSjOKngizPVG6WEAlBUvKxmZ+7MY2eMKYFBU
eYyxZKYVN7N4E/cboLkHM9e9+vFq+3wIS3Ed5yji2jL5NwGrg6CVb90OUubP4jNsnt0cERsHiYJp
5RQns+0p0VPtFkRCWb6qxSNMwDCZfIEeCXZLopqbtJ7IQ0SIoPp1wRvDI3J1/witwBAK6yS676+e
ME7qVTMhKP/125xEvEgJrfX/PjntoW/x84o2dGca/3k6PWg1TMIEmXEpSQdKQe9zuEyzLdGP1jtf
iMK95u5mJRfeGkQfKMZcsBd78Of8F+DBhY4+F9RGOJ1Wg85JQc2TE7n0NsHeb8yV8C78/b6fJ5lT
CagTziRa1HXF3d/WBLn33vGVyCCAm+lKDliwdoayqq1sSJdwhEwNRrdingWkSvj2Fuy7chYCqgx9
kutcm0ksyYKgNjNnP4a+cBnHG4NMQyCBfPwKvw/TU6dpUojxLA8S2hGOZjc3XV407FiYYUfzlJD2
rVrp0+N9pFJTGBEBI0sFP9wy87BBqIQLx54F8xjjJEcSUtw7J6O0GS6dhYSLzPaZd8DwfOUFPlbP
OrQXFEkpV1QKMJhobBzJnuZcqLtEDqOayoYsPbMuqUvIVfkkVyhhH4vi5ew5S1IWb00jiHb0vJKZ
i2I/X/fEXlus2comiy6PkQ52fO1NN+ahtTPfUjY8JxlyFaePJTxG/Ds6TqsOW7PobYVpcC9jHqFQ
pixnHV5U6s8FZniSBS7PxxaYD7ZlFhapgY+4dklfwX+te2Ntcie2qpHko13/G1/fl4EzZYmcJhdg
+kfnMVY9WFomb4EAiyrO6OOOsYxVs8Esy9STDgxMVlGw3OwNKHtrWdqnfBha5/5P5mW7ft40iSvQ
TNzH1yk0AGv6IRsg284H3dlf4ZzIhfEcwp7AIY89jlaPt6nbgnOiI+yjXkOfk32PCrQjoqivWGWb
l1m2QT212j99vjwsVe+GElimKV0OWcR9G0ZZyYoQxGLIgzwtC2xd8gq48/gJBLNREsQKIqPuTvHm
5p5nnHql9zcalZNjd3kJ1aMN6kT/EPXKXpdGivUxwXR0WoxmgQyO9KcI0aIhrDGAQBJyBOkegBrv
dK/IP63L7OPWcQZKDZchxP/CLR1k/ZyRQ3H9hz+NS5KJOpFFaCFp66Gbta1CK/8PoQypVq44cddA
JggbY85VWa1xwPQ3Il3nMBBfF+2x4uYUOlXpZuAoSDjRSpntvfUJV9NN/zkhXo5Lgltq6YHvfyP+
c2As9hOMbYNoFM8jyM3h3SeEnQsGVL6Gij3fHanEi0A8/kI55ykgu45ZMDkNL5thhoTtI7xeNhJ8
jgiq3qIjCRc0xJKzCEUp3uTiysr/uSFL7Vr+KUbxG7YIarmEMdjw2i1r5n2nwfs5hKb4HUMBlDOw
bhvgnqR/p4CS1FXjLwDqVJLYVL6gAQZEmYB+Bx/IGqs6t5ioT0CdSi5goOCPrdDv9Sg06qP3F7ua
D/UlQfh4XtC52IZ86QIP8UCApTfeF8Uz0d5pSJpmh67nyq38k0x68jYZ4sFsu7V012ShZFSV2Wod
ST9J9+I/DzqL9JxHAJ8tBB2ID9t2fpk9L139uMVYC4PSe1TpZbbJ1kkh0w0sJMnbnEslt3lXxwSy
bPCh1XsIhA4oEhzljWTM6vflLsnK57KA/Wmz0XuJBBMSOdwkeNoHFM4SO43HP3/K3hRLX9KYGEeH
PhNunoN9pRhr9trU1xgE8GAj0wOvpm5ANOSpIECzToErg9rNh17o96mvn45Y/TRnAADHNCbD8ys6
5GoAfv81b2zVkiE5RNV3vaBFmIXDn51VWjWRI0jVVjc40KKHoKYdT4W99xcSuHDtjLXV+pftjruE
pnbxUqx0/f/z56Xe+x+j1FWhh7Np0H1uCAHvSJrQEjkcK+1LMjAfDnB1FxANb/Fa9Hz3asPSZ0mM
jufS5WIOCK8vgfK1FmWQunOFf9rpaM21mCxftGaPNJ5dU1QVIxtEgd3TE3fqFbP5AqWJttY929BN
8dVZP/2gEhvhL9216eph7aMAITB9gxVJL2bGkD5nwQlc8aDKnKvntMnbI+06AB2T7WQwSszL71k2
FtbcgCPR20O5t9cYYl9fXDvAP9nr0+GN3OwqNAR/2M8NLfkCqaFxaq+YoNyFHlq3VxbMOv/afCBr
eP2h7CQxTU2OWJkceZ7cQff2T8LTVMyPT/j469d95hmX1s0kHLLT4FFDXmmh3s/hz2BeFgM+U0B6
g8+mfcPTDpW34O0dTbRPuQyiolxu744DIbasjQaNAsoTBbAjIXhFBMCpug/fWCF7F8Gx1PQsQ2Lq
PyvM+Vj0uP6tvgUzwV3fLyA32Lo0ymETc/cLTf8gKKp2RYJ+JnBXzVsF+rs6mJgUuUAnhiQPqegK
MZW/Jh3I8K7m/bTWba63zQHKAVm+R9uRjzm8X0jLg0YVioN7RO8FVsQc6ULucWm9KxyHhxUq65Vu
9DR8Fq90ow4zGeSokQPbZHbc7aZ4oNXUdtr+E4pjyyK7HBztj2Wxr/4Rn11JzK0Zl93JuyLI9wU9
a7X5IJjVpdgjpnwhjz0iNa/GjWcIfn0i955J4pmr+WA9EiQme3LYVuDk5Zwp4mW4z7gC5W6PRnn3
RsaQai9QAm2CrV2JAbckPIpSvb7MIV3PU11PNyDgv8lzNme4YxghrxPSBtd2MLwaz3+hMHozI6AC
LIyRusurJXw28NLPIF1iEDi0egcZrJvSfAbWL6zJb2MIEjFferK66gZShUVuUyZx+/PC9mnfyCK1
eWzSL14gaaSx+uXWBL1vrw4XNC3rc4R627rlNMgntMVOhb+VEvc2xpkgnA/wWKLw7YGfcUtdZ04i
EfFDbAHag/N4Ac33TfZ9Jb23X1dXqrrL4QdaQZMSVpfDKRUDTWlp3Q+xFYCZNkvaoRWPcIs7dvqz
gkj9zanQHaS81yv1cIX87JeuTc30JWKcc6z2imsFTIdjvDvCSm+t5VeO6eGIr/w1hVKK1XkTDvWZ
oSOBun1uZpwE5g5VkyZLgcftiR/UQ+hBnMNGTLIULMteOIjrknE+6sMNOhV2qYgljeXDy8h6mF/H
JXQxp2uTezoauYhT70QW4libD6WKDPDxN5yYPUc6Z9uRp1OGWVzLcm0tJKZ8H4DUlPYUEzIVgmeO
MhKBd3cQ1ebHl35KzMqqquDv1qYk/YdjTLWEFOLgjRKOCnuKJc5GnV9zFNviMK1644dx9iNCTIM7
jpGGVfmbCUkPXzNjCANfcaQFWAgjBq2Fwr+y+TM/D5iR5CrWA9+4NYO3ggOP4n3GZoy0FmnuCjOJ
0OWZexgHYUoDBYg4+vtdYLOkBGQRbME3fB0Vu28ev3r+w8NPSiNmtmUrFLc+qu3FOEYYxR/jnKDJ
Tfq5nuTDGGcJtOoYftI2xJiAVOTDLJaDnfEaGPM/LyysSAG1+e7hLFWthyi2+ApXjGxCsYZGE4F5
/d7TOzj8BUQ8ofuEMhF/HuhdKg/pDoqULi370zT2mWlbmlQRcPrGFWGFVQ+jAVkkt8dwPiAYSSaV
jLDDToaGzfgFUmE05jFR6entpa5701jLhqws/VWbVs/ErZ+aVRWxvHIxtosA36n45zppIT3/NB4M
rCUaCu62tDvNcExRGMMLNTZV3xulAZY51c6gJV4JzdnSKFDv4kF0ITnYwrx8mGRxOAypQbQo4jKm
9LNFJ8y+X8oQGfIXjncYbYEu3pRrA4dzXpOMFUUHvUyhZv1gTgNOE7o6+MqGAPIIfRuPYnmK+WSB
571BdthHXDmLKQKhQLVTlx2BnlrWRJ9CulIelS6AJ+2j+eZBVQRTbtA2bJYCRk1D89ikOtNhMjp9
8nBQTi0KA/4RT2ULZzUV2zwrd+t7NT2t3fBtFaFDGJZKPGHHX2UYdw2nYhzFuW2JwtvAy8mopv73
2+jISOOsAXDbeMIN28Nn6KP6wD/Tyk0+FilA1YDsthZyBgIbZxGBGIECS7HTgc7QKU4BpqlnrKia
r3a76iM7fm8Ppd+QIVozlTJfJn/ZcEfoEsDaeUGCMBqCf2SqDext+QQeo4VtIzqId5GnPSP3Yuxj
37p/21ziudcS7R/Yhn0mNdkP7ZD70FLlidOOI6xoFMjJCnLrhfKjfqregVqnswQP7fa/ywF/AuiJ
mpKfyKQpMipBj4+yXkkQWXnm760gKOSAJnsEUh8ds5oSwU4y+eZkkxpc80+30alFhdx//zoYrilF
kuJ0jsXsdiQJ8w9u8cgOSzP6QUj2rk/7GCTFjPp+BEyjv/Q2O/nlqljA4BuDsibSdbkfNx24W5x9
X2J5jigJDpfpf9H5PhzMIeNWDwlKhTYfvsU5DkddbwG0tV9t6EIWGbcP7JA0c/zx5a7vzywM9Lw1
hQR+SZD/mAr1XjDSmmGq68TxG4rgMjO4VBlBIGN+FxVUfY6SayO8DIrezfqEWlf5i74pB1OcYJo8
YxA2ZIVj0/tBucKiOmcU3uixkp+KTNKLTIJWKxrpKrH4TTQra7nwtUloHEX2DTkrDg3wM8DgmFLv
aHiCER5Dyb2cMH+VOuZRycjQwAeY4EcNXiHQF9lambsClgf5aBMv949AWTcfW9YQhE4sC7Im8mqk
f8EdKDhq5OB59YS5suzi46bSVRayUE3IwOmQGbvitVHcImYMZTiRVmjZ1IOZ/GR0NkLlohealClk
wATrhIGCU70sGLbd/0MSAi5VxY1MagEsGzdGJV8IkRJ6iQuKXn3zqvmhM34xZZAFw6U/8h3PtcAr
Xig/W0C0GB1Qzblr1Wvj5j2KWdu6vM54Amp1RBhOVDvKAUWOCp9CTvYLzMk5v5XR9MGPaQWuw+Rr
DVSaO/dBF4ZCwGCDQtZz0tAEHanMT8GiyBeszA5WrK1h1LoeBALvmWKV42dAq0Hi4aKUbPp1Fiqb
P9CKvb8QxrDDRniNnJ/9GRNPSc9qhmM/SrjknAd4SrMFLRNBKex18IYH86Ue+h9woGXJNX+75KvA
wjTczTXzoTiFa2hVazfFOUW7aReSz3NFX2bH31iOAPoU1JqQTvWqjFcO/4jrfNJzKG14d+xN6IZH
KZVRAo8q3Hdh0e63gewym/y8ge0Cqatjx139oBP13Vo1U78ayS+Ejlt7sV+4MuL0ydhbf1XMijhl
iaVgjWCdLCG/Jr2v76VaxIR8w2RFzqwVGKckNiBQ/Wv8hVUpEKcXmktXYIEGKOCwMJRSl/4XG1IX
4ZnSFWgbyeQhpdYJNvYR3o5I+QIbWPmzNrqcAIBhi0ATh1G9y8WpdckSZ261m0UtQxvCcTTuIGJ+
yo/PsiRwaAtN5EDwiacEbfLjM7BkgFNhBoHDVXDH6GKoIvjC/9jukVUhbPrs+EndEP7ZFCDDzuT9
9m2FvOsuv3tRO7ozCWu+BQNom8aSOOOgi901W355egv7EbxxXtsGv7ioKxXcKSF2teP3LiOC+ukZ
YefMbDUcCIz26pMwwWicj3r3nZL21cmAQ+NDZ9tlMsFw2bCXO58iviITmjBnrq4rlZK556xSFder
yC1DeSJpGW4RTbZga6eNyHLlrG/SCxShsFbM00vMPQzFmexyinmYtg6ULdwINSeX8v9v96ThsHLx
J/a1Gn3KLAGo+01gIV2nN28pkMhr+s5IiMJ4WjlQflgx/GKh3XuNBJRhtYiHkAcMkAhnS0tInhsi
S1Cp3ctEh1dS+pj3jOLNbB7bcoEJamwX1CuwvVa5CRoxLc82ty3wmfhGrR3rOD8tuCiTJORX/6xD
ppNE9rjj7MELKmUHahnYMQgZNoZiyLcWoJ2VxTPxsL0vgV0Xazcm2dooceJH4TsgmcFmmkSTAmWE
fUg6sy1egB8NNpLY8BNsMkK13tvT32xfZ3rcRFFxlTDDQteed/UnSclBXaTPQRJkbwoDBuSib5lL
3vm1hRIcQYAJTBleIU5S5bUL+086wV+ZC5Z0Mju/XePU+VAqN2mLlOjO968dQ3v9+o3VfnmY0M2x
a/5YroQF/8aG9uS5cHr2F9lukAeNHh7hG3kMdcenZdB6wUyd3U4EihUzRGKdeu0r1GHyTVZNTD0c
pwnP2m9TmWXz5AqmUaOH138r+CdCl3nLJ0xlUSFRfkjGND3qYXH1EuVo3hSrAKSNhaHVOF+QF81b
509iD5CyYzpNgjtj/CBBO2VaaBYFfMrJEOHQlgVvZkU4iiIN6m87amEq4k/Qjb4t+vZfvS+EJqiW
/ovpDMQuj54oVAl2tufc2009B0kQ0Dj+VsZDE5DC3vhWC7QuK2Of1ksNRDxXekDze6JQgV1m4D1V
UuXDj7VzIp1JvVUynxHldbzCNr0glWjbMOqFTdcycxz2zWO+gilr0SO0FZZgInbVuoUODrI80uWo
BEAncn2ul8aZIaO56VjJjTIKIXAsMJFWLjN9ad6LMo8ho6m1UFA/UlftMXqcxrO0EcY/H9QFAngA
7THJLSEoQ1ETZsgwmHoHLN6/fprDzNZ8yRtqDon12QrQBVAcQQ1dvq9+NfSsQaYMlj8InPFidUiw
mv3WPZXOg/U9QNQ639u85Q1VG4h/TnozrjzMjFsbrdF4Xen6LNT//xDXWyOAc3LHhjG/agxSsmn0
kJHLApxqYT8iw8XPvuAodVi0Y2LCulFiW80ltn4y/d1dD01MXBwIp9pQBsGo2UQhHX1QzvRk914a
aWrQEYyJeV3crIcIEA9TS+qJg/Oi5K/+03sfVyetkRgbbjcntGvrULrsne9q8FiFbKvk/SqzdS7p
d0xscW7ho6FTd5MUmBeu8fGrXV7feN/+o5jSBRtA1pvamf+e1wtGwLuOnUwi+jmaqtv8EaQ+ZRXq
rPKP5fpywOQTj6jbluL+aQ5Iphvp7UrZ1Ddftf0JQz+bjjO7z+onUAeNsg5HolXdKwvGCQthjF6E
JXn3av9SNjR5ex6/Lg6c54qMqZYUcgX0SR+zQ2mtkZ6Fsf15Mxv6OROehi+pNy5AUxVes7wyTv6c
z6T+ASGpdex/mmnOAVktIr8HnN5KnbQsEEZbeRk3GYUbwBzE5drZRXfDwgxf81ur9BA+/bJz26Oi
6VEOOs51cJFl1TfKOw7XatpQLcyDslbbP703s0/udQSvmTkAhjfBID+T8p864p71kbYz4QaM41OD
kyj5xoLq8CvbIGmLsXkAAJDLV/KhrRgjdt6CfM8ZsYHkspxJHhiVI81lvpbUFnO6lcXJCpSKTRp8
zyUITkhnrWtQDJcC6dzRvC9RN2RfFnZhoPl6T6Vvej25mD0wQvJO8ii5A454leTEQriZA+kPmkxP
qxR1SwDOr/irBh7BUoER/GsMIHWzYCjbBI6NG4L6D+mwQTtBQfF6bInMycgm9DH/Nff82WqOZ+vp
ApHU8SuSlhi51/amQw0KDuuOTRFrX3QcJZDQTQtCUBNKlQJg32VJfEFwAkoA3Y681TqnPLFZy3Aq
z1MwqorM0nlpgmcmqbkQI4rp26Q9Y98VAr4Tx0QMpeCbOjdhYmTWI/iHfsvONelsvKxWXYysfYiR
6QUoH2SLVnA7/A7lRGyTzQID6xDE4d0CQkpLGNeSthtr0CBrV74mGSuQjk3rtsqHe+P1/bANl12G
SsVq8d/t7h05Yt8e8qixGI43CE+/InA+9a57FG6iyE4vxb9+LkHl8D1KxAS0ma+o3NHRKzQ6Lu9T
PUhn/5xVMGbsyBQ9rv7bafK+TghGw6khE+Zko0yASFFmqi3tMo3phZNBPt2VV60CPMzZzzPWs8f5
7C7fYezLd3NsZNS4wA3RogmVOrkudvhl6mDsZ8t1o3jVzn3p6Vsh6Mvxvy0jmAGiw53GWGpe/8xb
ZsAMALvrBuWQopTNJAF9Ms1gEPy0XmlD60gvplz3/mftnUVGVFxdsoU0eWkZGInSsrE19jBGekXq
cP8kpmXMO9bvhD4L6iviHDcNHQ/INNeEieeMcPseFjHociURaoMF585XPR583AvvFr35OUvvhkEj
KBfOrp9JhJ6nZpTPS1d2Q263mXwKfnszjY+/zoELWjBslDCAVAFEXdpv+qQUsK7HOmgEcnQxfPH3
u3Ml4q0poIIkqPZ/Erw/5YNZQR/2I3ytDRE2nBgG8pJt/G4DmhfOXwKjGKdiVurJEISGE5DISdO3
FD8NgcQkufRQbN0AhvY1ghaXw6WzG73tHYHedF2dIsuBUHB+EYPFktlm0BNonWmafeexPSyegB0A
UluIQofkbR31IsNhqult5eWs6OUWeG/JZoxOp95oaXjEwUG4qickOKm3FAJUozJ2662zSCTDL1l3
Ajx+GOw2lph7LsOlWpGqKhn4hqiL9FySYvzV5GSTG9nc7D5Sfr2jwv1gfaDxa9tdn8/NrAwxyyq3
MbbSRlPOcqoL0O1TnhRox82om4RsQSxMqSNCjK+4J78oWgTyfUM0Wg+JaQPvInrc9bbL754Jy+yb
woj0ikJ+r0mPav8CbnQQYmAZyPzVc6JvREqZYjKjTlp5IOehWEDh4EuqGJTnVprtnBHc7DVAlJiw
0fJWcQg18sCMX1UPvWh3xMZ564cQUaYi67wJHXRhxMmEi+rNXWI1SOoSXYzNrRBEGgYhKP1S7nV4
2qqNHMt5EikfbjANiYZTUfWXxXlSlCcHj64I5kt+58EuG1yuE+dgVKQ9oVMOCGD4SgvSsxLChxeD
TMgGN1g4LE5VSy5IcJYOVyxLPG8JcQ1EVV3K8GyHjw0+4BCBv3+ji+wmEKfk596P89yPxsfFvhzY
aTJ3W6PTqmZo4hBdPfTyCR/34KqotR8g7qbV9GX0cPekyVwJq8LLUmEaDJR7FaP/PEy8w9HKgzkB
RJhVwrgi8w72Fh0s3iSNYMeiCd3KsqMzF5jjkcdPWzl/Px840uVXA2RAW95oNhxrCg7UHTeev25A
BXzqOIPIdOfYMXsxXu13kJhSI8hFt0QFeDevgZBDWcHjocTrdQGJPjIreFgf0lHzejW026RkFFV4
RN5LOOUy5s3YV04UUQeVB+onovCzkWUp9GtmzeLPd0dA/jvv4c1poBwweo0ujogl9H3SMdDXjaly
oOITb3u6s//DDUfoOhFoRsy75YebXeHDHARmRYcRVrD1VOiLBmJjB7DZ64zVvUHxHHEX/L+/aqWG
ogMbD7UUhIC7hiZgvrgaAbR8QLt9iIRhrSb+ftpgdc/+TbfkbO+JVjGVyHu+GUcV7rurqrSNXW76
HdmuWwNmG7XSMOQSgfCUWO/OduV/FqOPBkTZAOapDuVkWbqYHE4K/xd9YLqPen/vttwqfJRz3DnE
m+eJXn+yXj3/4PH4rmCRQhb0VwEr5UrG/1VWA/f31uS5xC8DEh8Nzymgz4FtBD46TS87whQDPAEr
7h0BBUpcKETE8D8wDxuJqHX5MbbG4/vwqJEP1/6H3/QY/M36HliAMlPeGNH1o2UDypwFG89FGZxw
ysFl71unvbsEuc8nsjlKNPD17QN33gpxL2K/lBV06aJcvaDiCcI/aFND5mJiqJZ2iFNVuF6kEwdz
NZfWTA8VB2Rq0BEocXbuijdKgKgz6kuu9wKRXJh8oFPKV9fq5jMYAGpNMUFzP7V++Ka6oEz2GH1n
K8PS7qb/EjN/84fwzp7E1BP2HultR+adDA+n6XYjipGNX91ZIqPfJdNiYBe/3Opuj945NajzyVHx
qFv/DOTCrxBTPpCqGdBol9u0C1T5UpI/7ayHAJFaddIy3MWpfYkCgsonz0d0gsh1DbhsyNM4xcGC
qZrF6Ah39E/xudMiZTPiTA76smTFwu8A3RKRokKKis7wgVy6iKBvKr/pTtuyZjBrXmt7ayEHT4jx
osbi7TOTint+KjTsW+QnmPb86THRZ9Tz5blnGdQ3GN1Bu1ZXgzwWYze1kBY9vYJn11DjER7a5q/3
AlWh84AHZwGPx+rpav7qQExhcejrLIkYB1qMmYRib1zNhxPrUIMPikB9NLXP6mmNEFIM6SFhze6b
LGO+g1zmim1hS8xggxPZ2qDTeJ7AbImXiWmLzyIbNuAsZHjCmvg3fxIO7zb6PQ11iQHjp8KgSdsZ
azpHFY/vI4pCY5E6Xk6VP1RM+Nf/uR32nbmbVryhs6modCRnxD59cBW2iZ618kVvEzpgWXb6b/x/
LnoDHq5nQlWpTWA5FhRskKOYqRvGBK0wP1yTajzZi9WKJrnhgrMh3tO/PeDMuX0qsXguYhUnGhMg
/oky229TDv7Um9zAXSpQMls1VFrO1kVoGKOBsTGjaOUeae/AsA4uBSnPKuIz6u1WyNbp/Y47eBvP
UzMUnbHms5/HGeDRkv35ELvzkf7aGO7jUZhk7BfMXIMnIXG7YKcjt1PCyQKNhUgwWesU62uzSM21
WiH293+QZLZ+8fEsXz8GFKqKXUAPYC0oD1h7M3I4AGRf0JZpuQXxccix9/mEtYm7TJGv2HJWf1Zj
Me2fxx+YLfRP/X55bPSpR8XesaBVL5pQ0Ueg7MeOemMqKkq0PmWhSO1Opyar6QDrzVoDGDbC/W0L
/qZEW7smlOAchP2nYBypMGTOUKyywHU18gG3wW88Q9qM43+0Ntt6Ozw07iMJTpX4tHek+7ElCURP
Eo3g4vyf1eqkztcB8P75CRbuof063EDPLUj3a5Sgeh617IsYChUTiJh54K9LRVF5IyAcJga+3l9j
76Okqzi9GwX+h8+N6vZwRQ+Vi87NMtp6fEZvRGN2FfQKxVDn2rox6ELNBPyQUIKgRjUT7B2c8lvk
oidQrg1CxmfG2UV1ybXnb+zA5aBPsYUfOiwfog0taRDd5Tk67h+5vBQVDRmp8hWGEB2pu5FWRleT
NdbdWT1jrRCicuifXqMoNJ/EOwo2QOHIAs5op7X0AkokIfawydU/iPbzKOYEXsbXqmxmAauWS6YF
oMdn7YqLBhLIVNFajpHlpWekY2u9+1/vHXmUUQvCWrVyche1CAZrJqm8sq/XKOHKmkiqX3HisVKj
qnrOnAsIYjCrpvQTc41bxGuQUUcV2cR+yVRWQ5LtvEX9aehx6KPuv9oLgxWFFRzHzGrQWw+Ug433
yfX1wWFg8/6uVxbxW4h4J+Oosiv56J8dcwpkMXOQI166j6ptm+dJ1ansh64tIEx1hDtTZn/bF0WB
+ryvK9Mb9BH39805k3fKqngAA8J93YPSyQXZXpSVmM9RV2hyY87EHFVJj0qxSnlmP6U+RNzVAA4r
KkrwK25FZoPC916O1LRXObpue+EAqyl6A1FqJDQJ2VX4jeG2jrVeWV34PAHlBnzuXMxzBn1gLkry
mHnca/5jcDpQXcg11saBSe/Vk7L7GStBNq2rA0M3i0T77TShKWEd41AJpi7/g1TeVaR6DBdhZAn3
8NgWlZNQNSoSbOmnB/id8txtVQf/lEWjGec87mcOiuD9842vAqqA4EeDy/oTC8sHs9UGfPgLECHC
p0NPQkz450EZVsCayxkkIh2NugYFFjPlVqoIQZ4OSWd0lbJYkOZtU59UVd9HQXjh9sUZh4ujU+Pi
CT2dtT4FBemcTf1ewdnjw5T8pQ8nu9CSqiQpGlsF6FBLdUFfkxGszb0hpK1HR69vbBKZ8X5+IA8D
3xuTuN0EBhVy3T4FE3keQE7pDWzI3DL/yif9zsx5+zfU6w8Uar1gSEaUo+CWyTgjwXiHl+b7C2nL
/l8MQXY/q/XfVd1ps1H4oTFqjO9xtzdo9e12K9QRAlZKou/1xP9+Id2N8rWVspFvUGIzLQ1mrb3r
CBRCCzOT+WQ8nKCLepzj+DYfdbCzM5gJ3SmhSS7qmiJxcOIIDBUs0MMOGjfXo7phfgAiDWOs1ADt
wXthk3qQ1sfdj85RoBUgK1AfIRtu2yKxO1YXOflO2gp6LK473Z6lLqawY3SEeXr7zgXn3oSOiupW
8kXjvcgreTYfNRtJR6pTuYP0vFQ9LUJSI+WweCQTVeiVym2FFghSmMJt8fgoQtknv1E625m2JaCj
7OMu/P527pnyVpd1bwod+U7/uCzVLAO5NR+8T427QvUuSPWAFVEk9flWgTb0RD5O60cjo+b7HXYV
yquQfcbijAJzd4M8ZPeWUFS2zIoC2Myp30/1tgRAXrkOw4sKspi8A8eMskqkqVKE90GgmgL4/fSc
tIhdxeT+1GC6SRXYpJkkXuSu162Fez7OqQnJb8LXnINvBlb9rF2iLrljtA1sjBPb7R4K5HghkdoH
IDNksm7011GD0vxLTUyAD1RfmCT7XPPj0CPbNUnQo+82a0BJQVnIMD+9RjwRHI1L53/BNsH6qfla
QgE5Mlx5SLZ7KIYKvIQK8FHRbqw2bzctewE8L5gxDil6C3vFCWjZeczfSiiTrZChX3fKFc7W/OU6
5xqUan2i9gZDzqY+cP98vrENZXqFoJmf5+fj9XJIHNeFaXvmVCVL/cJt1h+wVFwKxIvIZD4jtJOw
dikA/FbhC17a8p2y1dJbI4+ejapEZ0SnwcXEvy65aHh0zIRcP/oW1ZduUlUcEE/kdN7hITkAa5u+
XuOo1NsIBQyDDbnIQ4XE+QPa3Vp9bRVOhE1fuU0s7rcsarPxZnE21Us1hal4xnj/NYCDvw/swYqK
UsQyZ3ea8jNCIRwbOm7rJ/xSrIEBvtRKZdipUVc0YC1cNj3gN6NRxLJCTfj+KKlzOuEMU4ATpjGx
fGPmvq6Ly99Pe3xIoHT1iYyOvQOSZ6EsjmkwWWh54i5cttiEnpIIeR8+FAlLrUnOWi0L1UxLsl87
vPcfejFpZtFGUAg4aP9qg04u77MO2ofwzkr/BXWMci4ugezxgJyyjKDWlo4ovGqQzlEt96PstJbh
tHIAqf+oQFZTXoIpb+1lmUWVljfNJEa3pAB7dUwFaf1RQTYCfPGBD1IeGnN6yM2vVc2uTUMf0hbL
YMQuHnzZzbCtHY6Nkk1Gn1KXllxgXv9efiinmbUgThk0rMXV1E4FsQYrNayOMuNBm9got9MXZ1jl
quzU4Wg8SGKjH1Z6suie/tOz36gXLzRrnWI/HU29uHUHLy8Zu0N8L97JOtlJCCopALEFDDPoAma1
RzdzlPJ/zZygeTH5LevPGDdAfjXzW13eAjFBG18r52lvAwCn+0WPrx/SiUvmd010xEQEiB6xMueA
pddJOFrV3xXM50FuEd7be3C4RtuVwi8sJZdy+rFYfde8Z5yYsslDigYtxWN8gdTlQNduo0+E8syG
iXTARNl8x6jeJv2ciYZecgNxM5IGTnzQsAvsqwMWcAfRGqllXD/snVU27z+kF1GpAtQp7FbnC1/q
YClXrxB91l1p2ly/9HNloc2aqmnt43BivAiipMxVZDLaMGhe5GEYO6z4mNz+m2jmQEDLCBQjZ2io
SMMvacC2+ZVQ1L7v2qq06yx5bmOFyJkPSX154GJW6FC9EgG/TSvbU14EYYG272oYq11fbm9fiPYG
yIUxssm5vDD+dkmVjkUBBTz0QOKLvH/WVzu4Q1nVvdF1OTHbjMUUzCZsDfIp7zIL1ECeOO3CZfFs
4QzIwR7G1n+ueiatzzEaaWaeUmPDBpvrIsDdRcVRVdDsf/bQaeYpGV1Hjzn5lCamoJNdFhghLvIw
+6efkssUj/TyLChkhvn3jntYpbJtEpr7UaPyuwHu3EfZV7f7CY121PJNtVylnXxWmgOvIijV50RO
1Mdxrq1tr7QqKFKYWJyGDfdwo6EJPQ/0i5OFTI+nhpsx0sQWjYq9WwlfcbqRbXv0iH0efqRCmtD/
zDYJ2bBn6Zc37c70CE7Uc2qWTd8xoVwTZnnPxywwQTXZ6RRyGoVGWxYq1KIx/NtEtYTJNtPu62ct
xtCVADG3tsj30I+feTXDeUDoGQDWu7z4Jw/POhjg9qUf4I0RKswSjRoLUJ0m1PdHEQ4kSgERN0jl
faWyH9K6HDXV325RfbmRbhhiYUoCFA585PkH7uzG6SLUAcjW6qbRMJfXL1GYPxaihTyQhUi9aKCZ
de7tjlngpsUjOmj0GvHdSD8s+82M8W9iucYYfXVhNPQ5WrqMKzj71WnX+lafLMQG/IfcRnLBIqk1
LHBjZOn50WxT9FJhudrTfnki0SkPDlzJK+sutkcTJpQv5NyE4JfxxPvmC20jWkco6BMFwgeJe+Di
eg4f6bsTbWlXhBYRoRbWfrrYjI0X7YWMUheocWkTGoQ01tFsOOcscF667kqrrRf288/JLk3biI9i
gVSr1JZS26Kj9vrDnsZIt07XKTL2Zq5QT22XplJceGoRyjVqcjZUqnKy5rKrn5GtYuLsEKZm1gmK
qhy7r53uLtY/NlxM0zH0RCz7CD0vrlNliMSOePnkcMxd1Ni7FrJDTadmUbD+7+q4nkxFDKLUZQ+4
yUEDh3WHH5XlUV85Ag66uZfJDXgLqraqr37JiO/SiKbYBeB6/9g8+DqqzMaVf0LzrQvgthHImseo
7RYGcN+s6V3dsD8RoDexHb5vBaN5i5ZYHBSY3otkB5mAByjTc5GP6+iZaXqrp2QgCY75EiMTp/7P
UlU8aAirxK7e4AiT07YRu1vE0WgBw6zNjMZ1iuSIqxhOpyi8eiF9w5rxqYK+jae28rulxgvACFbZ
TThuR9cQcVM7DR5+WzSMpXfAQPayPg7tOnnznFTIGEAoxq6z/6wHBZ8K/fajT/TP6lQSyzdmlZBa
d4je56NgR8Su3fX370L47f9elrQSS5n9O3kqtgdBZ0bNEzXWwYL+7QfJBJ7ap+hLxL80I7OcTJ5O
FD6Zdxpksalx70c7C4NUBd2AMJAnWBv4uyTlfXX5an+nf1AZ2/L+Jws6yKWNmNut5cd4SstDVxLr
jlC8uUrkmjbOHiw4apTejy28Nc7M2x4F942RdltxYT/dkJ2zU6QazFjWl6gXPt0MAubxnuivpx9Z
HMHDe/MYDKjiPjk8iFZuXKM/F/uaSZwBpl2EitsGl3P5lLThqw9tgbj2W2lYRVckw6F72aBvak2R
2i4ITigWCFNC8xx/Elb/UDokkCw6Ihdzr9CuvAUUbY+vzkEJMsXCPNxg1IfpdeazSckzsiRJNi5k
61v+tRGoB5ijQchREJZ5kF9/41Qzj5tVockn7/1RM9kz59USJaM2qxLyqXIzazR9ebKiyxpMZ7t9
QZY/U9bcl6vfXJiuXcRrt0arOO9XBAWpPHZzLEVpk3MaIg+bPuvIRCKKYZQ4XOfSCFL7kV+wBQpR
yJ9BobfqrSKj10IT18YynKFc4LpUaaNIv1Rb5cpQ97Xi+SUdZwmwcmeMxk3i02B9JICFkbR4DBaC
jBnMnc0Im7PuI81yPusawTHi7+7MBy1Ru9DOJOfD2Ael3wYcXzg8B5fDjiiniJED+HeZTGClwYWr
K1E8q1orKD5det8QhcVKLrLAG9DdKRdLGp20DMvi6neak9IeoUayiRiNFkYgTs5fZ3aB3q91ltqE
fzt/Vph4cQco2nufX3YDkNsYWOezw+CvsFx707spKshY3OnIj6rQZjFkKLV1nVW3xQjXki7K5Gtr
+FI1yuaAnFnXbyXIhH+pWqGqDt7iSe2A3AUT/DLBoLKDikN+fqF8LvzWS0ItE8GS+RISz1sHluGc
PGVVpgCnph5jjXd9xmIKVEqJpvEE3iaC92+TSnA8gH3GIuz7D8DINjXQVUGTUY3NL5ri35L36Jc5
+MWRsIoTyogMegKDoB8i8lwTpuG9BEr5EyDTCzpO+lJIbjBdsVs4F0pU5kLfASRK0W4IY0W1KaBM
Bpc/8YQkQyBP6vlkrNUGaRAvmWCYKd0TUPNGZB0UA+0SNzoGfgZZ7+xYuOzq+VxEHNOh7cwIy6Gq
wiWjMa6nv0lbAkhZEuBbswcMyzNl4q1BcH0kXWgmf7v3uA4ZaPbkLCuCww+hH/l5LiknE0S3lApv
hpuXHFCjr2Y8mgFaplv/wBF/GQj75dxQ38LUFY9zCJMKEzviPsDNM17vcBrWwoAc23s4qkYu7bZ1
C4XdEkWCmj64pJVcDKfrCeiWdX2ajIJCR4XfL8p2KCg1Z+d4wuDerqeETMQ35LO7ADSJQN2AVGCp
X3dTI9qz/QWiPUr8dvaCeP18eWmNQi0bGnDNdqpKhM3vKgQ346lCmcVKrLpt5JSBLCvaPs/5Ctsm
JwSqzgqGcz4SE3IpFumlhYkD+Drq57ylQT2DioHYdVNce0wIeOdXMNQRScSzuBGAEGwI6gb8KObC
fEql1TT+ca/jxoQo5zvni87kVoifu45aEayRHuE4HcVtZ9IROku1ppMqFIrj6sSomUSHjP8UOFvn
ivZDWUpiFgDNteoot4G6VEH4BSSCa758cUmIfyaJe6rRiBXHxw4J66smgYMjZ0pKZw7Mou1cD+bD
qbRQ+MsZ3AjCeFtRhd+WaaifFQMg86b6Br92q2HIGa1yGNYXdRPR33PqZPtajx26JdXApO9W7fd9
0Nh6LI06YsX63n2ORsNKR9iMW2VuVJ+WVy8lC6+FD2shDhQeOvFDwrsllG9mGEY1U5vTedYOY0Qn
y2f5HvCe0ZtsPVD7BKG0e4XFYfvDU7+gqANinahHKcqHU2twcyNUAgKXTyPyQHKdJZH5Se2eFXf+
Z4W8zjNNrEf6A0hNwVgggoNE1bTuSS2nHyhwqLdxhQ77xXE9gf16LzBFrWKnN2jF5HrNKW0dpfnk
qnXUjgvb3C86dq+y33EYRdPxVnj8yucWGFJ8dvx8Plk696eIOacwl97pj8CWjNnEgRjsp9tJKP/I
uYmZQGu4rl+5O3/FgzGRimZjhr5AQvsIDIaM1jbpjaABHNHCnxeiCkfIZ9pLmowE43RS0d2o3Tl5
5sDSNCrVt7U0NlmO2wU5W10BqC+Wn2s0/Ldu5/o2HwKkxl1P4KAHnUsAD1V99mT4W89BNVnyPsLx
2EUwMzYPjgbPHtal4tYCexTv9xFTl+CPvNgSSiRzJk/VU5wL4B9/A3vtQJ1tSb+7La0xTfGq0qvU
ej2b2qMjb2ozIaPu09wNiXjBcsQjq4HpMLBUMhegdAfIE70khSYcru1QgVp8X+swVtwTKkcTmy/a
pkuYHa+j0ecYkzUQlKMfWu1SvG8chs2EufD9cRhzy3woGlbtz2w2zd8COdEABwdcTlzkfTiyOQMz
iq4MUWYoSPoVOKCRMsINJz8sRqIvZ7vrWhrL7YxzhzooWNngA9z7o3R15sfiKS/ngieRyBY3Ew0I
z1jX44zh1LnTCAL26yC8xgZD7KA/tJKh/2iokCwIyG5mq5B++D7pFdhFNFgSITjUyagqfSgofYaT
sjGb5xGKEG6gUdgK6axZliPn9LpIE0sO5gTQ6FVjFlDDCW+5G9p7UsUSpMoOwzPWatw54TqsbJEi
uXoWKV+sK1GQlX3lOTPPJkv5ou/8uUCyitKvlBmDCmVTyElOMPEvLMYxX/r9NIy5dj2iUuBPVP+n
3brgRrsqTkSqXJp06QWYzKgnNzVyoHn8N1P9VgYidTWHGZx8hTPWkPnKQqvQc2TBWumWtsFFIeto
ZgN4zED7B6hn9Lf11I5PP2g4vcYmCL6MnA9F7i7msCCEI0cLw1Hzc5maSE6kq5BKfsftKZUYbCOy
mpbLRM0fP/f95YAUEi7JUp7zVHN2KI2DrRuRU/iS1oaEZ1JE6zunMeibDJGMdnMtgTi9JsykdQMh
0EtV+qGYlRdChQhDA+8/lpd7NC28VOfOYZwQ5uDDmSLN+VUXqBa2/q/HSG3UyWho7VBbEF/T2i//
x6e0bKOyIyqhd5yaTfTjcKljXj9gGH+SkyJNf4FHU57u+giL8jlVPSPJxEb6TAEHHTtLNsY4q66Q
CbzRGTiSufnX7CVgq2b+K5L026l8rgQ4YL5ur5FO7SqL5C5wkHgmnq1bzVzkMTTnsAs8PImPOYXZ
fjuftiNRYBGIXh+u3KW+byL9uoPVwzm1fGcZHD+QL6L4CXcvZ8DNwV5WSn3nCHScs1TiPYMF6h2k
c62ieeDVU1Dp5KF7iXBrPng/3F8IfZEwQlatJ27xYrHcOpXUliKblkTHn1r1Bz1JBEBGS6hav3sy
4pe1cyl2W91uQhtgfbYy0M9+jqO5G7JtNMpOchNNfpYR8W5fybny5JAy7fF9TRZLzGOIPkeiAgX2
t8q8mj58HQWxIdKhS4/IOCRpIr1Ch+0tBuUy96C+KRkdMz9vSgzL2wRTiS9Pv4JFAu62+xkKOjFK
Ch/a+g8Xyig56JLL/DU3Vc9xADtt5gd+cCOxOKvLpLyDNfa1KRcGys3TTBkQRFcYGKTf50wzxJE1
Tfwml3n7ax8OBYByHqaN8Ag1BFt8KxxSeQxjVYECO194nhdSzRi1EBFLU+DTunKx558H7Bdmy7Jx
+R7Rk9HaV/7IeE0aBKqz4EcRFf2/M/bszS1MPdDnTpNWj92UQkxl7aADT5Az+afhMy3XXRBOkGOX
M7iJyeXFMkXvuv9eUVaIDu2zl/QZuMOeUs2QDSJh9Z+DjDG3ouBRgljNx7UqZ4OYalUzrLyT5lvZ
Dg2cYZF7lWk96Vcb9Noz8XmdTWH8FaPwd2TAzOdVNIJFUxt030oFzU1VPf4qt4JcSM5bwyQ549+/
4HiNvXSU+fK13JI+7hve4a9Y4muWZJvDIPk4oy1YgtnJdMmMy9dPM/Pz0KoQpAutTaCw3MOZ93vw
he4zL8ERMpBzV7l5E/Q/7sEBQC5GRm4doBFsTSuRni2x3adUjFYGhstaZQ1wDjtoNQNLnlr0mhG4
oQiM5rMKys6kuhOH1+C3ydyxhiVyhSWv7CbnwgmAxmgNStd7Os7VrrlktLnTNDYA8bQHkVuiMPUQ
GUo469evJ+n6WWuOEbP23aw0bHebwjRwrzIzAvQzLRu61TXMshAQ/bVGrka7ZtgpyJZUQFNV0t74
UMyEgKPUiFRfj5oKXWfoBP5zyPg416pd3awGnfub5pZrJi1YYLYkSu3N6SXtobT6TCFeZckjV48d
vICXSHFXYQipmViIjtNwTRTWoZyc3JPPU2/FW7KH6ru119LKCJuDB2vuRifaiDm+LK6bqKkV/Nsn
Qnylajt0y8D4biXJxUj7zT6mYbGCApk3tpaY+a1btUZcgFAbBWquAK6Z6wvuS4pTW7YrNxc09zPB
vbkYnw6ibwB28H1m0Nm1hVRzdakv+BYPY30EqvwDMJuEEcvA7YFKhqArMWYrWCcTy/9uMS2DWzzW
VrL0vvR/hlIwOd8trxHBtdP82UXWdGFViTsJ2s+KWASc1b+9pMKVdZu80VhYHQAFxtLp3XzCqUJZ
EU2vOvcrmA7P4/MSEzrhBSmqUJooKxxuIYH5knuGCTpSFFyWKY8YPfHRzHJzvZ/6+pPeIKyzRK2f
yG9fKRA7+CG1aCx/atbPTNNVqpKILmPvwc91zy0TS0iMnvJW2vGOrNICLG9M4iNVDtb53ITQqpky
susppVFbQhVM+j8aB/+jpPXy12U4aqhm2YjfHz6tQDCC0B0j1+edL/k+XQq2L6GGuK/nlP9KnB9b
+lduBz26V6n4zfSVOdfMRJ6sqLQF6nuuvtHNCXKI6KFvDjUbpyY2erFsgCLuCV/JUqrlgzphTB6o
Gkol9af/MvLfPJIxiKCD8KkVgfNLFoBnrRkLugN98hBFhbCMdnCx6cYA4TamJiUARc5l5d7GpqXY
yI0sy8v/C8GenEJq00mUsA7OFEY299LxZh2KhVP6HSh0YMkXFP5ES3u5m415b8776XK6ZG+v6tEW
9FQypqGAZzARpD4b5WuBp6nigi5BuT1ap4HyNCTuuqU7amh909otoS/5Bgt6SD/W5VmSA0o2rjCe
CNRrUBaQqhWlLb9xXieEnEPMfy3VP8In9sqjsmK4XiNd8tOUPDr45BZLsOOCCNJWMQQO7W8llXJw
ZIcWejib+z63pqTDJZPkqJHMupeTDcdUyEg44CU6QJu60gqLGLpgd4GRHfOAO7jC0dEI8eX2+p0i
mzRsPQXEa9R+TuZ4UZPcM7BLvJWO10xwMdZy80Wu7z0pgUq6LtzycwdWiA8KrIHmD2Cl439m38wb
AupANLg1r7f6f9ImVcP+A7vUBoi8bpXgOxGUTAlqUX/S6/2BLqMRObTrYh6zlUgNbf3KZ202L7Ap
Aqv1prLK1dn4bVC8XA+q5X8tN3MzGjsHLqmH31R6oT7doKnxwNkEMyEmMEWSMZ1eocZ7KI3NAyi7
N7oyjuWczYw3CTDlY3yANqH7UbOXAkNlbJWyhIn3v2Jn3VRI6Kbi58wQoj+5K+uxsDp0XYPbs0WJ
WAFSDaV3BF8g3My2D+fKYL/xHBvB2jC4OwLxNJDetlxjitDBsnXLi0cukzgCdbNE2IQ93+N8fDSH
GliDwsAyx6J+yVaGSX1sKG4x2mGmEWnyZMKs32kSjnZcLeo/rJw6w9vj9kwaXMg0mYXfFNgnzptM
J03WEGLGndIyHX0IZEHXR3n/QkGZapHXr32llO5UejRGUj/lmAik9WAEh6vC0to/OFrimw5YJBHq
1iUvKiTFUufJ+uscY7aKgYZpCkpabXRdywLuWPEWsiaFWMHFYMd3I8yEs7u3AzP8h2YCNqVeN9Xs
nDsQ0bQ2bO13djqWkKMMcCmRHEWrgVLLp+Ubd3tKXU3z2CYD5mSlp0sV7WHjpCO/xpop2lZvuN8l
k1wton1UWFquhwFS3RsMnz7G1RgPAj/KzMpBN467NLiWbffhGrgmDm/xgrMRMgNiVAbo+Kt2uCWC
LKfnu4c/UrUnqtqKtu8arKwliB4n2yBeLx9Ept5j2RdraPGNBIKnVyzY8nVrtuLfaUgYykD4ds7Z
MkWKMtviMRGPhctPsQRlWOfT60hSQOEr6xBVqXqGJpknks+Wj6CekxjIE3b9Mv6HojFBNVbeESEQ
jeZj1WhCdjkcG4oVt6yWzMVopt8jt4K5q6z04IgccqPwO5CXKdsvUHyotTfkbwjRqjIh3/x+7dUK
x8GcMeeA6L09GJT6ZOnT6yZoVtIhd5ZcqYrTsVNOUDKVkHC4eP16dOF5I85vlwrYc6HKbWf+oePk
AnQtiExzQreQeVTW/00rF10tf44MjxiW6hxpoy3qjlX8YkGVq7b/aIuYyvSFa0TYVEg0cRCM1ZJW
2QRl090J4HsGoTb0p3Wa4lA7hIVQ45cnGk5Z94fqISHzYtLFp1nGsXRvtlFOzTLlO0PCWkIfqlh4
zwVj0JdtNIp3H9f7MFSEtH+bXNuno9nQilcBo3l84+UsRO1+LAGYRODZ3N4arrJ8WsBb2qEFVQ8Q
Hwj5Wo83V7Ymz+Muvrr++e/Ov+GohpapqFroKkdPvL+jfJCp8uO2XQ/VLqLcd/fjhQi0hbRffu7q
dwgbDOi4RsAFFlRiN7oGA1+MMv0rRSDwjO0RBEZksmoW9clez1jHR72Mt2NhYPXBz5MnBc74aOvw
VQP9kAcomph/rmkhsEOnLM5vj9VX8H9j87Feb7ha8BHI7yewzt4eLz2+zOJ43L0hs/xAi64OhPoI
BBVygVi7ldAVRctvQqT8J4+mhlNGC5BOhu86pTOcz2EazOIgCdiU+sWALcFqz7T5R1PJemqi1N/V
xjLX+PqRt4VYgwexTasm1GKY4wRzByhF0gnwnQy4jZRmDCgacqTqdi1F3m7SD14qyGRi6GFe2W38
QgtyCcf9ZzGr1tZWdIppm60vlNNJwKG1ptAISfUGhBDid2QHIP+Br/YkQ68WW6IHtKnif1AxFTcZ
zGewV54K6JodEXBFprGtBtws0EC6UKJ4cDgSNo9itsYE6p8ThXCi7SZVly5VzPU//6KYjOso7eoH
Pt1x+lE5pHJVYQNR8l4YK/WV2LwdxUELVghNOrryIJ8qEEmmYSQ08kB0LRMFz2/4GOM2DlkFIn5/
I/0vqkm0Emy5IWqoBBKDL0G0H3or39J9KGOXi91QXNQf2ZsptmIEsdJwVAiNubZaxuc4SaG+AfJV
RouV67+Vi+3XzdXLi9ESAa0N9MdboHw+7LIbdYBjh2DFdPip7Ea/i0L5iPjgR6gBUraycVITTiJO
3BfKI5UZnlqDTA/f1pwmhaumiCKwFPEJky1NeMOsjuGKf5uXuRlQYi5II1cvDP9oIIUq0r7EO+wT
ETsztDAk+FPlZBIusmM1fL+mDA9Ql5/RLCyiabpJ3SuqcYsySCg+/Iyebn2WLGa8teIOJzAdf6EO
OZQBeLCdq5d4d3V1rK6IAdnuFMbQTdE2IYtn4VkNhDNNSGYiMEY8sE4ox62hWfw7dJIw6fXHg247
A5Pjpm4IMwryAz6axSYcNjOjkESyO2qs1SLyk9DXpsk9sJ2+yiJp3xQheIoiDUBu0oMRo5GyqUWJ
fi1jENVylHtZb5z5wnmYF8vhimIE2ltm1JmFLqpD4wDiPo2nwho/JMHNLWo61qtyNgR2FTvtCQtX
pOOOEzmQc9AAv32eE6yfPmhYyNhDbrk6qy1meRSugySqK+ojiLc3R2MosMhzDSI43oTQW8YIaSRX
a5V/x3G8sZIsKRKKnjSVb6OOVXf13b02uggYUrjN6OqjKgSfioY0HlvtscFvQab9EFAjHBzX2Zc4
uf4K7cCvldf6uF1RIW3cBKlLdPPe/ys4/THcX7pqaPLRZEhzCsymJ6u8VxDGP6ox61hbFvqivFyL
0n/Ogc90FjYyJxu9H6rOvP6VNoGRKQKWjPUEsgmyORgRGrCq8MjTscO3ET8oTbchAJ1vr/QkmEn5
yOrU7mIkNb4l70Ay8DFvnpIC4LXbM9ImPgJiBx9utTslDdc4EUbYm30THqt1yX0AxAeuYFNDkFz8
wCj+Ep1K5sH7CJEwgYwzKItvV5XMKUoaxVxSOWhgp38h7rLnICsSaU6B7BPumm2aSrHvs2Netsgd
zcH+QfCQSDNegPZSkUWo+1Z4grNShTJZD54ZTzW9NjDthYFiIZMDimO31x+ePm8YiJDpuhxKgz8L
FEYPCu5x2ppZCiOTtXgv/NI1DgiYvhmCuSeNr/KOWf94nK+IO03sEbTwIpU346c1Lx1EV151xWAI
fAkBrW8/AR10Vy5YXFTw0R6qOxoQ55RnKR48bo+sYqI5nTqgb5W3Xncir9CR/RzWESyUFTzNO17A
Rzx9enDRXKR7sT84iwNV+T76fo6aRj+z5aDpBxDnsvdohlPGetsqpz7m0GHy7bo/mitOrE3TgemB
tQiYi5NO7ubexYLF5h7+HQ5ZXgRDR2lHQ4flFe/+BEbnl5yBjP7gURMbXLx35e7UI2mDo0pYygxg
9LVtLisH+MTlxrFXhosP4NNQdsXPkI6htVxaGQp7vnQzlxesp8M4QsCZ5lsJtBspFFrQWI6zy0iE
+TvY6rRRaPONrsqcSUc/yagJ1kVYQPaqPbrkyysPvFMBDJQf+ei87nnMy/pnLUjr59gG7TXBPuFm
jLjilyhqs7gkCzK6unp6D3GGzOtpuKYJN6JNsIKzgOMBfQhqHCQIWGJnZqhW1WvuEnKqCHSg5iki
EciR2eeNyFczBJ+F+bkJaLq4k1FyA238hOlgo+dQoQ1BVq8hbJa045fO1PA+Bp0EExUehYk0st1L
/12itSC/NbKvIyEL+ubcCzU3G2Y6iQOFRQIraJZkb5VYGKzm9kl57HokZbvA5YKR5i7aU/HL4FLi
SKq87mzZICB+71nCxq3Whot2SiEsdV4qlZYYd9wOhCTsHDIoabRojrVrWxZdcrZLi+IG1lf/UP2l
/0ESaoJjSU8iaAxwNgZnuJc+QhUBPT3weKkqXl2Z88voeJGzOW1Obd1RiXSh5Do2+ekfbM2hpX/o
r+tB6K2SNjYJ2+PBQmXhgCPMHgIDSHsZBCK2bYwbCfXyFZ0ceHXlEVKM0EegdEHlKWUTB8gAdpib
Sfl4jYffBMW4aQri6z2z4wwBaveb0eG/k+oG4AJ1CvaRd32NPCeC6H2Ia/Yjc7rcBrh+CbSwqGmE
NnBwikdj0OjBa0TK3YWC1Ou60EvAywW9jdfGyvJk6LtpfmEyvmpnMeDH6vz4AL+GIvyREMJkl2Q9
q3P5NoZQgJ2KocfAvWxazIbNztsnokXb1TyZjjJtvJNMAXpG2g3LjVQap7zJ0pX9/UETqw4n7PJ4
xiE+mZ8ri0bN5ZrA6RJwt7XHNHVf6wGAkJGLNqUUvnCdC/pEuaQ/4755OEmz5IA6+DbyR5MNha03
950b2WcXXEcyeeoQB+wabG/Gca3drULQE9OQZmou3elqbIliEkVjQrueGoho4hkWdrMIA7p12HLk
d3u7h2WL8Bdb5ZYGmb9qT1jkogAnlMAieqKGw1B/0vuS9U2Udc/Aa2AQMnpzWb3z2zsIVMFSGeka
nWuFgiT0vuXpZHlrXQWpm7tjLKlnwzBCydp5TS93t4SNEg+edGF4BR9sr9NBQHhhyT6gpLiEXM6D
x8faLPu/SeNRO/OcPPsZ9NR5laugSOgPGl5awhaYNAC0Kp4XzO8U8+T/Ne1+3inn3gfoqYvWucdX
4jS7oeWuhSjHEF2kXjJI9aKV6ylK3hnQt3KG+v9vIidCuIsLaS/nv529Qqxi6Vy8ONYUgtW9xQjL
gctMgKESpumhuEbF3iTAwvS4/jdedUKL+FCxSwTKbZ0I+CcM4hyQJnOi7VRLVSRaZdoAYQgLACmV
KIHq0A8WnZfdx7BfNjiRTRVZ4FH+OQ0/2Z1KDQwgbhgbh4IEWpbZfbwCvAofDqzvEWxdvWlPhlWz
CQxcLytWb+lI5PpIyqabwu+EfTfGxcljDvZIEVTn8vguBIBVLjv/Tb7nR5s5JTWIR4Lw837TG1FD
YQUx5zx909XN1dOK105JxY6URqTqPi9ozsvkS5v2crP29I6P/7+HgtlKs9G0ykoJ+ezD16mQ4LrU
ABAMrS9fxI6KXQ+Dw3FtQQBBG10jVVpMRLdGLgcdi/ATb87G2iN+5fSqm730azK3mzwvKisR7oDo
Q8kPQ3HAR2BTSAFtIB8TFy9zlgit5nRPvbResFNXKu0CE0d0P29c0HUTBD4UNvR+tOKlQC1XxPXi
hYSIE5fBTdhT5g4+c2UBE663j7mOKWozbMFgIVAlPL97Xs9G0mTZMv4+U5VtctzGAqZ3MX+QKjTs
6dY6VTMAwZmzg9+f3cLXl7sm0/qCi3zqIvrOzrwkrHbmot/CUgfJ10yd3T0cbUE7aQcE5dr+yPVV
iHpGHWdFenQ49FUKLac33I1REduhzT6i8vBYvFXNW7RT9E5isAUVgHd40t35jWc1hUhwcsQGOVtE
vFUDmMeuKhI5jGEhc/guWvXQotVvy5j4VYu0GvO9EZrYpDSs2Crh6cO27OBfY8mUYF18nUbV+P4z
/TlHoZ+WtZYTtKa+GxFuDiKautUw6a8gq1mTwM/mm7jhuBr1VGfCetC84yHEvmJPzAwADbGpMlOg
kkJi3pueAi8sC6aziuKMa7hlkIYWiqBxZrvFYjmF57PONjCynFclGHFNMESv+clc0/5XdxhZo0ab
fiqRsA8MICrmF8Ym9tqWZuDU1pBjqx4ocYyeo9XPbTStCJCnjfra42GHSmsLncA2oYckr2zXDy/V
TAssN75X8NNRHTh/jt1ECJRmTevghdy08qUTf2jOH9nKjU84x7hvsbQa1lg1KVJrBFxeOvNQIp3+
w0sPynzJd53tGAnpUFVRYI5CSwsHG3z6MODLh8pGv7fxKun+Obd9QBCq8q8qFuh9V95s//AetBbC
27BrXQbJnkOnZ1Q1lB1HxxOWbe8PQHJp3r50Lz26X+1DAujoc/+LcuhJP3m5V/qaUAyrvhcR0Toi
Yw4uyF0++V+x9iHeAjz3+e9Woc6UNdl2UJTX6jEuWCfMKbawP+SyDZuMfVzhupacU/XRDLYH4ama
yj117nEb+mhBqSm7OWXJvlM9zDkQEM+Tuvd6qs5U3awMkLn/zCtlkaGZlaOMRl4i587T46TPine8
CHJ6lxiq81fLTMbOsvWGcHlZEKy00d76PZKuahpWsQDxB1MCAftaVZFYs7c5bGJREe9y+/Pkj4cb
rGt4/lgLgTUphWW7LAQP6PiptBIZ2iS+fuxNUmdvkHLhGK3R1cJnfWpYgNremHxUxW8e8if3cDot
6Ui3HbjrCTQoI+UREsTjebWOttHr2RCQlUSwYxDR8QfDazXcXcsr0SqK7PhxpbB1KFsD17rTw9EU
RsJciVBgAkLzHcsuNrEqQCEEqrEl+Gay/IDPKIufwJZqnYW8YZeQDw5wSzdGDjC9dMVneclUqRuV
rkQQ9aC7SRXuDJLAnwTzooMpUg/Pik8bdd6TWA4YElYHzeYHUbZSIWm8HfRUFv1cmnDYpN/jXrfb
WHIw/z1dywEDvYvnxz+vY2IHTJYG2zA65viYQn7GFkjfNnxLFkXFv/JfMPG/e1847jsX92HUBHJM
YfvvL7NRyoP6TBpbV/2q8AVZvodTMDl/2DIazVVLJILeYGTXLm+U/+VaF8W1aG0F+Usv4UDiMxnR
z9/MQBMjjOAg8S+5ZMG5oIZ9I5CdL0QLJ/50+hauJ8NIQfcU0mQNo7Zx7jj1jMSMCmwcNOJWlfrO
kn6SIL9XPTevQM38bl+R9x35kmZhvwZKxp7C/5rdZaJajsnMTew2jmhdf7wr8sePsiQmbott1JRf
fgDUCvDuWVyCY6gXrFTxhOsim95c3osupYt+QFRndX3msSQYjDVIdXu2iJRu6is6CZ+Fu6o1SYvL
ZjnP7gq91C6S7kcVRv0VMK9xHPryEVAaPwPKjw5jqNwOUX5ab1aFdpe9X9Ja5fTOpRsI98OnZwh4
kJ63/9DZ8cxGawjZfwYfWHI3UKL2bPYDgnyyjczFUP8LabKBkfwh+6qSGjDXHzdvR6ZckTVS4GC9
Pe3WVwP8uuDeDsjQDb5/UPzDVGCBweacBJ35rM77lJS6CJOi7HaMDKZKSRA8l2X3HPfYjMDVUC1o
nukYM5fN31CkvKcq24cxlDvP5u+DWWqL/1m1ZZJW2ITG07UjeX0aX8XgO1xcHj8S1WIw2y3b3Xin
Pks1Qyt8CgsoAJCH1XBvxUJY74WM0Q8vXK0kjeDLnLmDxprDAmgyb9yOl+Yrtlj1xIlVjJ72/nDD
T43B6KPCPZYBiWkAxM0BE+AfALRb+puSnhg8pmu2eJqxBIyGWRRXM5Et6yQexaCEjoPeAxE7OWc9
d9ZKvvDq7AIMWaj5eZHpFpxtukGQ/50iAa2jL19y7oSle9Pr2JTpwyPJd+5PJBaPNb9NhWqt/yXh
kusXKSO+JpWiCshCZQURx2m6p0HReAGTXuKltleGUfhadNVKGzleV7XPMYNJX37AigeN26Ocq+s5
64znTi0UVMyhnNyONvrrDgU64BqXQC8eQ4AQ+Rv4ILy47S58qUFjv8AWCsIGseIEQfh6GKLQXNB+
x3CXhoyoN6kl5+DR1K6h5C6Qk7eyo4wFiTU4cZcyg0BSeAwMFCLhVCCrqUCcwr8FDBvCSfQngPuZ
JjtC/5S/LrZ3aRL7oJngJFZdjhurMI8K3gArt2O3xWEDaZw0AugUTk01Vkm4LodB2RPFSro/uZzr
7K7tbgidDuQSQV39e0XV99QodWB7+9+ZWtB7PfV3U6RdFxzLgNrV50DebcnFWQK51cA42Svrmafr
uP6nASs1RHzp2XixeZwGcD9UWDbxHkp6W88tV7NnlNgcwzL0LKDvziIFytsSUtHvrTnaES9PIJ+f
0aPThaid6PTHGc8uj0qh0a1y4WF8Q95WJuXoq5/41bJOkEUvfi6GRWDU0b18mpY8OFkUGyoGuhHR
sysYQzuvWSgWBpAJLrGt0Av/PgzHmgBzrZlM4ILrVM78iTU1oojcAu3bfMcA1ZzJodY2betFcQzr
hjw3r/XdzEiFJmKmKYgtHpRQeT9z3fgFFlHq1Zw6wMG+2EWjEPuYOU+4SJeB87ATlBB0xD1507Wr
4whP5MKDY9kf92iVxERoc8E55ta5kEykvglcO26oGBb0fBLQupN/W9NTFX8FR4bvfR5oI3BrqxG6
sZAFunx+GNAW7v2x2a1duR52+B3demMWHBBzbOy9ZLFGCEjCjmn7N4esPqqOf2sXcpVyhA53ssCr
H4XFK3FTo2qVA5hNExW11ZUowSxgtMFVhoauK8eR1s5yxwfSCUKlMLzYfbImgaYJlU5x+0AQP+VQ
5ge7hvHkp+x6lkziFAqSA2hc1VG2CrgDQxcoDEkXSn0eLB7gbWqZWdxNkvLt9KUKm2hCVyHe9lYb
KRzk5VEs4HJrGFTdDh2vf4mRKosWfG6Wo21D82+s1MoHBiKF2tDzTGWx3oSiac9SQrl9XYFgyxPj
tciTAR6ZoBNv1AtFzQ36B7/MTwndavElh3HEPwr1J3N+w9xACaXSb/+tnrkJqZ7/bM+kk6rHuoRc
DY6UreWWP5zsUAIFsWjKMQfmQuF15i7CWcTalds0cn8zMmnRkzmameRfUJSMgpmvIVzRQWempBMy
9zPvyzcUAygkmkxOcpAu0draVZPtwLOH8iieOHhbUgQat0/8VaypWp6lpPMUbgRKz5f270pNdmrd
hNiYHQ5izAxpABiCJFE/qynezSqWx8PN0AoppT2en3cHia2rb93Gqfmmn70Q4PDdoRietLFDUzAF
p6M+NwrpyOQE7+gE8Ohng4DDGpRswdmYhrUp0APDlcTLjDX5Y6V45nran2yqHh6Bvn4QCWMpCqEH
GlBRHvr44QW7A4obtHD4x0W1RNhKnCtFc4BJ5mysAwgLshDyjOqpHG2HDIChHKV4Ed3jMNAC1YST
R2zrTy3G1psYyXsM8zwE6LCVdWqRLUYUvtXX4HsXqfbt3NzpvlLyc7Y5W0fGdeSzchuq1gVgkOkI
0xQAOkwH8Hv6B5UuOAXe2exGpH446u/xdQJGCnxmlElwroJ0hZLawl0WdJvo5IPt2KKsYnqUXA17
nYtQwAD6iDfVycZIPIM8NWLSw2NNJWl9Hdtd4BeUrozI1InolNwvbITQGdPYY1fFP59wgSOHIUAg
VMusp+xx+PBOO6z6r2g5Edp0nnTu1YYsR1oW0DJ7a/AYEEspcY/RRvNSTsikSWz24a/c8pn1JOJJ
AwqPNN9xOvCnV6kX3pR9kYjT+TomgvY4f8WQZN2CmEG8iq5Jv/nx1N+aOvi/5FNPjLTP4q7c75jH
N/AL3YvzNa6CTr5czdUQP7hN9b3JUJZeCJcHatS+f8tQVDxn14Z1Kbo/5LAyAIuGkmnM3LWY6aav
xwBPm3xsFay9eCtaaKZzERJC/X129jevA2my5xd8mqjf6/mcKZRa4ydtCuk+wU/yym4yQHutOgQU
prBTRMlAfsokdQg4lSjt8wbzYhU3IokV35IoID3YJvSuz+Ws6A52aCaOGToUif0TY9LmMc0DpD6w
o9VmkNaw9DZge+TaJ23MfjEUQYkbskTl+5bBBUzPmvLKlhTJsbFgLSKAjERkkijnlbeOtaGVJZ+x
PaFHliy0g+r3yAE4BfO//rjd0pIMxBzt3pvMUCcA4rzTst5qUpOnp4IxqJ7byULq0J74n/kWg3QX
fUoIvR8KljtZPyVSoC1u+FxuQuTEmolbDwemIaB8yDEuuyQvjIh90xbgzAtsNPEHGnZAynYp65Cz
9+5+TLfn04XgDejCO6UWlOKuXwr+uvXDEPNpM9QHQiQLuS4cO1J8ASbna3HY3ploxhFmC5P+Obhf
BO8ATFrZjQYMnKH0bPMplNkAabh2CAJkOMym4NZGNcuwwxyS0AD5A6UEBIWAth7qCPxyrtdzBa+T
F5l785J7ir2sT9ROSBhSVTq0rTcBitjOolH8X5JjK1nvVNa3KpUOvV08NI1VuhmELHoluCZJcJG0
2cI3o4YvfsyZmpwvHrKxK0K5Y1HuIBztY55YQ0YfGattRXAW2Fj+uPMoiyiSgnntdX/HZisn0Z0p
NOlzITK2+WBOGuSOALnuf8UkwtJcREgUCZ3iNrIepgqo5El/Pg7CG0P76q3y3Gh30w9ux494Fw67
ST/aAB6Qzbel4dI2e8NEUMyHqDTrbzoVu44+HsFYErxcH6ex/bTIgNjlVMEXPm4tc+ULgqYAn+na
hYcl0eHO/Ut9CHu81SkKfIWvfUW3IF6kILCZGIIWxBArsyElf1Xeu052jFXURVAp0IHutENB7E5z
HrLKI8yYE60JAo8xn30MmZNrKuQ1e91mzJtb0DuXVp9yqfdd1TIMtcwEsXXJFL6TNwneh7BNBnyd
8Tt1sjq9JJG0KBbCnqSO5PwA95TdvqvvrUDQDOhZT3gFy4UnJ+BSfEb3gW/ej0LhugYEoCXlmEgW
Dy3FHbDTdRjOuVc7Ap6yUJcVMv9dLKugls6MsC1QurVz7DLol0TI6fySzwt9OkuaaRitLtHoZJbH
vSrRrLCgABYgEIeujS/TgVs010PSvoEgvZjbdpZBacCPq+Q7RvRqnRna5+ZSc4Rz67eANxqLJzqj
glfACUjTIcyrgsbAA09L4RjHrcz3Nq24y35ngzN2em4l+1ayphqQhwfHsgM6x2AeRz+YBUrAMCvw
JfxOZNm7fgmQO5x3pt/M8jW7+i5d05uf385qazlGGwIn1L3wWD9hHDlwQFbirNoPkQheoXn6iY6w
bCgXVoMWPrZDaR+ckbx+Ct1+vleRlJl7PMUOSvaj2fzEjMx3UnRgF5zenbalSG37+y0/h4UFrx0A
S6bKw4tBAzj09jKXrQhOgIjmOBqeC4jAjJpTAgZM3qcw6wUMk9FSU3XFfV7yZ3SJa2RgBISt/jzL
jfVl8Qto6awuCzJRiHul1UzaGXZCaHUuIv5FmYcDwiS4qJA9sexDMGAwUOd5xCayW5FHgDNMSxsf
2r0qWNhORAEu2jA1xoYc6tyel4pC+XiVt8S2XvZvhNUEpJzATTjMsN7cAs9fwQ46je/ks9OqtrTH
b+AGFHcE3x3ZhJT9oFHWU2Ldws4cFdhPqAz+r+FeIywSmRWkY/3AMWRWNx2jWE4st3ZKlR7dJFh+
nsu2hoj968AAwD6PmtHL1J5xJKse9GwI8765vs0V80Fxb1yRIm1ZkGq7gs3E85xcXCOlJcTb//16
WhTr6NRrEY3Lx622kG9qoKsv21Npe48EtZS1LZywgAnEKjIyIpJcAJ0sKvjWGemIO69Ai1FQk3OA
paS6/MzTlTRWzqgNieHEHsUjaglwlaXDv2SX2DZ++0dcpeBf+LDADt6Q0vmzxTehDcOVruwcsSMA
S2Y/60YUAGnaL7BOIj23uj1NCCBs2sHKKMVvjue9T8zomWVJJH8brfbFkZygJr4/ULD4H+0RtxyZ
vUkd8OlrBpFtiOgbwxy38LIM+s2aExc59EJqW6GAS6Y03ZqCIB5qlM5pPVQ7jhQjdH3lzqipdtPH
xwm++rwG7GVPrleagjVd2u5tk4i2eVUmmeC75VPR+NNWsHKULYVq0w7wM6Sr7H0OBGmd/Nr4B0Dd
O11z0enKk1SrM4VN/F3eClO2nFp8pyS1MC633jeG6uM5sEWYpGyO3dPgl+XpQLcAYcBHeQMCarBW
bRN8fBX1FZ4UvLKId10/Ov1j+K03XG04aGP5slti8crorUR0PMg9zJLyYpswurEXguZBkKz+xIpi
EBWb1jP34ra6gGR4bBGIheMuuHWdX/+6UDkJctjzwesY6xvHj9kQjv8h8m7zbVGXPbmmIlq/bOUR
K3CkxIgp+m1TqrdRbqhji2hC67CSSladcQNpB8MkRMnKt6bsVymCkdHpXGf6bQQQNaG171CR3Vo2
tTl8kmG+i5ikJ49ji+5D4yCgRgbrbck0qecqXlFYVsCQr91X9j85mjoNVFt2JkOMpOA2qEV+Kfoo
fCjKjBy6LnOKkZieMDLWsQ7KQbx6A/15cx+0x3Bnx8SejvGAAK+8dLioPCikLHjJqDrKLasO4TR9
nZLITuoW+d5n4XausnmSoDgmzj6PBAnVVRJL4MyJoS62gFJDthWuWW6/t0LTs/PEXB11hDG6TgSv
TRByrjKPYDfr3a0bNnSqeW6BZn4ITONmt3yjsxH3NUDcbrLU6kHYn5XBt/9WhouEtE/TWlfXJ6By
DrlrQEbXEoXuiZRpS6nMAyGpeEfBBlRXgr/+Y5KYeJmPi9wULCtm07HK6VQUEQ7PkQCuEXY7R/T2
B+SaqNAOjs+oKqZVz2nJ5EydpvzlZaDdlNO9wT3nHtJ3eFmLY26Jqxs6GipEpZUvWEpcmCKLik4k
lTXmJm9/2KrLJWwB9Ev1Can/O6TT5qx2bJP35QAJrJ5SuTB9bDH6HERQHDoC9fpSlJ65hZ7M+MXF
E7h6ncMZ8la2ZvAqfNz3NkoBJjCYBssU57zSHk+G5qXOlvRU82YsoTGBjHIf++vZ8n/2EONtlH1h
vU34zedYVCkG3fmjvYTj8FPqVDWqZz+C/liNRRwHm3E/2LA/I+15O/xm9TI3TTibuxTKI5Hq5fmi
HeK2Z+Y0/Y8GOmJc/8KC1VZSVsME8nnzgMbwYcnNgfpwcERK9ZoLW2G8Hw+Og4zszTrW+exp4GyY
awdh7VzgOegr5cpbBXFsjqo9OkHkrkkb7uEhbrQT5N54bVQLTfhFFZfFQ6SH9hnfOS2nSMe/Djuc
jnrZiOxKfb46WR/z9eupZxTeS5xwV8YmeHeJMoP0ptV5u4F19j7G9ifSukovQX8tdOjQoD4W2Yip
+2cxloT6FE70m79dH7zacdV74MW5DtN2DBX63KF1AgElxflFdzyYJQv7Y0Bmo3DqxULxnfxGLPdj
ZDIkX0rkEoYsUp9jIyHTB/iEMtcwIqnhgkLEE3Z/h4QCqJ//N5f6QMndDt8yLUhrEUxonP9Fu7UN
Gb1a4RNrely+eId06d/PFj5c2QFK4OaV4DGraNLJ/jEmPg+Z0ETkCK2IGAkQGOYom4qKXIAlET9s
kLMQfcP/uQSegWhQ8QZjX1Maz1M7yAC5GZ+kp2QKBb6kJl4+jTz/FzytiCUrGHHywWTJPLoJY3a6
DMcc4vLb0k4irLKgYUehP4ICE28V686Mkl/mCt39HLsXgHPssmsmqnqnvLgBgpogWBEpLwQNxBjS
7ng6B/B7VnmoM+vvQYB02kXZ75Kx24XO52R33PyO1JfqGgRo1GOvFxrYDA527c9jle7HpX9qm3i2
Yw0h+Rk6XkD3dn304TYuzzHA32Asjq4L9u3z+ewyTE1AK2CODNQ59o1YxplqcVoyXEjTcWDapMEk
6iluf/BPP0+Me13teLqnYQpW1zLbiYxH3TpFaNqI/KSBIyb7/PQgFl6vtnYU9K3gUrRFDQQTfDUy
BxtIsLsL7tjrFKK7sN2fkrc9HvdZ5TeF33cCHNs5XFBUjEku7X916lT/Wcir+ZTJh3zKINmCUMtk
Cdj0LR7GDLRNIif93Wit26Zr70kLDRpvWPOt1nol4cJHLmYT4fZ0qKCqAkL43INRxq2xHAf5zXYN
JfIitml/phrECd7p7e9MpMaqaj5ZDuUVgwYVFMKxYp/B7JICqeH4B3CrnM9uZIOoEtlGljzJ0S7Q
XpQQU/Ue42hkYTmCRBOZ46NX/foGjOC7vZxthd9f6Q0loOr/9Up5BTrQjnVgkx61yhMh5GfA3iIP
VgiwanRHnVSLSaGelLitZrwLO52aPJl5kys2DZ3becWjNDLKUpgVPgA9HcbNDkmks3Px6jkHmojl
ydxGe77WyQe5tjmBw1j5HYXktq69rRjBjSianh9Mi+0tT07vqLAoo1f7zy8iFsB8T5nZ+e6331sk
Sm3tyigEgcRtSXl1dynMJt7A01UTFd/TZ0Ey7tDt4TeUYAV338HgkjbRtgWmQn3lwvQDLKtM+Mdn
uHRNbi4xO9bq8Eqzbchqi/Q+dlwERthOksiiqX0XItjP/Obk0c2n+y57UndTVkkQzg8vBS1iwDxe
2x0GYIUYG/QGoZlceP5BonDk+SJtObzxIP1OlvbBxWbK5ssiobONNQOXfsvJE6THN38cI/WqtoYs
UALptikfWVhb+WcESdN2KRmYGRBBO4WEj7rN3MlQwW3EmWJEbDwV6Mrq4k/EzkaxPQsNpwXI8qx6
EmVN5hrGV2a4RloMjJIW/rGN0xidD0z/3D8nE8nCFQDC97rljRYmXSaXiFkCpzm0mt7DzI9QwlYm
ZTRyJ9X3XbZpMXJlzCg3TzSIvnxjjGuWdYbODXIF8Drwpd9HFK35fEv2RpK12+Vj8b5JJh8Wc/FV
hArXYpPwcfUOyEuuMxb9l6VoZQYx5JHZuX8u+8nvyvB+hMWm2pPmXR6dBoe8ayrAYsraPDcXBmTG
HaiF8TYGRc073U111i8RitzgHbGhDnu7VeCB9gt9MW36V+Cdv9NosgmTpbMQEOx1RnLgf4pr2C5y
1XqfPK+GgGLrrxb0YvmrLMlfIoKe3ufLZeP9plbyAGZ+kQFRxMR76C7OG3M+tzi/ECJ9jE6br5aH
v2motBuI+60G5rrlOs4nSnEd0QGyxg2xNXlezUL9PyIEAWT70jUQJCGGabPeAGFrmjKsqr3c1Zlh
sd4FseSaJIFEWn9EWjq1Se9rK86/XTO3xBCI/Sc+V0FEHSNxT0DMy952gGrVxw/fWze2PJKG7Agm
tXlw1R0NLDRybB/TXNxGU3hcGr5bWhbwUK8Qa+VFiBVN+49OK1pTh2tGFUEuab31eNQzuYhBnfye
rw9C80l/UYT0WiYx6hZPO4kWAPIyE3P4JDlPM4Nzk+vJRHLg+fgCi0oIhqetheNojXMpHRxfgwp5
b6iPPqIopBiK7JmFpEbO0YqngCMbOX2XGmT/dd7VuGq/YFRT1NfuF7Qwj+dwCEQsdvcJXF8NLvxh
TfyYiBvgXFU9JYE7SmHho+w/1KDEpYb28LAxy/0i7yIs5l4dXB/E8fYKFI+PGYFkrMgSy92pOrwf
lErEb+Fm2RnmKP07R6Su33fkBW85LD5TTFdMHJu3yn3iBHNpt5qixqiMVTZfSJzxQnG2CGpa8EZ5
uJAH+K3j3PTP3b6oTrdZ5Vt+He4zDF7vk8hs37h7zPe2HPSE5ll6M7vkjsLC6hkHlbvn7PFhhjfz
1k5SNapbHo8wzjaJX7H68U3u+nYud3ZFJFLm1cxq5Xu/I7qIc5UmWLXdnZM7JmBGoutc6NzWQiZW
Pkt5N/koppgGeDJDgrOmpJ/wmYA6OtMk7UCUT4MvCS28gh9PxRcRr7JZfIQStzUM02RmPqRhe97v
bmGwtWskVRufqfhOxQJlu/4SMs1ElgaJwvOzmPn/M3Cie1drnsRmNEZOrHQgRE/yBeRtUUr2bJmv
Bsl+k1pB2DODwOy8grcF7LtLCN6QROg0agXObhtVoUA1nS27P7d+CpRDHLeirvndWyTHOla4AGwo
8n1JicP4XrcTiaaF6qV8XYAB0EGt/kkoLLGaq34ILURIkg0kw/V4bMhNu6PAQ4UYG0aguaNTXYGB
EMnFTeJ71++i3FNAJVD4KoJ1bSgO+pxfVqQJ2Cx51wWBBA2y2/MCxapifAbw8x6Jsabs7G7Za0ck
tuv3nIXERRGx5xpI8kK9daJ5l6FSsqU3hJwLG92ZJMZPa932O0kMbZe5gvaKVeLI/MMoc6RCIgPc
6FkNyI9nUeeNz71pJxon+8VxSPPTtmHpic9Atxv2+hUXSYrxBDKm+vqz/EzOXkNpginw07S0dVWg
7qC06aO96XietYRGtJl3f7NZQI4ESj0APzsqTExh63gP2GLX6y4ha9SrMYJqITWf02CKvBR/87oe
lbwBHBL2QRs9n56YauOJDsi8+21hpCev4tFy0iv4LNwofItv5jnlrDGok8MlGxZTZiLJoPe7iTeQ
d1HD+gT2HB03hA/usaXTOkmLsfe3tstRSCNVksHvF/cTHnOt0kYLyCi3iKhBJilNW3RfEh2iK6Ek
JkH/R2WdCHiglMGlLBFBllCLEqmwi79KvYQlF0DFi6XX2IMVLLW329ofHvxJ4rcLn3JLYxf7PCyM
PfCSgDfAxEBoDLOVeTxwpZ7G8qoMG6UpuVETG+UvTHoU5iBX+luKlyG45VCsce6uwce7BakKUkQn
jHC+ZikDY//kRlFwraT1Ex0Hvu/KwlWp+NTaF2R4k28fPHIR7kH52BgbeiuLvdXazDTofl1wJeMn
bTSjNNCBzeA1sRMPbXdDEkjnE0tIansicgwC6R5NY2np9oKizsGoUvxO5K4ticvlZrv4e1HGYXqm
4CXN99tCtwSNngYI8ZojzCDGwoFuXWz1MtEog2LPZY6MZm8otyPTI+q+cMSqj4TN3AYf+AMjYP+F
avoosamePNFwjJTOT2PWnSRqyVZZvsT0I5SPSOcm3VB4qlSZOedzUnBJREXqPc+hFVKuHWJmzcC/
zSrYXmV81G6HsGuzKwAb31qLVv7CiTYSn//PYC7EyMQT5BThT+cvmODqx9q1Twgz0OCnLEXIxf3Q
xWAaSIMDiQ/dH75S9RiA3byQyn2vj8kFYwsleByUJseLqgHox19HWm+wlQnPRsnP9MsNu+7dU0Zp
0M+S88fVsXgCQsFxVl/IE0srmvIFFcDa3UPk7mqikuV+7e8dXNyXd+MfkRegDVgPbaA2/qgRS91l
fWezkzqvfPOqacTCsuhIR44kFRs83FPRp+iYmqWAHYy8ApdHbocDnxmz/SDlTYVYWC1qSc6m52Qt
fU/tvKfpAc7vzifsCru0BZW7aYeDdLD5aVT/7CdnWIpr02YqkGVQeKs7JnYCa5VD9HwpdVwXOZq6
y0KWydU9TwLD5xsFyXbtPMNV4I36XtxmnDlK8ZW+IEjldYggriYlcsl4xyW+h0IFROy9ckWGzQOl
ynGASeeEUnfE6VKj0Nn4iix5+leI29+xeaGSMG2Mt7fnKDcUPVGdZ5JnY4CK/DZKNiwPvtspo3eU
xgjBS6YNiMrKtgz3GMitimToBSKSN/rKlnxkomqERHGgs7b6++nEuQkpwrDOncbbZ+YIxUi8imDm
5HLAptO++7svWY6zR9TGTbVK+wTvf72ebfVyU6hKxQpsREhG4siqJPorhFdd4CXL1IInUKAEYrHl
63IN7q1u4+nTyipwEFiaIdF8ONxF7xseQrKTWs1WYOWD9E2ncPYcOTUcQoLiqi052DAnFjMO6wt6
lCIzjMFsGRJ+Yq6ZeTOUwJUrDwz8M7qQMMQ2XJEQsCfo6cQKMD/hjrq+K/rvKqmUq7sP4/JbOCE4
JZhowK0a+HajGEwOIwykxEOMN4sSCK1m+TBGse3qHy33D+hM1IxQ3O0zLW4bJanWJsvyejOZAXmK
UqsD3zvNyDQqnZ67aMbOqA97Up39efC1jf0+Gx4UvaGURydsa+Q5me8lUHDJSwIu3mOJnJhpudCx
7c08YLV02oqcGPKIzMqyWdz0Cz3kZwz9S34qd6eSSgzazW9WpR+A25EPEMRZk92MsXTPcub6Rbjj
2eEgjXJqxXT/tRaHv5zYHLZ/V4q27JrgzeYJwdk3ERQu6a+ynsayOVPYfLwi1B0mGcLYg7ZcYuds
5k1fC2BJE1P8z+vj4ZfFlsHHxiQX+V7uyY+81QKVa7qDqsTty/JJdD7xA0Dyx9Gutu967VNzQ0EJ
kAyDTlDuWXhZ7vedOzYMTT+EibPc3ZHS2ek+UNv1yUGr8oBuNX3iZLjdPbC0uOCK30TWi2rQQ42c
9QV3MnpdlKFZ6r9yVZJwlcaQ2El0wr/5i/wKMPOUbH5n3maweTwI8pAcyumE+drOwt8hxFzE7cE7
C4zHBsN8UC7Z3YFRPDvZ7ZIv5RqvJf3vA2LEjpBfSYuBp/sTa4NRxzcFMgLDyM/8aszxPbQ2D7Dc
rQKyEajNt3jHSzCQS35cbfaERGeYjQR8rbU15EdTSkvueR+P6UKM4pwXK7IYCPjzmFMDJh3YfPNO
1O+Ui0ajzfOtEAmD6n54rdtzgdhgrcfvOephAwvAN7fCQXwr7i8DoE+noTmybJgeSh7Bxd6d/6vh
8VFCjS6q/XiCSOZY2rquEqhf7+DjJ1/xFraZjEIIaN6YTYa8hJFz37PL5+sArcju3E54ok7nGR5u
hkAGnWKJhkEGBUP7JWiDOo7kpAbxyrlSgnf1a8HWK4DbfTb/cmiBEJPf9Kz7hMK9LOSmzUQbcJXm
qOSiAcn8yG26Rkx6VA5ZO2POJTTXVS1KL5UfO5yJjbyaOqtQy+X4BbhUiyISA0P1EmhcqAATwhO3
it+jmiSfwrjTSwzL4sq9gPMivLKV0cjqFAYhj0ce2rIHoNLRzJZ9YO/hxSra14bA3D2Kv9BhmPiE
10MplJ7EiPl4aG/g15pHGYTpRqJcGaEOZEFPROpOODbgZfFwXQFMjJ/plIziSgtUVVMw4L7wgG0b
VfCbr04l0QrEDtFfq8Qb2c6uBzIbBU9y8t+f162bZxG4fXr/CoAvDGHQhdwCDtXskouQUGSilye2
sCY4jJ5q0avL+p+yfYfsWzvaTOB8g+P/u+P0jlWG3X3jMn5EJtcWckK9ypq9cQaCQKRLHxOSJJ7w
je/zhTzl9UnjvgbZnDAgtM7VzK6oNx+AZKPhPOLiB9680KLw4gN4+0yZRL8uGxg8IbM6rCzcqqUm
TyrTtMbMeW39yX7Mjg6I+3I3jQ2fUpHJbJOsuRw4jBysvyTyOoolHz4P8vHuD2iHOJuSojId53/s
zR7Tr7tLiUcRngeCkbApNYkuOZkVyxa8XK+BdUy8Bv1GAr+aG/5gwZpDM26H9WdfMb1x62hZ+JxP
VwJNH54SnimbMj6uSYIf1E0qNTqgpmG37Xgkgd6x8KPxFVQ4dOZ/M68P4vPNUkXbPiJE4kVbfwDW
c/F5xOslW88o1/a1crS8NubOH6I/WKJPuz1yxxweUXy9FFDKu6eAaFy31nPJ+yyRZmxLyi7vmpZW
m1nHRc9m6Z2m34R2Gksir/wA4xk5YzDkdgMHF2PoRQvjyXEoQd+2rJvSmKWThkODzqI4EU0BVv+D
XG97CBGF/60yQi3bEnia2G9/YUkrZ4s4uDMUM7YKv40nuWD1SXrDKSO/vUKb6KFYGGOQT/1u2rhl
C8xFZjyHDhL3L8Mz26N3jwjOszGjbKH9k9LIRnt914eJW/beTf/zK1S348/tuhM1ZoYVcxsY/JTx
TlusibNuYeHsKm7sZhIeIkowFyzFlzRCqI7mD466bzTF2FJR7UzBKzAJgMtY+M4bwPKUChfQu8Id
KwhlzQIbJ6JL5Jc27kWYuU3HeKiieXCcfkawUrZogzu+FJl5AHRZSCQRIcO1AhqLYd1kJ3pWHa0m
q0CVLE2rGtJ851uyi3kyFj9cMCkVVO+zW4UNW5bmDLtj7aOLB1tdlEBaPhzRqf6X/zQJMFBhKKN4
aMqVH3VhpPbL4vGqZvEQq7f2m8Q58GzmlfHTGdUX1jKWCr9KHNSdBa+oAps2KoInG+nu9XhqsNgg
mjf1lkunyxl6b6YPR2ZzGuItPh+0/cLjLJLi4CpqpTbVl68Jl3MlMqfCwYimzPn/Sg2BP44i+G1n
O8gW7FPeXZVGgN1Q6YVzndy4pep2qCj2r0Nx9VE64eAd6mXS7S9Qp1J0UTemna/ZAm6rMSOK8o9G
2Px7cUPsRHNiJiAvZ9NKlcFCzHwc3YbeiK6yNqTI2lHdFyGK0w9EDwKVRAREsWyNSQG322TRdMJs
Mtk24/QEA27DUq2mdMEtNliw8iUFkmrlYE/dgR7Tw0OA0RCasPYWBiPi5KJtnSvB5cWQ2kbunuhq
CHw+m0B5fy5k8FPxG6CjiKBJJ4INxhBSZnFz6oXn1xlIM+B371OxSnqdu0uJymNrvqnSOx09+0qg
A3SHyZAQJkKfa+3nS7gp9WfkZFR8BAVorjY5Uz008Vk5XAP5bOZO6530LhH00ZHGbl7nxW6stQo4
PnBWMZ3WcDuGmUSb0viqH6d4aV2Mhl+wP8ojMRZf1/g+dhjb4LxR+GrKIDTPhgAXSWDxppyj/fde
hga2LMkuAoaewtBDqkeRhqzK9RMX1goPLbxmGfxDi70mIgiswW/eFeeWvRpUC8aFDrEIUKqoEfM3
G5fgD7G4+1iTZiG7ier6ph2qhV9EL7hlKoz4OE4TCipEcnh5af5CKEmtmWO+PaxsloXhzkjcSqeL
+nm0oH4m97Jdt+sA+Dy5drzETofpfryuQqWgy9VjYJBpEyoZqrTO2zHT3fD3d+M7khnRyjwZYS65
TZSyiQLiZ4HH7eJARUgPrJ2s/F7iKG//vJ6jLpAaszeuzYafOQMg8+JW16pX9uojsSPbvSjA9XTy
EZaIoVsTmIXmvsk8O8FI4pTH9+Q5/jYQwL86FKFun+/fU9149TMQrPNGX/o9sJlB0z+78n5Tulpl
ZYin/FvjtikZIpZ5vUWKOhp1aUBjxO+lTc1ErAaFGITq7CC+Vm5C/br/ybkDMzjFYJEY5NoPfTDw
uuyszfvd23FqtsS10D0T62Ob8YfdDsGr5b+WZCIObWcUt4trdnrEKOZfTe/MHIb0mv32io/Sb3T7
yQ161Fkl+O1WO5oYGpARLUvRLdCOMO2rwUv8WiJYhckul1bPtTZ/fipNR7a8GDHv04Q10cCF7DH7
eVzLJd2LNQBDhgw0o87RWd0TOtQaQ7gr/n5IxEM0M77gd8Q5EaXCG+GTtn5r4/fNyX9KJapER3ra
P5msfIrLXhygnD0gYhw90XdsHb+JK+KFhb6zgflYuqMPRDewDrBQUlY9zpE9aW+tPto+qMMCEXYG
zcLSGEvgKrJ333Pi6isXiDsQPga9gGVZqnq285jGDZFqNjUep3BzqXN0dE7dAZdBqr71J712AQSB
fGTvidL9Ph/75y+4/54WkX1kj45uSnBYXrOvhyAUzvVJ+QsBhSeWsvn7GFDb8j49ves8BMzVZZhE
phVEvTcJmrtST0wBtDLTizBQxVYWM9ZxC4S+7JxEhbLG/oMfokzNhyb9/JcJ5KLUrpxIbAeZnG6L
o1oNlvAPLmumAENaD0usBaqHtCBND7g/zzPl1PdPVUq+gL/YHlB5Lo8Eim9mAm5irSl/0qIDKZDy
bRS0Tifv/pOLrc0++aIjCXUkEKqVtvqoDZb1bl01ihDvlN65JPW17vMZhJz8o47SGLLm3AIjFr26
jC1s7xT2ctvdrsQvfRWzaTuM3xPmai5zizxcRsOwm/LbYI32zom1znWDKPrGWq/Zp7Bk/mFlnBh1
EUc7EFCS3n8C0fLdIqih/xWBaoU86rbtAG7qSbfE0glZbZLR4Ek9wTnJRSapUrECIvByTJQK8ASe
p5sU2Il/NPtq0dZtB9asHRkairNjXOuAcnPHN+wGyZJpVSY5ckmiLQDklj9nuZummyj08RSJoviZ
dRISoZ3ClXASzL5Px4JMrU8Wh3l2ExTX6kjFnaQv+w1CfDiWugxJ1jl3DwOOm9dLGmAYNninFQUS
7px8kPLXRnDTJ8CUNwgr5qeVHKwbZhARM2WL3joBpQ1uA44WV0PhgtmTPzJSADy0fcMNKLIGB0Lb
YP4DRxAP7QZWNXysZpxA1Q0h5hDBGlZ6nfFuhAAxSWjBUvHv/0slFwZlNcmd9wliIpnqRrA0MwMk
W2fxiBbvO/uhglUeOxrUprTkuiKa8VybeRJPrh22KWRW6uWXmDmVsKPqomcuNqNNfIqbFnoq5C+I
3/lT52tCHQ9KdLYxyMLS1gMX17jwerIP1gYPM3y7ZXK6dRhEIdr1FpbPdFtGS+E+Nk2gBSqBy+v0
jlKt9C+CmRnkF3shQymCzkFgmprjsPyvsXVe/xIc5Wne0ILNZFgCA/okCh7tknXpbVLh/IshyZTV
kxJ70+lObN1BuwC+4Q1Q8e76o9siqkSovFBYKC1Pw23mJFtH7zVsdcTrjM83TZs52otYStPV1cB5
7USuQSBWIJfWdJOmb22NLNUgSdq0kLKQ7wroUk/RTLLstZbXc3m1JI44GVdSSWlAe2zDvoW34mYQ
P0kVghChZEsA7pQa2lDi15P1aIzyrPg7SCNwe7yUVtUgzcuErxAEiXHojo6esvXz37dStaR7hFzy
Oqw2seHkyAzljm7MJJ5ZXgHqM7r1n+BzsSudJxibYuzscRphSYDEwcUN1dNgmIXV/zIwSuWjttpW
5QTgmEmC2togQCaU0T9vsrMp+MAXWJ5CBWHLkb3IUvsSJ7B4l17bWvixD75i+gXpPwbWmBXHC5Cd
uBwwR1wMRGffGn9So+6PPnr62l2VLLwRMoryWMexsafZAPH3y2pZxfw29F5b/3zqdcQX2Tch1Bet
X/4unYBsBDJ5B5oRvNXHkQ1Ytx6jaMUcBxCicyVbv3bqSEgLL+5IebB01WKuJgwzIwolurI8WmnZ
ifWjXonrZo5Mimp89xgL9z488AqbdR/LeO1pWylUMW3rwt2l8lIPSCMGZ5NNpGl8Gs3dlG66xdHs
uFhe1dJf8YkCoqq9YZnxJDDXKyxVwHdS9MDquAeaQr54/KmM+1eBZhXpS9FsW1e74kaXIR6f/WcB
ldHyUKD5XmvuCK3h3wu0thEvu5ltHoQU4Qc5CzZSks9xyOGgKWepFqZqIzQMPASEssTj9Bjjl+pu
yddsVzXVQv97uNY8WTh4+0BNgyPjHdNkW7tRem0Va8N0aF/MB2klusra12825PhIsuVlM4W2gFOF
5EHAehJD3/Ggv9Crs1Tln4/736F/YBeOMfuhUsQsZDOuGrNBnKAtBMotiVu89HenT3E4cdQXraqL
9FaSMkbHxceXsqTC7Gqcg4vpY4/i7YC/jCSaWRau80LGAwYvUqeZGM3mCFDNCcLz0zfxVvJFje6C
Q0NML75ksR6hj207W9FuIBA5lgSizOcvZP+rQGL9U5NAUFfX93bCSNSwTA6Pd8ZM0UmqX2BPVRs/
Zw+MNkGrrivGw/M/jbhmCk9tBfhLEinoUEha+euytRBpwBmPZfNCdrwJZvEekP3SBahlBKsvnzav
cLAGFyDw0j9orikKMSo7V9pEGdG/iHo2TRsWU7snaXn6XGsRd0ixXuRcJ4asRbtoPhWutAD/vNWA
V7BPzQlY51xEa5ehOX0TTZTPeywAWjuTQDJZFmtrZymNWpI7f/HvY7RVPD5NxyyH2p9jeUkDEu6Z
7KyxJTj3tjlbS4zx1BuAUKyN6yisTNvQymfPVRXgehqQmeM6LB6rt5BEtua92Qv2SeDjVYTNW4lA
Z05P6Z3WlXlf4lhb9ZNOokuCeieDzIKSDthLUXxe/kvGqyLMHpKFNBld9iZJEudjxP30g3poO1Z0
5i+UyQLivpINMjfw3IX4cP9pzgHB/cXSCoZCHTwVBpvJRvdlRBVT/+DskB3h7Etaa/TxpY0lMbpQ
0x0eqX3OLrE1Azbxr7uGwdFJ6P8/zyxlth2nKIZNuvq74jYnwr2hYNUSRDKliQd6CWwUk0AzkKk9
mt2wpZp8Igkdx8nK1CtLkdiGX6XdBkHlhwA83VFCfg/6TND72bLJED4jA9aJXZStyTZYbEh19EoZ
eDj7S1tNehmlOcZnH7vlp6Ubf409O6KOrtzASKJ8MqVVV/iZlWT0mC7hFnqtYxT/FYVH+wqCW5os
yCQFaKkF5DZyAvXZtk4CX3kYHwt6UTt1f9BvGTohql9NhwqtZduhFnsYlLviMtNDB76oqv0SybUG
NgzlrL8LV26VoumdHVzfXDRoWajbClddHi9Iqebyrzz49OKmV1XbvUodO8MFtvdcvTdOZFr/orb5
qd3eZkTMJ70xvi41nhgacpH+h+EG5kkRuTB3bv4+LXa/ImV6zFmb3s/sBGOtn/0WGK3XXjS6P4Oj
VgTyPufXXjxex4ZsBNLzX977dpM6YK5vmaBoTgnJI79fywc3go2uBwmGBaZlUeYf7TuxEyUJHLzX
dJdaiGII94WRxNkc/anbX7auIfFwbaPcMvD7IV7FhlYAY6+7IOGiqjQZIYxXK/STZTEGu60eX2f5
dsRbYdwX0HbWwZ6yU2rdV0bIBzUa0Feu4NLFJsr5v4k7SXZs59GChrPHFFK3Tf4ocSL6w6v54oA7
TGhzam91CQB6KHX/0RjsNMVdJQeIM8rjkSWZjhjAhA0MpoNDcTdGfMQaLzPcoA6yEprbiB8sZEjD
H1SJGAulOfsmQnkE13eL84kBKP0O8EYx6gumZumKjRp01t5Lflzy24O5Mn/UvH5gpiPbzz5BH41B
+SLEou9ZQFO2armBr1Ii/QNqzq6UO63ZJv016COJMvgqqPs7Pn26PZ/oTHP4kvmZdxe3dyvhgRtP
igcqXosi+tt2HnwCaqc7CxzJTP+dUyArxFVfyiZCbA4yDyTt4F+tORvw1F3fkuqSZyeLy57hIXat
pG/cuJ/HaopCJ77QUS8jdSsq8+v3culn5v8Y28RzBP49zZBoVLSwDW2oMLDLKDJt2B80cNjRPxXW
dXIXCWfwVzm3gfw/RExzYpRMB0qvPdp8gPpHxwG3bwjSw1mHOgl9GAPf3SR9L+KrcexYnO62Svwr
MoNU/zoEgWATj5mRs4+2hJ+UyclHuYzW6bHm9EtCXzXOKqfAOPY6CntjKsjlzW66wDrtyFq8HKZP
Em+y5Y7g4UwDzSlUD0v0PuPnipZ7hXZ61ggZP9UfcaWPKI104MJe5bl9DuKav+nK183ZK90z/hqL
zw17kkyXKmpwpWjYAeTy+BorvaKJ95EHeBlOM9Ny/aRd1zRV8RivOdjTt8YKQY3tgrJkPP7eRnYp
tDGXofBLSkkhaWeviwG+jAit3MtHes/oEpn2mNnAWppHtplF8dNGfn8Qv+2zrFZwILxU+iQws0a3
sYmDAjbHEpS3kQBlEckLyoYdP9mPgqipflMrfmP0/bTsaSxC/B0l+Gl5lxWdnlCxxjbVaEPwP9WQ
1Ao/JiAXTX6GajOTePQzsuRxdKNs982gBj6gdcLJtw8Kzf8TEjIdRXRxkpE5fc0VsL+tFoY+qhFa
nXJ4V7D3tx5PYPb68O4JRJEzxfx8eIbmMO0ObpSAG9PKxGQ+Gdv8SdwTyEhhAAzIXG8tTu3CyK0s
eUZ4f9IA3ZDQXSR4KiHRj+rwtIiIv30g7LRwQzklf835v4VG/WhGelQAWe0lP9GkhDHZ6phUyY2Y
HoIehrfENyk2JhTffSIWkVPIK7kxIc4or2rhJKexvG7hCWNjmeY9U7190hukYb/C+ai0CV//PKFg
Bm+cuyR+/TU/Ok0uxURwz4Mb+5Fh5pBDUJcMUHgvS2ES3gL/8syRQf9vjIKZYFs3oaU4jfKpYXVZ
SqtlVzzZzWUtZuNsQo1oE6Q45EP1yNJMoZbu8eAv3mhlETMsWQKxQSSt1rYzKjfAQttvGVO+ODYW
f4iwv8hWAWOjbvsjo2MFcY/gdjho41M4gBzKEoqgGzp8Gml7J/qMow8JBfQdHf9rsq773uH9uBRZ
25LRjt4bDvg/kz6QeOGc3v5gZtcsWGl5wwNhHDAjr9GrCXOUQ2cMGvwW/FP82kQurDAe6PVSX5Pw
B2f5PVyS6NynseW0WrJBTkDpxo/g8VxWVLxZOGr7Ln3Hzpanwvorf9mVA3q4IqCZ/fMqgsWDshci
0cVxly1MXdOwMvR/otT6MS0rEfy4GHtBhonwV3h9l8iWNz2VsxjPmKOb7HWHoJ+1n1Qf3MvmfNrp
ypIXSBRd3WMCDewLKOv56Lq7o4lGOB2r0yObM969M8QPFmdgBGFd6XWB8O175J+KimNWC4KJNtrq
hM6NYwhsZWeg2an1SptnGYKvCerKErjRAo82qscYGMAgKF+wj3PmDrr/+0BYKWN0GtEOMiQp2Kjy
kJETITXucN5PYdEJR70TJg7XoncktLtq4ktVjjK80NKdhsO5O4SR6iyCa2hFfBzMGHc4D30+owjd
Dp8GAldEJTaCLhZSr49GeXLQACv48IEpM9ojWbj1feug7/+6vn49Tkf3v5AgV6JVb4H5QOkF+VzC
8Gr5zRXYQKwK2e8rVyXXgqv43hG+3laDlmONHEq1u5TtB7JVndMhVQu/3wNk1F2VCHieeY8QitIf
vQCCCAogL2JDy9c7B5UcH1Xxv6fpToPcU204aQm7LUv6FuycK8a8ajrBLJ8M61cjXD8iAwMscK6R
GegpbUY6zdaOrVdDU7ozXN+td7qX8H+riuhiPEBKlsPGYlfzVdaPi4oGgeEYwlIHJbr/Ysjo8TNd
F9SCXOZ2HoVYyd0pgDzgWuR/NNPxWUEmCL9zWDDg28ECqqv6KVXMMuK/l72ZfzM820qX5oZC53j8
pSpt5SD7xBdGFQpQLZsLFB0U12BRpU3kXBTxai+Y7aOP2szojNq3v44s9RGhv7254SonpfoKhI+K
bUeBEXMrtGhMpm1ahobcxGx22fiCJIo40vsN8SS7nwHvZgXTfxhwmgMsielIbd+U+0EUc9oVhHZd
IOTkHidum27LEH86ZStL5Zm/bPJCtmNpoSB9PN2DJid5oCtQRiqm1P+NG9bukjCgiA59QpUWHgwx
iCscVy6H1wbHq2xmFmABlfrxK8P97/DT8E9VCauGaSH2u6iP962g73xlnXEa3gEWeuecUVBKNng9
DL443iq5dpW9eeh8GL8AIYVPZ4ipWT2lk/9BZxTDVG8citmVR11gj7u+LkVaXnOksOvZ7hDcB05L
KCGz1AfqAzSg6vHmk8ZidL6WkrROo779SZ/nY03oRM2gxSw4pBN7usc0w35saa99+lX64YjUF7Nq
YYonqrnEDaYCESvV1ze4vyQTKNb4Pc0/jGYTVMpZHaY8fwtOGh6GZQEVrOyDr4UVII5l1CZLzBgq
NhzY+J0EcFBqZCBE/0vCME+tC2JPjy2qBTRu3FUb4AbwZlKt2ssx/jbAd1mM45/7XsT6j18992Rp
MvdQuqVPjOE4ZpJP5Gy3VIAOBMGZBWJT8q86OiEMcm9ezgj/41MiLnHM0eWPNceNEAYivLB9d2OB
UnJ63trn3VMSkeHHgTnS9JC1/0nKe8+dT7+bGDZX6RPQyjJkbvwQpq4py8+A/7OLi1/CQ7WYTSQU
+iwy5FB8JmlOjwM9F/Lb2sZITkd/3PfKB/2uQH/LN5bHmqKzW4rtPFF/NrpOMssd8wW6GIxJ1n/w
smsb4+SeGKymmL4BuZ4213wWs0UFA2w7/JHxqAotL9PNyhu2wOQ3ONio37DqmcZnUVq90Kvwd76s
YxDuDi/wVVRBqLf0W1+oQ13ucwwY1hSwx2Rg4NPsOsGtkdjGD62xadbOTdSNrRw5Q6UyHVGE8NvH
z4FqKiy3Ct9SvrQnUPW42fnTWMQND4v5Lp2i5sj/RO240pTaa9IRoNR4vY/HFDVl9W0y0VXtv8sy
ZcsQYlf55I65TVJu4TmYZ3+ZRKyQob3QEKeMi1pYkCuWDa+hfpvtnOpsrz0WPOz0mhxSalIzO46Y
F+3fONps+TClDy4Mx8dl1GRIGRunw1MjT2j/J1rbLiP6eiumvRFi9hQ4/++GiR2aSbOJD4rDGseT
ip7WYGwyaa9w2bn5JJQNJNoel1P0uVM5W2lmNmMfY3+JLRMSsNdieovTqvYqetNBIRjT5CKvdA1g
PHnRHSHxNTFZGJIkFhfITiLzm54VwpZDTsjh2plGg8hRiHcHtFn/KVCKy0uSdpFjG8oXZ/PnakAf
+ME0/1kWGGt+NO551+Y3C8UI96egLLwXqb4QpEuMDtDRepuDIWBWEwgBvEu8j37f59sZ4WyWwWbS
1+Ep8omwm0qaCnqugVSPxCEI3/WsPODRztEhrVaGlSmD+LYOXb6VQ5ExXRFrrQ/qVumcQxEpyjYo
StZM5COYSW9iwynuzLqSG0fEIDvFbmUInqZovY35p4qLHZr26CxdGBJhjKdTNfwtSwFbiqLeqeWX
QE+HsOLBQF+hIYskuKwkmPMyp1q0dbcXIj8+mACqkAfp8RovvxMlsVTpB9/nPAzWfCesMkasXcyO
qrNKAKaDaZ7V0GKhf+IKcYBcUcjJ6HENv1Iy+6vFxM+14h4s0hE0LrqCg8dButcfj8xAEGK/2FQy
ZIKr9CsiVh2umc3DDIyu96EzDBPJZx+XQ+TvIGWtd3tCxZGqFeBuWfljpj1vVsVqD0Bv1/0mN51L
RK8bbAmq802H1pWfClG6+XFPVKU8BEpTJLHwCkwVyRrW+6q899WlMlaC+ztzQYdL+pKiyuxFFdeg
4boLuWLGsn5/h3A9dxU6N1y+6KGhUskrFViiB2JPMKDD219ygbmuckwyftKN9F3j+m03sGVUt3bD
u/vW7YKH55JSXYxv64XvyFLZlGTMZYK3dkw0ilaEUDhFE+FILeQ7sfDQH86N/O2tY53Zs+ARYKa5
+RDBwjkNyWrrdtFWu9/HbrRFmHnud+l+j9WqAQzcteNH6+pyOG0tytliz9IabT6bf6zF1XUsH0qH
HCtJw8IJ75QsdyY+PMF+BD/57MuIQlZcDrRgWMKDL+ArMxflna8+1oS6LNAUCkhRXvfqcdT21z8h
uhLom8pym7G+P7FlOK4pcmJed4QCqApjIW2SfZ52fZom5ErKUhr958a19g/pft21nwlyELvdMWtN
fim0OfYwzPlB409+ZBoNjQNcfVd7Q6fGdVwBMBsxW0GpOP1dJjcsRkQ2itMQr8qaigRWkdbugXPO
eS3dE8h3uuoku3VKV9XpKmF5aUE8SwIazqbVBF2+nDF/zK5Bj6lBClau42HGDC9A2CRX5+1xE9VY
1EBvUjW9u0YjF3OrE+k+u6C+ZK31G7Z3leDMfsnbh7oKmF2pUfmZ2YsdJB7lExI4mmmMz5MhLMAS
cjYeph9LRCiNih20/oyDVDNOeyCUjQF8NVkqCWuMR/TyAxrgyj0p6sX58J5XbNyr8WPdCz77LNqR
U6uzBz7HSj8nW2d5xTHzEdh8lEIp1Y/3/5fRhRcAyvNJhtCjuy9GtdnPJBLPNMhgJFEpKW7NMKZv
yQHNImqEwZcFJ7pMBRtw/c3O8h58na0Vwfq7WkaiQ/pBa+48cYZ0K/xk/hmHfKdcVG2oAUabMGrr
RtuYs3266t1u5mGpw+Qjg/MZ0HO2O8CNV4wwgjhXBERzJUcyI/XH4YJgzsw0ULoMi8G5jedbE8hJ
zIKJBIrB+Pk0mNnPMq0fjy6fM6Yjwkzbio/KxTKK2HYONUCbHUeUza8k1xUC52DHpZA8xyiSQx8x
VSVNOj1WMu4xeIATLJ78t2dftJelr1XXIIsqSm89c8xuGAoNkFHfJ4VojR3leXjHZVVMmBJXNopr
+SgalEeohmpAzVYPuclgFJZ4bVmYVYuAoro0p5bnqosLGzQtgGkUsYdcbSJx8PgUHa/BlATBvjdz
Qml8YFUMRAENnusn0uzdcsGCfdFHoPbIWtcZCkYqoPen5ERbsvOloCkhkV/Qg7LFW/T6EyJZlS/m
vmehLZ2Qsx1gEGiFb/wggem1ajMnFtXu5B+8rglihQe4PpeK7fpVoJNRr7YNO7NOgjPhDzoOM8oi
8uiQbe0DER9K1ZXff2nI/c2Q/O7o0suhx6CTj4NppaG0zVg7Y22WHXlq/QywrcAVUn+4u/HjuYM7
t/YNNnGUNsfzJ+4WrAXBd4U3BQwa6n/jtjXRCWTFx1DUnL+Xc+2Os5yP0/ruVjnk0PrCeXztZ9IB
G+/LL8FjMlVlvMxUSV0sCVYiFfAjDjp0qW+Rkn7qOdjg9tZ+ZaeT7RhkqHeMgpZCfPZ/2E/88MQ6
x5mXfllOUm8vYGBuE/rhY0U8hsln0mZ+rLTl8+HpHtuKgqJiofzjLXJgQTHHMzDSoO8fS2iGgGyk
28F6SOmj9uWnqix7f+Krz5gX8b1WGa1C0YIbCS5daE9yJoQzSxK2lTU7SeuoDj59Lisqi72R6a25
U6/GL5ORNIQIeCNp50NQpCHTE11cnTzepBKo4dR462a36JaAsNp8FJmmEeCxJghyOPib1jmJdOsg
admvnKa1k7HIEkDfby7Nwp3aBOFnMDvFvO6XiNpxutqXJgDoaWb6GEoXi5X4fdUhcSXyyF/i8+lY
vyA6SYBRE3POKCfq0UTZodGpTrTP0Vrd4RlXG1eYHhEDPNNik+gHBynyYgV0tMZ0N+Ihh/NWGlaG
qTobtDuZKDmF1vMf6mH7VhV2DzcD3bIhIasyaa6TaJEGbZCt3nGr2JfCnG812Ib7C9e3l6gW4JMB
rXQIiwvo5i/6ciA2TTCKTmCK/GG2B3X4cOZepjw+UudPHv7oFJisn9vTuwrt6u+1dMPk4ASrl6s4
aJM/xyYawTFEEhUcGdJuS7865Vl9wRUrdAUJtxAVYyZ6UlyUNidZMpcdgxxJCJrIjW8mYBpqFakt
X69t/s1I+UvuA1TGzmRQYY1dmB5Vx3clpRddoy070tNgY3UQ/ivIuH+YxaRy4FuZhStZ6gFzZGeQ
uq0qACGG75jDy0gMFW0YsHlW82Ioled7d/Cv5mcnqzStnTcKFsNmdxPmZz2tt4qI5di869xObWF4
3aY4N3MPay6lsAP8LiBEFwTG3pC7BS5WycLH6D9GjVnBLqEEwHMs4HNmCR8LRG7EEL4r/6QBhQQ1
g3J/Wcx9uOdCQ1jX7hPGTwiDnbmsmI1XGvwYdCsJ2vhzqX5aj5S/KO3eJF05OoCCuuqMMZ09cCFj
UUG0rmd5quE+pGOScSPc0vqBLYh92LCj5l3rmXbgWg55GUVRuCxWg9Mwnbhn9ukQjyFZ8ROgYkI7
V68FF+1ynsJYHHk6aO/W9h/hCCPGsAcaNpqW1MFcGwtgbbo/cPso9mjAVBdiVH7I3wexJB2tcRTk
URC13jbT2tWNGPzkzwwlhQB368+XYKwdsT4SjjSd6zqLs/5A3pzjgTfoyOzMp3Z/FfNLsKB2g9Mx
P9TwtSxu3gFhAkZvlom+YLyck434AfKkonV0rR040PIrvwQdpHZnt1ToJUCWAmZwBJmv839ZDrTl
5qRMdG7SWkot80hfLdS+K2HMQjqWO8NXjOHcIM4AiGPy/pWJWJ7L4FmL88CKsqVc7kqhXdferITk
rPSti3utyCrIBcCbDSvfYYPvRdstqTOY33LhxoltFq29ufnFTP27uohZd/5m8PfdTUJ9aOF3cZnZ
jY5WlRtxVX8AnpZWmyTLFffmZSrjwDxmKu0urOHvE+QbNLeRNRBdI4oUaf3H4Vd2uIMweO9pEDGg
e1GC1QhmAFDr/m36GA6avDsjRl8Axqye4o/StXB9FOwoNdjlElqio+ZoUojBBqE7EMW39wOM04gS
Yp3us6L53ganzl1LVeevpvOwedRIHRN1LAQatwiSFQLpSRz6MizPyIkXgSYZXWtnAly1ObshphP6
rnYJFyrTCu+ZCh7GO6g011c8o6pnkw7ggYXq9N5JxUNgXr7aOJ81UgwTFiv55AbkFuCesOpAVhzV
4XihFjjOLEw4yCJ62QXpBFE0B+hc8oRiD8PDQHQL1lpFxvRj0DleoKQ0TGw+0IeLE9srqJRWkW42
1MRH1b2PPrTleRD7//flxvs5vxpMoenbal+PDg5hHMxAKIWP60SXlRk8SwrnvpUNL59GneJ545OP
YfxMYHLVoXgHwB8ysvEUJLqGSbP1ih/rKRGZO0S4IfGv7cMxGAgyll/v0o9in99R5qxlBdnO2XSw
ybRndqgXGIp02DOa7tglLReC5nIg4M16qabO8cswlVQwh9dnm6oybX4khrhBYHjFtp4A4Ft2Qwdh
+NxPYyczIVEtmP2nndsFznIv++2vR9ArmMUIPQlX9cEYHsG1uQwrhr0rzYxSOsf+Y8ruWyMimnAJ
yjWGx3kBkEVILNOA17AHNcMIADQD8Lo/vg9c2XzqooMuy20yg+QnXrHCm8LKFRoW5eYgzDjM6mHo
RF+6VwKL5n+w4Mx1Q8ozq5wg02u6QAMKhgfuQ/lSjhJ/oVUD54Zc5BlzpDspA6x1MItC6yZrAIYC
8JHql7vYlsXQe2RfJnvSi7wuV9p+KOIeYci0rtXFkdSnJRQ/OE4N67Llq453tSBDqJFPky7Gvj+Q
InImzOFsC4w0vmGBzi4UzWhUwkXx9huUFlFyryoae6cJ1gg7CN2Adv32qtv5dn2PRMeDKL2Rp09w
G6xXEOJqny87dAyo4TCT7F/ifi5MoxfH7JwXXImofVy6nMxnX7mLoWFOjF1hBgJL9sAMaj8EUIaa
hKw4UeS/VNNyFr9HRnk2oxfeSfKbGgVX5EuMcjhnJaPWosU26f993HQwz29bPo0T70qllFDzarcZ
cWzsS9xZUj155FVTzwWo9t/OoHZWCgOf9h6BI3TQKNl8EE4Opl619ir0IMcr17Fkz1T6299n1wyG
54pxY3gtSV/UKdBQbt6QXE4aSfONtiRPqV3FBR8ZiJdmQgQbRhgJ/MW9Vr90MVueE84vadGGMxOa
4NhKYGBi+xmFv48YXhkC6zUymO1rD+Lwbet+bp8NgcW3cFZpWql/CD6FYs/suddspBJCCkvtv9eP
hGd5Lr25oBqzI6wOWAhoTibiKvL6mnzc/SfQjwXZKi0Qgt0nvJBbIrJjlibXANuXOc/CZ2rnZT9K
CKTbzNNzcmRtR1RUkMlkt3nCHuMwCnNtekUXVLAP3GygHN2kemzr0nYcKiKmEk0xAKKlOOVv7VgV
sB1QH/M/WqJt682Xt/Oy3noSFNpCGOyg0u76E1yPfBw1PW/b0cThkvEgNSZLNRs4kQWn0dSPfax5
CwI3iwI4qOvIHbkpRDiAuyfo4yDGhzSQAI+E/5GjBKggJqAhWzHEuHI/Vvjx5GR/9bFwQvn8d5lp
iHYgDaPJwQDkf0+HENVNbKpp/jhV0+zl6ww/ZSoL9G6ZNGcwAJROyoZzyxpy1EfZy2Lc0tDt8Zq2
BJCo6DgtQBAkExJwKB4Brbg2ygFAZ9zpHxX0aO3kydLj0UNIsiqX7ky9Z6wURJsFtCka8dy3A27e
Vt27blPfGXnyrkINwahOyGh2V29TnpPS51mCwU29PJPBkNtqRHlb0ORrHSZpuzOuIIFvVm34ATts
OTeOtClMMudRPi4FA/R/v7yr1zV3qKowlcWQJBY7vilut4blwA3T++FncXoNtJ6UBaK3MO1E0XZD
IAS6iVAzHssTVM2ByUr3Pv3f4zoxoWGsdnXONr4Td3qIebEKhscKyf6MTkn4uIj8orcBR40AQ2qk
J1nH1Oc49CaljUMFSiV7FGor04HYuol+l8GzJCl3OffPuf1Px55PFzgm3vzJCtWVCHHuHdYCRAfa
c9MENOb27AF4qikRGvQaGRdrxU3nH0sSEBJxbgk7UJP1wwdtCLfwwhF6+IZpYGEkeLyRE1m6aNSC
gsMSRTsJUU41AT1sIOhxzMJGCAsdRHuS3gMSM8Pige4oy8WqLAqzdRHng5PLhN+Rf+vBaDDJJkLn
Koxi/xI+8NC9thJZDilYGomiwf1talADg9CzLF5XsPR+pRpnH4rGu2gwgd///RTrF4cyVg3BPoRC
l0JnS8/LpjZPyIrTsI311XRMRvcBZoaTO4hzXvHB8vbcMoexCemRyzFbVuW/Y3AekYWbuXlLHUG3
wAfQ6OjXVkM7NdlH9EBhZfgEyOVtx0RvyWg9ixcTAKb50Wl0FnXtl+RPfMYLXV1Rjy18P8ehwc8H
0ptYYOhAiPyA9PFVSNdNgCS4d45+dhzX36ZVq7yePCgYew34EpelDZw5qpwzzZSKnT727fbpjwqO
79/OvvO5QZVe0nZ729tuudhjmqTw9n5V+nhsY5UoOAhthk8cJdRi2kpoyMqRpgr5R0SkfNFbZyI2
7AkQ2YjCW2zgQJ+nBLdv5XeSKiEq5+NlUCOeeBV6obzDM2IM4u5Ktc6JsrqAoTRwwQIner4xxHlA
0L5sAlbNeduOfZ26vj09W5EbB6IfdE0VmGNNFkPofROzW+U4D/kEuZEVkMCBgrMPHKZM/OJHvLSR
/VXIrplY3sVFLmipYfuexBNrELwHu/40nTDSdcP+c5Q9LIR/wup72pS5NGD1s37+SGXY0I/4VOMM
/z4BlJioWiKFIEEVNyJrOULzSPIe4IPxYdsUewdjON+ALoVM++ZO+sN5UlwcFeDTRj9syByTcOzh
aevpCvwdeBNuX0AN++GXRnR+Cngbw68oDf61mbZ/XZTHWEQ5qn9ZnnKXX19pVzfXbudcvf6qBilE
6D70xHLgWlVCqXQNAxbLmWXtSWOCjI3IUwCVbGuLk8ZvzcFGkQszjMq/mceE3KZxIDr3nJU8dVWA
s3wrfhxrdf/y9Bnz4ixM6lWfUrNanPrP0g4Y6QQSzZjeTndCTBWdDglBPAiLli4CW5k8SrW9AL+l
u9TcxZjVOhRpgDhafULynBbZ1GNs3iHeNtjPC/8UTfsyyqNerFx9spLjW/b9DgJ68NUy8efuUu9a
x880nZnj5Ooq7x9/Mye0LyH7I/PHP5KbgvpzdkcE8eJhQAQgMX2qdXE1ZTLsSAWzn1TdjOODgjT2
ctKxvVJ3rKiAgh3pOewiS7U3NwXF2rXhx/gX92kChZYTY5Bw7Yj3ZJVrdILAyIIUdc8wGEgbPbuF
oYFoDg/eCR8UEHyxmWD/795JJKcG7kwoCKBtVbdDk1SStCqzUN0cOENBS/XlVclXGu4/2z+FRKhY
QOUh7C7eDoXjtJYyyhFbknO/77/bawdOX667njr93ofGgmZrJffAZaUffAvSJHk8G6XHs35uVRRa
x/l3Fhw5X2+gqQW2njyAK2Nubmz/9K/NHtMy5eFx0jx0OF7I/9MYm0+tYha33uG6dr2Ref0WZUqo
g9aSb2TEbeycFZS7X6vliFPUyFDWJWd/MtnCSC2dQTIasOjAWGxn0WT79zybWx8zNlVmx3B+W/ED
Jiwo/7EmZVGBLIAHgEGqS/3jLWP8WQ8mz3h1OlVe7ly+VtHCxp/cPVPHzlujj2Y92mOeFpD4oWuL
0HDLcbgAzzzffZyHlVOKiLqpUWgc9D6HSGKrz3jRYUQkzbKu/dpOHwjjpPzlgrlrVEaiGeV0hHpl
GmwiEc/YOjWHQvVuDbrpDXonWCpa7af6wAcsg7eb40CmjExjpM3xKXUsPgCQph291LcdLdKRwMBE
CbwbDIX0zFGOftE/+FN/4tctWz6xoASS6NX6GmiKESZm4u+sNEhcj1TlstxZk7m52zdUQV3Fuo3V
DjrABkrt13jIKj9uXKjb7qY6ftfsHdiKKB6JFcYtizVh/fgy4vKwwaOMcFyotBTtgl0ZSnnRytfs
cDYaK0YvKHFzMvDmCfaQUmWU5VCtDd4rvnGWIYB414X/+EAGzrpDHTYm+5V3stCbt4wHreBrULyr
+3B5Qr3FFQCmmw2JV6qHRWLExa6DCnZG+CAFH87n85qyY+QlZZxhnWbqPmjlxh8+qro+ejm6fQj7
RqCp3TiRfdbD7PbpU2Dn6pFD3JahJU5wDVKgsz859TxNaAZDa+OXF5LhHUqV7SlYLUUVDbNma0ZG
nTvdX4pfw/cV1G2FoHnJ19KKIVfeHmuAnZ02ivjFfj23YqUxmyJ9Uw6EII5AHlMXVfo/UmvOe/W8
ttNDwQlcAb/2vVtSsL/YccKTvDRL6Zl/w4yltQJDZr8m8ern2yIojYGTWkEUb2veKWTyaebIR0bA
Pq8Im1Nc7VkakdU1Q5CzlosMXrLJiYA6Ra/uvVIvKq2b7I+/YJqcTL/dsqfctVX7rWSoOPkBCe1D
MI7dHf8y31ZJWvkptdDYRLCYYxYwrjymv1PAYF8SymhM7gaKz1tQGYeBY+CgqsUZ9LL1mfB0Qfog
jvrWSLVxkvuLUQnBD2XjZMOItaLVlKi6cKIRoTr9XUkfovOYEr7bGkVfK9dfhqBkyXSRjNytzRbN
3E9HdrGxYyoEO3Vi2qdWGnqi9tucUlnKIO5KllR8gkq8SbOpyMprEoXuVal0vsIZ2l6Gul5pEKOa
418XYFRvz89KUdfRsOAm9R4jmVvG5Zvkzh5bPRRPoVGA8aF3SUD2IOIrz9/T3pW8hOK6MCVays4u
5kRiOPbDCsmX4n6/EKO/SgqMaSkq8SttUElYrSnCPKm+X3yRBE8om5W3oMNYrG6JcLOs2DfWqFjV
ky86GQFkOA3jfC/IVrYxM9XxOkp+uKxzYa/UJTGUf/QNBzjxFystsZm7xdYg8M2Ory3jAx3lqdRi
Ro+hJerQcNlp9ag0JvBJu44MfWcxyHtHrY6tKKC5r9ma+5DTMBfXgzk+eu432OnqmaY/Z+3A+WL6
eTF4S5OdD7a9ql6W7sWCNWg2khCkNCZZl9Y1f9nM4wWh/VAikxP3BUMQ+xPKn5xKSaCZwLm73q1f
WpMnO2wZYGq7Yhw0tfQjXYn89LHzKltG50iTFSXVTlX9F2YdQ0LbTmL3f8NblcrCzTnz2zThgMk0
h34/6qz3qBPpuNGXPInCRj9DqMWSRiX9YSNn9GyeXWiiwQHTxtaN9C0ZXFcKzB+HZnYelhtLB6ou
NICMNqgGJEHLoXufmLi7BCo48nVUXLJX25Shkm1k8qVNupjQHi7ylMjtUFAujS4yE5ztNy0kHKIS
TSeOYEH30J8O5aJGaA1twlcns911VuJpo58b28J5/B8k2tfJgWx3GG55MQJErXAycsvhc4JEQxVF
SE8eHw9Ialj0lqoCkGTGfF7Vx3+ylrSPwk0uszpeyFAoORophjMcdTRQ+Dyh2Cs/CjjIsEwpVtpm
LxGOCcHIOQrQpDZGfZBb1mLRrVfbHX93MFCwabmoQ3TSxbTfidVZ845IviSkFE0B4jW3krU2eQ3R
h6r0lQ4xHwzMcoljBfB/9uLRAf2V9bybcqt6068ERjVpikhZ9vTjGV2YyHCfPCNaIgXIEHSeoECO
+onvqjtSO8o4wvkClKYmd4x0fBUwpbNGTTBrLY7vIq53kTt/Q5j5CcTVNm54ZL0elhdeQ7McA7s9
KPT8x9NciONGGktE3d2x3HlmO01oI+Ko+ZbIDygj5kc4f9ZFvFDTrHV+EOApcFiBEUWht2jjlEWv
JQzofyNDYqv4H6p/J2j6Zjb1fg5lrwKMEb69Vstx3AmfF115dp3+2SIcZf36AjHO6gqD3YFCerbl
Pciy+LCmf4e6UqNe/AuYp62Rf0zNbolYF+GXzrFbiqjGUSaVIoJ48RN5ZOTht2X8xB/oMbwT3Vx9
kElmmgkWyDbK+ht7VF83jkkLBl+HIN6AkUuzv4rcltmfl+iSMKAL/uQ+87l2UtO7jps/agyolHSw
mWIpk4AfJaGsJt3jw/5kekskKQqIt5vLW8FfmpgMzkrmGjV63+3m8sYoM1MNmSMD29VjkDkizz4M
ZxuumIW8HHDEjTo5Ot2lyhG8uaLKMLRHR8mZiVZbYGqHYTVDvzHAald2zIhgc4HKZD2QV3V5Yzxz
LO6Fx9+DCBv9CYpq52ohzZ4QokAhdJJfuyznd8ip3hgvVpohWSJc+i0JD4qsKjQ1qChASRxzXSFw
4VLiCDVH6J6AwPX8Za4NjLEhfjLQrTXcH33X7CeXE20EYc8YrGqvgAEvVpetBk7h+EAmOi3cB+sH
G2fu7rGJdRiINODlJu/eGNf++AREo4RbEtU5+XoB2o+1BnkukC3iYgRsB0Dpf8Ba0+ZBtXJby8P1
BlMG9X8fee961gZpfZ3zfgO2hOSWJkNDror8y/YePYOmX4R3So1ja34F4qPI5Piyphh5oZHYI7KI
D8d10yK31ib62ATiWGDZpDRKu9v+qPXfxv5RqIdr2zzzOCzaL0hwAlEfSI3FGQzEh6/A5rT75m/8
8dcUus+1ah0tUqyC+EbgJuiarwW6phStv+avwpFxxuO9SP7RLWhMoA/Y5dU781k4fkfi7iLt33vp
pv4Op/DB5edi13XovkzLX2NXHFVoFOJ8ShUyJ9snpOAf2EByvIUJNNL+p9mqjCWrgPUpRWz0l+C3
VihxsfPiBIgPABZU8LU9VHG62Y3IHuFTIojN4nlx266V1kquE+Lnh/dzG652tDP1BNpQ2ifPMzLC
Wvzp9OWF94qFRgn0CdU4yyvjD3x18HMG8BKP5dJ3t0npWioA8Vjizm0vowc1Lev2zOUgLz8hw7UM
xOwVeZJNZDEwLUG5IWEFszcOM3BxUR4R6+ER8c1F+BtIT22LSeByebTUXG0y1exlGGxBtjiFLmGB
A6hCQ4NPVI1kLMSE7yVgKOn0n6rjcOVWkJseBgSer+hztut7GqmDpXpZJF1yDkVLpslNIfJJT2Si
w6VTGzec/Js/2k0RLyeyYyYWBjY3rfC9/iIF7AaSW8UPOVNf8UU7soorMvskroqnnpBAzxais9pu
JvgI0BQDO+bohMi7KYvu/rHTN6xcFz66Xx2se9JfDAtaskvlNchkzpmVPV4tFJdj3x+RtojJ0Kif
HInMtCKe9b70wKb7aojqtaEKLzvI41xnamcjq6D2hksYDvAvK9S8JFCVLVq5HtdiPC3fAoGTd/zG
PHVg9gydXczN1/sKjM234IjM2LLkBE8CngTxv+SibeMg+T6vhjYCUCM7YPxtob6W7yOO9ROFhOlI
/Y8L3XT84J2plYWmY9l282BRsJkOx2a3ika2VnsMtlgZ5HWUQLQhtrrVzsKrIF/rtS5L0g0/H8Hg
30hqKHrreSos26kyCgYhJVjJ9L1SJrumY/1kum6Eqcr/NGXOIMpzH8oliDy6ufxW5gACopR1MJuS
l9UXKSK2UWsQUeHMqm67RO56nPhX8o5JJvKqH0V332nDekfBJOGwx7VVwpLSkEQd8scspvr85fqc
Nwx20TfUncSYH/O1mRq/CCxBIyaa6Bb+YBZgA3CqZhRyzS5JHGsEq7o3Y8LpcVjSgHsDWY1Q0Xe3
TnFppxxdsbNPVzkKU84LC/+25GwdSFsNuzmc3w6e1kcGONoHurluRj8zl0V/AWT4Ily5cOM/C13a
LMe7ifDClT1U27hgnZ0yFLGvfDPj0a/cQnApcBZAaMXWMnCah7JwAX3LY6oPFndPv5g/RovpMVjK
YyZE6BWu81b8Ed7/VhvlQFUgW0gkYRWXbLHs05MaNay4jaEiq8oZwwdLnjMYhEpqiHgrxBNHijzR
ee+QVClgtPs0QGByLxtjomku/t52YcEsANdskew8BzXoyv2Ec1O6fNGSO9hsM6AOzvw3W/yRJPE2
9jnnb2yYm0VdGasjFBPd0aHLJyCQNzWiB25EPdSA2VIJhKe9sdKAnvDijXzmn/qVMqUiMzwgDz3V
Md95h7Ks+YY8/Rw/BTpU9MQKLE++joy4QGwDkjgmCOk6q4YgxBaZOTMg2MP/SLn/JgC0IduNSq8z
vyWrUgLX6toszEAx1Et2pmDQdNm/0eImdMmlnHN/mQAD/UlDYHh1CPk1ac1QZyZviFJX3I29ObXq
9Us5DJO9568D2on89HSp/dmJOWIDoB2b776Ljgkv3njUDVR515gWgJZwqp8nu5X5KFG5NAaYZiw1
o0Gt/2Gl9Z5N+6pj7mdzM5Oree0qiOjmZt303BgHSGiuNAX9FbKfssRzEEVB+P7GiYdvh18s1Piz
DnJm2YPBJI67cs3H6EOYk9xY9tYFfPZhgLDX/arF7NVGDubmNIR32iYxRS172cqT6Erc4z4hZHfk
y9pflDtP6jcAkOYxUSPegi70QtPzVGUNHl2rOv8sL54sqjT/A2DkVIlo+p3MNONwbBjTCc7iO1N+
JZx7YWQJiOnLrFaC+uxgeTuI9l6dPdw0O4aLDZ86uQVB91EWeJuwCOwF9Gftq6zJM3QeIWIPn9rp
xODkAfIFTvA0y7KYjmdvcu6L0K4eOkMNtVgfstmP0OBFr9YWZvzUpnKgFR/rw64OOSkSkc5eC9pV
zPfZ/A2w+buJbwcZFa75p4rTYDjAIZx6TWq9NhutFQReqrEV/J5Q5Kc0nDAMq0k06sTu3iN944rf
UieF5eKVpVIyZgGgpGW0y83uPuGAfvWX9RHLZYyH9h45tcQE7qL2TgkkU3sszrDuMDyJt/nRnm5b
/1xJegGVEc4e6UmkQ8e74DFOKyBAWqCZaLlhVg1VM3uZzh5p+RE9bbWZpar6II1t+9Eah0gi0nsS
Xsm19oJfvzUXF3yxN5Ra9h5u+Y1qmemIkTbISPZCLNKXdruBwd5kiYtkoigfrwqabAZ5PlFZQv6h
pF5/ZTNQ7Zo036g6o0iQHQs/1ZcHE0N0LWxRy5GwFkiCoNNaGSrrA//WNvB0q5HSC7gKvJkEDgjC
Oh3mLR4zkXMSfxNYUDiCfcYV5+w/SZ9B2uSThE0HrKx/dVCatdK5zT8dayRTMFbZORycDVbJqRCH
MEaW6efmM7TIyML//QxHtKZXC5o1MW5x8pgthaYP9GuKxn9/d72GR/a3FfKb2zyIMyBbm2V5rqvx
zYEi2FDrMycHWTGDGs91pxYeNCyE59j1NSG6cea1ypiTUQ8a/Uz662sb9/izQ3B6oRSGWs0UJFY6
2GOII+9L4GP4t6GJw4okkZL9SRJqxuT3uoNP7n9WWE3WsTZzoaYv0nFD52hBGJUbfnVUI/6sTyPt
9rSI1mmV38i57M/d+S4wjACzWH/ocxH1r7E0IFHJurQ7r9nSVhLfRS4xoT8/NwNWOUxi5yzZnbq1
gJY+QwdkN4/8mNo97mEYfuIXeFuGCWLy08sO0CwmJCPO3Oll8CesE3BzOk90CTJ2dskPJ4MKII7k
ham8BdAZlldd0BJbTl1xku0WjYuPS7zbcX8iM7F/4la769uXLc73+5Km5cyrdFYLxh7r6/v+jJCL
8WVVwifSlR6IC9BW4i+7upnfeR9JuR4zFD+1O4SUOu2Et/auEmYcpjJyefAllnYnmZlgs/dthB0c
wOuHFC+ynelFFAXKiuQblfSmHJrCrO/tiDOOcRrV3dbB/ZaXRBkL4evnzD/En92rhMOCZIRXyF2X
CiaUfWZ12JSr2a2byGcdFZ46fQM84h3dNOo4yjJRjY2jdM5wWyWGj1h0vC0r2YdawwbhEWzpE7PC
a359DKQurMkWV6iyWq0SeQt+Eihvry7kbc09hSjgXgAOF9thhW5JqXDzTBz3mLFVk+cgavF4mOKZ
iaZYd1dHvRUnnsGZKPjK2GduI7OwpgrrVBlj1U+phTV2Ynok71FPnfRGZewDGC4tX33lw2gs7g++
echvputkmiQzNhiwU4cCP73z755DTBVc2YaMmioy2Y6GPMlLIpvQ1ZSjTAH0z4+4jIvjUUf3wme4
39e45wsNvCa3Blvrn39TowVAj1CV/mY81QiIBl/6KweQycXqLJBYBkGwlZJms/2jyXpOgCBJsFJo
0YUqzCl7YjCkcG/PwBnIQgI8+HSGEf/SvRl8HebVeVOKwb3T9ciqD8jlGG5nGzaav/7woPdeTDdS
CKOZ87BSz5A2ydBkIh1zTx6j9bP5qLHYxpV/gv6u8TemFEKKkZnw4Mv1IdWHItc3vfyP9LWbWlWg
IncwVAVcUcYkyhJ0YAzVkzJHVW8i1Wci1yTncn//Ohz1SMaseGv/5E/Ye+vrslFolSgYH0DvWhA6
UkXxWBkUb1odz5pDjC3yiEu35D+cTJnfnjVC5nNxE/xqQ9XglPyPaDYNaJjVVS7HXXtbJndUTowr
2OdYKSIEeHgTEPcfh2dfnMn1nY0FF16+9//gjECJON261UeAsqH4yz26x7/gpzS2RT+4LaGnEOto
VJU8L32PNyKER/xS/6X/kYIq5T6v9l22s9YW+Gik2MNNOmcdCKWfU0qn6hLYagosgZRIW+OQZGU1
gKk87bQqVqm4xL2EKGVcRs/lRQIwXdshhUYObvApklKl9najTNCX/iazdJNHBo2GJ0Nv4vsicGLY
4q3+z22qqj9+bieshflzOGAxcP7fWTxQDcmHpOuc9yWJi8e5DJ8WRP4oSWYcOuXQqdmuTQkx6EIo
j9UV4t311rjC1gndzKpaJF+QVN73duqeejgrPm0AwYxCtLTOT1GJGj72tPnytMlj6B9/SQvEGbkJ
pt6h5WT3KZLW6nobx/pBssaDt1bWsvCnP6zt0kZu6tey9iH/ruelfQlGz5UHxE7QL4r4so5qm8Kp
EqqH0jJmeRHW65G0ALuAz5f98JyK7LtRgq18VtdJChSOS/bZonlSsCxHtV5JoDUNUwle7+Obt77J
ihLounfD46Rb6WOBtdpaoQi2WqszwXxQpN6rLtNrA8yOcoWTfKAeojHprpKgPA0Y/U2bS2lYh24M
NuBuJDpEhUJV1A4fEi8eZ+cxHsqvJseWBdfaeiY7MHXagmrLV1eQyCEEdB3OOwiGJWggi8Ab3HK9
FkgN9Px3+aOIKxUA2uosfnXiayGWDEIrpdnPmZurHjbRiUyuc/gmYlHRmOGm4xiE/UJozhyX1LSS
FBWHULFfWtY15KI9k0QyfVf5N1qXYGyGRfl4vAf4AmdDa9SFHc/JKW3qBnAVFBifwvkRYLkyYWOi
Rcp/f6sAjFUzQg98jhT+XU1Dymht611OdKOL9UFXkZbE2SysF/x53e32i/8eUqyHcn9myIxGHKqb
yMXjcVmhg7kld2MZz9sZ71n+kl9hDzycYYQFkFKfQSm+kod6EofJbRGxq/ldCqU5sbe6GlwKE6mJ
ShfFWH1IuAILsBR2BchI+mgVqXS7gtoLMEGz9AAt/ZN/9U2x4Qt5A3e350mJKbBbsHARbFHE41N0
9ZZ8OACB+yDo1+rJVme52yYH/RRoAI6k87+yrFw1p7iM638R3JFXEBtyHniRdjXC1CyFVrgYp7E/
ZHCM6kZbRoXd8z204g7YzvAF3sT4jR+Vwuk19Vd25tTlFMI1xC7FDdyBfQyipPkhDrxUWkkfKozo
ac1Y650I3FjAKwrfD8TMOhd0koum5xCMBFZQtrY1udULCY2O7AtcTQX3UVGBlCRGBxVrvlgGTIJD
RHxMxsi6Zs3dSqxFfBFtc40W+Zf1Otrp3bbIu/4VEy3AXIDPuK7uamedKhBmRVZJOpo3CGgTmCVX
az0did3e/rROEJ3deKGXZ0EAJvMyHV9/CgBYPb0uk7j+FhJGeaiqlE7Apa8k33TNL6eV3cKTMvf5
TwXXbKrzlMij2Het+j1lH+ngKDsUUXnhDro6/Qib9aqMxMhhuZBWaZ861crV6OQYmBopR1vwx2td
9+n8e/qzxA7bKNksPNEYgmLaHzdfGmE3DVfNt/4bnpHojt6gPgb6jRJqxTcYQKIwRZV5AybClAu5
kPIH0EKP3cTMWFQG1PelyM8w0WBb+RXlxM3gqaaOwXqzalrwzgKFS9q/n+Sypt73GZtGp4n4QaWW
dQuy6RX8LacniRwZpLmSZeBzxd56bWoOT1LmnuNXfN1bh5vtGv1AZVF9d3L31HtMJ8kibYQLMYt0
Iqszf4acf3flpsG4Du1qNG7qW+izTZCX+7KRBxpV/EH5nRHWPUay/XF/dLT7dCxZ1SFpmv46pVD7
/nP5DkYR7LBpjTm6JWZjlUbNnvh7tl9rFaTOaBzmDhMyzfgYVJVoTuOTx9gTYwf6MsR9at0VW+uv
ih3RORRZXQLIGB4Fyt/itK6nPOZ38fsH5/D2nrb2/Au9iCFaPRi0yC/bSLKYu/ViQF4m2LXeXNOU
MzK8K9/ShwXZNI5azaJeGHOOIMNCcubj7PD9naVTqvEp8e/p1IsEzDDbnFJOnrIoOzEVAYplzNxo
WQtbJVHoXFSTjPcqHpcXsp47kNHvBe5+FWZj83W+aSN4zGuQcmctxdPClDn/F3yEEAavQXW0/Uxh
W00Hdl5tp24AAY2vWfZXVtcKZfmJo9qAZ6MuwLiTW6IIp0WTHIEC/15oesaAvLjJGTJaWfqvqTib
o+8eSr6kOfh8w/1jWA+ulfUJq2M52viMz6gYIs/Phxx4yvwkmAtbfD2Apn0rBy1x8nXC3sixzKaL
HLp0KrZfk9MLPF09bZeDc0v5/eGESlQ/1GIo0SIspJHOMIXm8e61J2tzbp+O8F6c635ZJtqEgzo1
Sdh4T2wVcCWxlLbVOzRgFoEcMqUyougwS3092FCgIevqRLbhQNANrLneTGJn7PUVeBrz50EjDqot
UY4qNV73plkt1ICwm/1sv0Cws3laID1JA+Cr18eY6ptn0LG9CFvKzmRaWy5zIu7Kqt2LrCaOsFum
EIr7CEs+okersvPFNelXxL7ZDy2+BC+0zoczsITqrn5fVfsfXMLEQC/h/5F0QHb+jaO+DVqyTQJE
MrUJ0fsFWsHa3RfeGHAnAsJpgF+5yYYC/cx6YolD9HNH4C0vx5koNhT7yd2vtlGbYlKriBqwjEJr
1Z/PqWc9nGTUILHDdUA7gkuY5xmLpi3AvuwYM2SWDsp8BOw+r9zkzzv7wPx5T2Qo/+aDeuVsY9ou
14UcS3YoP76BV3VGXgckMIfgRREgk3dwNO5aYMqpbvluPr58B2BKm0hIaLkmkjKA0wFt1eoRdAHQ
KwI477fUTrQCVAmu85XqVbXZDMPblY+II/LZ9y6A0HXIrWQfUecHxabOreqp/0S0BsVN7WyuUdoH
AyVU6PredTcObHnOYGm7GTyiR9M+RN0s3xE2EKjb4MQASTyWDAcosPZY91sWAPd5oSGZLIfkRWbe
lpDBQRfxHl1GXTtB4mDTGcxIloMmrYqzrfMQLbeNIbaWGAzs5o65hfRoZpXSn36DcYyjpsZZ9rXn
WimRJW0d3RuQU4lAltAavTk+5OyWTmbWNPKws6rKE6m0NVh/CI+d5LfV7jUNOVEmCkKSlJg22ARt
e6pR8ai4JzI26QW9vilFwVnLZxts/zQJ5N9oLdK6YjKNeMe90Lj+K0d0nL9HSSItP/7QwaWozndL
/1Gx8s5H37As2E3TP7HHheyMrmeJ/DWoJxOj3WLUO5ESyQNpO9Mci9SW2WTV/ljeHYIcdZpn0rAU
81Cth8FLwZj1LtV0zcxsztMZtK9PRpT0ZZ2SVlUtDQG4CkXmsVoWFt9TwR8bf764Xes+Enbf2xPz
4gsAr/q4n22t+wV77NPcWjhkjTFDUU0DB/LOCwKq1xyIPw5deNvDVTeCoPw0DADxFV/Ipl/dAoCj
PdbWZmYhkyRr0Hb7u50kaGS4DgIE2ZBeJ9t1ixpkaHclT1Z9fpYcEcJ5RGA/gUdarz4VywZ/6hri
fR/zgYG1+QMd5/67YUytdzJt0aU8iTGCWIfsq17/jfoUZdcFV4aWh9z6essPGcjyi3QeolKAXsjY
PEVHJD7rIb4FsAzabaSkPRUt+r46d6sfygsQa+zUoiTiOGayzOYPgXz0pStt74+CajXdkTKtmNEB
3v27Ff53H9hdFGEoAq5hxlLVzZtOJWN27ueqkL3T2XXckn191kRrqcatkjTZtP1v6wCIJQG01jjZ
hGpJjsWlQCHmpiRa/YchaUvz/lO956mL2wM3i6qP0exICHqF/BKlAQyrjU48sraEP7Bak6w/wtvc
TyitEych68m7Fmo7FmAnvx24i1iLdG2XMM/Og/IRNatD+CQRbO/PTwh8/ZEcCWbzz4+r0uLY9H9y
7kZhF8lk0P90TvDQPMOmVHCVjNDVY5IFnFwYQdaOOMlM5Xqx9ea6gJgw814uRrGv8iklYQ/GlPpS
SEGm/r6vK86iswoVVfkJWsQH7hb4theeOuZIXFhzXBumqrrp4LZBuwB3vDPhrB74m18Vbl1pNZML
STEG+wWiHxoAUsfwWzKDkLuFTUqiekRoqX/vp80xfeNgcpWZm7yxpWHewuiS7lTjizlXth0J/SpS
WZPQfWIzahNeTflvO3BLQiajJFiRRUJ2/qPB58QIgsN+hKbEnmQ9GU7E8pEx9hn3OA0Oy08Bp2sF
i2JLWeZ2MdFJWjfrLDB9PBHPH8g4UkZxOByN3GBRBW9zsU5hItdDV7kjPDRxWoJ65jx/cgk6zFW1
tIYG5I0S46R7ulS2i9wn0P9IuQWlFysNiWCVWmoX4d+fbtAHt9qIBo3+XiBMsAofIOjp9OVsJooJ
wZyvAJc2cDIvXLCKpXkl84XIfhIwgdT5qGb6KzPSss44m6BPn0FLF0nJhzrNZ3KZ369rTxZcLKuz
LNdD0gkoefUKzdHGVnuSuq95ONyQzYktQ9hnVQX5tVi2daJ4F4XbaWWdU0iJlAgbISO72ByD2p/5
GzzvIPkq8j+ItbdMpEo+1R8xsTdUnpyA+y4Rgic1pWieyJyTURwVrj7rRuAwbbj6IQ3+vYP6QqRK
ZvpzWRoqslfaaQre/wa4cfz6h1mR2V2MI2zXsMDsjjcPrjLiFg3PooM+E2c2HUqi7S5YdQegfNRB
bFqWJ1HwLEoW8smjRNt/nyjiqv01zO0aziUzeY6Ls0wxJt1hVMBL6uXlJPQfQw5E6lYeOkcXinCr
F37Sc/ovbElCNab/uLhYtbvSHun1AAHp6QJPf8qOKVSFYmWY3JT1YgJHEsEGjjRPoeX6bWPDNxSp
HTbzFEBuArhIuhRaECAC+Tyn2HrLeX9dTCuybtb4At6TYutXqNAks72elfNj1CPXnAVHERUsYUga
GDtYuPlhVKy3zDCRqfLN8Q6YDxHQYGjefLhU+/cLfq/O8USag8dyDPm0301MtsRnV+IdWVdnKIPW
iXYHlje0CTc62qvTGiHjlT6vWGdIL5IZYTEXfFUORx2WCcKXLP9cf6+4XXnejf0xJpcGTrOLQoF+
T7Q2Zs0sEi4itNNFaTwNU6x3I73N4DLt52MI5HqbOTmOPJb+96QnC+/VRo1aOeGQwaCj5vHoUyoq
TrgayjNSYCJ9Sa7w7GYuPsvAOwlY4xi1+phN8fjGBhu9x0ug4sTHywiqbfjyx/vp9vBMzXf5/De4
u/LIbH9xBDlqaj2jSRUzwug2yj7NxZCX4D1w3Y6m4cs62GYeiKdChdchJ3dMPCZZQnwNF2hmK5zr
d4jHqQya8fJWrknaTuce2n8JGP9Ww9OcI7JxWygBCK28SdieDdTAwGEqSrrWsQQDTL/lB/g0WAgc
g6Hx5S/CVg24owGEBoE/vP+7KMOYj0QIi2gegLOpkVcaws4s/zZLwgFVTqZSvZljQIEKIv34+3Ex
wl0j4C7dmPeqFkQPBPZG8vVnxA0c/wJPo/rd0/DQTX5xWdiXAJ6SaCAWhknFuiXNCrL/wU2IgFy9
uLu1Zg+oR7piVo1eD652Z7K/k66eaCSvC47FGdMYMchdOgnE+gN+Oa2JAHRDSYbzi5o2vadDt89F
N2bHq+CIDdwinNAIJP/QvJUQ8JF+kh9qmtG8FDFU78hJvG8buA2LtTFq1ZCGE9fRVImoxtopih6C
5t5wtycUo4ZVvg7/Nq7uJsgpT10ikW3ZlQpKq5EoUCgfJQ/DJkMMpVfj54aiiADoqhg0+3Nm6SpW
t2ahRxqSkv8qISUWgaJlZBY+SNUQplhhPnEuSnEInsK/MIru+t7tfT4uOLEmXbBUtPVUvmMw7w3H
jjXREA7GIkD/kttVk+Yadddi3C1YgMyndixsHUmnuhLw3wZlRO2whIkePMzTjhVKRwnksrpq5pYx
Qc2/crzKPK4A5SJmA/ai3cPVxp/GaepT6MO0vXeoNNspZpunIeE4y/SwuVtUDCz34sja+sYQ++JS
pQjSD077bS4CuyaHNuvOH6pAlc02E8dF6NtY6JBJZcraiOEsQ4Ny7ZoDUmGFtQDxQ9iojKAXfpiY
6/X5Mt5LB0+pGLSDazMIc7WG9iIA0wn6lZIb8WGR9vuhMTssmePPeM99pd63dVWgW7sXI1tH/cqW
WzVwK4Jf/GWORblqMQIma4YI/TsZrny8AxqZRoLEn4RygSCOhTI+21/y8pv2i+EKLKsyycyIzYz0
2zGYBKnlZYt5nymb8WFpMA14jW8MUswQjTMsu2IOJzmpyTCcfbpGyVvTAXHmLJ23gMRcIZ46LAZs
9t5YxH+DJSLRWgw3kn3imQoUyySkBbDla1K0cQS1lFjrIeSB+t8Hj7RhsksI4rRfG3UTXa2SC/gy
H9WzK4WGlqRZP3ltSY/Ds2Mcj6FvXmRjfp7LgeIh0r+BC3L8uCI1GIdKc/tQEJHcTUTohoEHdfvT
/NQ9jjZkqv9PPN8S66JEAeH/+KKL4MvFfGM7PIcFfkiFOm7PbjtF0deEosbcMnO3J7nGYF8tJ60H
p9lHQIwdas34vVdpVxrNg5zLl3UvK838ydf7+U22rpybw4GuVIhJAxU633Jmeqqw/UELBmosA2Hl
7NdVSKsxV1e8QBVqFxeZsips2RVpckgWVf+6aKGgXgxFu/Itu4mQ/x2uJo1COzT5cJrncdZhr7Cc
xI4vWnoMN2CbEA/42maORjwQqe+qXYTI3aF7CmLbB3PjpzNkVMju/+56CrDmxfi1pb03tliIaChD
r2XrOyLI3O3KO2s2D6CbDgGUNyGKiRp60e8wMc0tbTNigobleECyIOq5IXGjXkAaFfS/Yt/MqX5+
de9sXjYIw8SuXPwgEb1F+EMjRPD9hR8wyawOd6kKg92lL6moDs06CYaNaAWCDcecmh+RH4WLMDAs
hAAKd8TIi3aUADmuIo+3okgk0fuc/AN3xAiLCtL20FQSnWCq+xTe1LKQZyfNMdySN3KQlJaCyVaR
YPuTeiDYMxU29JNd+HoozWLcWzHcQATwz20FbihYTqg54cnyc2AZV3cs9CJp/oR/TYrnfM1naC2v
ADtdzjOYbjkeYQhzkfQNVsnufY7q5/t3alKfoW2Hjp2YMh5lwJXB+qZUpYosQLTRazrgZPPFLZqu
+zRm2Ve7plTtiI5j4W9B6J3X/rTHFrlVyCSQM+AikCLVgpvOqXAf7u7THOCbIIXTVYtYB5NI4k9c
hLarUkqbpH0NfPHUkWQnp0eXGLMMgB7w4wDtsYlcp0V6ZpQ0FbxC0DEyaLr8+czIV1J+65FK5U3C
bvzgkEYX3OlhDUQhx/NPUgpNaxLed11w1CZAFLE5MYEN/K+9q1LqYBlrrdRzaFzagGdOoAml6ljT
ZwBDsXERupoh0FYdN8LhLrIId8SiQeIetIMHn+TLGOQCLomi+ZkpMhD3fa+k7jyUyLQH7SCL6UXa
90slksbHlNT0fdUVy+d6Q7OR8KnxZe/JeDXaY8Fi3bhvZoODdP4MxD4G+gwIDwlw5pBtOAmR2B8F
vP/DJuBkDUSDAk1rGGmyg0meuXT83/qn9yYGmMYA5x10N0wGl1XQb2kndym70SyTdihifzoPOzR+
69GGo1u5BEny9dz6XUiB/dfqv/+J6M3K47GFbD5s9M2iNvDc096guWZJSujulXPBlWFEAZplCTVn
p9sMnaXby8MnnaIS2qqHXxxRdQIabYOLgGRoSN+YQN2/YVl/ExihBpOM2ydSREVKJ7VDSZ4dnbMl
NDh2OLN69KGZaIqLQ9Vf3xbZp1QtYGcQB9pK+CXo/nWvcMYULOzGjZInOO+7Hl2rnITIwWTduMzY
T2W3WhQX8kak0FzKqgQdCsy794LrogKIfAAix/fVjvBwx0sEk9R5hV2N25km5syX/7S92rBUqlLC
FNZAH+63OInsFYd1uPAiyIvljpCvZFO3/HoScYmEJCDSN4vknYKmZtjCTbmjtfF2R9c+LQ5Fwa21
5vLMF67tbRsHwvUKGEHK1Bi30JBQkKAnxL2e4Q8hRUpoI/hFOePbQD8dUbtn5PGAJkfJfHbjBxc9
hwKIqitc3s3qZb0QUqIjOkMUXjipOPZphrdmjkhsYl1qzFKBZ3yrAxpOtwLI3Is0oGgyTmyS4P52
RRObTElrDZYuC0v0L+Z/27x/UCmDcA3brT3T8iKzYY3lz7cMuo4d3ijwGFhkxcZRvjQQZGeNp+8S
ICBlCG1sOkv5MrHaER/o+hMr671J7dyAnESg9P55XW0thlCW82cMPYUKeyaRhFLbSTMbdeM62eU2
sbCE73mXdgMC4sq1wzBWgoXux9SBZK4HkuQtY1SCheeO7gihx/BiS53va21aNXswx6Dk0/4Tnjei
fibp4T8tj9yhXDCVSLH2akEKPhBg8J1ezsEPiP8S1ijxeDGcu4MgcSKcS9FiTjEyItHmVW5K3e28
W1dGl83k4d8MfDMAS4+7V1BL4y1DN5WGMrW51B19kmldr9Fb2blgQpeoqwx4hygYDtWC7/BFCVTd
DD3OGip+9eQDC7adDmQ3l300EhkcxZKgxeV7N3c+ing9J+xCLPdjMNxAnHBJcg9B1IENAO+1jWL3
zWPOdyN+iynlZrR+0tdtN504j18yc1nUmF6xv+c2dyn/2EHzaY2Wn6SyJHVjqA+BTFUWvrUsFUEN
DieqKtLXEqzOQEOqV3Ko/qs4mxkflGPe2zXytyAZZGKsdVG0gYtmSAwze36UhqVHbwbDlMCtXROI
gpOqvMKfY/9vGLz+bS+ynhJ24nil56pdLjqKHxYMZb2ARGm+TX/cmQESk8ojMWt02XwJ/lXZ+Xyh
QXddQr1KzZ4IgYgpHez3ajZjMNaa7rAJXbuFAYQYgW7L5SBFO17DdB+1P96chZWGESY49tvBEVuq
ehdnuT7Ix1cC8ieU8OCj8+Bo4lFkJivAPegcr2QVYPK4PeOzj7A69LaAvJD0C1Q4wic9w53s7N62
JIzCmbcxuwXtd/awkL2wDv8lJrb3sDOlkaquLqTk18Pk3hKmvYhDBvqu3+pdey3c0tecfWOkmaJe
D9lkuVZVg/p76gGyPU+B9uKBz1sN1NgxsLurfkyUI5I3/yKGtPG0P4cZBmA9w9S9kLQS/nsPNiNA
AV9WNYn6911UmVbGQ7NohCscGGBFB9WKn87F81oOj072PBlVXGzwvU5hC8nPHJ8VWuOiLVd68Vcv
fqoNMaB49UeDsc77T7t1gXPzxL+60DH/EdmmrUpb8xQBc9tqBQqlkqdQjbuivCrT/L2nDRrusTbH
4DdnmElLq3qfTAGmNH9XZ+n6aNlA3kHarHhmjUzT/jbhwhKrH8yTfZ8cBfcDy1cv+dLEK06MWDCS
8/2k1O+qBqqdkA9EN5g1nMIdZZC9Uky1oZH6VwdsXZ2YnCO+Prymt75HAai7E0uMIY7sqB8EmbWs
yiiyKghOHqy/wEL5hDXNUTmbkGq/vnPYHSzq0AcBsKPrM9ZquOeJjo9jfy2vK+g9QKL5BqpDOABj
BiRRhN54tBtJ8qiN7LOtDM3eDGZSExG65nF0N6thcilV9bVPuqPBbyV59w2hXcZyMSDKLghYTA7r
7wvSfMAIatxMstDSmMWQtqolzpavoPr+3bgY6J6HaFH/ERb3/uvU/sSinMMsZXJzRjooBYxoHKjO
7fooWhlhsF25QOb/yfZpjjR00acFMkgEPB6ZR9QtY6OSf7DK7EcbbUgjJusq9FDg0NrGhHTKiThZ
rQZYzH0CXGPEgEeFsVYlu0npLohXgROQghBuDe+6FseFhUyTW20WqXQv8V0Dzzc22iOkSV8R9iW2
fq7/AlLbC+WcRLeqBSm+zkZSfWi6GBpUChSryYv0BU8aQBSRuTiWvzxmhZw5eAsqprzeugAQaT7x
B3lZ6MWWtB6GWvm2PubySu3xMLkN6dfonpO4pJZHcGMsNSEVPqts4rk+pvrMJcQR5jIZoCLQ+GUj
87WV2Ou91jl+ASz71VnzeR0F3P3c5oiOs77OfAz/kuEsYx0MmdpZK4BmTEWLYz9CrC2kg8mvhzxt
TMcT3XymMyWsYLX06aXUgNBxBSfJpHKyEIWMkvfRFM802JNFB0FpsdmdiD20xTCTUwyOjG8eqyjt
H5JImwI9EAjgQ+y5oz8QF08rqTXWgQDTgayiYrGZl1ARyY5qmeX2B2IXQjZPak/csHE7q7NHSGWm
IYKoXJKGPEZQka/rzTwfsQMlKCcN7JsgacNOd1lwC5n8bRVVJI8oJYEleUh1974KQ7n2h0AfMmmJ
Feu2lPGA5VqK2aAnz/RHcHy6Yf6YH2+kCUaS4UrXXR7vJrRDS5ONMrSTrdHmjCNxKl9RCmYN3+M+
re+lu5zTOn8dsZo63QTlk9sVgv4iATVR5LtU+mky3Ug5g6N4sE6Uh/6Tb0gFtjmcrACgHvG+gWGh
s9YOD/rTbtwKe3FXjp5RQP7KgHZYEeTEfS6cYd8xSoacEVE+8MV0nqNqpqisHDi2ybJfJ6xigtGk
nC/kuI67JFEzdxZx1GPuwlpB+Otbi1YdOXZKcu1gEJ0q04iZHh+ZY0cVR4uvuH8/1NittucPTfm8
gEPQLOwSlmFGi8v+4mA9vIjaozLbgPdflelT9qdJ5txyT1dW+6GulefbgP/sRJ+wlwuh163D18+L
TpnERt5S6RfWgBzMUwWDGMLp+rCzR6MPkVugDRGnrg7FOzpLqhnrimSIM9R3GKVI2jjLGyphmkTs
xfNOj8YO5/Mwde/Z7rYmaZwaUZWOJNBWv+eVHSuYaGYP/8RPMyxvp77tKcUlkZEisYto8IzUVyMk
Ugc2X6gZ/606nA4HoN2Lr7MMxnW9ar5cdOvWTvPjY2obEDG7MBuQ8Siu4mZVy4gF8BVUitEZZfzC
aI6yciV84LDgi7NI3bGoCJeW5bWd8+SpmJcD2+ex9s7jjQHcecLHEaEMCaRD8PlV8U4f+gqRrNsH
TR2DEsDE3U2bMZLO7TvMwJ8RSNO5A4UKTLYB0kUD6TOG6Y7WnT5IjBppKQecfOLMboKGIVVmq5/L
2XeJ1XE6uj/PuiMP/znMlus+cwX0Dqtwh6kQUq5PRKNVlSS7pTldfCQJ1ZVjc9Wu/ljZ4OWz5eWk
QbV+KxO7/WEyjkuvD0g0xnwPAeqpicdQNh3vy4zgh61IO0LwCw38KrUbsQyVmXbiH+rEW6atVJEH
KemoH05TSDdXwz2cG7RsoQRI6PT6jluqd3+JoHvjbkDQFYp+yiowm6cqIlI3z12V/ikaTwzGExk9
hPIu118cPrnQsob8wqJLy/CE5QcE8muZi7baKRrvngxJKAyJb1Kdiy3h0eEenM8x5mIn0ABKb0WM
fPB6QiLK0fr3uQaR6HQ7KfaWWULFV3PUpqjvnDB2ZLGOLXVnVfLDxooJxwgJmiV+gPVjZ3aFS6VL
JtNdJb3qGYLjpq1XHFS3gUm4+BA3igol04uzZyhxlgMkmpvc6THACz3bBykfJIl681+/e8Pw4h1N
SARORt+yTgK9CRiHYM5tjU5CsbSDvq0JnlsyO6ZUaI/CR5O/xlCFbJkdgsXQuxUTOisauShGRZIc
Kuk7/VVJQlYC6enbtBiCZrT7fHx9PVMZ+/b2nUz+YTqIIElu4JMRhEXh2byPteadddgCuLq3e8iW
MiJRFvPhzuCdFFAU2gt3w0ETZ+wA/UI2WsthnXIuiLcKLSOdzKb5aBzADDICrqe73lYqXr8biOq6
lt2ms2Ij4RaFvXpbYMHwdHHTqpgVp78BkMoOxDb/Cw0DA0BvIba3gzVR7A3rNlP/3nYqYxhaNXpH
iRGvgPiVuxclPvuwjX/M8mXvhGy4ZvSAWi1hmidGR95TmVGk0dZyj2+VM6utiXzGE2/cuC3JsXsj
ZQQSFMSatsuqsW3kuXCHpiOBHbsv/+XvxSeF98apAk45k3dpwLHO54FPmD9V3ySWABp9pjnHvMuN
mvxFrwZF8M4BXlWdirrUEesH/iol9hHAUOtE4qjebhexXsbAomeIYg5Fq89Oa0D2VtV+yoFUJ2fi
/vrzZDUBut8tRfoLQhV5froppFqtZIuz9TiPnDPXrR/UQdF6x5TzvC8+LDCtoL2tyj5tLlj0Pytm
X+lTGwa0fJCSjbDnDyXuRYX/NvdbTz8bH2Sv0vDwC8IFZd5SGgnPegdbX4X8s2vVEBQweJlAUelb
bt30ZElV0wryNu7yiaUz/MLdtbYqPzx3jYORyiAw5h7I+sAPjmt3UyICmQ4ZnpynAiHYbsRQrpBw
XK5ShtTFajipEtMQLPdZqnGat0Sut/AHh1QWokjm2+KhIhT0y0q1C1Gv1YpqbhoCMN34aWjVMcCx
NbkvvBRR0A/u2KiIIt8ZxhoWe9PLQ2mdpbhytZy9niLfskICTegPl2+77xBq2k74cpsATrSSjo6I
tlgcDu07FnZvnEdA7m86sZF6gncT5Cy+T0fIMjilXShbIGlhqbwgeMLcs3EV2TVLOA/6u/qnT1lj
reuve2lzIhteIuwhL7bZrEuJRIWTLF3823WiB/9UAClUu/VfDUGSV8qGJHLnj8zxWKUTsUiR/p8w
D8RESB6gPQS3+uBkAc4Z5i9gFjAdBCF0nJFnDOol8l6sTmVp+wUPGFWWMjFa52AlPDlyiJOFEFjK
mChKFMwg4tdGvTxUG2waN4SrnoBsCpC3bdMvoGHDfPv6RSGPt9TwUk+4EfOPznmYtSMgbeSRhkhE
o5D5KEgtAyDIJw6iPQ7BMPAlecvnjTFFGe2y1iqWm67kbOH0Q7eOeDdiEtNFvik/+vlaJUFe+s4B
jbsAwcz5UJJhuHAPx/cvJgLBb+ql82Sz8etCq5ldK/ufX4I/hpCT2ccjeo+QFcCm6xTr1natJHmi
WPhgrVhOwQls1ftKn1pmSSMwHmtr4w++UdnaP9GHnpbG6UIrejWw34uETploDh/G4qC6Sy3IjuMP
Ox248HewZfHUI0zTKIDn0u6hmoAk3eL7KrA0SeMaV8/iKKlnNwmMuUv1XD06wJsny9yT90hu0ZCZ
9xuWXa7j2cYnn6pBMx8ZuzT6M5IZrJFqPvw65ewsboqugXZtBNKuTNj5t5uW0gz7js9Ui5KvoCll
eklvF0pDO3ZzMp7m/Y02c3D8bLSdtMAKrWJco5gcae2U5U2ddRLaOuq3EMutV0B8h/0ai8WIISsX
EM2fIRx3pl07ZWxvWTBq1QcigKIe3kszcij+riOLgLqDPz9JFtwc5a522frJ22XqEY4zpeGJZL/B
lsqa+b1JDj3hpUqEhiUz8XQPYuGXA46cJ0osfIjcsNI6hGEJ+wIM3XIYXEbpSlpZaaJSwI/ORN0S
f2ZZqFnqqBKWbMFlIX0rNoe58/zdxcDEdbgk+8ZuZ1jyJOtff7tN0jOIyYqnjDEExVvjz3ZcUe1f
gX/udxJG4aLPcPSZF6Wvy5mqQG6EeTgfz4miVOqeLOx5ogy7mQunmR3L0KaSjr2J95NBc9XmeVSo
0WrhIt0e81CPiACuYqrYb7MRoS9QkvOjq1EiVTkPMUEuFvTURvOFPYgZJ+h/Pmhu7Jhvg6X6uQ8C
g7EtbAFqEvmmb341A7N/3c23gd3aLaO3XUCLbt2Rak42MmBmXMBS99z14F6zzGRKTJVqg6t1UtyC
GUNvfkMDKzYC93e6C30fSsW2ZGXv3uaRDT9uF4c5FEU/2DSVAPM7ctdcdMV+H28HfdJychvbRoIZ
fgBEAlOsazy0dd9cR+hxqtL7CRXXzxq/WGgiyGawaGYFP8QB+vH5hk4UTa6hirp719HIDJ2WZqVC
mK1GBwfy3nqQ9enz2Hh/N8jIMnwEPGlY8IgDPFsGeM1habQQC0WC/ypS22iVMi6ByJ6Af4BYjdJu
ci1YLz7nXyNVwAWHyQ/RkpIEh4DL3MIMvf4E0zG9l/hPodd08ArFugjvb3EvYR2JwxQXqrXgiHl/
6XnCV3hxqpR3XPhmBCIwUSXxhCbAcuyZdD3So6+/nOSByjyNjz/JojHDPss7rvMYoMq+sYR3vx6T
i0meBJSQb7XZx5R3Y7PD1Y0Fvxnb9uveQ+Xnbb0fJz/a4M8NpZU+P5Mzq51oQTwj5W3BcB7kVMZ5
rSrFONlTmQCVUtd4/LUMvfNbQ05pmQJjVRLsoawFQtj6txSNwneOpjBhkUmbMJAAysVhj7a7o9nI
sVzu2Doi+WBmAZWDmnl/WsI21SiJo7lled7JOajq2Ukc87rFKbMTNsZfMRb+fRc+1kukqG31nZ8C
SQHEeFkm+PSVkuAQ6Y3o2uEJ+zGiTUHTwI0/fKPteUkrQi8uuKD2ltouQ+8xdr3rfYTHdF5rSDiN
AWyPu9ON82PR9XZjt5PjfrAJR4COuG378jI6UrV6MVU2G/RdbV7vpBPVbQE3dsXrsdlK7NnxFDGN
0w3RgPV3NDH2j9ZEOcM/keEbQdDhVDSCRggm2UsZRglIdnIo0zrw6VsitV/tAhgoA1qhzcZ+sIRS
kS9L1UBmLpMTAGY+yN3AJxgErSr3lJ8uJR+aHhsL3eaoSzxnB4Zc+ml6O3BN0D6FPY2uzHqmIxlN
Td3+rFShLLxc0q2OUaGFhkjrMs9JlSYjT2MarmGkJMtIjDP1dbuzAmwSmOJg7q+0ATYguFS5g/Qh
jq4UUpQHMNDw4LEBRVdV3X1cEocDaFvWz9KwQjh2qfg141/35/mkDmK0IohYZG3RXFlBFcpe1CDQ
nLlKMvWsvypXX9h2yR6hBAdOcAWCapzS19ZKd4dMiw1MOFVnx3pc+jCKYH9za4QMs/DcTk+6Kh99
cPr1GU7bclkZr1J6IbKF9LeCxcE+PORjTWqmRH8O62axazxh2l94Y1XzXgCgWUaaleLP1b0NfpZg
/mU6PT37YXttGmN0/VGf8lHNX2EYB8qohTu1HGRK9CY9Tdf2B8fJ7zzJ8H8clnhpicklSSDG+Rcp
ESisZuENX9gdqdShm5dSa2eXWEOMG3up+tD3v5FBpzJZ7k3cVv5vwGJBGrUDod0MB2jwCn36CQ12
N8wCB/gSXavt4nbW8adFGqKUJdo+c1uoFnE8Hjowys5W7o5B0IB0FMAV5O2ujCrgIynNvXKQ2Rkz
itaCcXSm9spZtgE32CcIH3/+0S6ggkodGnBhTEmhvCA1RUl+pcEeuvxveeUb4vA8ZrxMIgYlyDlE
QIXPy45EsaVj2LeZsPfLHTkgkezgRRnNQpgDfGCD/maJT8dqHU4zEzso8PTIOOR0v0dYZm6swRF/
tGpko4DUFv8QyhC1IDbxHb8PbGTIpFbkvHZDgxNC/MuuD7dLsIVr4vWi5ycVqJyQ0m+vSzM4hFqM
ekp5mP+awsjGlgn+6JnrVuq+eV+WNYVgjnhxs7AxIElk2X5Ew9TuTyLx6DxVwyUgoe9c+LGVbG8e
fK8nBt9P2EPLKmGDpDQVzWWPbb8ELC532Fu7Ds/LOZ7l2zcHo7uFKXeH2I0E36Pa2v+AUEjEe2Oi
M3VCxq5DTVVCXWj53hw/SnmN3WAuq477Y6H6KZJ9oriutpsX3Lx0qPOKgHc1AHLIih+9vxWHB3tt
9jf781XoNpJiEUsWgABwQAljkiUmSIE1eOmtHbvrJl3dZBtpPyGab6jko3v8SN2ueG7Iy3/rexyH
yTuqE1b70vKez07aNaBVV93z6pfOMsfRZ4Pepd0CBLF31MctEkqlchTDSDHOUevSehdw/bmv9d32
6RxJMVH/8VJPlwLq0MsXcjMhLBhjI2qEKbK7XnwlBcv+Hwf7Z7yR0fHEX9p+w/NOR7k+1E/hAUX5
T9xtswJeRCm7esCXV8nuU7G6TQT8iJnpbeS8Vqot3AwPcRAxKHlSxS1Vx1bSjlmMv1JcJuYqVVpM
12UPGPUqKMT7rz6N3QNSjGZpEGC65QUTLeJZE9R5KVV0ZI/vPrIwAPj9gHDTWNLsulTUUp4E2cL1
Am2DZdHSYHi8D/YBkm/Z2r62A0eRLegnWxasgNQHNKn8Yv1Pcz0Pw31VFaHPjF9VxgwInovbOmAn
iNjuQswgHFNZOZO7N1TpGCyGPD6gbNbxEK/un5hIHVV8Tx5wOKoZagxIXz7F+C7Y9iCKb+I/K969
TkcgrIsUqbH0UubszT1dfJlEtAPcDwSg+gWzNGUqtJuCCRQ5A0DgDZy8BRVTbnQJfiHYaD5LIMRK
g9IUOdEhGxdzU2quX4lRxKtHX856jDYd+9ZQgsUa4h4Rrj/Lv9gkYbDQra8EqErBAJFEYh+4Ffbk
WzC46fE6IARwiBDPdOUo3CsivXBsapm54fvgmXaC+7fSf8gLCsd58ANvpyOqeLavpTY0XVh8aUZg
ktoKhRgZGkrnqCZ8zoZ3n0otvonKqUq1dbrLaeth8VRWkXNWp1e3L7WzNq2y+Uq+FTupkvceJSuf
ADs9haIWskV9mk3QPPOhYe6JsjCyMjx1DKJ+TZGee9nEiu87bg+bu9M90QUa6JDCfjduaHFpF9C0
39arxV5b5wgWbrhBwqzPFE6qb8X7VjX0qoCZtNSnRw1hJVIM3aJXPx4pntift+IL+qiSLh83vvPp
utDDYb+Ih8/Nt58ubIO5mQwoho3CjoHlcbifLKou8P0dtwIRrqnktZb+42RQhMCLAmyNWcDSUPfg
WZ2XDQVm1uNS7Qbwuf1O88D42xO6OA3lMbUJjnr5dVCi5fRhwJNek6+Zl7gYl/TlmFvMPaEYSQSy
nOhFMMeD3Q8OsILutrbITfQ0lbNNG8Ao7vIq1RZwYMxlSeOw3zUYcMf3CRpW4lLKtCTTKCOMI8xA
8y3NwU1hLV//YUAKyVow4ZC7JjMnfPY61jDBX1HgpyItO9Hr8DDeA7NIKtP1ou4xZJJXHIrx3Qax
IzEXSMqrYUX7igMvg5c8FK03K96qeAhb9fw95fEpCFfQEzrKDJbaeJEE9T5lgiccnhW1AEHN9hKA
9C8RwoQ+airfjF3HwNrkk/208UrE39zxst53l4v92kLxADWGf4ozLd+3iNk/mC4xGr1dJu0VjhlE
I2jIknDDUw/TK+b7OQomIHzjFqORxHXBQgiqq7++BjgkhmWcMMEk7M8czH3LItPPXLrWghb74/sP
uKgHiWixKBmE0nRZm9UNkTdEcSnfessnaSmFU4o5L/VIvt9P3ftWBQ1Z494Hc7HyrBSidL0c7+V9
UH24dVyGc/mXh4gQRRaPZjOVPXNblZ8RhY30uoU8Wr0bWnT7riQipgM4F1I/fHhkc+34F6K5feJG
Mh8Ug8tr1vC8UlIgc9oJWxi0DVBvIDzcdHE/N/skhEDheqnnAHPvnIHgeclVF+d5DyIk6kihV79A
BdnKVOI++awE/w6yakFa5u9f+xnX9tERYiB9302KUNNxSPrDWKURMuzOMDX92m3a7/M+JMerV5/V
s/pcqwIF5ziI6Ep7njJ4gyQqJmBc/J/tTCd1AjGjXJybRGDxMH85BvARGYJQIkU6/QKTRZT0z/L0
XUZTQdncBJhNag0SM74wU1QcZAonkOpS9vzUvN+QmBjkSpF/e2Fr1B92liTUzauO0xrGN7+uM6Uk
iKiPUxOh8du8B0q44VMlMIruUI74ZxakLarO632d/RUJEAraBOf+rT70pLcu4zAWmFbW8zZXp65I
pYsFlZDzEkeh/amrzzPAZXDBiXA8+K5NemCYA3bJKSdMF+5WVAlCYSjzYIyx1utt1Rex/NmvtbeU
8IFWqFFhRP4BoQ0JhYmXFHj09rdylyoPzVJcCUruWQxnOKNVLSFvUYJ+ejOCrTkFo8r/bljGPHDR
my3LL7HwGO5wUpTpAtxtGF8GHCMYnRFU7AsrzQ++HnByhGc0dWJRT+QI+3RGHCTfe/sQDok4vcoD
c2/U1Afl/TdU/nMGKzQf7Koc3/qWSnF+3NrsQsKCLPfxJNz7m7jjfwBJw4RvM1+7uwZDcL7gbazr
2pa9k0VLpmK0wkWOikewz5vQs/f65vbnb1FCxuywXFXWmY6cvCnEY/8HWNdRWj6feKlx8veHN3sM
uSxGjJqQT/zT/xXeU8fiaTtvCYaRiWfg/ZKe1B7aO8HTKt8p7qSWEK+AT0tJYaK3H4fBsIU3miWj
wUhbpqquXXQXOzJ2jNWzTRSor0oPMiZWbN3KNMSZBAUIb4YMnzDX0UGnTRmqFAQg7RdW2cPfx2dF
aGzenlbOa2Ul8S1aOB12NeseWOpK2a6fdzhfEoOzGCD9PWTtEhw6iJC7DFDxoLVPrQTIWce06093
VjKmMkuZ8CeWEUCpkv1V0tKpqCaX1bOQW5JGODg590XQHMC/s/JRYnjgzMUonalPOsGjyV5NVLNJ
4cdhNGxDHqhtTVLgt+3qjcRFl959RdIUub9PsLTe/1P0F43BLJZCItPgSp09BWh/BN62qvQhe1+8
6/PCdUy7UgLuOERxWVTVX8v2dtMmQJoekrIEXmZKSqSXKsjoxxq6j2Ba10wxniO9764N7cLa1oz7
/JC79fRv9q4cP5e+6KWbYKXLdIFQQ0nWecW/94Z6YYSZSwqQtiwfySYCXjRQyO/yt++ZYtnPD0yT
uSTWmEuWAxNOKgvQNUx0aMsG1V8OVsjQ1cptS5c+0eGLRuTUJ9ZSH0XlfajmvCQJARnnPDN1UbJv
4fsrWJuVyKHCTR0QJccKRyWxZykTiRkzRdveG7eeWTAHO2hZjgU8ZUN7lDct8apPw0G/rKK2+IQ7
a6AwIGJdAiSdq/Qcn5YATUHF2PxAnOwV1EJmjSvBfpfEVvH6jTxLNndrFGSUx+CxVAqqaIyyNnd0
IFN62jxWgeyHmHZog92jk6SlxKvf5Pa6TWixCEu/kp8boyWc4ldzrJJWr5j+Imeqe+fNoj00X5gu
0egLqMphg46L2nqiYo825+88lq2bNp3nuJtx7weec3MqKKgUrsm/vzg7+9/8ZyxtOdsEx+EC967i
H/8OrxiIvTaT81osRiQkodROWVTW/pwqfJ/Sn4dLfUrXUREcKNiT1/a+SKUpFyq+qkxWszDrc2Ps
w2szM+RfJbL0GjyMBkn8bPf5SH2hNDVZMie9h9+Yke5F4JbblEPUX5mFaNgYq58f7xcADqXdeVeY
uy+B3JhemCc6nDPbB+JACOEk29k4Oe47KSwRgm1Bw9vM5UppIc96r8RzZ1lmy62cTKQKTDfGj97a
oeKXdwZWiys/JuBKeXkcyCtbnqn+n0CkzWp9gMEMI8cQqEIz5DH0l3xKIlKi12pRyKDRKwUCwPty
Jvck8SnKRveblaJDifGBtkZWlDvOrwT7NXsQUQHe8ol2397Q+Lfxtb7cwrX/oct7xrgO0/5ydqJU
GV6vpj7rUNxz+yznP4syr8wBf57fuWy/tFLvHbv2jUaXPUwlEaf2qgfDUQvfhRWjlaxzWKjEn1Ym
1M+518BQ2ARkTmMFNwjJW1Gic2Z0PUP/i0MAHcWOygDyRTVlvN9e/x3msKVQNZQnpTG/scKJljVN
28T4KRpDDAvJ59onaiw89qZB6uq0BO+ncshWEZtpgFqeUpU0+tWxqJLjWX31a7C354750h8/AMy1
6JdRdAWBy7Wz6NF0tXu2zhPnCcuCt5L5tuV3rLxtFjQZ2TU50G+Sla7Wor51GvEf7lMYNfnAokdj
oq622WGr+ehH6JFpaSRhCYDIG7pa4Kd55nQ1ZT+8EaXHy3udiZJ3VVMfTLbboFqKm9J9DHHq7ibu
S11EoiMHhylBUE7kSywYieN58CPXelC58owysviYBlt0jjIcgnYrbLImX7c6pLmxG3gKZcRER8TZ
soey6MZJELh/K2K/T3MtgN3PhReaRT81FAK0rPr9OzDlIXMYutHH81dLTdRdlc+1dp9Q2BXEQTad
q/kadlDBCjrCVVQsELqDhXjjdXDnSCBiSmtCwi/wWxLp4oE8G74rw2hSXX+mmn2V87jtBJaXbpui
Y8XA3uZMK7onVoYcJXydcVfAfJZ8eems5bOUtuwp+SPvAPNDQ6dW5qNe3Qzkb1cdP7xGZKxt6HGN
UGwrpCk/iQL/2GSS5JwjZq/PkzPin87bxGVdBFBimME9dgYu7OMdJRNySTY3TerlXNH8Vcbyp4Cp
yV2DkITmAtm0bBO+OWPl5wra4hbtETC9IqfpJju5+FceNMgqBaBUfLbAT+rIrj3ABOoJLDYxQoBW
rEjy+iEnMR6OJYKMGf5Ga01ciUvw4M1avhRvu8CYHYhByGJIOMS6BnNUzgRSICYgZxO/vGL5XjSG
UpTDRa8erc1EMVlG3IOq9sNfiR/uO+bGmQuvR53rvdn+XczuaapNzNRM1KeZ7bbUlDFtkmS4EzLd
jM1w3dUkCwmy7KTommLI3cOxiEFrKTsf5C5JI3E3oT+G2ueC+eyy4NGtLapx431zKJk5Qvzb7fYU
++P/2J1URaZ/aN5XP4WOrK+pW67qhOsqboedUsXUbTO2MWIKb+HqbuiSzZpiaeh6iF32Rq6b/lDU
GrFBwgSr768KBcUa/Bx7QCxUMPXOVx4vmx5j8m4kb1bxcWXscrLJIdqeYlCCc5r2XhHABE2s4en+
0PP+jO+HlbEoizfc6pnSYsvQafus03t1EHaVOELhfScJO1JBZkBn9i0w3uVd2Xo0X4H4zzLhrfUN
/nRUi1LSfDBrBNZO7VPkfoAUd3gJ9mrwxhGjrWbqG9n4VLFILxekRjBZMEpzCObCaytFyaFzZtZg
P4JnpY7iCOLGDZH3QDaXI7CMdWex2TXEuSFRwh8I6xA2yqoX7mlYL5gEh/4rokOAK0O1uKfD24fj
AE6nlcc/kdcRhh9dEwAS2tuet7DjktTjiMWeFiqI09PaKj8cO53+oA730+7g5scJn9wUXpbBFZXc
Ex8tDFRE0fW7bzMoA/871BJ24X3+znMaqATeWTui/QJHchgXyYhRaE8NoaWYfPlLjRYwZdJwLnGh
uxiF0szHsIefcNYr8/cBwD9wtx3gwu/P/BXCgcWbUjGotSkMzISkQZmqpVr3l3tDGGKU7P0QroMk
IQJUXirdKFXiN0lIRvBtX/BPgTz8OGr1sXnvyWG+vB3GwFCFrva23mcDkWGMdFzOuhUG3Se348Fx
+edgRbHy52C97UISBNWk0k7aECNv2E8zqvh2B/y6ILrL4JDxSzBcb/DCwfhWgrhSftcOujJcnpqH
qTxGu4M=
`protect end_protected
