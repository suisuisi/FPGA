`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KW+uM6VF1w2J59GnW9nCNlQJsGixF8tx0hAZ/rW41/3D1CeVZImR6WnUvaQpDzqyukd+6NkQKbGN
gExWu5ZqQg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xMDBrDpWBXBP7OHGwvc2M0BkXvMWB7ITv1UnT2qOe4Js2r2cnW7oeoh2VyCQnRlcD5/5v4x0ilk7
SYnxIKWha86OQxyXekUUk/FfC8gHjHq1onEx72iLRF1IJyP2uvfzkkf2QBdHOBx47ZQtZznsiMU0
L5XsqhqXEYz4PbWY2Hk=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VMbRO25j8i3mCoADFHnJzVSgm77ZT/5C2IIvlXnwpW4mrt7S7wmSCmqhiM5DFJ5Ws9THQGN70uuD
KB05OqsAw7C06UKw3jqk1YuJneFlrHoYK2eUVMMqZNujHBgqiSTTD711I2UkKNn73Uez/bVBPpd9
PRjWwinR5K0A5AmhD6Lz8wwwwyOskaapqXMew9NRR7uq0S9dPu4SLvcVr0bLibLH+N89ZXa/jbp+
3RJFf4um1ETeDD0WiPpKrrM6rZFF4qVHwl9ud4x+sUm8djP0zyMiPTHUKtPtArcITp4mnF1+NkrT
wDYneD2LHP0FAOPxvmbjqTtXFF4PGTOJ1oXxcw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
d1GSv9oPpaKSilyeux7u2Woz/0x9kjq4sTDzalfL5yaZvCk6EoZCUPWJpU7oZmRv/Ax8OH3z7k1z
METCJ+8BVuY2CDJClX3XgMiI5Py8maKwTNjYV/dHYTYzLkK3mXJGbg5csvPwrCOeU+M4xHazRoE7
wb9weTpiTDmjjtkQxwzkDhueZstExobu+o1+4M1IlkozLe6feFl0cjI2cqPbUwbJTGrZZF/k9SHw
3wyjv2T7mQEH62Rg86xozQxnvcfMaL69tqn22/3E6/vl89HetxqVzvvqRP8tLywmT5TFFIT5j0sm
3c+IS968fbpBOZYIrEydYNeKg72LmSE9iPpPdw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dQr35UX/fMxQ0mWuO1AobCiYrdyLPWPk0TWHWdk3vLBJgl1LfE+6RDUnWJRXUC5hPVOWFqSZYqsK
AJZf/+ZnqAGLivhYyIF/5NZfCfoohZ1m9YuLSsEh621l020TqGOoUQpQShaWgqMoYKhxj96b2z7+
YdqoO9I6ELgg19yegcw+dT0uyWnqMVz+ht86aoxRRcTfrsbsjbLWpGQ0zFrjec18nsVisJ2mDHYi
vyhn2bTpQM1hzAHgNobep29SCzR4ti6jMCHejbBYVwUfAbTgkeEolUz3ITQN8T4EyIlw0lNjyE0B
QAFwREf6JPt7qAJK2BEECVwApmjimifT9w8+gQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qG9+1e9HWsJbBpwAEVNnIW8T31cZpOW2uXs45hNxf47rvFTiBbFVMhyd3zCjPtIaPRmEoBb93+cu
0EmC9pGWL/bVJG/EU9c4aPAamJKgILiFaKDFwef8LhWgpBn4Pg0usZUhKWtYKS4kecURd43d6fNV
O7c1lUHnr6MhTqMm/DM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AdgnITHk/9qVO+h+BJMfl1a8jrneXRtseQcUYD2qbxt1U5m/vJIyMxzOcspnr7kzQAy4iExLkHYB
i6IvH6c2vlU1/DTjG6yF1rSHS0JWSqSp5MOc7FFGeKXAmrBbCl1GijRvlhH5yGY15xGlRfMQ2hX9
6dhQBGdpLmE7cGcjhrBhvlOlDglLxPii3XLx7QLF952WaQBkHb/t5ErWcnZaSJtyb/nMeA6N9XSX
7G5mgb7LS4zWeIT0uQUaOCyjrWCSTFpzGCi+rh30sIf3XVyLgJLu7z8TGE38ljKW8e/zuDJtowPf
8ed+mM+eBRp6Zg2PBp1eLpGzbnhBOjtBIUf7pw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 67920)
`protect data_block
TgmIO1kWOCWWI7/DH1ias3gj1rZDjBJHFI61bR8cQnhcdK/buedNqGcNLnqV+0TBq4JgAhYP4RWY
WwDY4oTWlQCTFsI/mnBZK+dyKusTW8HtOe+SWiqp2E2O6/DmfCc+SqKkVoOACZNNGtdAOfmmR4ly
uArSnJpFppA8q6rWW+ETTpylB//IdMFCa2s9fhmWDND+OIxszxAIha00xKwCJdN3yVErTR/kCg+v
o8usycUmOVSCQBnSDjBB0gaKh/4gurYkLAeTiRmXp82JXa+U9R8+e6wl3JB5JiZ+4+cfiMFVK7Cy
zqUw4Nx1aGNFq6C9+oGkbz25UhPJ6IzO6Jaf6VuiUibzYnjncMS8elEZK/5bseg+3mlyQHWA+CS8
mZKp/v5Hl+JEtUKMskGpCtquiq/LA/YuMnQnHm2P3AmewfHVnkHeAn0PqTm7/yCnz3zFygnuwSVt
470b3oHLs5r+yTDRdUDa5UoA3Riz5nZQ1ZFtPlvFL4g3S7yk0z/ZyX+Ppt4Ra4r/GN8RoVKiCg1g
ulW9sq7TJFyfvAZNbrNkltlgVlweDLelae0938hkXp6hbIU3ObCnxe8PfpQsqAH5owHmOiCwxcek
Jg0SwvQnuFbKeaOV6xAlpkHi3kQHfmMPny/MU0az4f4lZbT8lm0xHGbtEH6/AmG6Tk+YXZ7JHCr+
dqpL0Ev7sA8D1xI9fit+1bQg/QqH0cE09a+v5RkGDPH+57Bz1wSW+f+yp1WDmlI3IsV1MMLMFKHL
DClVWV9s+YMQ/eikrXFkwv6oL5jHyVIr/tv5yU8pksU4I34XRuD/4geRzoRntPSxUJhctQKL95yd
yaxeWbLk5QExFw7W4H8Y3ZRRxyNCDBarYF0Hn62H0Cv3nUI+kfUE4yDOtoSV/3CFhVzwOC2bUGMV
T9ibR3fv4bmm41S+99Dnd1DJW6j37YFQ9z8kNjEwowi4JuUCVMfO/VKNn7Z5lFtOtO7J1Y4pgQ76
GNvttxo+FIdKAlE/uVw+fK9JEinqWNH6h00twcCatwA/3l/NuLWn+DIQYd3pMEZvlVZ5JkuK8eYb
DZY7Lim7kzTaHNc9NK2OPF3KC7Gr3p55Dcu7DcxkC7nvuce0ULArYgizNw8JeaLVX095rqLhlaNy
7ko7NWVi9f3HbWxE9Y8zmPDOO/HPxx45Ujh9/HyskxJAslPDCdVXPJ5GVUXcj1l21x2E9aep9+Yq
8mY4CMIGonVnBn/ln3v7riHNvh4xIccCnsKTof6IWy7OA07hqNNHTB0fe80wqigAMjRYtQmRweIz
fSWy2uHlWO9XZuwVnrq55gh7E3E0SNoTLnzcliSma+JD/bvpX1J+jKU8zc9VTUxmPAdDEmsZc0hw
6Z2896EYeTD5f/8PlC6pdvXy3wEiC0GqlpdyAP7NJvinIOvokdngbEgsGdj/bRj944JJX7/zKoUG
8y3Oa7exlBEsbjyuryzKuR7A6fQRHVHdQnDdRTDGtCyTK69NT4f0SX9aP1IINDVPSmeUJmM2iI2a
mPmtGqz6EFSWsnEOJpqZ3s6zs2QZzS7Ahxts1Lnx2KEscmnVVouookM2WKE//mDbVzX5KoI3AbP1
ZfCi/Gu50o6/5dutUjzaNiCOKPV4gshGQyJrCZSaUFM7GaOL0hzwnf/luQ5ysuOisDV06hVDRkUv
9egUN9dKYlB2nwx8BRn5If/Fk1feCqykqor7DlHSchl9oa7vm00NTSy3dGaWWV2stF6NfbJ0yLvs
wknqrC0J77CNtzDawsM3C/OEKYbbVr0t9TE4L6VkqoKuUolGSzIvsXqOgWNDjfs1xn2qfcVJtz29
uRfa76WmJVt8haiTtjtiq3VFwlWShEKJt4fbvjPiba56FSzBx5af316OzvZch9PIiuB9LeFDkrDw
/Xp75xqlJguJ5B/MzFZ2RiFPG6JXdCDmHeO6gepo9OOrmrs7kCStY8RPC7Y0l57R5x57gnSbOVOV
h+CDSA0Q846LnBmZ0tKgT1d9RyJBaJOlx8XIn5oINC7BuB8q4NK89RMZHg4S2iyGGwfGO+dYFe+2
MzMMlTfydsNusu22bULhbdykP5+3uCYZWpvmZILoS9n/bCWLFggdXdvt0xZXYMpfK5L7QThLS352
KUbG8yfL7enTpX+KvFMKdCIGCkduEjXkS0m322c3l54c/9ZcLZi0lkicQY92UBQ8HgkzJ9DDx7Xd
t+xo0j7ZDfoy4JJRm7dx0peSUyjk7i+RY5T3HcYoNmc+wR+UYgEV4bw1zoqNTCzWHF4FcJXVOHCO
4Frmk8/V/pQi/80jtP32SmBViiwyUIP7SW9lZGemMtPkwBlMKmSRGL/3GwNK3EAQSK9e8YS0OsD1
9aut8p+uRfMysIy0YvrZRoVvT/vLXOy+5ryikNdKYyEQ6mS2GewR+aPUrxqPfrhZeO/dXBtD1uX5
BhRzsUnjMZPSfqdRypSxWyGqrcyRqLy14QJhFAjfXsF3ciJ2b9S2nOpFnU/jytTioVPNRK0/uOeD
xmPxEUhqg48AN/9v85EdcJn8IJ5aGNul+opbmtlvaY/bTnCbokv4kljQOeS4ZP0camcVw2Gs2UEQ
h76xP0JjqClZSKAyocrVWZvw/gWCBGV98S4p8pvtn+2RoXxuPYDQwHTG+2PQDIkI55YO+AFXFJl1
k01D6orj1ELRhTOOMkYyy4u0qxPbtRW12MQeJR2jJ31kqAYBfAc3uzyNC6mYWBUZ2Kn0oUZqGqrp
ZRegiNCd0OM+ce9Yrj73mqmBn+atvtoqC545W6XWe+aWV7YVzt1b16ioxKk47+lWSWFJe/d7sZZx
Sn2i/Za0x5zl2jAs6pYFdUV6h2OL94ICCfMG4URCrVhx+cBX2hfSs8wFZwCW+3FpJYRDPQZJR2wt
bf3ZBKVt4RBZr+tcrjPdr6CSuO3k+CWDtVcE7MIRexUlDTEtzY9d904apUOXDc5zEiSvwlm4/G5y
As6Cup4+Xo7ouppxmgzWPd09vq4YAs+dJWIPTYsG1R1J1VMLp1PrunFoA8H4jGU4l+8AzgKMrJlK
AkJsBLM/kW7YLUnKCpxCq+/dv7m+R4F3BqLVf72PjfwZIV0kh/5dpoYGhD5AOuBDBvz2UGqC6HjM
9t1XDvpaf3hHGYekbtF2ccJSuS8J5hodN+arc88x5aqvJ2DiHAjcpV+uA5567WdzztrqaV+KEvl6
xo+/ge2rccPYGOE3Q3xPWP/f8pB/I7KS/c/HlXxLeScTNxUgCWuVnY2IZBls1ZVUM++v5pRUgN59
Tbj74VXXaYKryqHw5LftwzaIvfNpGJJQ4ea6jwzRgMOre9zaQKqHSEht+ZVU8iJ72BFYi25HtrG0
qLi7apG2hXwwpRF5Vf0fvGdYD8uWdkfRlVaqnk8M3KZOUMTgk4KpWRUclVqOYE4EyvrePjfEYFdk
zw+uOKjRhEbL1DlzW9rXM0Ryp4YRcnXpRA32RFPZ/kaL4TnMYnX3wZRkPiDZafCu8mQtKTPFDxVK
w4ykwSjo+4E0FbGpNYs7ihOyA/k1gznR3FyuD+88uXyTIJNyrrCXshG9696axCVUvLJrOCOupwIk
+hi6eeEBgdNpgl3UO/TijeHeMhZTwRTJvvpfvPfvXXQwq8ESr5UHYCIG5KdsTupcUZS9FnzpT1R/
mwW1NnyEj4cAc/uUGLZbU+YVuz2vLZVhhrz/psR45QCUNFAG+D2pHtWBaLdX1l02NNPVbi/jnegH
ZHyJd01MmgKANCXu77WrkMdUohbo3mLDmkimj57sS3nKdUWb4bjFjZEf1PHrXFhqDgvjf0JR4Siu
D7ZRr3sDwn+HGlkWo0+OL2WP+20oS5cKWo9px/GQNEg2SUOkYdCWW8ReQPSEK5AXPV3PlCrrAbSz
6d4oiyO+YlAJhW22l9S+Cxg7sIIObC1LvijD6y6LI7w8ljAVb1w4Sb6xlIvlxCM7//4GKF2I2S0z
7vRKYrR+qOybe57e+k4IwG6deGa/g+ERBrgVKnAjH3LL7A0aMBnIhBEH8ML/VGIwv8m9bpK5jtz+
FBFKfsmT0eaX4Q8hrgNfQpzTnn71Qcv3XGokNJFWF2KCJBjKyZlYuRf2vSE294N+YQ2U4dkaTM6l
m/ekreCh+65+AnB3ZhxlcxvNND6NP0qvaa9yVscy+5vBjxZnfMp90oGr8fyWIDCSTdn6GnK3uCOZ
u9zYiKL4rxUOp8/xeG3CENM3QFp/sUS4VxiJxbvshxDtZrm04VIWvzAW2+Vm6wyF8UgxUqVrIJsm
V2d92R2lQ9HjWYuRciHdmurFDUGCNgkjAsCe7qpF8sQIk0voXT8yiMIlDjIkXWRLu8u3bLqbIYdM
L3CbnF1OlebQVY6D6CO7pmZq+jZ8BEp5avL3hw5YKoP183H48wJAkgK7EsgEJp/pKIulsNu3rffw
w9VK/UJPmqwwcfRd32TDWuuqglT7TSPdZRusEYEwh8VjnlJ2NZe40BjHre/MLZa8eXNkxu+JwtEv
kZc/QSct35A9/8Gg7FdaaoMTgWzC0LZc8fkR1NmXCPWB5t+/qaZAuN84TZZA1/5QOUc33gVacs61
HeoKDkjC2oSq7M/fPGxjszfaxiLP2T2ZHVERPfZwxEGCgilAtwzG+mvCx/MQllzbAgTrZGk9jJm2
dvGaZ7dMQo/qwMvzU+XE7shlikmaJ2p8DumlD+KkcowXq7eFBFFZ5GXbTTa9pAs435NgplSFB2bj
8RA3GEFLrjc4zN1ZGCw6OJaEnVrS9nbZqYLImt55wYqTdO9D73O7Khcbi49f9S7aKpi5fySKdukj
5YJXyidPP02mx3x8ZrED4yU2/zZfNW1bIBkUGwQpO/IfBVQ+TYbRi5ANfqtN6VlFg1pUNU4PWC0k
8xHf5lvF/+WnIZ+PaSeUIDnMR2ZifYwP6rSeVCIx+HgqFiWh8pn2JaGFNNTB/CFR/g/MW28En53I
35dlvnCMtTwXjgXxCe657re3tWIE90r7bFlf47p7qhus/vABtnewD5hlNB2VKVMKHwaXeC2TtzZT
3OInbEB7hVHnIRHqBaucHk2S/YboQgpPzyqgPclzXULzIMGitcereNNPIz+VPjGZitwO6ZhFFNbK
lKwKsIdXSrb1uQac8B4Du6POJy4jnCp6KtTwK4jiQ/6lNUjO63xTxltY0q1P+iIyHIqAZH+hLh+s
jNusWfQSqi8NAgtqtiHGJEOfv6H54z4gdVfcvrcQIDvd+Vz14h37M28IEr9+kjTXKOAK9Q5HWhrZ
61FP9dD22TvWP4DYiAe87CSvUWEkbYGPLdYK/IyQSnU6EwpgmT/7Y5QwgrppBIUXCIAmAFn004GR
Jje8HpwKSOETVZ5SyLDv3UDXrPHPYwr3v41eTB0FrdzCHe088OMejZ+9NqoBkU7rBFKQSojGyrcE
lYO1nNiLF68eXcT9TdOs0OjUcciNv0XjqVX9uEnKFhES3YQS5oxydiuIHho+jykyE8eFVNHIk9C9
ifmFqFlXs3+QiAxrK+KolhmR2N0os6FYXDGhlSFcpQdkb+jHBYNynn43Q62SrhRCovJ49M7zoTk8
RxYorcIfysSemnk/LMvvbFzEK3wRMHBxOtQmyK76uoVOP9yt1gPzwGk5QzargagIINBObqlNmbZZ
wMV8ZK4SGQxr4GTF+nlpoxKone94QN7noH1z9DhcwuwVHzT1EtqYx6AsI7+7W0rnbvWWS5QIhrrz
g/ZZAI5pHfv7k6or4Q1+gklx8tJl9p/n/Ugf7cf19q9GZUqZpLY5TmLpS8pLaR/Zn28NpUgNB6MU
WTbBN04nFsmOc4jAJylhILiav5zWXQAOAes6/U8kiJgx4boG+IogL+VNDE+KM7eWSrgHOdL76ALG
4F+VP5NlnFuuFaaAynzesZy2VIpagHsIffb7ZKnqsIh6iAKu89d3dlXPRH5CGHKUwT5MeZBVlo71
2sHxoBWVzv32NprzhMhubvHctdDqr7cew4ANDJLIPyWNJzfvcdJMEI6K5KMTWHq0eoPUUrIfZI78
oZAbXC0898vZA+TJZ9wcf2oQpiUd1dsQTfCnp3LM/U3Pjyp+nemfszZXvCGnUFGb5/lJu7D4rUDi
DRcDeiYvG/RW6EHgSKCa576SRX5QIroqzx56meEB/cEhEt4JIWlUtNy3gj98UQz9Y6IHiRrNEuUe
w8HUef5hSOLozmiNphBh+wE2CR2OqQ6iFBKM6GWV61uDpNGfdDbbB29cbjAsev91k3IaFYJAMAwD
ysdLrK7dmTBbVOb1HzAroaGY+qAiuaUbRWOHkH3tp8VT1YGe3SxF6DLZWqP87awIThgmSTCVTkso
6rr4aTLLLq0O7nsPvcxaNB/CKAwmS1XHSTk6YWIMCQJT1xkJYOmY5TTc77W16PWsq7R52BRfhWkN
eMpBL5+SRQ3NriXPbF2hlSUj31OFx+LAWuXjaobtipRkVwHrzS0Xj0qf1ZjSqZ997CG1DugYsVmk
W82GF+GtUmcbn4tMzfnhLNnmCRS26kzBsJJTk0vkaSUOUaoPmvNrcUX+5BcPWeiXfumKhft9EteM
ASLpbHAK33Bwt7wS1TddP10hiXaC4qZlX2z7q5rmpZfF8HDCJAfJYH+HNxUxLuASEvwpJ0H6NQun
QXOdwps7g70hb6LzKvctIMk72j9FVPrxnTurFhVyl9QywPFAyT7Dm0MRoonBCBmlADcg2ouDqenQ
Mc+/DJjMWsQnbQ3feEM7R7SCErbt582gWz+Izm8xfF7ddbC88xyNWNPf31JuBApBrU7rTSXofLLf
O+oM5g6jhL73C3kMFsklYme1pjV9J4zWErGe4VYTjpEGDAO2NiVBWJTozciuIU+nwHX+/fiuix9m
8+XXGevTZOLyFmL/g8KZX080/IzaEA6VGB5q3ycJhyAfnBkjbwRyiiozr0W1NxZLMQr+UGFv4xdZ
rWtZglLN9sxVyDu3kB0FYKGgakZfTMnr1iP3ZM+8lu98INmrRAoJrHYL8z+j4ujEriQkrftLgaV1
wFck6+vQU3sgpYP699b1ax7q4aOKc+6+1A6ZWZW+PyEb9dJgLHYguIn5p6yrbKO+MyOks0Nguek/
0ZoSc7vGEXLvfcRfUgBy3i+5vJDPS1wu6Ne380GICibHtqgoKSyszJBAxK+HUcsDKtuU3TCHYI5v
DCsY7JKFwpvtd9OH8RxFmFm1QCA/zzfNVcJ2LjKlo4OggYGMymbNJnNiUjz2MrSJ8OLrNwFGBwH9
OzfAG+ZIrXIbVyDuXUM8i6vme9RssL6QWTTSG8aB6u2B/KJmpu9pZEOFQXIpQoiKn27JjbA07S9I
jpfNiszXVcT7/4J8PEeCRxc4Wk77UtaKfTynzGw2EKyvTK2UYVi8pCWbXlYegZHa/5UWUnaLNINN
FnpvUZVYvDCKRC977+sUZmXODPslL4kI8re06ZnX4cJR1JIdaku2OvznqxigLic2GTNzzXy+7Rt4
VJ+pkP7trWhu5SthW7YzP92DOLrJpBDkXXV1+YJGhh73uuSjDdB5BkcIyTmrJAAHkGemTWgyBrhD
67aQPM+HvGW0KVmk80q/dwx0MR/gvmBw0BakprUgQNFG/pYygGt1Jt9pxMtkXffKyXlx6+qNWisR
2F6On3tZ8JIK7ZZ39mxUquFdAylJxbMt8PrYwa32dNbxEztGo7bxOxfiVeu2sUAtdeudtis7JYev
6tH82kxJnS0NNGXctzPVHMd4O5gRoWi+cIk5gLkfIDvYLZK2MDcxgBXn6nkSlg6RPikdYzxgWss9
wNk4YQVGqRH9fhWE0A8Z8X6W5TC5ZNO+/R8ZiVQ+RrAxCHUGlRbPZb1csleN3GBTpozU7KIsJ0OK
B8GT7K9PpENSZL/xDSonzZzppTPR4ai3Oup7uhw2C3wQX/wGVHXuRZmpepXM/OkaZYkY2ALQJxnz
NjOB9tVBBvOS5oMCpHkq1KTojAwu4A/rn9E0R09Jl+95f+IwcvrYyLT9FffSmYFOYmHT3zJG/qiN
njTJb+dxsikD1K1H/LoNGLZiSf9oizbmpjhp4lY1AJCPU3QCQIGl8FgEAZbUlLrkdKXMqPjpKjj5
sdK77Ag1NdSpMnaqnUEf1BBJUxcz6NmIlk5j+zheu9xlOk6pX8W9J61MpDB3zdyNnGlffUb+bOAt
MY3EUkalGWiwEDoz4P3OKdJuL+LJiLv89nv0EqE+u83rlmn9MkZegUiia3isXjKLb0sNU7+mYkFv
fJ1S+2bHYbGV3r3i0wv1AOTRP+o7GzPsRIukjV79q66W/q5vH6hNDkPuawFeYFGsm3qZaxKnTOkG
y2PuNFd7oSWWq6QqP9QBySB0tKxSZu7H5KY+M9coEGU3x9VKJ9A8NtWnWGzdFv1R0a3QYmfxP0nX
w+SXh/HbchHGz5pf5ZQyhpKXxD7CrMINplB0uDUE5gL8e1e4BhU5yJQWgYIxrgCDjP1loR8FhERV
7gDnmj67qUKu+xCVm6ajBY4pTC9hS1J4hJ0KQ/g21yVqLVv8+vbfCiG1h0DjmVrZLk9PwTSs+sOL
NCf5k88RhHCmMyuzx3xecr+pfBxklHVtj2IfyOWzWMwYGtJ5Xt272KwauTs6VQYI+1EccNeXIfm5
bBFcqdg5ExDV4/foiCBSd6k7OmtBUofP0pEWSplr+afH8sqT7lRv01spAMungNaDhTzU0Fs7sSrf
eAQ2pW2+0cVciWPjAGqk75bVtX9kj0n/mbls8lnRS06b7qgZaWUGSijPZgV5NKHncjEXesyToDXE
CDMzi7m6qpPQNxWxa+wTBT+6ARJNRy5pdQGe00QRcYK/JiLtEVAxe1GfjQ2jNcL2tCv5wgGn+teN
tseyU984507LRGOsBBvo7X3y9pK3Gl3lVfrz/gcLBDLYQ5OI2eAiqI7KZVby35B9u2TOkHyd4adL
CDCzQaQE9wS9Ot+xvgB6HSmpkIKwz1gHPwivjggUiMPmBh9ZXwrqRjpxyJLzLp5b0YgrXqWaleD5
aEMGl2v5RD1/edon94dQ8+Eg0Ack5yTv4WVb6ijsjZi22GEKfLsaE0DHIe4onYB2P/n5fzPLa4xl
y0dqWXlZlssnrMzXSzRK3XlHAk/qujwtOnorpByz03jfdewZotnONi6Cu9SJMxHwUNjpp2VxXLIn
xwQQrxb/iRlRX5rjNateJRdcd5zgHe1evHe9U8Zpzr4q+5GL02M7B0I0wyckBsuN5mEQhNy5RLyL
4tvXKKzGKims+r6SZD/MwgtQwHdhPkdkstKzbBMMBTbJ2LZIueSudMcCsPh9YXAQeyaitEXzWk1K
Z/829/qxo4B2GRcMDC5HdSy5Fxu8TajjelRnSZeWRh5g8A8PbX7El/39mNyJna7ptXv1+5b9OpKM
hSPeAK0z+4+W3DVQ8YLgszZ84yvB+rfRLIyYg4X52GOYTQWk3aXESD93eHWrgv60m3DKZgkNQ5WY
nfFLnfGo5FlADROc/AK2chDldNoNVJaFsZF+QrnkjsKxPfNJiVdK7XDTeIzU9NswH5r0o0hrYojz
SCxNJQtX7ciR8vadGZDewAVvIhvnb/FZ/qEko8K00dA4X+OdFDvYppdcRmpLjUq/6yMU05UGFdvY
BJACW6e3/7d5TIVU6Mut46lYvrwys5tLfgx+HSMdPloQlEtVWe2DfW4QdcahflXslS7vt1y6gIdd
G9vq1FJvagT14aA+F0cYCxyJKBVH2YsgdxCXVzWohpQTyZLSXV2OS8REbzh83VX6h0q/9TBssvMX
eqbxo3PezelAU3GjYflh15Uqqav/4W+G7StPgwenUeDFE9KDlPxaTO/s10N4XGAj2fYRDC2P6nz7
Hga2uIqzUz4jl3DAeAp7LaxAyaTCVOAcTe6JM3g2OmAxBaaWekXw+3a15Vy52bI1QppzJ7IJHlD1
tlmIKEf3+8g6abRivPUD2XNnzFQxL0EuOM0ePvYG0li9mgwGSP/cqbR6P7eVpJ6GjQu4ASR0Xv3R
rRy3LxrNyXfDiGQY/WQwWpnEp83XQbGjrsggTp+8JK99zwGT8J+c529IuHFpJx7te/QkdHlJSvkB
nHvrmnligK5bdyJHyWaGMEF9gyNDJ9Iuq8bFaYKQm/2WADpFDxaqqDm3YyqutT8yvNOWe5H9X/bl
pyv55OCa6AZGFppux2LtRd0eoyKPRWmDkk82pSYRxS8cVXQ1Y51OexNEXLL9F1vWosMwVX8+9UqG
mBR8YKu/TjPWDfpwGlCt7+nG3FF0I8aWm+2ZlSGJFGvM9lnqFk3r08fTQ0BhOk/SU5RdYe6wthQn
Xah7/ZxjajYmOL1veOCLeb5vFaZM1qZjMS3VPIJgb1ZF9HGlRdKAFBxwtNGXEFwQYlSVeWHv0bNj
h5nq6+d6V0lS9bk6YDvm9AUVPMsar/8jnxCi6DzLS5kWOozbXIlfcMMegybCE+NFBoQgfu710xbh
ZEr1zrY1cYFLpPc6vSdEB0gUldRRzCYiHPiCFkzGYvgjCgBQwl9f1AF/kCLeRtJGQgDjnUUtJBrN
BN6llwDi3NO/cPMTpb4bR1TUfdFXTp6cP2A486pW0/veiCJ0MTdL/V7WZqsSN8Q2Qc0ULn+EtML7
RmiO4UhytoOvccRHzRQsBbWEPUeh0zHIB61BpViJhpHN7SzRt5BNKNiekcQTUS6WCl8jGgduRKl2
Fd1D8vvhYrThgBkbmjyXYWVGcPGZ1999bo8v2SOwV/mhwcXoVkNn4hg0FUXcoW6A2WfuoZpgdypo
Qp3T3npz2QLHApIzbZM2sKqjoGIHgzpJMc9rwL+FidEH9YM5mSjpzgEqR64kioAOWKPQoVSdPYDm
grBsi9mHQATl6AXNFDSvZaciNipCqc7SFnov6MLQqpCFPHTYG0xTLg/Mgl3lpov7T4W2oywaXe4+
+FnoQ0W/WFQQbe7PpMMr/T/a0eSxir2CtnswWn47yEp2FRpE7gbvNjUECksmmVfalpv2aRBuTbAi
ferYsY4Kpq65pUtX1RaiI01RnKq/HarcuW63P4IX2j5wJ9TFgcgj8o6xtoypP2u9Tu/s8JTEoFwO
GTgBTt6iGHYoC4wzI+ArXlg7/98exsxPozb0qu9GTHuP+33JcbjvYNUIm6MSuCMBSUXVQU7PpC95
H3IymMY15cTrj+DnS5zrALpvuSC+z7xrod9SI2Ety6fkS0ELjEP5pxe4NAWVhgKEUwTiKrSz7VQm
FSr8Hei3YohJZw4JQG7I1Hj91IiXtindnE7dQIYedlDUr/X+TcW4FrOJbdo/vbxlXNZs/+ODSt+O
g75+fprDrpGW2G5BwdNz69aYUGtIKBIVRVdmzd6dUzBQ2pmu6A+06SemVRiSJqsKaKZ7y7ka/+K2
aXPp9VzOOzgf9WN29X20GHs/NWqtIZ9oAmUDV8iv1JBe2K3AOXNwIUw9v9GsWjZAssgosh9NqE4w
q1f4hVX1T6TkbaQfYdPe+zYyAb7sa9BqsJCu1QSCsFXEhknuz6AUkSK5CV0PSTkgQQQDOeNvEzr4
ZCfEn/GDDxE1+Wz1ngWtIxTX8wUUW30X/cLYKiWzfLrczy0O3E/zefIOiWcFSpxsPJ8qXxNtGoQ5
vpzyIZzU1ErF4qxOoxgTuFoIWQJ1Lktmq4BJ/Q3lwPJpdWZP53Nyahb7V15BtQX/Ysn88SjS/GhV
Bbw6U6rltEE6clWt0oS2X6CBoEiu3JZUo0m2UvVB+XO9CGuqFoVidjybQ2reBJM6P+Wk1SqyoSob
myFNBuy2IHmVLjvMuA0La17cETuZi/to+ij165bn7PVLAyN2fN8xwz0MoyUnpaT7by4ZSwL7H7fS
ntiqnShcDH/8lp37t4eFDAIH3eM4OzoPrCq6OjkU2Z/tAS5t0hb7TZw8IoNCEjD3tiRxpX/Io6NC
diq4evfUlat+S7RueWAWf56Hw8RPWUbJ0MHPMlY9PuJDQ9RhgDmOHCY1fkqq2mxV3/+MfkioHFnb
eGBJYNhLoSUuc6NsbwHgDWI4rbTtKaPaTPYSt1ose3KzsSgxlicNeTRrG+zLSuOv9OuPGjEN9TD/
TF7LBoimVBKJsu/5fYPwxDfLK7a7oGflNL/5K47/bR6ZR5vBwDIcBa27vkeYX7I5IBzED9CZ9Ydq
uLZLkmDnROU0wU4aA1+RAbpxufMRZ5AcgeGoK0JSIvOwz8FAL2fzGETQbQthloFkkskG4LYbAi/l
cv9bySaCuB9jnJiaPYYJlc4zObxSf6xTCIX9xdfniN9SZHtJTJ/coHezVb6x0+lM2I/IqfXTVEae
GKJR//FoXo/rx5yiktVVhh5JHkbfMt3bMIKZJYOiEY35DP7vksteaeTryOj+2EYG2FMweeXnHSuq
1CTeYOG8SF5PIKxREbNY25FPLmGGQsaElG7+IQOlgGts4QDNm69Dp6blBd/C0oqIMnqf30d6+Scl
0oCa0zDhC9/+ahEsNPNaMKn/eoV1XkTq+nQrsOD1dp62NTEShPdXhgaMbjA+wbExA6atzXDPaCJC
JegC2ntweagI8yxcBML37jq+eJj3ENIH0IqsxBoUyMbZkWqThsSpPvNi1eylyRT9aZUM8aMcXz84
OUHynNzwlaiNHlvs064uJUgI0Jw3mmoJyynF+UAqGlbz/OtIz291yitwaBrqCoApIrSVlvTa2Z0n
GbemUNkTy2+4AnCjmuMweCEFSDwnUMpQj5LOvJRjQXCdNw3FBv1Tnj2PFgDh5i6YxC0BPtkHbHnc
165QlP3uLijKlqR6nTMbzMh+A0JjaNM6B4p6YNvekbk1pGT/Ft5HiRkbzp+rjzStXw/U9RNJYb0p
X85tPmPdkfwodWQjB/BlKeE39rdIOo13KpjdmppjeKA8pBqHkG8pSMgdmQxTIhYCxOEU4Lm5uOt2
kTsNYBS0OwUfO0W+Y3iSbgi2YHBPyy/v7w07oTY9cWQIBXXjZHne1+Y1nhDWAIa53S2o4VxrdxKZ
uQMew7OF8ZpQdKW9yyyidhJr+VfxOa66h7CgmrWO/L0Xl4syb88ZoZeuv2AajUjws76HWglNwT6Q
amNCFkUW95VHBEBnrAOygrXK8OpMa3MXHWwQO+SCY+WsymLWVIJuCNr79DUhb5MG55dX84BIlrq0
4bNhKqeDSQXlmSkASfFL68L1qvTlBFosBCHW+5D/nZ5WL0Ib+/PoyyNRITri9wVMhsZQAFnFbdO8
KZPErHBXlpwiQdjBGZHuAHqqScoJSeFdKgxZ1nOIB82SjK/KDzBjGBSYOxYlCnf9XuxhaTKp4c/E
pgI06cczZsaf8AqXpO3zkngy/jBNolCctghNJcsCTbIq09TZoW1GVgdQFh2B4cYsP7Nkmmn15yW8
80iKYvXxvW+XwtrgnAagO8+ERy4spy+KUUTirKWuK+eGV+cYpADgTBKUJXz0ysY7G1cqnjV9VjLw
ADy/laUXGa0atDbrZ6nPG4/2oUIkLEZOv19W2H6yTpwJarM+py6+hPJ1dr+XtFTIRwXzK2ra52Rc
DMkDFfk/8wUh7BoOJMhhWqygZLjiGZICbtxk4sYBXcCVRwcoDPapFPQ+y3pD20EOm8dpxy9JS/UF
FX9HdyxfUbniQYYuwXbcJM87z3uuqLQIuEmltWmX+Lz4VGOJWC6CA1VdjwGsiCDtjFru7bOoilJQ
Eb6Dx5MRyOFdkm+PFg05OmNm+FlbxkG01RwlnRk7f7Lz8h66Kn8+afFUJYFTqk4VHEKFBP/2mU0L
vRW9nyXOencS/pqos8S3+ggtMgjDVgbOAMeyaK75+J4Nj87+68eZGLceGCDIdjO0EipwK46M5lts
WxIe8AGJwZnHpA7UW5q443pUWiYpK2+YWdyPiDPjyQZ3T2BJHtlIRO/dAZu39R8kNiEQOwcjbZ5k
0HG+d82OuT9eV65NuVu38APXFeO5DtOGgotF1BX53esp6SfB4tnQpvhEvigXC8y/dwIu6CuTZQkD
Ogg63wrt+Spo1y6FxREDV7dVWZ8RZGgts1UNHmkElnQA27DQSUOZu9byVa+TOMU3yg/PfF28Czzy
VahanEjUt6eMmVKQSxq5zDNW3Sr+Yy1g0/HsLZHwaIR0ZnQswaCtXUl4/LZH3UsE7qLYQdepk0a8
o0mhvGmc1CI1JL88YrC0kOPnXSs6zS6GYQsYadVQDVVTSdoRGkSO2lmSSmH6RLjXvfuhy5bkx0nZ
OlT+JZpT3kwJpbHyZtdzZDXcgOP2wozhd07QEBgEvR4UQwHKqJxkN0iy3GcbAVlATHQawG10KMnv
jq6Xa0Ox8+Dv0eDqlUsLrAz04MV7KT5gnYeXGs6HBxLHsNkGwi22wm64IoPkV2PfCKi/IuqKpGIF
VpmbZzHiU8ufCy+qLcriKIt/tmf8MJ4WL29KWTkMxw5NIHdnnuvy1hLwczJjm16lJyobXjFfo2+m
7lcMHJrTGYblhQPm6OFrMMfkslftKcK2ozo/POTdMZU/2P8/9nkZs+pOyjdMW3pdlkUwWuFU4yNb
+2sUP+rcQ6dD0EtoIdMhP/61M8AQ5P7m57EwdOI/FVsJ4prUFbmaZXVj6eyQibU0lTl2MiyhCSe8
ap9sJEwPT4oJGJjlsMlwIfbHc5BESLrRrYUQmRiGdk8fY1mBukqSm+07TJmp0RCJ9EbVUhYELoCw
vy0BUOhJ1/Rqh/YP7hawo0kdlHf8u4brukGvYceV4I9FiowR/EqO2aeFFw6t9wXpkeRgS3pCo2KA
yqcgT13VB6LCQ5MU2DCXXhOcjM5ImGfSuOYVhcmYHXkKhXX6tKKzKxzgaonS5gaRcgiEjukZsNOi
HXN2TtebUsQPhHb6peKutVrYp+Ycs6adTeg4RUOOUG5uo40RPj9l25gwCkofF7mhpeTmBWBmskvI
xUzlm1hcbxGSHKdER+LQR1uDqYWA7oVJsnZ/kaPl5hprex4wtNr0x0r9YJSNjM64uJFBJjalptNP
KbnoR7ke5hrg5Jc5if6eXwD68tN2fjlzJKsGkIcL2ySJYUXTxM4JmWp2SjxYQPuxKBYpBRFythOx
nuxoJoK3ixeSBSCwRBPzmAtsVBnD7K3A/VunWG5DlbWeDZufz2Hs5mWvifBjr7TGd5zlR+IGpCzi
g2saWNN4wu5Tj3Fbs8tKXrVxwypOROLTrdKo3EElRv1MtKodFlnOK396l0A675Jj7L27wVBnBK2V
3nwmrA1zDH6HviVUuff/TTG6h+CkSnUPZRCwPOxJUFbFo1ebRDY+KPW1p/w8zDtNlLdM/L9xbkbQ
yClEblYWlvNJJtcJWAuUOL0khodW2oWvfMG/Kmuoq5PkkMkBnA8CrrL+GKb8HOJTEEAobNLRECFG
WLLjryDpSsaZ75d38bIOTKbJfPN2qM5eEQRH9MyGnrpcc8T/mwBXKN5p0b5AW2k0j76owYdR4QG/
h+b7oxwxFwt7WVMO9HehQG6Py0IHEbyc6D/F1qx9rp38mwegVAJsKhbFcRHSANMlnQA/WOT0ysqv
NphxtVBCBzgam5aTJXX9uRlsyzW6Qq+PQVY7gbAJUfFj6KYWugEs98dHsELceeE3cmYL9X9IDP4G
aLZfcyTwTFrV7Wy2U3pZuSZ/Jh6teoZJnMaw7l89FQYG5druQnLNTaMWXU9cnSaiyvOkZhSknflE
J5o84h7agBkPkyRQ2JbWH5iVky+1GG6aQTS9ctAtIlhG4lil38pAvWw8Cz8qjBdaQh4xrKhuWvjE
SF776m2p5qyUjspqVKjp/EyXcMSQDPhSOF1sWHldT/sVw/NxEDE4udYgATUv89kw7Oti4CXeLrEC
TdsDOuPkREr7GnKjV6P2MV+gsm4fdKq/okxLxFJBI07/Y9K6DOV7QkM4cPm/ZtrShmAqyv6kOshg
OSJI1xZoAlI1Q8/71q44lccJaMtD810Dm276GjibOBhRIgZo4idARP8G1hO8Gge4jaZ3rHD8Da7Q
RbBmLEJVJR7heYlfL+KhVfhEN8m2UzR4tcxQSSM6kBfKmQKbQTzZr75UH4NHtyfZzZAhh2rYFtqP
eT8amd3Yeh8QF8DABk1+w/E0Stx+RHypVmQeJEIlUV+zUL/g5LlkwAjb42+QV6pNsnwoeMMSGMdl
TRD5LKDEkXIx99bZ8n8CcnazeO/17YPcS0OZ0pk0kYq3pdDyBzvmhteBlIHJRF5gjaz8E4DgxTcv
9tM7JjxUJ0/OSMLNLfhtmexkHV9hKm48RMLaOrbB93FMDw1zdu6x+aDB8nlyhrZ11g0Vg4VTv9d8
iEzRJFO6xkcsziE7B8WrAW3sucmINW38o+zem7kY2wEE8IpfcW50l7oooc9zau9d5YUvdvgWUmqk
GidhEll6QiOIIMQm8iO6kgoDVi/lVCaKPsRPxwb4yT7f2FJMCpV6YVXiFOd/uLVyE50+rd12J9Ei
ZgJM3utAVuIhFsx3IEwXe6GDfpHIoJNzoRym25GcMhqknVZxKeOHzZIqztO1A4DDwhWgMQIAWLei
RsZgYQcpYIsFBC/24Fiy5hJA2qkYaCeSAtQ+Rc3GqzCfBcTFIICj23V0uhlOiDWZeErs3+Qo8EOm
qfMOwSXrdi1dubTEJGvpyLuIwjyZ1c3MgQnraNp7ncV3fu04f3B614PKxB4gQDaauwvKOIDhu3ro
pBR0JkFLHNzuj9yn9F9rcRoe07wvi5wMxwaS4p1FJgTKQWF0g2gH3k61FTPqtWpu6eRDFc9ZbMyp
jCIhtydQy4PciC3bPLSse1mqAQLQ6bECnv2ZYv2Bh3Ze/I2xrT/Dhwt2991bPnixQpUPJ6BA5UxU
0tXV9k+j0cbivSkMaj6krV8Ej0ILqnKYeeJZYdhAlkDo/XVWg/SlO6Tc8oat3hmzAMT/ukXAAVKg
eBXfLLqn/SW3i+dWROASqPTBEBDLqE+v6qnGRGWSEZ5bva4zZEedNoR39Nt06yluYmhXE44ZIa3d
RnF7PWr7Rr+woVr9/E78968Fu+DNQpWla+15vcEIR/zVcs1lZojOJQz83dG+TH3YBs7u9njqzVFh
K3owDBiagFP2YXyWLvFeVN4dKz0B4ZOOJ2lZcMOWOaQtud/s1IwktA8TxVQZrZWtg6reBBaIWFQs
IEy0rrXGYsKkmGxmvsrQDYJoex8RSDGgt/+Vspkgucc5MUkfHrMGvDPWOAKhy9DJ4M6/IZ0gynrX
dLRFVwvZhsn3LLUxFf1o5bSEGYBkj/nSFP07expIyRcCxjB1ZYhkA8IMHUpcvXmmSpX1WK3zB4UE
2/D52ZWb1VgWTw6oAGtgeQQ3YzbSWpHiy3RDtWY17HHemyF74zYD9QvvEiOsMQQevWBRQbiJZBz2
ftG/I0sK26JIZEBhhyJZfnziNueodooxemxfoL+AC39yt7uu3PJxwcoGIpYJF9qyeXGsM8XoBHXx
fcEIDhurrwPiBFV7gfqWPVkMYm4tlrvvEo6KbUdvTBBIYkWXQlmgjkWXbwsnognyJzfKvj8weoNS
hnyQNWw260u8KEkv03xs3aiBYxEWKn4EcZwEM/HLJLBqwtmxJjeZEe6iWxXDqKP5ZGdPN98tnD87
GjJLIQZiRpmK3URXWMPUlFlL44vmMm0JIglZRQIaoWFS/i1qulgX/RgTmO/n5rDFYmlkzhehbCtq
9U7GuT5Tm/D/rZ4/WZ8ON3OgliKYPO0ttUNFJ2wJtQo+g9lsu93I0b+og0EJQ3Q1MbBS99ujUfaX
4DZ5pXwSacjUkEUyo1J+pXn0FG9FcF56h1XkUAHUePtd6RNcB+iIDNTAwmSp0I4EVZN1centrtuU
6dX6InMhkd+jrKSlnMOK+pzjBeVGB/YE2y2LUoxSY5WoZai6tWmJO9uuYRMlKDrZvbzTrtUsYr4o
JnZLnWAr7d+KvlQ2lt0AKqk0BuJVSO151VSt73qpAuGZzkJ4mo4VMnk6gbDLm3svAO8uCxj2NLLS
G+mXej4u6uJ68I3Pb3Z2Qj2YWoXClVg8KNT5fo66o1m7kLOj7r0ko3Od1TNiTZTFJyD5mdWoytUG
L48wwMqLQ+ZyFXKoE8YCUy65dqs1VTHFy23E/Tgb17rhHCgbb+XwsFaMvdIMwTeAhLe+OSScpbi7
uDmcBkYo/TpUbcgVVvvhvs2JNBWYnpG37gTQYcbNRhtBgxIKuQINmgAuRw7OuBv51DwWtyyQMJp1
h0MNAPFFnCjqBcvCa1V03JOg9Igp4+Qq7P2gJbLJCwrXZ0x9jSCGdyslVIOv+VeTSyBFlJjLy886
4R6v2lxiuG6zwl3rE88vMAM9huEfVxmR/h93QODeQRvH7OOfP9FF9/AptmBMvcpT2vdkHLJEELsy
10wCqnJ+EUo2VDvclEt9mJV+IwF4Od2wVMkYNHeHXKj6jnXExhQmn58ZEKqq1RRkTfAVqSO0M+xl
hb43qQ9DahOKhkHBkFEiIHfGnypZNCFQ0mPg2jP/y9UUy7Ne3GzVHa3wYsopPR6TkK3iYD+LapIG
NAu4cMN5HY2qWEhjQI4k1W1Ho0GLJRC4IE+bHbew2ie3sQ6FzMAWUK5eIN7m4mx2+x+FlEwci+jv
tgBlVyU03nn70dIaYksJYON/AylEeBxOadILR+8741ygLIyuCsOFiMP7RJKJxfsrq928OiSxXOfO
rsJBFvHRmXcKe6cebrw6rFJjpJMzKcvJPQ/K+Ua/SqDRvOv87QsxLWE7eAjZKLiCa2Z8+loy1BYU
C8rKof90jXqHrUFggDtk8OLnY4jX3kt+fh/5CTP99HRub1q48mQmtoPM/U3l2SGy7Md5IJoOtmYX
X1Crsx+Ohs0n8remHiRQDSMStXusVGf2WPpte2APVt7auUxu39aYNm44kx9BwnxG7AYFuOAzU6je
pblrI0gHV9sb6KVimbbfece+DzX7oTmiwEiog2FzVz2SpJI2ghs8moZax13Buhi22wO0w1dTcTak
qCYJNl2uXBm2NNOsmxcsEzQ5CTsPv6oPjyCK/JjZ1TJ5zk9tFJaULbpP3C5V0jofd38K59srLmJo
Dcmhzys88X5Vf/wHOiZvjdIzPjo6EWPNl7ia7YevoGwJ97VnLRujGqYIrtWOVPXCjZ53itInRTC8
TK4dOVJ3ELEgs1ZSTGkXDAGdg6UBEN8NRxKvWZp3eHx3OXfspKxWHEvkeT4rMyU+S08cLwDQQIBn
5F/ygLmXBAFVtkU7BNzMmWgO/Wj4K+XamgXqCXzQpoABRKNagX7WYXbyJ6e3ZL4jkMhJsIAY/pA+
N4W5gIHqQ2fGlAdvZcVDiKwGUJ08EGuT+slstTI9IH8Vb2it4aSWZYcNoh7gznlvNDBkRuZL/Yf/
Ko4+aTfYiT2DGUciXPrKbt+nEwEQnqs7AY4HMSH2o+qGHskAfXFovOG6wQL3A0N2L2aEw/p1rsrB
nGKj+mth+HcJ1IwBhiINBx5SGuTsBFJ1V6Y1tK4jC3IrIHiIp3ojTq1paZHN7WwlUhNRKb3ggnIg
waOOIP7vkpP41w1U+dWX4fAM5sD5ZrMRg4ftDTdZs902yLt+CPP1zeNbjiMGjSUwFq3AC+gJeqx0
h2AbduPsCjoA1KMNDGCZWMlutsS0PgGWqwkOTyorOB+y5Lseka8NYMbRJb92/9XBoCVDr/5uzznQ
enOvNrX1XtuTTTUyy6yLBsbNLriboUZJh/wBjbDcO+RUtB1MV6+plswGAgR1bI8nn/DJXfHATlJ0
YxRacC7gqLX58aXmawfX9lhXrgkjLT71hOldDnM9fHwuu5+nWYyUQmmwEj/odqdD/38LPLuFXrfZ
oLRzBGFwWJ4/3CZchXZ07AI3PVRfoNBtPkkKT1BhHfGKDeNfXcKzFmHOdJGY6hg9ZbRfePhpXBqi
tmyB0pGJuGGt/gDgSI6IiysFYu3xwEOKZ9I7Rjfkzua3Ea8/gWRJu8s7Bo40uTFg3pwto9VYwurS
zQAqLVVImI1x4AuaIYs8Cn8Uab7JGPDT5vA9OOsde7SQGVjWJ5LjGPIWJBsh5/b+Jdt307m3GyE5
OemYBsuibgw7QLu2i0BqypWuNeaHik4/sAlmafQ5XeXZtUEjEskOX/xAD+R5mhKcaXb5ZjoX7P6P
Q7P5k0WWCEhfY02Otc8P73r36TA7/mu8Gzrz7Lh8TAndWo/VyhPoSSPgEzcxj34yUI8Vw/ithaAe
N6WnrTQeHOMRJJayQhm0k0oPaZ9wef/STWc/yvVIkzOv+YtJwD5KuaN45bhINnYDEysiZORHB37q
kMMysv+bfxYGHV/soyfK+Aj1hhryWQyDfTlS7vo8Oj4gylT4bNMcG9+GJpmlTwUkhSx3bZ/j0h36
UePFuDT8SXxUk8cv0EqRuU4q3ld0h/PnIT7+gkbKwTQAR68eJD5QE3uM5l8dFaG3ud7hZZhiTghE
UNEDb2/88uH0OgUixy4hZ9a/8ufgFOsiq3Tl1xFjkwc2IbpeF7dV273KpdWzvRIzsu4AcYYnBelD
C4DTcqhU1CXukxRTXotYoFOIbpuodXJGI04LBEyEIg0++ICiOuFun2nbQcGKMpxMl3qh3a0KkuWm
0UomhuMrCq93btAeNbj0uEh2VC7DA9krAJnvUJn2KXoZ/dhPrBsYtNME1EP3KxYRzfHlldbZan91
1orIvsEX2V1eNfL7dX+1qE4XYshYYkah5gZr/76YS9KbGrgS5B1yLe676QtzNsic+0pNRNhY2J0i
zP//e9wh8wjzcRGizTshi1RA+zXlYO+S/Szkbr89JzsmNxf934D0daH1MthBwQlCvahW42Ym6ATV
dP+C8pg/qVL6OW13K5aN+7AX4RM7TT6EMo5lWFMDS0wPegBS+jRLlG37fN/BlZkqgNF9H/V9yUg2
S/FfmbxuIM7zMKQ6r2u799C78jZHCKVtN8YbetNi35irtvVjzW26/j/wFk6Opq4yImh3KRbuyEi7
3XGf15RYGFMpsQI64tlS6qgPG/B6yQLwuX4j1eR5jHTK+la7/cLlLTHwtUE/+TwBn5rcKsAlcXs7
zQoNe6YbkwRgrNMVhDxqPOgE9MNKUSZGZMFEuR0xnwwt9lbOTpq/oJaM987XVo0KHVUdnFVZAWEc
8CXUg8L5ebTSY9uflov5Bl6obwwmq5OldkIJCa6qJJt3UbcOoehwZS7ffyNMe//PaXLmQB9Eq2UF
YgsTzp7VLOhTTvJTd93/FP+1p5RG4I2J/ktPBLsLvrvuATdsVxu8PlTcvtFBhY17bigI1TH1nX5t
NThQMo5lyX6n4Ap6kU7MfJ/Z823lwcPzXpc0pMF1kJ/LBK+OcKeFodQlPw1YcQKGNLFOB7wEJQqi
oKThXcrfo0a+9X+DgwnH+nxUI3DtMmZ0uL8sBojTQbDY99acQwQSVWtSXK3OtfnXj9jQCdn7aTuh
VMZvzFDKLoU4nn1t5Gqy3cNwEvtyUpVXCbO6224w7Dw0xuuk4z68AvKdPb47aZwX5iWm3tJ74WHz
uY4NOS1etCOHKUcBZ71HcwaROaoQRjChA9v7wE+Z63CHR0hHjEvMTdXaesw713d8HWVNPeUdJj6r
giz+z0MPmjlF6XWyFMIH07Y3XS3wdMszonnXc/0hDV/StETP1Nm88JqM+8jX3bpH4ouZ4jMJa0Mk
xF41nxejfbWYkypyfg6XJPbhQRhVQ1X4N+RxgwLbU9paYVp1O7vgqz3viojkZD1jx/IwEcmFHn/g
vOxXYYxX0DC19sIchH0EeHXmiOhT7vg4g0QY9EQ2cW5/ji2sTHKgSt7XMj/guSm7QHAcQ2KiM0tl
kBcs5IKDKmgRxXEhqMRzzAA5TfO1BbZDKdmT0yUO+UNFeevYSupbhFL8b5XhwywNRwajRsNvS22R
oxqE4iLJ7foroTgLM7ro0COkj5lqxWy9XPiTgNZfNKQ6FOc8mXfYrAjwTDgsBg4z/md+KqklJQz1
eyzF1/piy7kSLky/l+UQ5Qfz8ecKwCI+QqSucFZYsz3zZnwDIK/SNJrHzaoaNDCt+Edk1hzOA8gs
/c6St91Vtmlezn9xsOZzPPWvptXzBEktMXn8c40nI0Eyc92v7h+8nVj83KVXqrzEAemJST4YaQ5a
5n5hOxRtn5rr/7cYn/8yXw+1FnfOBnU3KO8r4LYEZRZma+txbAbqZS12HQpHyN1aUwAo8faVQZwa
x6nyit8apokH4BnWL25OO1UMqvJBBE/kQyUQMjCrsZm/iP5MrqIjFCBcEnmN53yuknQ7OpTtIQ1D
3ogib+g7iTsfWiKXVMCxXtT1XqonQ4M9xW5qNlxIKBJLlm+tbBCxXfDD5RQ8fn7kQ35xh855s+FO
JrYIgGhqF/ReG8AHqatnR9+EziMJyq6JcFQd094xt/F/tnhE0jn5QBXPifP+XSF6ICmteHRzo4PR
AhjlpUuZ0OUsCwm/FO+JXJhqARrQ9uNa2jmFqpXpWx7rPe8DVzi3oJ/7YQSlGfmStBOLu0wku847
7TGWZdzafczfrZnw500J27doHOLaeKoXu9jXyhzjL2iqdWqR0/rvCUqEvGul87C1wWjtC7PsMWUI
vzEGJZRZnSE9B3tcQcGiAMvU8xQY/Ab1T9Qpbs+LaCNxUBATbCrNZX6g3Vs3jpC1yca7IMmS/rg5
3pwr2ljl11c9UeyN6CXvOcRbqNd45XHXfe+mKCjlEvzFAW/gl0fFNpP27Zg0eKFMY46zTCqFCd2K
teMtJ/gB7N2xD3FO1wAHt0CE7GdkZTcWEThcSg1ONqHBPT87xzzCga93aWgVL1eT8Nq35Rwe9KY/
jAxZZDEb8qEjRF+4lBfx0KAX5fMC7RObmDtkOogBjl1Jzv4Dc/nC7NCJJIEkDG0KdguiLoGv0p6R
Seg4mEM1RvX0BA+GZMLBRoJih1qqdqlTD0zracffsZRtTeVCi+K6cXABnXxWxTn+FnO1LN3xSu2Q
YkLxyS+toVOgd8DAM353s0tdb60ECK/GN+OfNi+MlUtZrAeeRL7Kf9kDMYLZGvvAGbhNVKpCjk/V
SFwSc0ZR7lYOWiiscgVq7A9t6AxdHbfTjF3ZtgoptS8qrGTXwnjDIW+cBDKPp6O+/Fk44mSWhpkk
GYLmw2uBdIWx3jh06gRpThswLte5unRCuRbtEa0UF/BP5Te8b/2Wb/GZdAsHkKfrvTmZVqXDwpa4
qe+kiTWYU142omGByVF6vZZUZwSol7TNPuDzUoh23o6nriOZMCQ517EgHcwLv+1pu3fTojzBL1r1
tMC3s501qZfq8IJpuOcYUX/dZEODUVRAreRCL2/G240TM6JuWQ+ZmdKPBVUZLjbtIpn4o1ZqQ6XB
01U1ogNCpe8oAaT9IFbCqEwqhBPWCycqvS/t+/x+vEV2P2fH6+MWbG/j0whKH4quvK1Gkw5WrBK1
8+GJ31OrgM7VzhUG8R4N4241qDEMTHqzIeOeAsetQvMhu8MarSa5lrUFjiDlkcwr0XzWxRsDZgC+
//Bag8YvpdFmw1mUvW/6CBzI4CfylC56upIKXjCfwYGJWzyE9bO9TFtd9CA65EtZnui4nqh8hUaL
pY0T8+MyY5XU8BPMLflnwrw94c+ts/qoqZPzhG0nU+3rbBcPv+gFQmpgDGQ3AI6O8XFiUjk+C6aw
xnqVz3VWSjDbCXteHcbrvC+JH+HGVov5SB9OXFRWFgxoVAwtkCQyYA1G1zXpjnn6UOyZYQa5mfLE
fNGqtqrsfx3OTSEcFQQxu3fh9LOSjv4gE3Qs5kC1PLXvqTL7ixt/aoXboY2nPs4RDG3alkZP/cqB
P5yNzjxhYh/2NvGAmMXWOTuWeLwpIWm7JGe0Y3fgHSqxlRiGhq6JOfuHzelciLxSBcAPdEY5dRDn
6+gKhCkT1Eo1APV3PUNw0n3gpXi6EHShEKAyGH6IqK71Izq4xJpqqKRTWobsVrku0hSb3rHTrxi5
eP8wmtHXiQOYeJ0DRrh1h+s9VnLMNh6RVneLk/5O4/0WiYKyx+A+xVri1+4eEXoZLGl2LT6vxRZA
ubPb9nNjAg4JonyLbRE5amvowpSEAt2M2Rd7Ug3uoCL6EWwHI0BaSKww/Vw+1mk/9LyfUav+wWeO
sw6j+0wvt5BMtoB211egSQ/NnAwbo7d7NJaTUbdb/7e4NAmvn8q+BnusXOsn6VnzZZ6wclgnI+ES
jdD5Yo/a9+x1i/k8mdsGWgxqS9v/jPL2er/tfTyxZ4Ax2RsDOKwoHsRCbmC/8StiE57XSTwlcqC4
NG2n4jha/J0ZnDUym8/uiRJKVH6I0UGe/gG3NPFyCPQff8kK+R7ZbfQiItEpQ/rR+0zFhCizJ4mp
TifnkKa1UTwqxft2vMLOx0za07KvjEyDBdnjCjg2l/EAGn56pskxLr9O639mWswFfS2t3vL0KnwW
+m6Qz9ojppwvl4R6RYS+sJK+NfQqjS2021AqSmJLefy5phNkPjxYlGyarXs9AJZSSXLt/qq+AEYx
VORjwHteJN21pd5wQvJ0g+suUiJFmK9Bk0DVYDMvW6lTgtt4e9kQI0fuE7EpyW37wDwES8IsHHss
SN2gic8f0mnAHjooEGlZGqdr+pSvBtRVcmVk76CvxSg+pBMus3pwSSeIiybWQ2n0BccHRlqq5UO1
D13hF+jD8ILgBnRT6o+z2HChBXkK3VQ3L+ooDKdNazJMhjrW4Gf29XfkfNHQgwRnFEPYHzkLCK6i
P8EZtPcX6L8NbpY1BIRIN9Hd61e9Tw6k+AKBrAHXJenGWfY2YBk4S52nZSLYmrC4/v9XovXfe3eG
Y7RiNP4HC7zHqDuUNinIQDNzpHpmh3A9pVyWrueSWMOGkDtOyRRyskwZ/vXvrhVwIVdnaSlbi0d6
K9DvtRaLnSZ8W3/Yfzzd59OMJOoK0OwaVloNMWRnzbM2wTsciuloWyvsOOKcIAqCwH+RZXNxgRqS
Ep9+C2X+XFpRTfhEV0QcKjP4Zd4uUv+4GxUGyyGrSoGJrvkKBkp7g0lV00gD7qGsmwbNKie5UKSX
Bu8bYFD2EUfmkQQEXwQObXfId99d3LtCZXHjL16We4cGs1RNp0HQP782amoFIW94ULaaVEPssrL3
SDp0KGJ7h6cSlWXZ5w8mqpDG7IP50k6Y0wiMWV/K+ThymhH8o3f6TVj0yHpBdniBFlIfrYDdk3DF
0S2LkTbg/jEBBO9c/B6wyu00O6MQsFLP8SWh/+K0DQ8RCATh1yRUE72atC4xJ5/cdcRKLFqMjcMl
WmWlqNnTmfWPlhgnJCVxiGctl6AR5oeOL5MZcjxW9NciovECAU+W/ggDPHsdo3sSLr6dB1PgEGmP
O5Dkrv75FJGyX2DzjsFIGTEhaZcmWCovPWSMa6Ult9imU+U/B3dD4A69n0Po7i8kFgAjoUWTqgre
LII2lMRRASJ8/pf98Z7JjP40J4eo3QbzcxF/GNVsYRSHOCT7CPmyWlHK8awnBea0cnmIQF2TpokR
ceIbq9W/uJRCahAkbs2hPAoGExTaLN8wPWjJBoAcoeIMVSsOa2jFroWThnVTZJg2CN7UPyW9f0xp
QOAwFC2ighBhjL2z6sYsf0SWtnRJaui4zVvs3EjYJxbmUESNYnO6mjEA3sG8pJzc4DmjBnxe7Bi9
pJXXGyTEK8rtTFOQI6dCXMZpPaz6J/oH2QkMplxVr5WMxf3iQrXpJ2pDTtE2WZxlhdu3MLD4ZDYO
3kQ9D9SgcR/lxwY9EzBCLi90pMsTy3NSwna04vACM9AD1abjOCCBc5AiXCA9qs6OnW5X8jgUGzJE
SaXL9wmhPfQnXqCZy7PRoRRih6JxbuiaQXdHgrilVKYm9qmRV+xBkntyFg5+D1l7pjUeUWmWYLr7
gyj8WA+94rCqf4rK7uQ3ey3jyNPy707twg4FJQoYXByF3jIxjYjYoDg3v0E0IToY7Y8xdk7vYC2X
nGVgT8Qog95bjBUUyfxZEF6T1Y8zhYjX5E20AV2zojIhms20dz1U7b0Uyws1W+Dq6LyxmITtOZOr
Gg0XC0OyhKJZDXz31DTGUQbpFbhJ/Y6jk2dz9yz8Infl3v8DWGwmyockt5DMEkM4iveIbPdRRuYH
JHKtpOvf59CTlIcrkATkQSTHasrtvU4dP3dZ2OSnr82x4Zeuxv7oNdFHoELto0s741myPqeMzC51
qMfr8S+ds7pwrrpiQcMdNO2G411JDquF+ljJPKPa4U6/uiw5/cfDVVwGjqmr29qY0v60kSezLFZD
nuUiW+h7nPYMuDKd5Qcgl4+pGu6rdYd8t0OMwkCY4DQ4N9mioFv/vCgWmAs9ON2f0ZUv+9/Yj8fI
A2IzhoIaqu9/Rm+HX0PgvVa23OcslNJMKRV1WXT2KiwzG0JWPNjb+WqFZekoKTJZHMDZFvi+XlhL
kL4nSYRTY2YN9LiJb/msvcaX2qOUD8BmHMp4MF8pHoRrcpthfdAptA+0n77/+q+VDo99AyxWZh+H
1Yljb3PSsvuhHCd9Ws0lPUxq0xxCuD9s/mqmSbym0VBvX8aN8dOTOoOBFD3w/3tGNwPyuD8XWr81
hsUaiuUcdgLBcZBYxU3LoZP/hBqCy3pmWUVJNo1EBs4QPZi0SIq7aN0+K6PPl+E0w8rhsTAM/V62
ZSpoX0m1YuF/yA2CYKYxv/XPOCiv3P7wKs2Xy9m7sJ5UFk/zW+SpEYKp8E/I0IuScIDfY4euhvra
hQXwaIo1vM501/5COBEsq/qrtdm6EF7ONtF6ouYjdSOZuQPa0F4zOpT+bWybgvbg0Ogiknnpho59
QZ4BX2rzvu8DitFAP6mDkMZkxdo9/dI2WQQwXJDp1PPIFRcoI7e5edQMjODiMIPwvZPw1sr6G/Pd
xrDB12uqXiy0SNXVfeXR3Yn0cH8AvIV3CkvNtgc9kbDx34EVyx3gOu9l5t5KETy/k4tKMH5Xqh40
8jIr/FAbWAFZ8eL14KBM00djYhp+zkn/jld0nNw4KQp7mCyPRX0PfO3GW1JxcaxSqqUGHR5ACiPm
e49ekrL3WT6LotEaluNrDPmtfjUeth31Pt2pUFQGH2fzknKSgQT/4KGotnHBY5qTfiGPHmV8gzwK
sqBMAKSK/xqx5EPv8XJdjcWTuUn4d55JBszV+2tvh/CDgK7juaiU/2IsTPmBpYh0XVzXpvnlqpLU
GJkyux4rKgp8U64iCPX9RQGnDoLpNStwTaNaZnaXBu0oOrKbxYY0nIhmDwcla47YRcgHlaewTmn1
/WW2/QTbTh2f7TapJQCuR2p0P3Z2ob4yRIgOG9pwvzbZZtvF+1OsKsNXIQUpLcDjck0zEDp3dLmM
OWw5jxn5JeuouW3CoPOosXF2c9xP29YQg6iablZOQcfSVz3Lx/+V7O6SHpb/CQWwVLX/R+sErOE6
2Oa6gNEE4uh/9RAetHI20Ay05ayq3fFN+ZoFmnoP9xbI0K8MaMxg8LSwIpc1FS/pXqgA0VOm3Wav
KeOzdXhCFyLK/D4RSpBlw9X7IEjJa9tOaY03se+IeRsPxxiLbgyzxsHjHFB0M4iUWxB0qU1vRlfT
NUikpqDw2dXaqCz/8kpULf4JwPZ1yfMo9LX2vKIMGa/+DdP5kb1QerZk3qcw/rxzUA9fFdo4+JbN
6dD71biKchCngfMpmGqFhZSzMXV/BATKw6Uzw+g95XP63fm8ejQUXfaxagQVCX9kq6na9nmlpp48
c17RRpLbmc8ZH/Dy3eqpluN52OdyJEEAjDVq37sMvKCBbneVrLmrlY29X7p/91q/2WXfBHvDihOc
1t/S/e7HJJVPnQm0xfYHnJO+OBpMoHsrIdLNB4Ys4erEqEoYONmuI/rNxPLKbMUnZjetJLnS2Ya3
nFu2lR+GXbPVMlQUi6EhPcQf2vq4iNKd92KUe+DSm3TxTLrRmOd+t2nap80PDauFjrS8YlPakCtZ
9CzQz09ArmDr5AHSA3X8QvvtIsr8pfNLS2mp0s7i+x3ZJRSA1r8Nm5MmVak9Jivd+z5mK0uuf+EW
0rXMdcxUVxMzp7VxkAJEzRQNyZVKOn++t+jKJQGPXfoGcTlq5kHmJB2n9PlSAslz+pJ89MS1TiRX
g5haGUh7mytNV/U96EicrJMWygmVtIiSICfy5wHcBjzGSxX+zfQ2JK0w5oa7QrKDnNsIQpIM5A9y
N/PCejy5aIDM4pDoMsPzJ7dAd91Ofw+FGUeQN3Vd2s09yak3/CwUgVpeC+ZfiWCK5p7sbVWoIywf
vgC1rq4AFiSRPqIsHCjvDXxJBQTKdQRIsGpT5NyvoPgTVeQRbeOH/Z7uyc/5+ltqpIFrcmI/NP/x
dEgydEYSevH/CU6U/36wknH0ZixGqJ4HCkwKJh3NUfzOtAgS8RUnkn4i8ImZxDh3M9+ChIjHtlWW
3PF+oQkW91GKQKGQsPh9FOmMAmb4jvcWHn89j4ckmBe/M5Ptd2sRWrMNqKp3ykFvQVpy+ByHLyyu
phlpMeXQfZyY56FszrTZhr52QJlbMSqlyEPeanO416J3SeySSeEBBOBsEDA51ryhLPzU7IMO/G/F
ejPKU04S1no82FpDgvSlSAiTypbmLMC8Y7utAoEAXX0D5isV8n5OgfoiuHbm9xoVvgkMgwWOx4Yg
m9w6zvFc1CjzbqHe4zKLOo24CwKwjCTCldQTTYlsEU9x2Oel/W3MqM5yaxLkPHm6joiza+4dXNvK
PYTRCyTaaifVO1PvJ2EMHu9qrAIQKcYPK1HUdmD6BCNSad5KQYzSM0nS59cFvHNYYdK6wA6lY6MA
fVyPZdZxEf9baQApwY6ozLp1BgjS4m9mCzzikWfP2QZphK6NLAhtN8iR3PWNd27Caotc5ackBo2v
t2ggkEFMUVxbZQZ/s2X9FUt6on6j+uDiPUeEuIv+W+Y8V5KvcT8xzgB3GbT0WFFqITm8zFh6IiVm
c4fZoPmRX+4coCPKtumZKcKMnDjCkpXCC/drUJINxIhqqGTxSui8nJddsqr2ATZStgt4ftGQEkMf
fASTvEQAXn40N8MOe7bvUp8WKla5aqukowo0oMxRV4sZ7sII7ZyZTY24LqKIp0rkVuJX469xFbX5
tQDVUaUIuYnaztoNMPmblJhILuiYIjsGXWC44aX4INNlbDBAG33miwaORXzN9DxHsVhI7Q+BNE3A
sVpJcxv9+aMU286brbz58Ifm8W5toUvERTTXINgXmuv+Bjn+pO7116Oi/TxzyK+1FyWUnjlU5V2N
r5CdsLB3wwmxghwb7E7SukA14oyrpZ4l1TMGI5K6ojj+i1FhlD2UM/dDFCzMuut1sn/QqWlDCX1M
DWRkYwHXwLIuHI1IodAvmg91wDsioDy/9TqQceD3LvRObjpcE9nyGgq70UZha2pJJxhc8RbJs9kO
Ica6Aw2WKRfjKjNIEHc/tJJWdjsXWbko5wIAImhkBeiCsQkFJ5mgLnwQAnhCiS90o72ZvZ+hEkYe
u+vXLyFYc7nt4IOZy7MeU0ZdVd7sF0chS5pEjXwdordvtNpN+7izFyDiHRYzdSeUqx1kVsgXrrJ8
f8aXKPv4UYALrTQv3QKIjPEyeDaN3IUManS1XSd6oSmZbgyH46EptNCpZJ282nmrokmu2lD5dW1h
M40vzQyYsJUDXpFhzjt4jdyBFa45UhXCNF35nWKOw2rQ3YrgMyjqrY67o0zItbx/o/wAh5u7d/rB
WQt8oZA5oWrpGlAY4AjNau25GYDVk1JYEAGFiArj9uGCInrK3F0e7QZGRhhf1s4yLhMVBSWTwHOk
1rBg2NErhlrb4/VVCbZJZyoOSaURN12LvVue71VZUQ1KphhddxnOhisgip7JCnYBe2umVIIYGMbj
1NxPdLL8Y4pYvHXv/k6VLJUs9l46kM0b28JwoaWh8rfwHC9nSEIR4TjX2jCqrxFtG9XIMmbhcgrs
40KFQ1UzLRvCTqwrYAjlgGDlAdNGD4vCTaR/MbzfVEDFCLp3AezoAYjZSk7guYG/a4CHcN62pd7/
WkZA/NSKFoBN5/lr7ZO6vFoQbHALLo6318qKUmw/A8naCc5QImPIsCPCavPiGK8bweJGb07pq7PT
J0cuw/GMsBSD1/Vkw8K4eE5NVpmDNIZ0GT8kUT/heOOvsAiiF2ANBem1pPZ9BsK5Kn0BQJju1VYN
oJ+64L7U9I/2WOVm8VSCCw/pN9PP0QJs3GS7oerAoDGiu+jcxQpDQqWUE6Cr4zV0AtX0lV81rvHa
Nzxj81oqiggxeW20xXZQ+sj+7AMG6Lqe2vDDE169BW7wLzXcQa//VHf0NoilIylyyzKYWm8pXz+S
sy8gHyfNY+uzbzwYIQqyqGlZ2XLryQF60mD8x1awe7AuSs1ZWOImMv8/Y5OIw0YZdmzE4rihfITJ
CWHP/Uxw7mHbzxcQjM+NGkn/sTWjccb3K+qkzTydCiTraTtXcGHTzj3XAxK73ciLpIskU/CFAF0b
D0REFrwPvoU925j3pePy+1/5UMiXABZy93ZV9eav+xKrb3z8vB7aXiWj4BbeG4inH08DEZMoaMeW
UMalpCS6NO5XpqiVo7MzdnAid55FE0+orIdhAfKEcwzRphw1owSPJDem0HOwzjgsLXSHT0ER5m6m
xVxSgHb988ybZUOQ4WoDyR7WIqFF1N4hzquxpKiiPQQrCXzFsk3xd8cjJgq4txt0ZGNhki529cQ/
ybtzJAFMRvS5Gj7Fc+rH3xdrQI1GZHoIy3skZaKUXDKGTFOBBWkYpbKJIVxEsZXmdEtQjDOGUWkV
7LqS56yBYzfkD/QvkbFYMd+5lFHwh0AN+aKLJOSTl3hfEaANEG0/TS/HPXZVpi/dfGVZwbhF2+iK
stUKuhOHze3ifNJfXABgwfgJXpzCbrb7gP/KvaJF3bpXBsVwC9GBvuJ/CyA/4L3ICYEnvooVlHz4
SZnfq0W1YWloFie1GcRNQsj/KqMokw57l0Dz7q5nV118dotnm3CND1+2kt2ChihmQWlOmBhnAkIY
eRfT9nds2PR3hxKLK6MvA1JlnqSTC62KDLgLkNbIC0dVNz0mvNbkHtFFVXqzI1kRp2eod1IxQFkW
oF02xg0s/+w1RWd33w5L8IYZq89gLKiAB0rIGYPTcyChmergFMO+WYlhmQBKlqSASRJlMOFFdIeZ
Uqfowag6nKtb+M3E/mo6ptlnIu31ub9H3UK0LxFDGCpdYZU1UUjZRQAkydacv1dTKvLslY8CCvno
Ulsj0LUjDVp4IeojoUN0m+MYOgiCohhx5oMiUX45z3JwZUxnplHeBesOq3OMz5JtJ+TN3LvHCrM7
trnLBhrTZ9mnz4KZmbKYIa3pZscknm44cO+bvrRZ6r35fBJCUmcuwnIQBq0lKWLUqBBdqmUDQXmf
rx0KzoDYWKStrwujkuw0BasZU6EVTFEj4kpmhyl67OOLbbRXOmNj7HS++U0YZ0dbuzU47CNt/gsy
Pz/eiP//Y1GgKDPsBAppllZyH7N0O1vH9VIViPIaCsQaWN2vTRwzjJpUyhGH2f9qCMfO17qvwGtx
dZkww7x5fnzC6WvvnbAmxshqrvOU8QIRF3kjQQ0CXSgYvbCEuy0zva61pwOZXeU0tXT8KDNPGgex
koW6BV6FTORnC7ypoMZnaT4jCDMxe8wp59IcshHjU0N3ystBX8uR761JEpiO4OsPoe3HlURQhXW/
V3HzTR77wHIH+3hB8w2XwbM60hyCstzllG3N0YFsIdRkaNCAIEAarUhIaB7omg3YPQERwgSLJWf6
Nt3/RRouvDPM2uATzDCR9BWJyyerVy3KeYSuKRw+DJfK7Y96+NcvpzQi4hI3kfNL3xQEkRVWuCJD
MKoq6pVjeFHds3yRGAQs/v9x8/owrrYmTw8GR9kkdPBSN3hgl/IBgSIp47nmZT2/6rtGGOJ3dING
oPdfAIvOKjRggyQBpLFiLr5mFFSSI8iSgkTOF+UgQYQQ4Nga0Gr+ieuVBnk02NkQUeWAHFp5kB42
SeKc1kJdMSj7Ya4SSNpH838I0rp23gWdsyciI5ZSUi8ndCBvUhgjT15P/DlXicbP9qckmVwDpIRs
Wh0/NOyMEm9M9p31jOV3+19oURAnMM0pkpCvSatC20aSwJW/bRfANj7kxTgApEaFqeGJ6GylLV0I
Deo306RVLhSZq1yI6ZZ3wCYbnielcF1iPqNztjohkgx9i9Z+qoMd8+ZENQsVlEaekQWZqRc8uJZ0
wfUgsp2B7S6cS/wIXLKjVKDRRHiI6BDWz/h3d2SR9b2clqE4AoNV7asyLplbcmyubWmKJAXhfTgP
IP0jUiPR8TaoZDUyfImjZPczbrqhlKSczBWJHLnvYVrfCq2LBNWqBS7oaf+eGgQABjCxu9oBPM4k
spRxIFFUE0XwbkZOcNhl9qxAVP+uaU/HJ8MVMjcd5NMuY5WCXUDJk94bdP7ypPRJxczyPyuMqaSj
U8VF6ewlF8Eh+yB+S0TKUfuN2yYPA0dFbnnVU2bbZJtPTOUq0aUjT/SMQLicPzF/9PHlkkfdcMpW
jibJhYOBlW+9ya1WeUxR8vzJ3tlt6NSuUV6VENuhWZhCTnMKGZih3QkBg9CF1QcI7dTTZ2FXCnWy
aG5jYp+GT7hXc7mXyuVCkd1Vh/5+36ElPf/zu6MaqjjgACNrpwv6k8f5pK0w8Ab26MgmqtL1rE2O
y2pGTMFbP3ZqnJtj5PxnbSU7tGmdHhhyTmJyEFM61rVeLjeCiFszZyjcay2s4R9r9FcrnqdOn6tK
6KrVmsMAc2uK1zuyqFUimIK8RTXT5KguY+RB5tshl77nh7CSk1k9H4OkxiaN1he4MnovnODfZMnA
KI/WZq/T9WR560DAwAMjw+qcaNZXkT7oM5BU0Cpvs0gOVA7lzrCwpPipiu2koOPxkPQw6TRCWpO4
ajvdGfSj8wLOwvZyOT6VAQpua8uwoawwUtebC54tMH5RRYPKebz5pC539rr8oR028JRC0g8BFbPj
7AwpJR3v4m0WTpyHLygoFTnInchHmH5JdIsyCpKtZOGNVEU7ACKvhovuLn5Kj2Ekyvw5lZYAKaDj
F8nCn+2TulLO5qWoqnaRtZUUSJ0aIyA30FMxE978l7YbDhQdh0UI87ePMPF0QKwlpnE4S1X7YEj+
/4yIoIwdlQMde66XbSv/DNoVTUfg6Cg9SSL7VuKIfV/e/DhBQ0oWJerlAw8E0Qg+ruQI6rs0LNi4
QD7qGjrX9vuc2p8Ymgqf3JV4IwRfqtLB/n3MLvpwqor580JVPSFxu2DwUYfkq0cWDsI1kRSOXrYA
Sk5V5zPp4PcUiKMDOHE6uzQWVQ/ZXo0dSv4nS9ZPKcWOwZ8O56iOd+0ICiwL2npiOY+smoPOyO/N
zcgrSMrZtGS16yPashN+Fo2sLsf7uP63pfLzbEUrxuMp6mO7f9yLD6OWnCTKSupYoUM3gcG+XwkB
NGB3x2A7iQDIdXaCiyxHgebInKUJVgoL1LWtAPMBcKn874rxrZtZInx2hAA4gsyZ/XoRfAFFtDy2
249a7VMbeoQQYGEdssiGXASsdKKLI3qezj8wDnyAMuXAgGJUfxL9SYbxPUECTj4gPY9awTr0wXY1
LDYd4N7+cRxGJS0evZwtMIcgqtEzqf/ElFtha5h5bUIfwBNLxDQHLpPlLMnhN5188nAeqRyjm6tj
+FeW+rofua09kVSS+K8gk+1lgr83G40nlSbQkhafrwqL0g2kFIHprqcH2SAm78RI3jtWHMp+8yzi
iWGfhiIFgsfMovZn0tp+odSQG3ENkwVirJGpSu2Ib2ZKsofMj7za6Ir3oESwHmsdEfAQn6fX7Hl8
DTucHMXDluivduo5VhU1afefznX8l5hWPKP1BxXZFrvcyE7dEsxiz1YPeVuaapeXSkR1e9/YiKO0
0luvraQ1QtumWyqOvulEK1DCBWSuyUm01PlTQHk1nWwrkxfobKFaX5Uy8e0UmQTrmAEIw4Uik8yx
ncryyOlI/s9qjKeZS0uKx+S5eGOUEn925i6wc7mYw09wr9zYpQOu5V3hdzhQmaca5+U+lH+j4IA+
BCdIR24nqyYrVAjjNPrRbRwOr7TNY+O7NdCHLfZyMTWEaV9O/ojdwfcBpxl3ERl4nHhe3pXdaPeb
Srp+nvZtXrmd046jWqUKVHDOeriArzJbD1XNG0gkbjUYc6qX/Ql/Cr67yU7R/iZTqKzfSPYkP1rs
vur4Zh94VoL5ib46a47w0uV2htCRGRRs3fhF9oWeR2PQztYi8T3Z9RHBufKgQ0y/Q7hV42ANKoAR
/ki5Fhp3ldPVbbAmb5VVapUch5T1ntXfzI3qufzjyqWK8kUz0FTkzcOrKPknPirJKJx7F8gKo3VW
ufb7NgPu14x8wHa2bpyUq1oh1bPbCwyLIJ65iyIVKyjHGF5cYwigm9gTJRRXsCqcSSasmunyH49o
C+B2SABuslZKWHYa9+uOMkf44WFcIGsdCKHnpoRRdFZ3Nj+IjX/aosxF9lIqtc6uDGPhRuuHzfUn
z9hIPBZSU/tBb+LbFtHdIpkIJ4TjM5xNNGHRa5TX20aqmz3G2cpC2xGHnL+kDhc/plgaZ9Tis2eC
FEWnLm15xniZG8sNpwtLbreMxFgXArys/MUwqa9RHiDCViIAOtA1G6hCHgC2lNGDUcU62dYgmIUy
fr5/WHiwD4afDKVWeQ6r/U3ZLOEoSLWx8surrTViPs2CKfSJWS20T06sybKULD5jJ7AGLc7t8Fjf
//b2rtP4gAm/Bhu7EA7W2Q5m6ZOvx8XOiUBfOZtbIk7/uYdVs8rnobTiH27an35A6Ujbn4hBSYnM
OpAYKjlcnIDSWxsoTLZaZ4Pj0vaQRWKVw/8aQDIvXy6PblJkXSM7fxEi2/TgEFG6B5MZ+CSWoGvo
G3sGPxmvo3Os8tCjcf2ogwWKer5q8xoALztHjOOTdX0yg8p7557FFlY+znUSzvvZKDK4ouqw3AWZ
m+/NVEVJaneMSnByEbbmrhxnglStqZqA0c9bbZD0v9jcBY++ow5cx6H6z1g4Kei4v47jsKBWv3th
3H1CMriHJUr2IVPtbGaburMyxheUgoZjk86gwHTsuUt/1lAa42fiCU3Lt/T3wBM+ubGBChXTg+TV
4TdLCskATdt5YyHv9rc1RqpyCqyhm3Pwdobq/rcS47uRUue+fWK40t20ABHtiOFiq3PDa/rH8629
rUhvl0PWVWfv/fR9xD6o+FYO2rUtnyu7xRIQtg6RDc5KTcLJlXo2MHPOdDrBFzyuwFbUhfGixIXk
qMJvHkXRVlBTfXuKy/LG9kAy1FeoQ/fJWVcEv/N2uxuhJxaD6kGxF1HfE/56TKVRWWWuFSsXvBq/
AQOtTCJm75G1n5/QFis8NdUr53D6CC2U2Qn7bw4X9VocL27HKIM4/lU9N+eZfSGWQe0iFW6uwpjm
JNRShkaXqCazLG07lYJzZLkH3w+YXTRDaIlO7R4sMy9DQ5huNWWoj/d5k6tdG+DZ/96ZqYFp00dP
N7nC2MqA56N7KyGVx0Gz5OSx5bnHkkvM7/o7mALpmY5Y66JrjIEtlWzcnzMFMcRiOdh9n2Xj7mgu
zdl6k2upXRH0ziDmQrGX/ZpC33bq2gwTzk1lEZXGQDODLNDI48fhtXN4DzJsVtXGKPZSLeqCbIDz
O+VGdHjyai0g2qvKtFzFSXo2qpnLZjj/qeatxoNqGns08qZdYJ7r5ogFsNnVngFNXEl4E+zByA3z
So/031h3z95XWGu2R/i4VRwqfOv4OYxIfFwd2vImL48vDrj6dR8wpry+7Vylt5Z/PG9WBRqjV8QC
1eKBYgIFktUpQ5kxDyfRTy8KCAU1pn/L8mZGOuL2b8flNmoO1bCIiaijl9Phj/tHFlQ0C63cY0Yf
sM20+PoTBpLOA76imq2VIbreDgb1G2H5xkWgpl3okKmiBkCM2lDpt+KOc6tmLDFNElQw4sXDMzgw
rojpbyDmo8zqxD4o6WiwJdXzzIRRVPhuEeAuK0TihwQDzdw5D2tWSXt43AIdxBih84RLcV9hCM/8
juIboyE/bXKLqdjH7/W6dv7tqvAf7AWiel4AF00+N4x2EMGIxm5mp5uOMaGuQlHVZnmAYAA5b6M+
rH+0Vlz/p+ZibpFYgRkDUaCwAVktG8tKXRhZmXZALXQmZdTiPs0mvtqKmxJB9raXeRjA6TfBfmX7
X5b0CF/uRVv4WI9Q1eFP3hYihpgeqGemX2atvzoklNbbqN4jSuzDEPtQyMDK6NepRz1yDSail3Bi
jPJ873VeEH16o7FwYhFr9ga2gk+Gj3Mf5s1MQ8Mki7RQytrEn447xojsVs53AXKQzPrJFaFLeFN6
Ao+FBEgeeXKkyypZeWOmrGT2Bm5W6nL4yNNWnNxvWL0ieNVNPMeFGorefLeBGzM6fdxURbX8pKNW
1mvdTx2UoS8uzCpA339gZQImt7Uhtu8tpIwXEMo3Ercd3VXMpqP03fxLi3rwXAhBd1kq8NNHkacl
GZycpP7FXCR5gm2UK+89erMjENNUZGpK5LAenOtoYmMgxBLTHCwhUxUd/mrd9iXhCPsET7xw0fHD
FKMocKJxCRF7BHWeLVttFTVw2GfBbbBNczR086LxG6jECSUaI2f4qVE4x47w8Ts+foXuSR+H7ura
78XckDwej8m+FhrgIVUxKrzlW1KJefXMYjJZPH8+z14zxZdSij9hBl++C/aqxaS0wcX5JweTb+Op
HLq10kstdQs9ym2TfcoUHvVziz+pGlAYw70/RCnhUdWFTA6ip8Lt2I01+Mw1RugaRMfkJS2eATvs
LOQMB/TbnScXGM5186ODz18b1ZY8hfIsEyMRYC2Ea90U165dlasitHLLKriEOWsvHc7evHDZthP0
V10ivXGrzo3BSsm2DUG6pHWuKB64ea+cW2d5PmEIvbNTf5Z/+cWWdk6KjYX27SpH8Yp92V5ScNas
chZ6Sh4z3JcKFu+4ir2Y5kXTgqiJN+Bs2uXskqCX5MzN74NmE11b76XtqlYRRyspQQCFfRabNGCe
zFyEEWaE7llJHEc8ygfp8sWPGC8vVuPqEXfwXSeEOsVX9zA/5Fhr/qUDiXxZAJZU0sANsEI/Dydh
qijQjhTTquI6QFeyZgZ7QfNgiO+NEM1b/F7T0goraKX2uXB4G0ufXHYUDuvk0grlS1UfXBHheiV8
j/9kTku7+c2R5JM6mEOTwhwlaFhMXeTJKPap32+OZsYqJno6EgxYZQXmrP5szKFEMvINt5nrHUeM
OpLof0eOKAkUQedKKm5gj/io4dsy9TGPooZ2X9nSFfAag/fIgMs3JBydbVEm1qRGuXXZ//cFJzj1
vd8rxBUrLsvl4iDGYB/da4bMuvaq//FoIvh0Nd0EHxil243B9+sH+OFV/1aUDQhRvmOWWLHZIpyp
3/V0zO2kBD26oJ+Pa5v6qgm/8XhN5TG17C/DRT0IoajvtYYzMHiA5I9TgJnX+zwAaEYXGbDNRlkh
KW14JvqnzDvstRK5KfaldBt/iPnTs69rvWWVxlM65PEnNPPs55MPorXQAugUMNyFWebZdl6G7CMD
BkMvlKDuzgsYDzpy7m9zkO97DJbjQx4u+/caM7YSUFX5M4Q0q+qlkrCGgdJhl5g0kO3es9J/RqHU
CM9i2pu8WSfLg1J8t+jDhAQa8XMC35j5g7jcwd/PsXr9YD02n9NGawQhWOh1mtrezv/HiEQnz9XL
c2+fprhAzcZpgZZz6vKY6PFHPjvTZz7lYnlnIVgOL8cdcrDVuyaXLiTWdj2bGZAVun6X5MRADaus
HiSg5BwZZQg9lEfy3KBeVaKpfZCJ5Jkr76vDCdBdkcHyswPSUp4zuUkRsVMhW59w7Dct8Lt1j82z
BwTX15rFAwvEg6htoXmCpmhzcc86Tp91jfbF1K+Uvpx84P/1ZSw/CdVqUmrqspi5JINMsztYRPoZ
vQlOOyoGeYpPI16/zshFXjTuF1WctW5eBqQeVJDX1G6SUawBsgAcxkh1w07z6dFiOZfEbY9uIH4w
WQuWtG7L94ep7KRBb2eNEmlTG8rDjw3wpLR5GtgRdcHzn5CIdwtsaPi4iPRtK2ifoYLStYc+UIvY
uE5KD0UI4iubwhQ8SGKnnHHcVxAkPOYuq6yIkP0uEQbc3wM0FqrnXzpSBOhVxiinmlfU94dI1pLk
WS/4NujnNSB3Ie/+WI1UWbLzpcB2+7PUeNqidPK/ONpVWzuqH++68oPNct1zO4CUXjbsEctrGFxE
+uc94grQvTNc9DcO9Cfm4ZzD8h3KC6UsttyHLTMhtfg0m2KHe7MPzvaUKkQ6SyZNGWoLKCWy5MJz
yO8zIlIg4ZfzttdKSHpoFE2ZxTO7suq+YTWUQFLCfmETMb2s7lxy80ACAc/PdQqeKubgX0Momr9G
KLNy5l47MloiX55P22s3S3Dry7Ypb21EORfgUK73sGg3hkxh//gdiGnq738MJBHnEmJRdP9pOirx
mlNrJOMFQVffoF2gEmTEZ8aSFvidyVOV3cYeWmGnkP/Vkn7LorlQE389+7/fJC/9ppdtOjYVXPSn
R1BOBhRQm47Oo6mjiALF8D2GnmgGwn6SU6qOeg2/5k4pR3ycP89Dx9OCaOQziygZpQ9pMm1dMoYG
Iq7Dj2a7IGCmCH+EKZgMMNn2O1ok9VZsux6UcAVb1MlWuLgj+c7HgMfA0yftdJTdBL1L7ZVENuJP
bD7UipXtM4RC0jtCObxUWVMCcv9uKn8wPB/lnzO6u77hQVPtgcp4byIEu5pylLYxqo8yvaodvgRx
TnGBsqJRtZ4NwCX7pb4gAv7KtP2qjeQHIg2xYWMzAwZ/38WDR/gZsJKcQI0lymVaILU/uRXJUx3a
yfsEn+UsCjiyMmW56DoDUBTNL1ddKVCfkO8IZyuqEZhj0WD1Z+j0gYgy7vSdIdwR9Yd4H8H9Hjfg
68KXS4nTyp1s/9Lw2gIThF025PskfsKFon3cqmu5GmtL3sgj6vQ+vQT7jm37SeNsyaldgRKluavw
IkVttnsyZEKFCWtZaB5S1RRNulN34eCEM8wRKQq0UV7dvV/5Yvv1ydKWaSGB1l+hCw8tBVpFCUrV
VzzDIOy4rVWhZji39Dgx+f4Riojc3rJZJEVCkkXZDjFdWpioRwMuOfeWHLx1UgOn3P86FTRNgR6D
LNL+cx4+xf0KrZgwHaFr/BaLTjzUKA5M0JHHD09SMsnSyLb7beMpIIWuVDNUhEMryyLbGnIuAIuG
Yw19FUm//kfUWmOIb9im1TbQcqvmaycfM+1HIHu6qFeMsF+U5ORDG5Fb2UDM68ZGk26AUzuxbQqe
mOsRI9uJz5Jly088+pF/orfKQ+8BIb7v8dqkEYsGOxTaOAI7Rh1d76gWhClgXi18O/4wJSNQtf8D
OGS0dGDRDkXX2rnnZU06Fxh6kC2814bwwWW4IukwYsuJyCn7ZP+9yfkT/JIWDvmOxmYfnUiTjQtg
RCzxkjJlf7UzTtSAUhPwtztuT0+vriA/5+dnfciUEntwfVPxKunA6eAWtsgP8mg+HZtfrAJyq4Fe
eN1YuNVfPk/dmL56ayuB95Ap/4PqvdpINdVVqnNm7Ni/6QKhNJ8asgrhcGpdP5t4KEW3FAjTjHOX
rXFMLecH89lOXOrQtECZPEZbsRdRArRH7eOXXaMJE6cZkLDh83DxUamIcXyT+VwQ+l8DBVVBt4q3
KnJIFjfsEPIu2qZLwSYG9Jp5wAUCh79PJZ5LutiupNGclcoIK3blOcQlIwpzRbEvW9sXmMMww/YK
GGHVbp27/4ACtCOcUz517EcOMFtlGltcWCFmEX+g2oRlQsyGI7U9AyDBWgeqz3V/lVjPxSBpQwp4
+N5RE6neaRKuxCNb/a1EIBhisqyRvAME+Po5BxMk9T1zzbwS9zvNthAJAjjz/dLmgbpJFzR1YBJO
m8zbI6kvZwD/Pu0PpopJMM/bnFXERAn2TYUpvamYwTqy3cafdkyDPDWdhawPUUIVHzO0XtUc5Ula
arHK6PIzzWYFs2xTpT2kX/FZ/f5L+C3JQA6LVCPLPsUnMgufpeEehvRuLw7pllo31LbMyZKFm0Sy
SxlUBfNCR6jQ//HjdLDoRHdm84WxLq6uHXB21kE0vKt6W24orWdGRgTFCPOzQcqSEAjhDMtMiekr
vG23Y3L5AMcEaai1ybONcfhsbf/3VYugday0UQwwdOoOpTrSfUasMcyfuy7SBBd/87nd9Sbfw95L
BiMn3fRSZV53efvY5pqsUJRLP9ZW/NI4iPk9eIhXHxkpBwLiNJFo3qs3Ygb7jk7hAj6hCB9vnQ4R
UMSHiyAVPtqXe/wQmryxHB8m8ZZaCDPm8xdBCBhrUmtzX5gOmnfdkv9O9zRvOG/cjaX7Z7OBzdsa
rjcn7jxwkDk/5PGGWv/gop+Oc5da23GR8oG1M5doBnjOiVzAQm8noJayKzmHGHyRxemipVxUiaeN
klPFTG36PlzEd39AjEANtYZWjHQ6wZOO3q1Qrk+GIvGDAecL+zxBcUMvGr3lhxRuXBnnaPxT433N
vIKj2NVwpJIgjcSEOlata8clxSaJBciCdg4RmOCsz2rqc074CWaT2NgcyAexFsewhyiOMKa79hLZ
PehIzUurAY54gjcz4OjXmZbJAfOfpHwHuMo3V+EHg7G5uLVou0Zd48PmhcayQY5BHIgA+VZHuyRF
eh6Nv5S26mTndo2G5L/V66A52XbBYqAIDH4vS060K0HSLCwE9IemFcpc2VH0sEhXAI5dtDnib91J
aJLkEBL12WLI38muJFRTJCKGk2UY2XNzkd5YiI3jDJ202YCPvWm+5/ZuXBfYSUYjIIn8YX3GPVUS
JxBglpRB3Mz+89f3LLWASUcrrW8i0kqGpC8u6mZExiXakm1I2HPt416JhH6MOOwUV8KEBt9dx2sv
djKMIIqe866cGNL5dIo9qvRy/AqMLvYpxnxr4KlnZFZ0uXYZtczMR0nvwkjky7fOWI0Grq5ZiRpi
jrzy0PRGHoeiKD7eOylWxJtgscBTdK4Rn2rLYJJ20wKo2DohOEfSsG/VFA9NrYUhDm+aPpsPdgKY
tUYLrBqF6suUY2XA/2pDcRfwKg9DAfiTP0quPAy4QzdrqpZInZy3C2/3MhNUYSnFZtbRpcGvaq45
xSZpwJZvAyg5NS9rdASkR9Mfk3rDUQKN6t5aDd0AmlcotrllP+u28CXz/aD+lgEhUTGqY2wSJfgu
MCvS0wAJSMADyvcbh/O6NJHqLVUx8N+BY3VLGXQMKlzZkwSKnSCCl5sMjBPDanU6L5OvqQHNwiIY
/fEbqbPwIKKIVZTAfH2FBQ/usmxCeKYq2bkUo4d1z0BxOyPaTQib/FF+gbO4X3IJj0kmbrYu6fqJ
Z2VpEjdF4rHpDfeWG7c0/DiHD7AsCCFeUthsOzmn9jS/sIN4mh6Hp+KYgPwogn860Qh8QB/L1cXZ
QUzOo5n9Ew/jxYBJMq0GGzN2eeXPJyxwpZMEn/kkpTknoIv2Cxc/Tp4hLYLIHK572TXYiAklB/WU
hpUZR5eN1hvrOtsYyQhRyftpdGBRbietfZHnlGc4mUkLRfEGIu7ulFtvAOxvyGDkkpg5KtuNOf+d
E1CndFQ1FVX7RR3JkyekBXHsC1+ojPpWn8mVzg3A48RPN5sfCYW8TtX3muJQx67rpn9XIUXOUQNP
/eLDHuFGU5FJP8aGFPuT1ScGHFk0+3mSpg9jOhja2sJW/A5ezcbtgm/VaVI44UX0YIKad/GO5R4S
xEJgcpduaAbxks+7RYWH+wGWpjSO+HKBf6ZJDmh8FJzDIDnWuWwOPNQT9FrFvds+pxcTlf16bMB0
iyE1GG/b1IS45C78lTeavZ19gqzRylJZ1ailted16LQnA7Vj7nfdcJwYgsgIaOAf9XWwSq3LKh4J
tAxLuMGl0sEijNHg51g7jxWh2jeIUcu9BwOIMr+arqUhwR7uztWG4wTgH96yh39HLtY4U2fZabkr
vzIVHD2fAnYy9VMEmwe/igMx/tgVAgyPYyeJYbPBxTteoBq+ashdBri6tHLgUS2naS4KpMq81T2/
P8VxgKLGrZG1lu4lH5Vu34BgjsjrQFxCDVLToJYn8Pq80PV/JLDt6+/cVuEUXScJGKGO8NHAjnV2
yibuArMzcZvuO5fnZMIQjX77/pGGQdhI19wowzb4Ixdy06XnqHrZQSYJjL2IzucBV3kAQF7xHD1w
YANb7G6EqVHiisHC8L2ZEzpeOd37FnQW5PzWQ5p1FVNxV+d2tVDJ8OPu0ysSckGlCUInbATPUwFb
oBIqg760ZZoxmuaa2YqtfUXYKPxV+0H+bHZj1CcDcG89DqnxjNSmZplsWf+dwLJWFUMoYEHtNe8/
tUkMLV7LJ7bw3Gt8Lzq7eb0rxziPiVN4NQy2t3bgnsGDmdbI/3jMLXlOYb+7PMq2JuJgqNEC/vbD
SSgKZgurCnrPnU7I2qWYDoWC04Zc/26s/NaWdeP1NUrBVMuH5GFuJkak/71mJEGJrZU5QVRlZVR0
nYw2W+zVcMGVG0mBKdZRDbctQTp3l5Hyd1WS84wLgTxEYVoTuU+rIeu6BFCzXKR8bCf/g4mr8z1K
gq+Q7X4oZroPXeD00rJS1NBnvuJs8ZzBShNpjHgVilsRbMJPvkxRL70fQzKk2UahUVL89UUf5ple
pax4ywEb2lu0T9SToUUC++KgaEOfYeM/B9xC+rCii/lwfaEeIz2ZbS9j5jkA+U/azkLVH1z7u5i6
GNFm5Jq1vJEYrvgNQ1J93Lz0xdFdd0yA1bh2jA8I/m3pW2xUHDTzsXm/gTZs6x0t6HMNUzUQJ/kP
1HW1D7/dC/bCmVrbYWRgEN3Q/JxF0vu8sdvmSVU+EIMDBq0A9EN7XW5qBqg8iT50Vvt4zpO+ubph
9p6ouU+TSwaKS9jO3ixQ/IX7sktvTMLLLZqYaf9vkOVE6z8rA3HsESsvmFcUC0GdYF9clYwet2OC
PJlAzyDYBRhzz8paAgY7kFDd1mz208WQ/GfQMOi8ROQt+9Vl7s8QYGXik+sYSFCXglrCh+ZKmZzt
WrIA0asqpJ7z/38oPOH9KEaolNGFqeGy/npMs7dcBmypMy4og8xAZf+UH0b/U/3/iET7mEMrIvtP
fH9vTHiws3BDCcOf/LPrO7I3ShWisHn6+oUv8n5vbEqUSnjXXP/K/mDoCDrGWcZMUvehLMtPYt1d
O9SfVC3hE5oZzBpJ+eSZe/r2evDItd7WH0l/6DRCUk9QYERSXTpUM0rxpcYJ2wcG7rI3XROqrMnH
rEvG24lj5LcGWzTTt4KfQjk3rA9thKnnqObt5D4af4b1a4nWiYBeCaW89IHDFycXrhrLRDvHu1w4
zO8EsHQtXlC1jBFL7xYWKwOTo2Qpmf7+QOdTKWSmwbQzuuLf2Y6lFZjbG87y6vwCh7lfQYbcwaGC
LmP31y4A4K/RJsPKvGL0pVvW+4jIBUhn6yGFw4mWrc+lhVSSmIwzAVem6sDEd6pXVxhEGo0mboTf
AiT1YUlQ6pwAgGhUu8fmCRJNu4f51+jvD6RwZuRtoZgTSvKI78HNvogGb8p4KBiG2kQzpWv3iluB
FopTwIFy92pB7FB/PmJk67bjPqM0voJaDJsLibVNilnwYT7p172dAZ6r7OTWxkErgWQY+QBdlCSb
ALbvjUX8ZWGb4p3RoNQnVEJeQ2xQ/hhVm1+4n9pUOYSRIgMC+B7TduSs+aQxu5qoyy8ZX+fCwWjK
rGuancgN/rAvmo3aqwv7qJSXPRWtciuU2zr/2z+UEZXcsF+WD+85UDKeq+W7TODlTXjtD3Fh6YIf
vmbX0ngA79XR/bi5O0EoZxYQFaYKGazr/D9FZ7LHh9vDK/9vstN33oDQTATHxCcb4gJFPIvV9UhL
cUl8VgGtS1/sh0WU0Z7zJCWSwD5opv+wFBCol4uIaV2MZofnd9uJQC5ePGkWkwrET2Ao2L0KYBtK
nXvLIrIo+D58TGZ5pdU5Z1X/gjZy9HrsCDosqxr6GwUZWxWiZ7N/sVAnHeAMPrFU6T2TzFuKOM8K
DB0+ZXs4rCLxqvcnJ8RrHxjZV/vVQrGEOh682pqZzNAXKgZdm1IEetDGkYqOAGXsRj4NVRYURHiD
v8b6JeyMpelDmzIL2Q+87Xa0SieHcJZxgC/0i5Ya8B6FlXgD7ml/wu7kNbjRRvrPUittcix+ZZf8
TDeRFuAYzV/qUjtPn3ViJdvx2yd/1kEAF7Mn60iaRlUxMVMJX1mXSlh/3rsF2EmyzsH8N89Xtisz
4ny6Obxx7qZiRybb3l87vpDsfB9MrFsCBBYsgbwR5TNDUtwbtZt2nKiVHs+LjzkElmJulWefsye9
EYguQJ8IOTHcgBlNC27G0kUu5wym1PUvdwtqLWBsWWfSPy19SbI7K5LEjr4/3wVWB82PhmEUA2DA
d260ySarekiLKCowgyi9b0lCmhZI5UmUTPCduwC39R/7wgyjriqaZd3jSl/lc1e08Tf3HBirV88D
4F1yMDLBoX9yMJDUqx78fvtjqawhbJBqM6t030qG5DeIA8QF4/4CLg1e/WQRiHtpBQd9DgixmcdK
qC1R7Xp49lwCErV1JqERjRmDiULyBZEDyO8GbMuWh5KSgXVIFDxmBWlIOdoYkgRcR1ihUBef1+zC
81ZI86F6AG2t3B0RPsPXz0Uje5WVoycII1lwKOfAzj7IuMeRs21hsdYeuOP8jtR81/pb9jIGCBv9
4pBWxjM6ffFNUwGnnVqsjaAPA3mmGytqkzA74rVfHw//S7uWSm3mmeT2YDxTHjm2SA0m7viZfQJ4
oKnUm+2cWtbNB6Gho6tBZPRsw1P4awChUpLo/MR84SX5GFAhO1LyjmSiEl0QKmmqBtbpqvOPAdp7
YjdmVYoR4c9uHhDhlInZ0RTLFuyAV3AzlbyWeyyWElczl86RQT4EQm+LR5okg6rq+f80JUF9+opk
+mpg1IP1NoZfO5s6xALPNI7UwxWyyW5n1T69Rux0HjK09OCWipy5gI1N1c8VK9WFTkZVajcSFZCS
I2LlzchQhMdMf0rXguLL1k7za9cz0kksar/y1Ae1ufobEt4LILY/xVwnXthRG7ngE5bSW3enClXr
MTzYBFTXwlmklIVEEhRdX2LvcJoe3yFWgxA3qAtqthPuy+CbFEWgycW9XCW3aAdfR+zD5oVHSVgA
kHwXKWrLHRYIpoaMav4iE4+NLHWdme4o7ojyuytcVMQVi2mLsp1CIhw8k3naGR2RUS35S5XfJXBf
71StMkZ/QkPN+ohSYnjK5E5v90VN1lOajXhmKooXu/YxWnklLoRgsLAUpEHnU/bHNRfGCJBqEoDN
VJR8lWK/DreHVMLiEF+jaPrADYVNw7O37q+m+cojl9XUcifyXLsYoCNkrtPUQRcsTM6RcIwO/EMd
83kL2PZVEwXPIZF7kIIzCf2s7Lk9V/jbcv0s/KzUK3MbKnaDV+LihJK8DqoeCVQsotg9iL3qg/5N
prbH2qJy/4FbWt74MfflPLF2yrAwDR7UBvgjdNL5xwwwgx7LapYhLkMXyAkAf68GV/9bWrZ5h85h
rXvzQmaRaMsKqkB0Rr0n1oa3hf32eA/OxgF4XRipyx5/Qg83WkGNuFZBXEtaIUbDAUXF7SY6yUiW
redxSCklHYRXAjLQ1BWDsJufT4L+MruH+afOnlgTX5ZPSskHDoEeuqbhY7A5rOgqwi1vzGaZo7hV
RZe0ScCUfJLyVdKROSDTdGBsGrZz3ugw7fkyp/XXf7SRSWTmbubiFzM4RNnvIOJvPpKT8HdNZF8k
Kdh8dmW26rxVvnCiGMWKTZ+aTfNm2Uen68nKn+idPy0oivDDWmI/dhBaYSukxXGp2QVXVHL1hHYa
1qg/GIICawoC/3hbK2CXzLXHWXcnMttfXU5gOy/DNy5o7LWxIOO9ELyZ5U2UF5VyvX5Qccx3s5Bz
WBAKHmNbzFJ22ECm1WyE1BznXV23MS+8HTOQZraSTUKvcOslULeesf/hCEuEzUdStGvu1oUV4WCI
8z8/X1E+yxQz8IIJKHTX6b60xMrAlc1T5WCkyl4Ev/fgEbQP5BZSJaRFCSboWHMJIcTUeR/lyMpb
7lShXipfKa5o6ZcfebDSgXBxGd1iymYUbcm/6uVY+z2208Uct2S+Jn8H5aj6/KAs3Ul8+mEXLyI2
OSVT8MWixVItbWIpb4HQDZFbMTMm0R4KEL5fN2N4ZYJCRR31zDbs5CO0u7Ut3r0jiCWPouD7dWCV
4p6aniCYgUieEXUwOj7NgrE85FRjPLCNkeWq9P5QgMUa8su9ZAxsj6oJhNjvP+n6okXjp1sx09Au
zEqnmkuEsN7ZU84CHab/7p39MH06sVpDGh1/oTqqzXVRCQTww+yd3sNiUX9MMAdE2GsConQn67AB
KWxHGBHTaL0M+jC5hBx3wonh5VQUnAIIjX+QQSEX0JhGiPIfAI8NtwiyRsQmHPhseY9xHpEc3CbB
qA+WOfV5QxuAcD/K9VeqJ3w8FDcV9+XJ+fIGfi13v8PUC8lhdFG17TwqQHKTOCo9NYn70OV6zlLy
u6I2ZdWFNlUDeRSMZ19WrJX/ZcBQnZoQ1BS/gXjQfyjOg6x3fQO5kRr/VVVUh5GBdKOtusDj82rL
cF7O8Cj7EGGqBOIcjl9Tsn0rI6wR6WkJW+z5VLcueADmkpsX7yQrRRKveTzsgMNVDclZJOLmoxku
LemWVtN8iTyHxeZG9e1phhFpHCQY3+x4VvEbdQeqx9Kg/n7xslk3J0k6n5PCbvGtTQvgdScRa57D
jFdWhbuwBa0SQf1KwBp/m8f883eIHMeg3HCI2ew3Sx2YsZPw+rKhY2v4xku89Z7x4G+c2KjK1IKM
XyoSadQptNWT3AfHKQHuSfW5fdP806oEGVR8j08XwLHvAld7Ku+0aA9u15OPilF3HS3RVBhd+cQI
B5ea2WIwyi0OvUp6XI6j/G6mdozAEmnfxlHPQO6yMQIMul6XUqJ64+iDQLGJXiYlwyKF/qyQk1GN
UfCfNLTD1O1qAxx4ucdy8GZH5Fv6OWPt9i/mSCmQK42KHPG7CR4gFGC0GOtqCtB0a1Aml4PSLTfM
4ZPpJQEb1Q7Cxz2FZJCh4N3Sjqfy9Afchs+Kec3XDRyl07VyUbgGG20qLbwBDVodbjnC92wtVP3i
jgYqsXtlSSSBToTtrhgEtb1kotUx9PlRtpyhUnxQHVab7I3kmrGTjgeHcR/yOwNmuqC9RpAVR4RJ
d+Xqe2rRdGLsVgRj4HwKhTLD2uTErQlzeUJdipFMsO1qUgRPi9toryHh8drBeNPzbMerw9kAvKxe
ikagZUDyGs130BZyR4zqHwFsg7CxKesaduvZ5qX1x2MJop6h6k6rJFajpLf7rhTOR97afp0BgH2y
RFuBvU0sbrll54lzdPiTc6aIB/PFOkSC8oc6ft8pnPtPlMn/RV+Xa5GI1pVI9uiB9ib1fgwd6lCR
cG6t/TaGkqXG2jXnfd6yVOV2ORsBSjSUL9Un0+Vp/cn6KbA4W2B9r/CPUGS2lKiOgR4hnAdxEq4+
LcqW2atswkF32Q0HzdMnM9/FB3ywQvGQHJkazoR59skz5CJq3nGUnzlEHwT04bmBvu2QFhGjFVNx
QCNxbljOvIEoHMZwHMjHX4qsvaa3IsLnMLl/AVOdfYLe+V+gyyWkme5edOMqVzJiJmKy0kZn04br
+P8Oga0/qLe/o/O40fufVMExrL9YIGJTSTdj2x2ePNF1+k+zy5kGQ77bMb91t2whr90ZTd3hw585
v2fAQz3KyZek/dB/ujF6Q8gs1vQPgUbZD6L1JQl7TDmqO/dgybyPyGxwSbfvov9qUsrOEy3sfwaO
YsOPVCVkA+IJ9/144jAMvH3dfOL9WG6AcwZZDxoswgd9EixBVpVX+XtyJwU/mZolo/vUsvQpafBE
BJbJ8gJ5k7f8YWcxpP5vaWeHCwpMxy62aoEl1OuWAwk2K8MSJGsmlqWsObK1nJMOCK5l93cHQXlQ
x8UsQ9Hxs2LzUFuRZjZOPOsInc9TA7jx33xkp12BOa8xUV/Ot5npk+LcvrgG3yXJyZXdJ5SwM6tz
KT4uNYwFY4OTX1OjutW2vgdbBeunnKbPNf4WUhuDOqBNEvWmfIn6ik1VTVDjnaXVhyWEng8hmtEH
FEUN5B7t2NYBmTqeW6OJsiTpd/qMp4kL8xqgP+Lhoe6hUo/no3zAmTUXEeb23c+TfV5I1f1V6SG1
7/hLKoQ3BXs3+J7F5ixkZxO8ayLyygOxjR+sCh1Kuq+AjX5F9hWfaycw5SXDe5R0XKVu87gnSCPd
ckCHteaUCCDWk54QzCmQiiOLnSnmSTuC3O1LgGU7W5UMC65YIlbiQod/JonNcbSnvPAM2YoTDjmd
EClk9AqglfOl7KbTcngrKrULL/j577igDrw94rLQzSGdgFmu6z2So8xJPEp8UKz34JNepIANqLnb
8G82CDL6M/Xh+wTrupmwJd5n5YCm2gfYvSzjkOkW8FsfFVUl62v9pq2W1LMy3PDa6Q3UwprlZbQS
HkV0lKKsVyI5KfqNxFlArY/dRfvn27BiZHifvPK5qD2EBa6tzyBD1yEbR+szbv6jKH6dKZT1/2WF
w5O+0XdT7vehBbrL5Q6zpZ2i11tjMnY/XSaOYPiV33IhXkkl4Bv0XVso6FsNcORAm+uF7M9+GWWZ
KfGIt3PLrRWJ1qjql4RQ1h7z+cOiiyWTUCWOatX7JYhgxYSREeAn+xTA6HoHcwraerY3vAbgqi8W
nCycbuO8cfW8Ut7+WuxnEQQ0bwjrhmoOqtVm5zjZVG8Vac/b83/lE41NTI29kpSNN+lGIL58Z+iP
Mar5FqDG5b5PznVbgKW3G6n+ZQHvoLdV40PkFGgfKgI8M5cA6XiE3tYKuC1ez+19N7IlhK9/f39+
2M1chA92i1bYbhwaeO7t+LIWntmD1s8ogOgPULMfhAXok0SOUqB9NqYkfPCOHFfXTm47kJUmBqkD
1nc6t023lMo11MMDPa37mmgvvLU9zRCUhA9aHs8TFd54YbMkVO2+4AT4k5rm0wkhSSZuPHYqLPK8
UVrZaWEHiBmd+nzvVQrnDNJc5fgn/MU4VDs5FhXS5YkKi8slP1GzmxoQ0SBgL+AwQ/qR+ZLuReBf
jvRR8C+MsZeo2w7d9jBWvVa6RnxZja9CVMFQL32EvD3PF/ukAZCrBlUn0m7dcmVQ4omLOPN+I6LD
/sKVwo4P+p2WXOAMZ3obc5EHBlX5uDJzzIl0JbTiwJ5G2fj/4PCm+i6JKbUMS3ZsjtoZuygPWTaw
q+tFBGvhQFxA9t8v9KyYn/tAfAYO16+4g+pSZzQf8/aiwabmcINvp1YXi9JYEH1em/ROOjX6XmjY
H63W81Uy6WgxEV6WLT/nsRXVr69vjfVwS/OCjdcqqOg2uU7Bz3rlnE3h8WFPaaVgmeQc/eBS7K/v
jQAqnqJLwvhqhZ5YyxL1HKu+Ghu+44t11OdLxOQbYlHpPm/+ffPT+mS/bpWYMQZYNJqCHeG23D9Y
CRQBWgvBdmIknbaZ1TQnQI7WL52CILe9EjSdfNpQb9FYXpluM5JmP0RklI8yNfyo4tQr1M2N+r98
ZSLV+iI5CMKkCU+Aj+nA/Tf0+T+Xb8YhOtafvps9/ExiBoSzT6G6jpuMK8vTABlsKbBvI9mbA+2L
+gnX7nrbdMn15rlVG9aaj8rmt0thQ0H0vPJaF3meZs1dSRry6QQHbfENf8gBj8Iq/ibDAyhlgecz
10f++LQ2cL6UZtngWRP+6X/uQ/KreAUFIItRHArLkQ0FvgNCpLrj8wyJDF14Ui6rV22aqkESLuA5
pyUnPIRkaLEwBcY537kln/BCtEm2KLsgJIZKmiGY9y0vAdmJUZBzM0EaEnnQ68cr3IksDJ8iF64A
N+OFs8zDo7Cou8fXjtg6N92PoRfO4LKLrE774V5vRUrHwI8NxOBYodlrKD4fwg89enuU3g8D+SL5
rCv40pCEx6U8X/UP3S8B4D599EnaCQ6kl1p9LLPlPq8eYU2OggCAiNYF2TDQ9kesSoaJCbQOPPJA
XP+YLax60oo3NclyHXBTlElVZng3zs3M/M02w1zjoPLY/RUH2GKcKpCh1Vt9ZGKkY3Y/CfjasJ5z
ZkSw3WDKTWY1Iqpwchqf38DNF/m4VwNOiUkI439plRK4IolRDbbjum+f44/lHygO+M9Ap5z9wn4u
liEEbvrQPV8v4FQMQK3M/Usj+pqROK2ZgEk+PaVHx/VA8p0XnZ2eQrvDYeeoPslZUZEEsV1/9zVX
ksJRiI28JzWH6KZdPv5HR1L4eUOGwCG/rvvA/GWV21vK/ZxVKiVli37mudh1daQZP6JK6f7pfmO0
n58BC0nxfUWWOIN+DFJChafl9PBRiHP2L4BOatYmRSXGztA3kvdsbJ1DFxoYlLBHXJJq1ddYTQSv
RsM/OC8fp/p3SUhslDL7dGSklz/icVgVSsmtTKu9BuwfNJK20SDKTzl6OngwnJiORVYvpm4dcFcY
Kp+xSVkOaDXHS6yJxYgQN4igRiJHzBeLjYgyAhQAIuEXcPLIkB8hF0DkDAnv8EC5CH/cN/L8IDf5
U90nFlPUs5bYIEmY/aKnHHnyJnVmJvZQsAjk3pYecBtj5GJhN9WScZGBj9V+PnXESKzAeMTIaR/d
2Khx3o0/pmAZxp5d3zRmHs2Hf3XyMOR5avsRSQ6lSDHunqhQR21Wa8s6fiMn0z09xX5+il2kj9U/
EtYt47GndMEiUT2MbrZKkv2DG/30zgO1+l7s9K/g4Rwf9CDfSyQiYjxIPqtCVIAMHLlXwJNTpv6c
CPrxn8WegK+tqrkSOwViXHM8MX9RFyQy1fYRBCctpMNc21eu0UbebOkr7/Y4tTepamgpP20ZLAzY
wF/uEqih4Q8w56ixooPTBNxagqskHa3T+VN9T9X43Ki3Rkl1fR22JYXkibIEMolG2y4qokFmDe6r
HoPszjo/UAdLtGFG+xM40jbSgqTFEBDLu2qLEjwetCIEsz5Vso9eQbCnNN5kLAKL0GfV/dZXYpA/
AYotcWu2kMsuKHz97GCY3byaSlYiHAAwTWioLaFYadsanaVN624T5TQBlDTwMRo97r55gGqjKNJk
/tY/5N0iFif/URlQQkpiIJScewe4QjKBFE57+xwYmsJLs/fNfwNfDdKKW6CBqeYy9wmUjkQHDoUM
JGCM/C2meiBJPQb+9RQUGKlrckr75nsUPQHYW2xIdYS4NwGAHgvRRUEfMmB4q/rw8VUQCnb3aeOB
XIWNNcDeWRqyxRXgFNF/SOAygFmOFNeNNg50lwEHVRSw/4PZfAdiiI0ejC1MqoOz0+mswU2LLXsa
AQk20UqBkV/QX0a116u5qzvOPwPmWwor8RX9Bh9x6dt9qeRaz+1dleR3zWd0h9PcRZqJv3fzDwpH
OgQ0Rdjc/9HIEgsb+vSqj79cfa8kmPUjT8QjGvl6xNk/vHNenmLGadhXqvd1looKSW3+wLA+NePh
XWspNioWRwr74sB35MJHmG064Froso1+Bfy0U1Hu0URWkxDpiQCN+hS/c9JunnoPhDTpPjQQIpni
ABjCas+5ynCjQ/dgwZQZPuHAfHz3S7x64Or5jBUqZWy4GEt8JPs+oUPE+mVnA4kd7MjLu4SaHTAA
k2cxonbV59V+0gxvcAVo8hZ9sZDdyiD11Q60WX8sYWcNVKp12pKg9F5/xFZkijefXromotBOB6Sk
R+IjSFFzvZx3XLOXWMRvH1g3q+QUxhEX1CUwH2pR1c5uUIBVogaTh1E5IhJ6logkGU0SquUfAqsi
gHrNwctd0lhAm0urWjrCB74Q3qVjvYPtpSXwn/Cz9MrdIlEFHOsV4DOl3nSpQvCoJfC8wVQ7XLzG
VDoRHX32ATY2m8EriJK53mFh/pUWP+Ne8D2SlPolEU9hOYDp/qC+DcJrUG7NotzsaDko3a0vj369
ZFJYjocclFsGhvt1+4SvbIH2s6av0cQFsAEfUxnblY1TSnQnq8cVuVh0uyDHUw/d1hZqA8fIneHh
p1EgEcONXgsYoP8o8f6eeJpCnp0+6ryiWGBR+AfV0KKftG2VERBZ1TAS7iOHFs/CU9xALjG6KQsQ
e77t8xNYFkph8q1aARUNEcpccuGrkBwHKX2rnLhmCRakdnNcxMQlpuIr+3HtkE3N4yTokfN/swSY
SE5JxNFfmZa4mr5t29RLAf2+jZEopB48SUSENSASmGCMI3QdAWrfdcsZww1RKwSUaPHKILxmgwsQ
aNIKLDnWQuCUiAapjfjJ8TC+W91yN+Hs/76M0VJzF0ufJoQTwa7s3tpX9+fZJjLalE5jNBQsmImT
1Uqfz/uz9p78it/fwsGOFdlqDumsIP944LV1eCMadxMwYSlmapJXvx0+mdJRIQjlITU26KvsMUvP
cSwrQlTbffpTvuLmyCtkbs9y13oe6BknqTheUh5nUPzQhXIgjgxJ85Jm7Kwoz7S1fGqlNRJ3xM7/
N1uGzQF2UMMmYtlvyK+iFJIBSXEhEFteFNg8cNyY6KpSrAJr6tp1tPACQ3Fq4G78GiCB9HegSsJD
rSkqotqZbCoSAZbkPpD/Bxx/Lx58QaBG7jvsuU5DeZuTpg+10qudkCxZgO0z82QZ217jl64PcE+T
beIaa8W0NhV7TTCyrQuAyYR0BshAYxq8F7UXaN8pNmOUdxlOZ0gZZKnOzy8DVDZwIJRSornCGcda
vdp9qinvFT6u+3oFDuzUDaPsFct4xCxWBy4po1UlJs6pymCJAQF5tVyCXmdW8ZUJcGLXfkL6YcZ/
VanCeaNyyeRPI5yErciirIRHapdWgQ21NIoZ/WURlgzXU2Qvty2BrGsTN737LkH+8HsFhOTyCbEo
x4jVT94H5MbDIi7ewEXdjqFplC4lOh8Tk1WEkL2q5rvCyFRGWeWZfte33Q44Wjkr6ewOqTDMo1Zq
rBvv2viUCzhI5MxjQeYC6/ot5MoUgvkGsk7B1h030x6af3zkKucVZMv0Y9umzLQaxXk1LaNqwGW2
0AI36biDN0ZUK6/l4WvQlrvD+rE/21S5DMYV3qUGlsa0AQSFxNMJyn/XjZHljMWELnSSErRIM4qu
o3glT40FqZcXSkbSGuutzywMhMywBOudKSV7u9f4VrBRMgdz5xFAYJ/NR/okz1osaDjhgT8MMkfV
IDszQp3C0xvdufMcQM45qgxGpidodRmvHNkr+VHjWaqFJ38ilAeRjRJ3AuPve2ReatF3viDQaI+G
DgjXzcjbKuqjQmnJNhZ26Lpge+R2K/IatYFTwQBnyKRiiB8MlpJTvLJKvXZI4hGE+8LrCYcXVpJK
XF7try29xNwPOM8P8FySpZqrG5RFcrJ83UdATaZdtNH0EAUuOuCsBKBYB3e3gP2JRMZDha5+N/zA
dD+fXS0NSZWld4oLKPMvJPA1xX+148z8CIbFuuWBslId9/bNJwum6KfOyyK+2yPy721Kf4urgdo8
yNut9AJYjH9JZpNF+MblF3+5k/eHzP9DbHnHrThqrGBWtykCH54PaHpJaeoZLCVHTvu7SpY3KPER
wrxJ4oCmyipj83trqbEYJFVsaJF/REUiy1rBgPk4sH0g6T8LWe5N9wUg322Ro1RR2j6T1Z0Mr8Pe
2lYZZD+mm7tWdgvHnIJ2iRGc1fPj1NE+jbNgY5iANJIIJzoQsoZVzB6de0fUmXNWbulagD5YlCHc
DUzj96IQBqvaDGvzkuGxDAYMETOeMdM8abIpl4/QRl9YguBO6rVP2TGWwLEGFWroZK6OMJ3D1RbN
NwzsTi4f6Wxe0FJlZL9idA5bVcuYkKv7vGlblSRbsr1emiV4YJfOmnY2QHsE7XE09cN9aoM1d0H6
76jqQIJrGBLP5Isq7HuaRRuGmdeVaKLKTqumJILKKUGoJys0VWqVU65fkg9Z+z5vLF3aAdFNINBq
t+ahYW5EiT/ksMqpNL4ShKyAWdC7LGKf59g2e+bJjnp/9rAtjlNs0J1MCE6q59vApO6ZJrSQZ0rI
Esrw4tv3Lo7CgM5wXlcaFBFRXSIWtH0JrLJ04/wIXxRIKSGPZqQOfbQSvrWggR99C6ozKbXRa50f
DX0rAA12VRtSf67lhHjs3U0QaBba9anAk4E/PSeXUusBxvC01bObjhLs1VF15gO0zE713ohxmUTm
wKyh9SuhMHVnrdhhASd+n5uhkgdekwXJVBRHg3r4iWJk8cBEIlxs4AnyRQnqaOU4Ck5sJFIdesY0
lRcdqiiogUimVrs1VoZ47qeZSO59KApAHffm7BhjZjLDW1Tv9T7f+OG3DbWdCtFf1AiVh9UxVyiZ
qij9UmluFJ8NNzBez/9utZuu5aDOdXaFi7ALC3iGtKcZKEpQrskM+mm1J8tADqZakHTI6/EPhq1o
CTCuhNkJ47wjBT2ZvsG5W8+6AaRfWEHrczdIw6Qs37g0gG2sTZzUwbrs3VpdKNof/yYxl0Ci0oRF
pmmCY4R2hAQcu6mlAkDtL4Rt+zQVkiBvy43LG1MjhSK2+D7LbuwWDGKGA7ElZbBi6HLcoUPZZiO4
Jg2chE1xOE+B1IRG4ITS94TKEBLRdUOPigMv2mnu8azNb+Im2+dD/ajP8rL5rC49gb+9yK8aER9f
UPNu83daEOMZpcH/sfIWC86zL/FfK48AqLhdR1QhylxuOrgIwNTgfVrri0LuThrZD8jiTU/SCN3h
k7tN7OjR5ayS6nqCh11RyIbu44zvKBETNNBGk4Goj3qO5gf0PmF5CfuZLbVpPdrbADQkMjiWq19F
0D2Op41cqrFyPkZ+mjQ5UacsPZdVnn5WX3m3rAJBc2VHckhQJdFX6dChonmjkYl4MnIYNLFhyThs
WD6cVL3Qo81jVC3wQu14gU8TuHj3pH6md2LJo5btDCQxFJsvjNKk369yTG76LpiYcZHyxi91FjUv
mE2oxCO3qItwbxyDFEei+ioHaFVjnhsu81AqWmav/HGYM5VDZcjHpau/5vFEwhL1UsdywKtrJ4Vq
0+/a34L4au+0E5NTAU+006HRl5uimTCoA8GQfUFi733y6Wn0NPE5GMfO5pKWs58AJlswIpQH/ZKF
L9cjCD+PvhEcte4abehr4QwAbsh/GGAdgNVkke+WTxDt1FwwT6cWh+76t1m76P+AVyCkVorw4j05
UuLokyDoNu7ym7rEFC2awCVo6EMbgsUFu5giMlDdBRX4H1yOdctxGaF3DvFcsccqeOSfG2p6tgog
+7AGGGSLw8ndJRYa7a7JeADoiZTQ52Ppeha6ICBVdMvh+nuoq0/jxAsr5zUZMmJ4ulZDTudRavqt
DOjFNRAxSYogCGrAavYyCGczarE2GxrlRdHFDozHscYrLKJg8ldixbwKastTeORaqXyxwrzNasX2
pWs7U25PJhqzfNdLqZQ2KByYdleGQVUOVSUOHctNyWh+ldmHsgnKS8SbuDbJBU5jFwARTofSXp5z
v1tL1kbDIwal6ka/Gubd9fR96UzF43m4UadchWYpF2LULKidI1btUDgnsZVT50qCXiwwbon1lyE3
DI9BhL4sODi/KK5Wx8kN/EkMiB0QuGYau0dEsbs4XzhIK+wELOiGvc2b329nmT/bw+fqOI+uWj4w
ZS7xvXULTesx2Gsl6z2D0QzKzCOZBjWOOjqeUeXzX2e8qBVdQYvTSoVWIv7pPXIkQxN1GR5FrtXv
y/N/NvDF8bF7w95YwD4JpIf+LmfjGK/7z4yps78Okr1J2siHnbdrjuNp2ivTUBxQzFHd7JsYw8CB
tzfS3kX+tasxSi9sHdalrjO2OSsy+TwyTgA15ktJhtjykby3E+xnPRbqqazFDEhY1gnk9eYomW8i
RR/HK09yOc8uQ5J6KfCv4ZQQqUAuiNziuCfIff7PMvmc/jFrwMke0CWFMdqZ/oDdV221m50u6q5P
zMuc17EcW8yiqXc+OKSsNDeEwkeAlJjdwhZ/lsBqJ+m3XWZp8UvIF7Vskjb0QUFUAVwpmqwyYUx+
N3sGE6l/x+QsHHI2EH15D0WSDRZkMrK2uRra8X1/ZHWSj+tRgyeNfQcElCilXn8wqTbw4fZ/Yfa9
0ZR1zlUmOpGqe5hVLGKG//aIadKNuRl726d7l9EsQ3wt2oRTpkuMXlU7lDZeHuhXsRzQv6MPdjWy
dSFYzu05+rZ3Xw7u2hoPXwqBykzaA2r5BQoO8DqlHot1JD1o+L1p33TPxwvaAzxPmnF5TL7xmuwA
q7VcX+bsL/OuORsr864tpm5+8nncbHiRcKQNDWlwK1CV9CTuQ5zDVpHva4BWmk61NUZRmao6ygzb
NT9VdOhmIOxrEDcrHhCvDz4J6mWdqNdssy+qMJlJo9mUPEKEPWooLfBsOnSL4h7BHUemwaZsXgXX
cDTHelExWaQ3fFqSWN7xKU8TOJUhJtbHH2E34SdXxac9FYE7L/NPUyVdqT0JxsPphWRZURtf6/h9
IcAoWTDOtQWNiVkFEpS9ZNf88iWECEJQRutiitRRJ3EtBaAhQUOucuEMy209ag7A6eYHWRkC9SJN
/WJp2jLY5gXhbcb1iDW5fa6ud9P7kzijisuyKioH2SuzN3nWVqBPvorGJ+XlQrlNskgxEi8ZT+f2
4OfpigChbJDZi6pV2jhCo497Q89WWAsw9HCLOZzqHkSgQcEkq8tXa1cyis5uR7Y25oTn8e6qM83R
+Smxv/0xM92PgLl5e5kzefXhs7n4Stj0N9CnKoTwOojm+tlQqN7BXLwwsxyobk2UqTC0Dei4oNtN
SSPqJ/QdbM/n0BHOzS05W8M7bqWfKIOencIt7bjWCMk4AzVEsh2x04oySo5yHCwnwOS7M4Ste4rk
6zlKjF664H/+OHvaPR1LIbH5/HX5tj2yDeWosZVTVF7qsU3+fLWgQf8hVOZGe2NLtpvVkFuknFLC
PEr/S/je8UdhbUzb4HJLBPB6dGujHyQhy79GuLxqJWR50rxLXIiJ6UN5n05u9G60fDOY8rvthyFh
XN/5zVXw8NqjOpxzmKkhkKcLGoZp7UgafO/VN5NR9caVWJLs95S3eIhz1Xc0BYgLDLCVnMudn/FI
wo9yOookvYaHdr7TakSAXiDVbat1FKFRS23IJgQpOK58xn7GDj7UftQvF0PBlB4nZ2Jm3/RbxXUX
KnTdXxefcLMISmU5CkSKtASkNnksz+9lSt6JfavOOLmnzEvZlIjf5yIwmhvQw2FASYpZGUm7dwU7
+fSaOqA8YWr/2DwZ4OqiRQzkUi4G8+Rap0cTekVOhAuRmz8UOGeFgoe3HPvvYTgkiqET1XgNkK7v
WIGOhhPr3/Xutq9Vm94W00FJbaCfLMVFu8vCWyuZZ6KSqzaCttjVDEyOjhtfV9VMkR3ZRwfUH2oX
hEujKt5HnA6XJSIHRDm9kZSmrrKcUKag6frUCzzNMq0LrEB+F4LJMFD89WHMzo4yV7d5q8KhUY2C
9zVEL0+8c26UFNyTg7p5upzitTHo+OwTgTmPBTmegFolh+yWPPXyOCD4SeoPaVQM+SgLymSYzZ+8
HN+JcRvFySfj5zJ0ywgrYM6CrgUzKs9aJ7Wop1OgJDc2mK6rTYozz5G72/W8fk8Umv6KKMlob5tb
0qvThSNPgSHvM3Mv5fuPQ1irzlvEcrYUQSYq4SUbVmvBbMJHKv2c0N92gP38SZmYQ9ZQ4FQfuv7K
OrSwrSqHliyoVujRnJph3B34POK361XHyFHEo2a2p1MU0at0N/Uluuo/9UWdh0lyfOTrlxFNJbQ1
SN/Imr5cIlwNNtX0XkmIk6V/2LenegLj0LNawhPXuzqUHvwIM4/qoxS9pPdDgnaJocrGX4jRQ/5y
wfngBJDFaylE+jPVTCP23+EpnhItUHStIAPm4os9OMM0W2Ej1NU0wLYMaK7NRxHTkgW+fDEMqdfj
E83naj7Q5Ep0ZROJhWwrM2s2D12QTHc22ztcSk9xqxzHQQ5Ij8HdfQp8FJbwgofG3NnLhTs6mQDx
/lel1YnFFxScdA2bVYTVEUb6JvZ7k6oQY+vZRYFjtROHblCHLpDe4xjamiom5R7qwkysqvHgikt+
xfxQVw7cOzvjgu0HV+vGnBXf4lv6rLwbmQe9RLqf6sFbzU2VLzuH8ijcL+n6AU5oSGXA8E0riHJJ
u1bghwXCdZjWDEb4uLT1/tPKmJ/yHHCvP+8S+JQXgxMxAjrIpWyTihblYV8xB6vqfhx/Je77Jnno
kupGtj5KfVJx7oHNFFBf/h3EkL6dL2RoudEcQqXkprzsG6WCueZzAzVI6V6wcZrLTFtpM/FIArxc
n7x9QSKv95CU2+wNmSBZvFYnuYIJ8lODkE7gM8niJohckxsaGriW5rdKdgkDE+46HaWxYeZZaURK
ggfFBkD78ShX+GOErl9c+1fX5UuE7qFiAoN59/YclzhCY/qfodRf+qToT2UprkUT7w0bJMTUZLN+
90/Tz26uuWUTpyJf7A/ocXxFPkhTAG/QzDaee5d/kRiLagnTEle81KmTJ2bJk0Yet2SIJxANALVL
K4IWEmMfnIpWWVYKiVuV5ifjmIOxjbaSNgSEMPSgeWHUrvcwSOCIKLFUGEjqmQfFKVGV6yVLs9zB
4VDjF67kmUoJNvVDt5aqtJ/k0sejol2o9vTI2Yw0ecdopMgOIaA9I5piuwo0NHrtoe3Uw18i0HbR
uOdzeSosXkzwFpG6AukP1DBAwmELmK8yNCO3/WBQ3CGq9/fMHz18GfgbaKoYHMC95m7LIq/nMYLQ
O9iKpAWHaswm1KCwQA3Y8zJQVoFNjdjr1WR0irtfev4LX1R9d6qsqcpIEo8HrdZPL1XRksei+jr+
QH7qxUgsPjBPtZGmHD/JiV24rvX+pnS2/UpXIXYvnXiR4lWedqSrqI19s0tL85vgqGbfOV4/tR9o
KDs8kAiYejgdbW9ekn6wtHCfxWta7gLbCCtmbz+XNn4HeRp+bsRxJ2bbZFgA5KA4j0hsfSIjDQ9X
Oowaszf2K8qI2J1XFKmveiF76Lv2cpulW20ryfTW5IPboarEi8mI1zH3XrQPJ76Zp1R+MCkPf7R4
SE7iHyG1sxm7VC/DDU5PrYQ9AdAQF+C7HCDjEOtXdILbcO0zZABz+A6XFdpfX1PKNWdRWaoa8R4Z
oI817XDO8PRo5dyLHitwbAaj+SPumK0SetTbTGJy6aH0YGKZDOFJz03gbjjwZYY6h41V2U0xH+jh
xA1K8bcJZuvupUelpRqs7RnzD3DTSZ7qI975pF93x7FCXUqZCNBaFxvhRpUgqNerRRdSaQVF7aVl
eYJrWA9LxfbSjZnOcEgaQ1v7NbA//XsCqkFKy1NFMuy19AysnSTGh02u22y8+VYMpqS5xkhyVoP6
lbWenoIRmakBeR4C0oarNC6v1KcQFHFyQB2GaHt0dG+Xmq91Aev63aBvhzaEJ+cXqO0BR7mNY5tM
DFlltCykXsT8lTDnQd3tZ1VgdfkOpIlIrrzIqKRYUZj2tS5mmzgP5DW/DWvgV0FxOFGBmx/q5yEn
fHbteuGkwomLXhovWJeP/dAiNcGBq080/ObHcJnmxAMRZZ+6Fb7mudqurpPNltn6+tS5MrFZywwC
3IKjL7I4qRuH8mHC8U61q7cO8bsFvx0cryPoyNWgiogumXiwOgVAb0GGUWdLVisS1BLo4hzcmXqx
eUNFC96Cl7cHB1FQQxYKvCTSSk791XyPBxWbFZCq7gwDSl6ksfVZfVH/CLWXLwLJ/DG7pl9nWANi
J/e7mz9LX1de7sQLW5O6o4Hi8M77pELdJkVFkypW4hoFw2x8WIJKA1ibwqpgjhzCTZLi/itpztDj
PmJ/d7En4XI1IIXoneVM6bpnIfXJF2f3Rasoqlo7b2w7AMbdZqhk/Jsr2kwFOb/iozalkpsZJslG
LqwllMCGPRQG0WOMmzcMK/o99fDF64vZzpF5cwNXID8/v9dxvjkZtkc159qYeZqsvc1YmTM3jbEs
QnBFhQj0R4lD1BViQulzIadksS2t2SE+JH48ieuJB38HOLVfy08ODf4XD+UueODy0rPDWKcXOvcg
bBEfPwm7cA6iQ2yhUQhwS8o6P4njlsvr9ZXZHz29p06zUOn/8ULNCGoFtBb+Bd91XB2XpxoePSQ8
H+KPLTfaTXcMBUEh0ssP268w/C7rKodNI2GbcUhRz2hnXf2zqT8SdT8rlY8qH/gmJ8yNxRRt3WMC
rc61ZMjWk1CgIOFrmswE2USdUaLXufn0yBqRh2Y5uYkmjeNDBbKez0uTbtdvuLMy2Ug4OhQHwSFU
Rwfoqt83rtYlt7RIvpAIpufcKgsusfSFdHdcdCQ3r1T/fKmjhaNsC8eBkxO7CH2cFpbcDNxm/pVP
ccvorPl0gTvrmaVP+5N+CwKXD5nWM5FlQGWVFM+KxFc3Ol3dxRg4BuY20x+00ESI+Cpb1dkIlk0n
REaLvSMhfP6afxBFOVgYDGXUbvfPx88W4lsz2EoWywAkeAoYp2ETgGV4xjjS+u/uHH8myeNL3v3a
Ev1H7oHW83tBpqRwxXjFcC2S722EakhnaDkEzwuN8KWI1iQjdx9BQU8ksHJuwqZG+Pys0AwtGkHw
byxclur6LwrX1oX1rhBF9TBXqORERP2/3ijueMD7X9JlQui9tSyk+OdYLCs865gItRv1kU21ppmD
3RZxIhCX+tTF9iHiyrpu4Iz5GwgtJJyhppqiyysXM4BmI6jc3xri71FLq0qFN/H+IOmgftRIXKkv
XRE5PoOT16I6+6ktsRvaZsIWKrDmtmersSHfwRkYO9s1mecU6c+uYE/cvc3PecaIkxzOf1FvQAqL
0sTjBlC9LVfNP8DXTHCg51aEq6JiJdhD7RoVnU1S421MdJXA6uc9HbNM2dA9f8EoTXpx5bmFguXG
7mqfbk7QKLPoEh2ZFKng0WxSuPk3X6jrQOqJfH8ZGi25BznvkJwX+lTU7WzfDuiGs8x08fXkI6OC
0lYizDQQW3BaDCBXMNGti/U7FYkHgP23IcoBOyPVVhNgnIFYl0zRLTsAiVeczLO38tviciRm/XH7
wYZouG+LXxV3X6GD5yjaDKpF8MOAtHevDuRIAFiPzNMlyto6Pp2ubiMMjUcShxhYnaVI54te4pvx
xxPQ37+dcW+cjqbWdea1ChLtpV7bX0MtZclFQEbOsoxczPPROnGVc5e/3KJUmkIA5IB7ArMZFIym
HVZzWT/eOYi6mbpww1JwY4Aw1Ir0zP2e+y6z6kkVciKII1UkW+2oR8qPivvk1LGhPJ8CZKXl2l54
gWvaF2hvl8Y9g9aVQQha6ZPsMPt92JLGl9POb0mFePXANKeDmMFK0SVEICJzqkH08sfFD6o5FXtt
tl09anZMfElxyK7xTmCjS/5fe13bGG8LldDlC7Tm04lI0VJeiiPrvk5zm4NRDYfnRxmekUTCS5Et
GYrIE4niKUCPDXEzOVI4BJTL7JfJJgXsYsrSkgMdmyBf2YROKPFRCX3ts9Z1xIU/j7gflHXWinO6
Q7I34vKTCHG4jFSeMo8dw61nSO2Boz9hn0+yw5iF3UrC1CFK9zsmzbjs6TYEZED6cxIxnaAT0JmC
wKU4+UZHfIxBIfg59yw7D6cdy3eR2G4fzGNZkF7x9VafLH8Mab4h/aETkTEYX0ysKpYK2N7H0GY/
+qwr6HWSX6S5OpVVMK2O6s+2HR4EoanJ8okBGdwuAf5+cl7I/tmmU4fmNwbJHmIEGvXQRXTAASIg
pZi7rA2eRG8Q68YjwZMk2fn0jkeEs43Ajmbsik4zgTR5+IHTC5m/vmnzBYK0fMKQBNAkPmCAv58B
TSp+RWK9ryIXdRPQaN0310UiiIiChG7tf7RLi+W8uo2JuUugPeDzu1rAeUbZxeh7NYsMmX3Td27C
TUEs1P3SZhm6AMjuVK0spfFbjuETJH2sdeKjdYn0PBvONS9mWIOwN2GpZaMKye/oA2xA8hBzvtuo
Y6orlUaE6O/JUmsf/hCHZV9t31nZMWQ2Xzt9OV0HH8yOd9FxplDUonHt/W9HMelyGFnsYCqW8PAX
Tq9GjlmKEC8F7utgifHhAkiD3kgnH+qNoEVLOJedWN0eEG6lHH8w84N7w9Z9zazfSMKffBBO2SQP
kFP3wK5UKPKgcSDZeON25OaiIMOvzq//7wvmWGX7dPFLgtoO9jBugqlwRaK4gbVVk0YJc5GTTpr9
I2j7gkxAYN4kzjIRi5VBlD6ZLHwFx5OzG1ABJEtO2jkWg29VB8NWT30dg6emOfaonO2UZhcCiL44
8UOBGYvVLLHXCwU25FPRg6t+W6BUAArDQDyBamS99E4gAaYpcEBoQ9abPzJPqH7hK6LssoJY5ASn
PJiiC+I8Zqt0uwtXFgDh8jIxRlAapeWG7YhMPyfEtUw8kTiyhHXiMhWgEXNHEQ9ff0Y+e0uc81Nh
2UDVvoNmp2r/TVbn/RGcv3M2tTDFw3r3t+JiDc2CsXcVA5lqA6GDMimnMe0nfUhPLiO+RFiB6KUN
XKqQR29b9HcE/KoSxHdJig5hPaZIGhuGAwiJy81M21dCsuzFK9zm0n6Olg72Lx2uiAqlXtZim0/Z
5OV+aKud7lUJGDVoKwquC+O11RL/7XBTNg4XnKuYmOtEh+kWtW7dGYnxyfYajG2MgBQNIDhGRoEr
PnPJ6yg0hLRPiYazUi2nNO/xlrbQXK4BzMpyWnoK0heZnvCXyLDcMtTHK9xE9pEpzUvPE46KGP+J
WdBocur+d0yI1M2cD6wlCHIoDZiC6DpG8iLQIII/6gnHmAeAY139mOt5U/Nh9bvNB0A4YVs8qf3e
eUkRjzitcVTDIeVP6KEG7uA1CzaR5CPhNxIZhRLD6j2bwMALXb4uP4Fbtx+dDLEIxuP/EMeGGoR/
Q9BJgIPENTiePtjVeevmUHMkfbtgktWXzFY33CPEuYi/CNg7u1k/lkVHxPPkns0Rj7t5Uzgl4KfV
JDk0cKBPnGD+BFQCa0PHUVDm75DB/v3LGSimFoTQUXXT+VQwuflLK7lSQKOZjM/XcAuZZ5JSEqkc
QWJ4RPyghSqQsletgUedZjzF1OTY01LAbYYe3WImYjKV7FKbLoWWlwqRndzzFjWO445ndOD6p2as
DTWNlw141xv6Nyc43vHq8/YoNbfFlxEgL/+y5a1CA0HhwrROze6/1c5krNol+l890mj3/NSUXGdl
XMFZrFtP+Rio7fHxIVB2YR+0QJfhpSR04GcCK6VJJO6TJE63rIwNxir92XuUaqyzgtc2zgqVW4l7
TvXudhnc2ALGLaEn0NTddlFS9vut7LoePf7WMboxKPhobHOdj9wUuLLoBuQjl4VLUAidZq+XLnoj
A9ChBSNHcHRB6UnoPSfFy5Hfe61N4lstAqeONVqMdDuN5BZ8W1+WaRHGsU+6dTNgEmDPV1zS9bJg
iYifDY8+w2Y4H4ZLOsZhw3AfUOUDdv7/+tyKjgS2oOy08hKgtUgG/pjKWaFHhltGKneg1DV5dvaw
VDt5575K0k6Ljs2d91B2+Yb3refEdoYkuchhFT+a6wx+Lopa2lYPov7DzGokLn/JlSfQk35uzSCz
CqT5HX1P5sW2StlTHrzoIyaNXBHFjqvwR4aFDhispRMJ+wOFPqeWohOz2JUrsMM17aG4mo41u6R2
D1UX5LJWRh0NDFJcaFjSuZBu5vw/g0iyBQUxGfulf18WJ/uw9G9VhVkAkzhT1gUZNEeoG3J+B2QL
GiDhDjyk8O0iTO1YKQOdeiCq727g9iGAZCN6ckem1cnQY3SJzzd4e5JwsHViS5muqpqGfLnPaHIs
gBko6NegMag5u/NSlojl5OWWU2+OdDuwCNjl8CHR8jEZ2H12a5b5M17Q9WyzHQmQRWkbvQU1e+Zz
1VyO80w4fH41PHXcvqbk1VzzeT2jnzJQjvwRkdRB6+fT71pJJw1+jelSD96d6Cg2nfGmgEOCnUbI
fCIJeORDSgwBfs3tZjIWIz94FFUbneZd3r3wmKR2nRHM/OHrrMuVLOiI3UT6UrqKKVvp/6bQBZiJ
ImhBuAgJH2QPr50jakR62TEoWcjrjU9r+55Mit+JcjWOmdr/IpebCiJcAUV2tM0v0PlHhtlCEpD3
FmW86alFmCR1nnSe3UzxM4LECTjQlmYVGmu3sAHGvy2SWTEmo/vGU4rnry7vdAqGRNMkX7jCVdf/
Jo6gYTNU89AV/POYj1LIBArKUwN3oRM5STNtejcPtBkzbgQjfN7Md52r4V7+Pr22dJggV9wwq7yC
NhpN9HErcsfHfWwyWQpb/aOzurdZtWlDqiYiaDc1gpl0XaxzGPp+klQVQQfJNcFshv3l7CqoI9wc
BK8C0M1eKEkdJQ5zyeBKrCh3R/XYNI00iDZ30W6y5xEXzBORPqmulspj/Wz1Ie9hLx7Y/HymEK00
G6taGiRTv8nr6heyfCXhHOEGsGDkH0Ve5IqQqx9OKIFarLVfxw+JLfc1Lgg7BAajiL+n9BEa5lwH
stcgwc7EwBXUVSkLbeg0dky7vT/Y7ux/f+VDZUyfKpJZOMsJzSgEn9jgzCMh3vZAGVpkXdf1V3bR
hEUNNlSKFBwKGqPvQHiOmmjcx8fU+OA03XSnQpYYTKrO022Ct9383l96aB9ltWQTHxhyV49eaIz1
93Pn5VwgAbSOreloIbpxzzzozRXoqrgu1YLm6w9LrqMLF6EzW/GngIOJk4pzxEK6bazLA2aRlxHb
0ZglA1pEGsjqJoh3tpPkqLSxzua7KMCMpRYGhnW1KwopV/vF7mJE9d6g20biReC0CIj/qQgaBX5D
mcBHqVD6BPlAoDudM5fCGjfT2BONKJxL0IL8a7nvIQrXiGDZn+BSnHWxfk766155IjTIsiPbqub8
vyQUZMTJDTTiIvjonLcvsAZ+zfQhGNNEYzB11Cs9hdZ97HjBQRHOVy4eGVxieqWgiIwnQgWY3bqj
L31XlrgHi8EBknMMWgjkUr7u4rUsZfpdUbLcKWrLtnmArB83+vTvDJtzoOLCOQrmXhQiDXHQS9A5
u9XZ589CnZaNvtR12VYibFYdTpFxjacWKiWqOxh+gzOZ4uP4JuLDxEsNZgGBOydsJqfZ0OshiO9v
jJLfJ3q3WFAjXcIUJrJEiytBS2WEGnhGUPjqiy0LljGRLQiZsLa0dgYeGevrVxU2Y9bgXFQ1wziS
EjWlii4IDOioW7TT3NCblC++0poLqHc9Vf6WwRmQNEHUTDk+I2PiTSb+iYM6mtwisolcUJ2n+vYD
zRlKUnqFycjSIr2KbY+TwHtivY7t7aMyfKVUlhy9P+FTGp42Uu5oaULtWtiihfDLwiLfHMsCjz7p
lq3VzuqXM7xEJ4eVEX1xh5/zxnyS5z1YS3EB4yMVID0S90AGOJqpHZYFlrpvsz0MKjkrC9aHh6Zf
z3O5fvbq6DsPxvNb5+WNFNXb7zQuTT4qzb53nl9DUTcqmAW1T+2coT7l5JabQGE+8TySkvZbFjfN
NZaiA/niT1twbpg8jOLeS7H+KVXAMzkN1XVmxkse/ZQb82CVYxozg8gTJCUohlruIKhY8YRva+sF
odyh0ws5o2kOUtv00VRwKy9g3m97ESvlsvxtgXuvTnxOd+bmsHU/tgqKMCdugSB6YM0AkNXbb9Cr
/1jm6Rr8iGm/yJE/uFD+rHRRvDKr4dNTWi9vJzf7DH/HzJFceQ5FQv3QkTMS8KFzlS6kEPl6YbuD
9HnMt5oIyV/PryZHXZn5nrnQcGwRhYX8T3UZ/4lupxyItNyipyGalxEkBD6aHs0b1q4c2PtoKxgN
dwIP0I5PF1Qu0b0tWTVFWlHiP+JxUW6HOnWWrTucqXVXLMPF+dnccxelHc6avjkssczx3HnxNcjd
kzS+D3TNY5+yqF+o5w/pqwouuVCP8Y1ZZvapLZwyjLD4Ftv5lsa0s+KLCY/xvhcfNxmW8B2+tSt4
ryFZ4ZrPiqFYDwH3F5nSSsDuG8pfLd3MY6m+RmvAF6JzNPa90y5slVhITANcCpB26Dw4uj+nF6Ec
aQv8GxV7zsHFS7VYGQRm9NrUlWT3Djl86c0PWSwU8QqdID7BvxeB74fV2BxYRzCaxFLYkmNbl/mY
FkJOHD/2m0gHERbl+KBzWuPQ3RH3ZWPlMGKl65SnDN1U4JFVCf2CyOS9/Mgwpe60QtUnbPLq09ei
u4J5RmG0lzAbjGdRcKqMTVOSZGbmK7erChtU17e3r2l5kT/av+pfkWsn2/LJ+WAuE552LN0+0HW2
4cd7vf6RLl29ukpJ/mXgfIcpxeAcF5UEwJxihC8hphL9bzfilNUzKd+nX3HbAKvyDy9hSX50kx1e
XqJEZbFKy9sVwaUGE3uGKx8PXJXsSgm/p4ATpC5oh/wXQi+WlX/8DTNbr+zZ4vDa0ZbLaHFC0UaW
J3WfWkn44fCb50wY4TyRKkwLaTher8DwMYk6RQV1xO4rYiJSjxol8dO3dKyw+N5j9/dIBOLoEJgH
XctEQyzP6N1Sj715Y7u7HVvOlDFTKZki+B4BdXupBEPwDBNg6EH0hL3QSBCZzXk1YuyseNA3C6TX
dlQNuoR3FOSdWOKqEYFea3HBN47OWgxiEm20i+woFl6ehjxcDNsXWysMxAOSiSOQ/+Pc++T0HpAf
3MeAjzIdfOGOXn5PSEgPUT3cS6ABhUD6KjyMFUQ3zaIKlzer3gVq+TPTTh0yu8cBm1IqE6zDHe0s
G53zYi5j6hiFiIlJQc4DOkZsBeMlTrjWAlouYmF7tfVCU5A+0nkEe2N2PGMgMxShvk/EL4qsqjft
e+aiNcwGeQlFsa0pqYgwXSrGdmBchHT+EFd4w6KWzU7H+9Dc8EibWFhHdetb3q0e/AiuQ1zxgv61
jMqhuqbVuDTz1LSlIg04iPcT6w3jU3gPb5F2PGRA4tAQ8dHluw5yIdrCkz74qYLLBk6CLGclwVVa
S19UeoUe85beBAHuo9ltzAjuS9P+aNVxtml60XVhhcoHeZJcfO4FQRCNu31G+YCE1nPuljFOyuKO
W1N3o/+KMi81kwwjooh4aCRBFr4onl4MTlYJeZpRh9ZOw3wHxUx5jZtrJHFpUu3TL5yIaJh4f3/D
jbeUHl494JwZo1Kwi+EdD1Pf2Uo1HGLToaBfdeI6BI791xw3OfFIYbiyFT0pB7jb3Rrbn9w51812
iYauReHM97jbwO6HVWBTWO3eYEI/AbdN9vh2eG6x4JGw60cPmK/kli1GQMbzZoawDTkZBInewlha
DPH7O5OkAOLiJvLF1/PHjhL/FjcymtrxYkolOrKO+8v/f5qKX6Fzw5bihfWbPBcnYBBcmcidkclM
9LDLRLEVTrASl5YaIgyLY7Abf60Mk0tNt1xhjZyhIgCGIsRihPHESs0RFka8xaAldy6zL7zwWJQd
tsF9JtyfPWyLNYsLzeTMj8iZtdNB7DdUeZnT9+/J+MI+PIvhZwdX1YvFUZfRkwZqNyCwxnNjmhAZ
S5inEE6ioLNdqDkrQLNtmB15dCOQ6RLaR/6KG6+4dVt6remewCNoN08EAgK2KoknmkyVbttpMxfn
2gcG7WC2+0lJ69P5COJ42F9+RR7/mEwO+raNEC7eY1q7nEz3GL07mSPmUthK9APwhysAv6wlZIGC
eqYx7XQ7mG1eXldS1LoGlrP9bl7KfrQSGnL5OCXhkxNlDL628SgzYBoI5mXcWXnCZmpHgJbpFKK5
CjFi2yaN65BHpwuk1Y8gubYMCkkLrsOIQ5RuImu4C5GZwILSVIP5jlcO+exWB0fn6dRb24Lu9QCG
a8B81bE33olz8hQeDFE4+8yFu1aWdqDv5XGYjSuMSVV4P1GGAevDhqXvcxrCvzMC3Y4esOwdL0Wv
D/4S8XIDgH9pCcT4C3PW18LcFNWyZFPtK16S+I7JwSYvRLAGTgCEc1WolExl69dsyTzBeQcjWAQH
1m+MgtVLjgI42RVuTJ1lAy1P3CmjY9UNaR9Gyv63ew+YnomJAuWbpRKzH4GhptWWkG6EKyr6RIcI
Y9qAqrtxaJxHhgMtaApBnhiNElwdCGakcwqmbRfhiw/p/VkHZjmFJ0dMuWELkCzFTpO77TshoEmi
Q7x04Gy5peogH+8YFt2+XEiLj2lYl7vu8mtDAozMN2nfebhlVLXnhkqFzJQFHdDqb//eHPCbowkS
TuaCFEgHAriIntoUC1vnFmukbCb87edSQsDu9ZSzs92Y4ToxYtO8/OqD1S8ZCIA6hFGZ/yxoNiqw
O0n7zehwNyGfOOUv/3jMg0kx9B+ELAmbWyIXkszl27umxnnJxUazziJOYe71IuaGyp5Jx/xihJS3
OQ4HH7VFHU4vMw/MejnQnnIqlvgfUSHzkDlF0DyS7o2sjLywkjMsAUueLK5XtfYVP569E7kt9DDZ
dwfQGmHJQmjtZot3wkvsYb9iLEoFiN3r8sVVJzPay/3m0eP3T3vQZSpY/MgfDA/GI610G1RtaZWe
BahogVGKQJQMFeYEDzm/Yg1ZXOaRqUQW/wzHu+71goe7ZRZZDGTz0JrFQ6p/xQ0ZhXlrT9BBfJ9+
shi8IDBdcPTySKuuZvkV7zaLXF73SqyfHBf9gps9IiiCBpQazElmPD3S2Qa1+NaxpFiqCLB+Qsni
UqOOJ2c/ff8rJSMK81HEQh9cm1sGJCDXINL17USSIUh4XmEtRwfZbRPMnZrTZVRoiYA+v1Cr3BEh
BFkXErlZ7/OlumdzrRoQ3Pro6RKgLMv7TcJLx4jHDkarHeNSzNSes59SjeUukjt3dBnVwAJ5md4l
e+Onnxs4cz6+gi2WV+KJQFG7tutmLW+WkChkS7Inl30difZ216Us+YaupUBpByHjzEq7hiaPYxfG
yoInCti5b4BpQgjv6K0A15cQaRDwSA7ft3Bn+5YP4IwpUJ6jFdJOWM9iFPNbpu/XS6Eocm05R4yv
ntFh9lR+wssVl/1E24pl/P8GVszmu+qGOfBvlWZkcmwONkvrUMYmtA1E0WE3kZr9izxRN1N7a1uQ
8bWCc5jLhTQAeCeUwekoY9kNHxphtpGobOl2ZxBGwCjBlfk5DnAPflZqcGtUZQ+YAIjmHYFNzBLr
VlcR4scITxcqltWOvUnywHlc0yWdYy7NB0pj78KJxxdNWsxot/0egXXXHXGOWmoKpDonYJ91c22j
SoZjm7hfv757T5wCYWISBCW4O4DX4vqGjNXqOQN5c0zqsJxvoiubckP3Rxk6w1OMWseOOvWHfHp8
H9nu7GoDCkGvOYsSW+/yfOOwLPY9ekPKHxX2Z4vpM1k6AbYvc6dSwrwqG+pWFiCkSyze2394qY4s
WFqYk1q6V9Zbplbvn/NheHScbSCaAkH9wecLfdeGOPvGwxMxgbKn0SU29ouhVri1FcxRwOqtv/zu
0y2VwgF9aEsKSyGMk5YV9EQZqglU918vvpqjBJau2lr1GL4kLJcaOXgimMF2o/lRbJYOUTmsPS/V
YOnOj6D8WLdQsBA1qcKL3YX4yXB+NIz4kqzWO94CXC75P3nY1cxJMzOpoZh8hMePSeK2ubMztbHA
ZVJ88CuSEORi/f91an80JGeLh/KEIVe1ferWaKq9KLU8nHKb9JTRxRGlXZtaiHhhkgi9EMPp4jWE
VTmv+JQaRc7/RuSd1k8Jdvts/Q5wAlYZVNBaRxt+u/VLIVq4ty6ObaPBLlR9/BOTZFDp7UwIEDmD
xhCUOrzKmgcNG8uhNvRZ6OQL2ZHRI+g4cw+PAii8TlwxeET7y7+q8+KCeBP1EdRiw2BrRhi+hOKo
1jKBdgUxP1rBnIFW2rgQHU6vzLZCaB6sm5E4A6CFYYxRf5WKS+sYugmEitNvFSC8sE1YLsEuQOiR
zY5FE9V+Iw1i9Eue/ZOhM+JNGCysQ9WPTZoaTm0h21XVVzWFzlq4z3GkIgvAhPhIXhoGnYbTVDKW
znZ79AxHOvHHeaWJLOde0ehE1DL5mdEWw3ZlYfMk7tZz7nCbRhDTuRlfmjqEtBXUdwTNtgRK4s9N
iseiCg3EX5m/5piSwWcAoHAYwUslbuPV7ZvtZBLohjXKcDH1EVqcStZf+746isaGyt2Amkb6MJWm
r3nmw3o7BRw2M8uZ332HD1rAXhM4rQOWbrUQIKfF0LS5wnJsczpSu+C5/Rc86NVwqw2y9SlmNZ3K
JXKvgBCKpcAB9YqJ8Pl3iSjILr91Iyd+v46+SeFemmqdpfmGrLikq9Z6OwBBlsuuDbG16TelP5pU
P+4aHno03kuEV5Sq5vVcOlN+ZETapAtySnfYcSAV+COk0uBJB5svr5VOrRgd/uAheSnM/WmvRrsq
0sbR1FJKxMr9I2jisYjq89ZMwfxwa0cNpEPWSp89BqNi8psKhnPlXL46INJCIWnGfsJgvPRliE95
sEZpaD71jTj/hCH7wYsKaDuAwCbLheDea1uwbWKV3XBZ0UUbeIapUcOi0hReGg2NP81in6UgBYgj
rNKxL1YZ0/8vY4ow8CD9sq9ZXr/cDZc/JKJmanRXV9r4qV78fV7bAJq1+9wmMwEG3WSK+YXhoo0P
zL/vzvataRz95cuye8rKC+oBXJflCxRtSwHeFauno7hBcBTuXQNPbZBTXx2ayj6nzAcnzk/q81+7
RtFuANSjalceh3JmUGCoP3czMUHm1EFC/00xb+RLeGwFGvJTzHH+vn62LDa8rQOf2aYA7U9o7Os5
ffi10dNmHm+HBEMXFXIhv8OIHwvJjpuhiGrmsfe4/OKMvistYncMzGjcQYu6lIo9Pp8HQLuxRi/A
p+9LW2Rosp+v5uQ35ZjhZzBq+pXGVlB2K8QmjaoD+d4jA+BtqwgIGlwON7dLM4I6q8w5VaQafeCS
vzHp8FTOU33zbkkNGjqr7tr8CC8gaKFNoOW1FwalGbX3RYtAQfGPhfeNqfvFUZRZWcqfTe+SUs6i
8BcTSuZzuUscY4wUubuNx6eL3+qIWMTK7qvZZoSVx7jVE5l+iNp28epCX0eWJ38j2N4utIbdJQqT
2124Z682q9hyN1Tu912LHnPIZl6irEre+RTf4F8GW777NFQP+sem5zeyMv6iFQ+iBnj4MG7ERxgP
qx0YJzBKDFrCzMMW+siEd34TMxsjPxijto2AiOoDQrTeMvSeabKufRMqoj0HuWebq19xccqPotC9
JXmU2Yw0sgmyUUXbLP+a8uB32HTwEHemlDGpXyirPIMe/0oNDcxL0HxPDu360QgE/rERjzWBL8oB
J0WYM3x0v92R7kHtZtxUS3ipX5f8KmAysRJudfB8fPX537rtowrYlDZ1B5UNT9DvPeuy8POK27mR
wBoZRUqNBtO+TOJqwnEBkSUamxHZY7GA9b+37QmDJoUQshF8NOnTymnjMgeKV8j6U4QsAjICC4UP
U7l85mPwUTUHXmc164SYDM3rbldYIcz+ZxkxSTN69sx+VbNfJKFaF1BPRvMC4saJaDY9lYZBeUur
F8EZf4McGFpcmv3ocaMimzIh4hTzhGSju5hn8u+VnxmcJ+VPCz39Th0xzjAsR/4xOWT9YXIl7ApM
lSv7fwMI4JF1beg4TCgKIzhlbvqjf0N273kz/tWvA6kv0MbYURSzThNxJqCYGat2kejn0Q84u6Z0
bUgIkcZLxNLt6YR8KHU7SjilYq8ZcDqSrrI4gAhoJBVSVKu6jJ1ijXBxhBdH+xBPvPY9dskbmeOP
R9StDR0DsTBMeq1dYusCdh5a1P9k0G6eBiw9jdm9T2ZPoWQ9DjSj18ZVpXXM/P1evwoV6f8s8g3p
6Bixff9XXcORl6hLBIi5nGjO9GyIHRdpidQR3WEi1lTV7J2RVDwr+wC25SVGep4U6Ysg49dSfHL+
+HhennL+ePod5tqGPs1NOFCTyJ+K6JDVMUzJXJMwIbj4iRxhtczwarAFJ8L03PACxaM9wNX+1E5j
7WdqxG3zj1qNjWT1RgX5UDYFbm4/PQuyoUDve0vqlwson9uNPZZM7Tl+4RpgRi/+3DFyPpMV5FYU
8omu+INpmtBZLehcA7l6OkOTHY91hRio1/DruAXg/1u+TbzB05PZRCBUDi8TNGgrBS8etpjZsQSf
8l8zRQyHtCHJGyH+CEk7lP640t2nLeIkHvWEYtY6oeAyPNlAJ6fsJw5cKkY3sucljDRu1iDfX1Ho
4SATM0PJrApvbHig+UsZD6/Ctqxq+CrqxFW1n+H7obK54n7GkndFPCJ4hRyeW3LIlHZ1EyQdny9w
D4Jr2SH1Y6C5Plk2PZ2pbrZfAQsgS0Ak2Q6W8tdizY4qRhbnKYjcjXmSo3cl0/kx+5P1e7pg/BKK
eLDGPfG7cpBF3Mih9Cu2BoLlwbIIoY37tYJAyyruHCH9ZJEQ3t+art4GlXKhFTPHOyOxtqChfIbm
pno/HcWILsHPnaE3sRPc39al1rUGZoWT0iRfpKFcCZ03k1NqZ9mcl/UegdmE8aAqaObHkf/rvhXT
Hvij7Divc9ywuwGy73I4MHjy8lQo6fWB4WAuoA9JdEai+l3ytwcJdHFZpoPpI9pavIWU6Xq5zE5r
xYh+4Yzq4PIsrZFXjaG/tuvhAeVo5/Piy5u79MhvxsslAJujVJMvvbHPVVjxipAyAhVaTXnrpiMX
JjB1zlvXP5MOoc/J5MSlhLbMdVrekRXtmwQw080odW3QzSDb6XYraGn85ZremL2N/mGDgCuF92w6
04uwCfqykuLI92CxQgPqwvjhGrM22h16ByUp4jSZzxaImhRRfuqhzV/js7i3L2n28lm8kG36M0J7
rXkmAG06gZfGkEhneEAGEawoiNl/p98n2ufKogtfPHJ9XIf2xIqo3XKJzAF8ijvAPAq6Yv/NLAhf
uM7HvnvNwk7JsnW+8s7/OHlMQEpd0tbyYuIS9pdk7qUo2ZM8kNNGPrx9QgIs519SpGPJX+hlYJz4
/3IutfDHhsHGrpoDLhaO8sy4Ovqi5kwyzZC+DBTP0nnadC+8jOU4f8/2p4zzxObKw/L3ZpTUm2fD
M5W/XQo6I8cCTwCTcEyOqTrgkAR9G8cJM++tef2WjpLSbY4nPSfsDYHfyGMUfV3K8RUBxICWlkg1
gRGNlQGqJ+7k5uzj3yuiaLV5XYwFyE4YfwTc0pcNF7AbcGnhWueJuuYnsWxZimd67+TrQl2ehqXi
IIvFOnkNzJGQj605iVUY8XAVAIj3fJ7ZBd83amPGsb2K/jN9LWGft7BicUaodj1g2SQBJwBoy386
8Xvv/GeQ6KpDys2CtD3eCv3EaMiIW1P6X8AkTRH7b8UMMhsnas44E/7kR0dSqzdf0vzbxD1lZuyr
youwnUl2JQOsI9QVmYvBt4Vv5IIJU+U7r+MkqPNj/iHifyYoa+lFDdQlT8qisLR1utoS+68vIaZ+
o0P4WIyP/Kk/PJxUkInLEbvIJD/ADOPcKybVR1y8ipkba0gSjFpQ94AhCB6LIhAj5EW7nJdZhhsA
Bi7w/yhNEGAQzBb1s7YMDUPlI15KL2duI9stZUq/KJHpPXDHBNnImP4LmS11hA4goeqoCHSpgxBE
BfTI8ZfpwAXvjGRih2ikIGwTJ8kvCVsB9gMpv2elw7cy0oDeFpiaGKyT4XLoXJ7cy2miuF3bpkeG
RA3A+KVyYZNsAo5CJDDnL4EWc9Z5bpr+isNvQH9kSmhPp3+05xcA6IF2kLSOfhjSkiwdDdGykrRM
hqN3x9K4bstzpDlR1q0AZZW/GVM3sxRSNFA6fZyiFesHbbRApRZG3iVJLs9nomnm99QLc/OweyaB
i20T716TgNj9I8/WTd/LtjxHHQRSuSfW6DAG42Hda0G1b52aFhflrkHBP2LqErBIFZcxooLFlBhU
uknq0oWJ1dcFjziZ1P1C+Wqd7DHNkWomzxe4+coQF6yoaKCAnmPn+iBfLrUKMIkBtni6SrKekIVQ
RKnN1p/0LRyLE1vk5YFSpL8sT/0YmI/RAbnBusXh3sPgi+zzSQLZFyqO9cWKun044BsNSHdFOrDN
2lnjh9mJB3tzZZzBRtQjqbsXt9Ef2pQ3FmvhmX3oFqJ+uldO80iWU7KnXKOL7LizhIjR13HeAQJ9
nipUeqYaqDJ6jhd1IiTuGrbi+XcSoa6yKVx6wQ1dhnbJdyxtAo+vF8lDpn+N/ryeG+b8/GOPrLVx
DaA3BpR/4Ub7itF8jzdNV8pMjraQnOgxMi3wQPNhdh7G23uq++m6t44jGvGVQ8zwkW2p+Eot6dA5
ZgqPr+yuJEVnj5fM5ocl07GUlA6bQnPi6hJLxgOmQ6se6pQGlP5SuZDizBH+3rhL59pINDLI+GuB
KtrcRaEMJA8iBmXw4kXM3yB8pOJIIEVcCeY/EIMZubYQdcqNuyWRwG+j8Urfp0oyXMTNsPLLzcio
3TDw2zObQvQhgX3rdvHZZXxsAioNyRiZfKr3yDHL0QcMPrNsWL1j4iZgm3ItpGO/JnWTfXlg3brb
w5uI+yFCxlfDLdXOsaHnpwCsTHUBXaTV+9liC6aOOLrubIHgluciT0FhWc5n0J7ieJDGiBtIo49+
cr9YrznK3IdSXa2alXLAG+4fRIxLeinOqGu9gVGV7vVUWfEJ4HPnpwzgBCI6GvnAkQotKSJKCcic
dOnBW/wJEXLtfNBCeuuxQkcNJZUC0W0/iSsf/WApQ3nsO9z0rtypM7CTtRx/u8ACOhBWRQB+dfUW
yUt0idXEg3ixM6i2FCmATd/6bKA7i+FW5gtlLnZ2XRaTzFWjjQQFKeXJt2iZ2J1jFGxNdQt75alE
cy2Y3F2thHkmjt5WNjysViGViAsA88sbfr/gplfJj3x8lINNqNh4fZ2/VpoK04yJ2TCPfsvgEvfZ
QI/Lc1PkYFtsFj+2LhUipMwhvp0VOLPhDhAgGKwsxlm9rtBKBMV5fXub/lRMg9sRxbHEhB4R8Jen
8q2nvUZtY1K4Ffm0cB+e/7V/Q3D+i+NSvmSnTF494evhtA1cEbaGPbQCuKTCc6DOeB382+u0zGzO
bYtexve1BAIBCZE9Na+FufU9W8Q+LhuSMb21LewURRRNsTXgnKfF8MduSaA8kuryyqLW//LNyeP6
SHr6W2lUFmkuTFs0BnUdFJ6V9bLhfSK17td+RMu7UJKg4E0X1VoQjXoFqGjilqDi3Q5rcr+sreum
J02ou4Er9DINFnPHsMdaBD+oC3pFEZNvgo6fc24ObRopUU1ewjZdDBTDQ08gwY4i+K0o46opKeW2
Q+rD2BKLauwhy1b/hGUce5GAt/PB8ATxm7Ug7pAX+ItNqHhuXvpdlLIuiF9CsZIntU4zRK0otBgc
VU0HwqJe74+XQkKqFLDHLFWfYxWm1KoTgFSFIJkn+F2ZAD3RK5LvGPMOHfy49XG8amF6gYa+dNT4
o5/BEQRmsPt9PIkeZyN0NkUOj0Jd21b/JI0yTiy++eNrCEPlm2E4+vZZ3w+7rbgIp2wBxKjaXYHo
FbnhjE+zJ5kRlxk7tmGEqprDtpI+NoQTFf3ZoDzEtCvb+OoMAV5Zpz/Ov9taoaUvBHIbSMk04Ccw
M6u3b6fOByPAeLM3RaYrPY/94wJNj0HTuKXtIOJZRGw0YsoembMbQMgrWNjffLa4SKWQJVzWr2SE
0HcQWNIRnHAj8Qme/HFACr91RgrNbcJVw3eQSgzDdRywPzSt4E1hPhatEVwlpXFLn18mq0RBdovj
aF0bx8meIjPo2YR9C7cJLLIRrZoNCuZBYsLmIRxxjGfHGonYRvZfRFnR5Q9OTOeZLsM29zoVtn0s
NU6mHdplDLdHZ9J/je51iFNuL/5bH2iiT2WaJjuOu64CPAys3cKvk7Mpo1kt0HylDyOX7B9xsOSC
fZR/0+QU8++bAdWj0+b4epiD3lRRRBFg5KqvoBW5e5XhXyoQRyFy00S77PI0XqvT23FxlTQjLSTi
eFDROL8jPwUDWXx8ZT7547QfVc+Q/xiHHzk5I4AGcTHMhZ9PPMIeeWSLIQBYpFNXZHGSsQABTe9K
z/KUawJseGZge/9iwuWWyWABzNNgIN8M7qGQ5CZAphrrkUayxZrVBJtRdgJhrEvLGuDXal3+6eOU
vrCpe+P4l94SaHExnUxwZmyilofV47FJEMwrn9VINFx0GTFND/+pvzPUZFQaKUSFdhgJ/fdosB1u
CPFFf+DmYzB7nmbewgRJT3O9ug3EMIiaZ6ZzOjX8FAtJ8pIgOGL+k/oa/Mxjz0fyagR1TIr48zna
A23q6LSIwe5U7o8tqMg1IJvr2w3ti8cunRqSHUcUWYF2vnjAM+b76dLI1/eQ5wFvVfY+x1s0/arm
h6c3RzVSEsX0sL4rk7i+niQPWv2U/oaRxL8jL56BainsKpoOscU/ZBmEtZxkzzX9aWh1ec6z5y61
AuwowFibfhK31dIqAcgVB7Eye4cpTDOTS+LXlfoTdiSylJE5FD07YB318U+ND3aTVWyiimXX8E2B
TO4dTpuFxiyGH45ZjMbTVX3jK1tiNN0SE2n/d6BNy1L3HC3ZdP5IFgZemLK4DmLZUIe3VG3zGHz0
AJab4ZsWynBqu/g2mpoiOVTjipFc0xpn9/SksOB0JLOrjJfXeeOU0JQOEl6oQAsLzV2ulxFKUyOf
bQZoyN7sg63FdjyebaEt8u2wJ20ZIf13PfjDuigOAVw+yOO9MPQmyQ0wjbcEhyrt1gll0XkFJ5eY
u5GNRQLoEywyz/gyPBpV8kSkKbRXFLayf1PyLbf+5Fb2DWro5mJFeSoQ51G6AbUBXPM+0xtRoLrt
BVL698376PVfnR33p4WOhOqSRAdoiJ8L+yAXwT/lZAp7pBSM/DAH0cgqVk7FTdALsqKyxEOWNaZu
AnXZ1bgAtl5nQKWspEhW7D+wvK74l+spCvNEXJXZyGLRBSkuY7w+qEqjs9BtaztbU2CYFLHwAh8M
h2Z/U3LrL2/o3404Rwq6lA9itI+4m7vVtAg2eH/qHE2GRXHqp4mgUP9h0yMXQLFaP4AGD8ZoBcHH
jUMkRCVr41VHMUa+F1SibIyp0uZVkOz5ke9G51BhlFLbhHOVTCvckBj+KNWqU0CcMLZ4L6F/opLP
V4nn6whS3O3HZ4zHLNw7d6PMqsXGzMUYdyJAH+QH+7bIDC7C2VTpPgwBAvwBOEufy6/8IfxFgQXw
MQCuVhVyvD/EHoXA+3OrWHtTSNvRP/MLl3yH3nqHnV4MFPuH6NfeTDtb/CVwtFSRqiiNwSmzd1Yk
WeT8KHgVWrT7yIw1sSgfu27IhB2xtxxiyAFs7rSr+2AVra4IC93rypc4+lm2GOBBtV3rkzK1aIrR
O1+txCh1TQ1oGXFAIZzXke9h4inIsP8OJ99xmjjOpEe4ZiwOn9oGMfIcRbLrUhJDsNtcSvYd5/1g
WfUGhwe/paQn4hOky7XEhRGuhAR0kjOnnqbgCy0qkM/4XwTKZg7DDLGU/VKe6DC9hssmCo7BUMYY
kZ1IWWi9NqPxp+SDrhdrrb/I3V6p506ZIwMQu864kpsYv1paxzonHhD6IzqXWNKd4Ulg75Byr9H7
DGlFKC2U4wJmtAp8xbp23z38Wi9jdzLR2NDJnIX9TodMyftSBo88+a+Wv1369vVMuPPZ0lK7yq2o
4kLsKT5Ul0FfDcw3g8wYdF3aQnSK3+SLYEaGf6HH017ylhlguqyPO3E4EkNxa9nkExAIR9cJTQhp
GQ7GtLAEEztKaAk7M8rfw7DNTez8K650464D4hJtFTnB1JHEqu/Oe6U/XOSWdMlszuH7Tqvnijbw
e4Axc9/wVbkYqL5t3ScYhkaAZ0WOf8beMYqF2Yg+YCOvjKdxtKLE93NZxAURCAz+Lg7i+GJ3nTVR
WLQ8vSDpXttQ0syEbNwPDS3i87cKnc0pAT+NxUxkfMa+lTeaiFs5kKwZBFGWiIlrqBHsBK7Z90nc
flq39TxtPwQciUmVOsHRnb9t6sAeOp5hfOZl9rL14pXeR605pAGs1pVYyUZb/8iBj7MjPqa0T8Zt
uYZNkyFoe8scrw9O8Za5JFjnqPkusPQzPrUS/djS+c1ahuzZ8D3XyObQJwlA6VZrsZ5wUhdO9Cwm
pKdNVPV89TRpjGDWWEdBRLF5CygdBViXUYMIAWP7+uHw4FpwpjCStbCR+oGIiF8ndGJdxZeeyLkX
iBSkfDYvZAxsw2QFt/Z40v/0tVGC9V1hdJr7a555volkUgL729pCW2mBv6Ix7bIBtlYagdrizNy9
I6L76E3+d7iHZCfWt3ncfae2iHXr40yStwvfyQnWAHj7FA5VUs5poDahirwSz35cXCKokWrAIVQ5
2vvoTqwvcI1QhNmR7drSxYdv2ugwaVfPpeB7I20OcIBET313dJX8VFipPm+tYfwqGe2+LB+gwGNS
pGI4avpUrgLnXZf7GVRWL6eBy7vbhv7uacjTV4/Ry8FPRC2EnNiR6fFTTUeAbE9iV0XeIc71dUiA
0F8XR2QE/FceeRMJQHT9YvcdUahqw8K1ZkQ48MQeT07jrLQ9HERFMHdjirjHwYaTXYPMW9LSxtoY
dTZxfx+Xpv2O4MVTyTfYzZvLveKdMWk+wqu3OQ2Lqo0YaJJBZDBP7CltAqaz29JoiGNuA9R6gzdT
r6/PMjBfEt7YxnNt4tKii59RRKWK+SwY1AOhcoT0cOqcy7zZekcuI6bsXm1zvX63yoL5GSaywuJr
HokBW7eB2Nadh+UIPK/ZyLMl/fzh7yI1jWK/H83Coa8HrzfiGRZpgCc8t/6E3I1MZm/8wfB2pMs5
P2txdlQ4yz98cnxg5KVC2+UqP4mkUfD/8Ep+0W/bDXKBcVRBI7YtGHpMDhm6ZNsbW1Ff0Mm2MQfq
VHuABknjAjf8vi7aWneEZmY/Vt+uPDpvX7xa9mPbkjKX5kCJcjWolVeAVpanPS8oXYiptNXjcBeA
oxslZC2u6fxdGQjm670U297/HPGETChkdzLCSVDDmNxddvMBoUvHaob8jz4OxDMucFIJeszh84L4
gBu62EXXMu7jweNJ+vczZvQG0zlURw9OO1lmlkEh0lSAdbkwCZRMAJbv5z4WmivWMwa0jUXnf2/H
P5AFHTZFatYcKR1fIx0FAOWoRhzClic3FXRgtPcqHGu+K3zIFBUeJeTC60kAqC8bSChXha1ynKrF
k+L81dqcH4yxKotPzsq6q/0h0dcQgLkQhrnL4qLTWISx+RyPexjBe/Ajjjv14FhFsn+LMjriZowW
4qZXqqDZJG6wdYG0krf/DMeIHXgobkYJHkc2HoDWrTWI9a0FZ77JWN2POJp1Y1HlQNJkrLSOZBfT
+NEFDmzFUQX7a/zMMHUICYjhRYYq18gQkqtg7lfTXK3U20i79YqUdh9J75mVPJtkDkKoQx2ZxcTZ
XtK12h26NR7t3HdY0fpfUnWqeIOzfmj0Ff4WMIhozJmZEie2oVp86b5I9u/DmmjYlz2/IgrYh62G
XyD90IJQf/IPnYFvFkM7f239jiGhG8lJt0glFbNSneOUfyNvZdOjWgI2WY8nqYVw64FuVpQBRF9C
W/bffkNqkYia6E6xWA89XhwhCjB+iro4OQwrb9P/hi59Cey4RKKZ3V9CKrIOSKeF3Cfn1mNUvvI/
1fca4vjJkw13O4bsCTS9BYZDC5tRAzksWyXTmyeLzrlQPT6IO4ok+cNwzLRHVuyr4SzVPTNk2j2e
BVUle0rPgv86Dv2/2VAhXLQUgaRvZ1B25cyLZ2mfoYqkz07S40YiR2aq1TJjGQ2yGMViTrEzLWWX
cF2uFXDXCfOVZ/bBpOUZfft7Zzm58rotXj0M+A9r2wSFurZrXy/0vt6CUXYDP5GBXUIIEaT0VRhS
FdnrovOx0KC4L3XaxyqRVnVAvgwt8SrBR+ZvYIXKG8fNax2sL5T05Dc3+lHP4h3mVulo6/XP40Jf
fjQoRGZRrudGfpS5/z2XSTNJhy2YsrgtfgTvoVfmwLfUkE1/awCIpkHgeGMOsNpYa8j6X3npDNjN
o6fiDCzjvd5R/z7s76PWTBLsEMq5RJZvz+zKRPzMTVw5jwspJJS9bO2Kd4c82B97ZTNuq6LpCKIB
cKG2rngfB5OP2s35N/0oeTyZT6URn/I4WEpDRQjNxr2fm5F0EXdh+oAMJUTQNVoFM0xzYoMvO993
Rr8GqRTR7jf5f+JoUWk2Pdbt1/1RAJlvYb+Qs/ArqwU/1YELhXWmw4LqZjEoV8dVMvnH+4vaImCN
Z89UgIWp37VhOQPRAJC5tV4HTNCo4sFxwCFIYUu2lWxbVxgQavMbLNSKfTw7njogxRTtuUIUMlmw
C29+IBRYKSknQOzC5YBaZVB2zykisnKvUCrlTxy/vYI4vl9mums59DWNvmrCiT3S6WZRsaszl+6f
V5PdOeAytV6FTMaJFSFpryQDUhNFbiP6rpD3mXmd+7F+uMPLcohMS18hufxuVsyji+DxxHBzTBaT
Ws6v11nG9VxEULKM77laOaTQm8frAiVqIwyVDbzfCnkma+Z5vgKidPLvJAhgF8nQoypml2uQuKAi
Q0JuoNISuKCAlVa5A60iD4jv4L1dOYxLy1SpVBxAzd7/uio3ZJF/pqueTXsvEKXJtDi/I6ha0LIU
+fn7ARrmlWRjisxT0iEgdHmTYMCnxfviVyySPA80UHaV+ZhbJDHUS5HURolF3bp8oN4/DYkfuq+z
0nTnzxPBGRUTeJsO3I2EmBWj1FEW4bT8qQb0635cC5W1+yUoYh3kzO3kaB/oD5NaBNXUfBzCV4R1
JoDgSqaipNvkd4gi/aankIwTG+v5DX35kxUaQtg57XtWfYM5mzcljCWVPARAyAWfrkCf9ARmUEdO
Yn7AGjrs8jkhpAc9Xf0srtZ+xap4/LnaeSLVYwWMJDdPdupTq80Hy0eWhllD6lZgdawZjimF0MYc
3LTOxsJjsTYXcZ+zx4UW7AfcA3fZ14TOrtov2/isJ1vdq0PE84mgebCOmnux2h+whcMgpFMWk5Vw
9/Fh163IBKWiQdFa7B/Vl98VUnEOCBlRpGmTIVZsFKvi7u/Kl2qS8mxifqSTL4SBaT34IWPRUAaK
7Mklt3V0LYj0lmVHKiJ6pyCQhtmxUZr+s9m8j0nAAFr+0n2E/jBD0014xCdXqIJ5fQ4BTQQpH6XD
vD8XWDPcFONMEBOaaRTVqZ0WyT2MzYPnKiuTOOmADI8jmK0WjpI3YT3BpUN1k+hzLrs4ywjZJHW/
xzGLifXN+Nb46FyYpz/MOFM0GoaOKGLARnD9oofX/ng885jcRZAZAExHsbbjX6Aj65aoJFgX/Qzr
+3bTuFZ8fmpTjLAYXpnV200rbw2xOPQ+qq8UgvtwBVo9xyFxSbdLJRgTPqC9JY0RPga/o1lVtOYe
+xcYGGKzp5DJNlsYmp+Wj2vNXn2XgAA8J3xd2VaIHCNOe2uqF+EitWHkpzU8HPJAaitSwJNNuHnY
1ty6E2TAcFKNtx5ohjQufVO6dU1IiP7tgIqp/kgCQbvOy/OE8BKkN8POXQcTx3PGQ4gixD8/G5nl
iL6kIc33fSKWz5d04ul48/u582N90cBfY8AoYu9DfTbzwYwBNN/91ZALOTbVdzSR0cWfY3ygu9cj
xSmI9lLuLsrWmcWF11ftodqvN5cXDZG8vOoI6617TXAkCIOzNn6WbQtSLcqDBr3iM1EESGCiXm13
FHp/JesrMFi7maaJI2U3efh7/Qwuf/eM4bsbf+jaLJLWCOI9hJSL8OSw92aGUR/R5VGwwPfibjpz
RR3KM9RzPvVIZ5xZAB9bIiqZaoqbsIdnodDQHXnGFaSgalejr57bQqTKQFL/5SDqgzSxaQpEAc1G
o2LrJpzg41HQaahDpyPpB70zl2yRf0KsHVQCcigPG8bHxvq61oLwkX4FzfbrQexSVSfXgWmDhN2X
DHHMn2Tpof/YJ5fvGjRYFQH20x6CJTJslRDpQnM6P5TNvPqooqqk0XVcLZKd42yXDwTQFbClDZ5I
y7fovN1lBC2jCadF8huIs8q3IbXQr4iXmS8EG8ffp0E/HpfIv+Edsq/JNN3PinkGokOFQ2jtuQFP
eM98Q75S7jo9HSmirJ6lTCNdv80Q+EgLbCyaM3H7XbzsFd+ug3yVNFVh3RndwwFmAF+qUQkQKZte
xKTDeA3HyG8E1hyMfXD7PCRW8LjbjZFPL4b4fQtrJZR3yewCGjjTU6HTizmlkyFWxj1dyyDER6as
6aWEj6EEOASWtk+eeJk7jc20F8tQg0f+svGl27JwFX5iGi/ocXz5eFvIlNNEMZNzJjnM/y1CbF3f
LXSZDiMKH1eWitmYmEAU0ZkQYi1If+WWHYGLeLSeLW8UMlIpfrKIunl8SKCn4neSbJH9JQx0KMrh
LnlrNP2AsQWlY+YKj/LNNx9JMNMw1Re722ltA/4tOTS2E52uJ4tICaM2TVdEqwcA8WZU+sgGHgAB
f8DZOyGSEBJzt0+Ji19EkQtQQC2DBPiqQLynKmm967ENSsZ8dyCx+LhaHRo49Jc1N2eK0/t+BLHY
iy25IhiRFAiQPDZP8ZoCd4Eto4x7Udjv2yrCbXnGJgc4SzZ5dYo6LImxFGnqZJAgVCQEsUbcaV/m
Z5hzLMZ4IohbBTuBUbPyl+fHzFXcU3cvpdpyRrW+tTetUzCOBKE4Jj4sVg5K/wQ8e/LPqM98fbQt
RFtbPOjJA6Yli00BKE5+LAguCm6l31oc8rSCAo+4kq+XNpHJhfrLHzUUp8i+RGJw98+EkeBd10Yt
2TdhSlGs8QEJifmaJ41gGNZeNf71s+xOdft19MNB7HwhB+RxaeELRElXwmL72ByMRPwKzu0PpdtL
Ahd1j9WaBNS2KTHR7bZymUazVYdPkX/H3nOO9aBdJfkO5p7KEEvtwXRCYixxV0/dslBaC63X1lMo
7iXth+08FlusZQD3NnsgI+pezksweQ9Yl5QFP6hy/28qsihraZRtl1SsCEPMKveLvx4C++uLiaQp
x67aSGvLarrmyB3O+MQ4AjqzycqK9zq4PoPvnr9De0rRI+NL4h8Hy0ls7IqpeJaCY9bWiTUY6UNg
ypTDJtDddEL0Xs4Lx/h3IOgm6+Rm/5bS0pHdVya1Qd4rio7uXOjo8L0l6BPc8w5e7lfkFfhtdOAW
M+wUkeYqBOWtqvxSQPeeUPgyYfsknwDdbi4w8MhGXybnP5//s+hFZfbH1g/jEer2yxKnogyXdNbw
ZdKk4F1hgpgbnNJCxpWPARpDs9eSDlhmgbD+qne+sgqANg/f/V3lVj3GA+sfeYQdxggyZHgHVnXT
x56dWtjaDUvYJVL+r2RPisCi/9JdC1X9KXOnu4n+waeoWZjt8CB3mqQaXOU0o3gsTtU/sKi2fmLE
mTzTVmGehFGwNYNhRAOEqkEj4cjxkKbXPXa3Ymk3nsMPCIyVQ2GbUYQb3BhLr3XaLSOZ9rDoSRFo
oYb7RAGMyLuAycxdbpw7P4mINvwPZRnMKMAbfaliy1WtTtK0VfvGjL3c/+kJWD2IdYtHL2erUGXw
wfdAIcnm8o4LV9fQbdYVf2ORPo6cfqUqlAf5/hfTeoc/clx0gLksPXxysoGLK+Usoh6xCK1axs0D
CTMFl0NUJtvuY/uU8CfmnjuxV1mKlAZlG1rOgKydIVsoHusHpdTsDaaiBW2qlOk0sxEzuuRR4MBw
rJ0PxCLrxP3DpyRz02I6GJqySL5UWh4La4FjxfBJNXs3ErqZ7fMTguRGRepRBzuWW8+1K395E3gd
pHncusa6cnGurw+GIWK4ViDmPjT8ez4z2DvI/GPtZh8Y/AyqHmM/tGCVeSiWBVsXftrkA6khEqlp
BETMHDF5dpv5PivNdu0/FpsbYnqnajJLnGQOnb0OCJeGuMj+FZBLN1cx9HSGPFmO1Jyn9kujAa3O
JTXDKDq8LMsokkEf4tAEwQsqQVhn/jDty/Q4Bhtu9oQCitZnWDjDMZK4kayZqe0cht/Bj3eqyt/A
CANAmMRURK0uvzNt0JIjKQ1491/ekNNUI899/84xuxvHaS2nI9db8RO/+KmiaEyZj0Cztzm9SDJL
zR4jsS4ZbcAkzK1JYST2PgTyYLWim7JFMD8Gw7tLVQ+MA/spg2mrzYVtH2qxELjrZr/+lKpazOMc
HofmuYPXSkeT3XKvRnYmq/ExCTXgHJWMtINbk41QPRsrfb8+9ZGcUxOsjyMkj3R/rATM2yr24e2R
LIgMYVyT4DWhxhGzECA/16QvYH8XhBvWLe/qyyx6rVDZgVlByJcDwxf8CwfFGpWuTjrjljsX4b5q
+wA6x/ZeoR3cvOT5GlLYdQOASE2dWrwPh4UoFzMi3WeZqJfGaRn1UpbhsEDFe1m7XidwHkSQHRYq
IRgTakKBqhnCfjGXasuwP/Jqu8qifyLc1stQxjBuVFrfxLLy4FsSF5zg28k76rZzlgixClvnkX8f
MVj5Ycfl9EOVnJhCy7eq1SxRSKGCK1sWVQQCIMAqItQl+SwQyhIsaDNC7t5Ta7iqjd07BNgRVkPT
ds7+lJ5I9tHbf7DgivNyLmjdBaYeJPOsDd2JYSToSefKwvaYW/q3ua0IhLy3mSovo5g/Ni4nQnE2
DlKoL3/ypwilQIOhKao7/On93WdhJyzzb6DcYCjgGexeMurqEub1LmEzGQn933YHA2vfJeehkC+D
TLjSHuXSaB0U41syqXerMUVRZD7QPYoZF9JX0PPP4ZcpzRqx7HMNX1zRV4Th4h6w4s8/F+qGIrq2
hHiw5S3/bY5wB9o6TfgvRIlyqs5H9nQPLmKkXOKaMJUFhahPsWzOL+FcwSmUpz3evrls2hA7PqYp
7w6G0hcpV5YbhH6J5B+ti+oXogy6UZ9HuGTJ1PTDv962UO5HBdzxKOvRBHqhtxCc0ydWyza5B5E/
pesm0osVtGWB5e8VAvIoIgAe8mOlY6dy3iriFHn93Dzu5XwqbG03SLiZhL/M+lIUQ7MGjgAIvpES
5F0MuOO/oqxe/dewa9dJGgTzvNs3NR0FiP4hMOJpBYd/eGEvUuUDWq7lQyDiF7wM+9bsE+vHicH2
JHaJsyJXsImMt3gsYaBNMwV5twz96AECTUuzI4l/wddgni6EovcvI4wHGwEqtX0eVJjkzpxg+jN7
49HATv5poADNP97SG1oXeh9Fap/uT3/VWNEtV+RAmDF37wpoT4gzpe+f/Awiz+qvLv/fuhJtV27k
sRVe/PihvTaar2fIOdJCJNsTgwynTecdC284waSI1r/AbSJ7uKwnXtfeivcqRvfgVZRb5japC3Hs
SEr6Yt71TVDM6LYCWxDCnNOO+rNJ8TXVFNnfGYqwafUaw5IlLXJwFG0LtWNCN9qDD/G7k+ybpPb4
xUZhN/9XxC/JKNCypPudittq1WNPYFwMlzRP1xzsNr+Wu4DtBmQoc00zuA4fxnXAeuRa0a5HqnoB
2Sc4FEswYRuG3/WfhrhGPy7kGPORDUyLwf6p+jcvNTSdgNgqf46tfWr09IDsJcq/XCx7EtchUQzg
2HO/mXtOO+VTtDWHDz97mdgo2/+IvyVtmR4Q5NC1M1bz3I+s0y+V+Spq7v2Qnktg7sZrLQrovy2i
0H78hI/j/hk2wFcDGk7ex/I/SIt0K8QVplr5Ht4+/CYZWcPNmiYIItWfKVH3WGPUslm9eHt7pwzz
rmBS2hlsY7Y+w4exYtd+pBwSswD8DY+jW28n4ZBxXIMYzx8msJ9PmJRa0zrs8cvCfOqW8xGGpeep
O9QkIfPYl2EQp4x0RfXSAbOpuJzVF/VytYR5CmAk8cIvS2M8cGf85f6FyjKHRceN7pNxh+JsjjoB
fjxk1LCzRH6cAVyfEsYQgqu4wLtN5MBf/lVUKjdJF1VDT2QmiIKtPUAlvQt/Gax/fqQKcZsqA7DJ
awQK0Rgr2yZMvya2R5SiEtupBoxUHWiJ2tQm8ehM+Iov9gbAdTUrOtX6eadhbxoOhejCEOtlvXaH
zcPQUn4BTIZJvrBSt0xYyK1M+BX0IIWZrrRW2+pu8Nilcyw3IDTJhSWb5G/9xrpBnyH1bHYiMgpI
Q/TBID0rNPzF/SqfeckQHZTu7ftWdGycYIsI7XZ78ffn2/Zdc44PhRZf8DFK4ft4yKohq6IliKGZ
7ElaMAI3ksXuu8SPpxxiSn+BM94I93rDWzEDCgoKgJi63XD1seWtohRIGDoFvjBFTh/L0t9fTE/R
E5QD3DhVdeenpAmwaEhgiHW2hjf81rDsY6NE7ZNNm4+IEw8G469iboIz1LOHlH3zEB7ENvTFvzSH
+0fVTlcM4rBfeUg16H8y1eTOAdbT+06VxUxVtqPAHUYrO+Ptwja0vJpPTCDtRsAvTvHbzs9ZRtd1
eYOukNnJtO+it9PEuNlgnm8V0Tv8lIcDLl3jKGJWuFBfC8RWnDZJFlWzmwCn8dz6bdK/BtwGwOv5
cthQA0KX2FAhOWTACNwLos0WgS4zY9d1EZO+4hwTvRHun9yM1YpAiucd0avniXPzh/irh2bu7Hbf
0qdUsUXlxsOTNKFBKfP/7w8akzX4ucCK0jyqc1xd6HAUfFq0CyT38Oy+StyTshiEM1CaFStZWz7W
8mmOZGPUuuW1OLE75Lx7vR3fjwgOnwgc1Rnf65hnPLheNc5rZCLuu2OH4/2mxLRLPoCcP4OlDoON
MHkBWW9BErqr/JC1zC2ov4Up5KJKw5BJbovQ2W+vBASbArD//ynq+TxGRmG6AvFkMJ9Z3e+dI+J4
6V8Nk6nTLPhSrnc2Z5Wj5NnVtzlT+r4hKdS3P5b6nBL6+EqlsU+4b7+aL/JtL4MJunKlq9oxCx/S
+WORupER9/PGxKdAsu5K0J/6MlgV7oOJx9Dfnruv9asmqJswmz+in3jpHYipEooTsNlIIvE7jKtA
ZX5L0VGi8Ul+S6AuSGwFy6UV4bMe18U+a0tmWh+FTzuf/dyRTkym4Elz6Tea7jvyiAFQAHoKNCu+
jwV/p/2pea5Ze7ZL0SfsoQdZVLybMYEiccVY7Io5dfAFDhMez/R+oL7kPdSS2xThIC/c42WvCYjg
SYZRnHyQ5m9gofd594neXc/yO9Jo4/hx580+cfywg1OMX+sajp9Xxm0aNt+xANqURxsZ+B7X6ram
OTphNtwvgsQYBffiqQcNIl53iEI21eswuZKxSnlQXS258GIc5My1Wog7rv8R/68/QCwhFsQFAqLY
iqcz+F/Qe+u/bXQt+zSNAePjfJOWCeSqhjVrPYW1Ykcy7vjiA1654eB+5xQNZc3p9KVZF7fx0ggF
ShgR9BMzAPdpxSOHmupJJRy1+rKaP7rPX/WoH85EVMJUJABoId1CIXjGFnAdis9zZhdKbLXzrOv8
Urpo0yRySqHzSenZRTGV2UlpPAUro+5NAmmfoF3BoWMf3Cu/rZoyBPRIij0U6QOE2TNbkIJ0Nucw
eLtg9kfogcV+5o5m0vMT/Bkj2Gmjn95bltHoy1gUsJ5qdNlwxzmJq6IUC4yoD1CNlgnXJO0mK79Q
6qsIx7n4VOFIzMn59a/EE+eRWXa3aaOveSf/2bCZRkvhJJobCnKZNkGlYFDat9BQzvDOoWx8DIqk
CzmGPnbPPERQENKbEDnkurgnP/Xe2fjCq7hhon2nGwUzV8s4p27p2Un3Gldidm/2KuMZ1b43fwka
zeK15liq936Fgd60by6DUKWfbr9cA5bJ96K0nfCdMrEGc47bdNY+7Zi77twu02Z8i82HdHIK5266
PqVqt6cOdSm1jfKEpuBJNTESl0fULR/0xLrGl0La/W5Wnfe7CpcRj472/FRA0wEIkhFlFrV7cEXJ
Wt4PZPXvK+hnTgzGGB0/iLtPjqdqnwxGdXRISM6y5GZMzFkiGJa8dUMMGN7Ah3qnUPr7CIP1QVL3
BBKaNroK7sjKzJRwIAWpZWKWU6w7sdsdhYFiuSEE8yFn6AFhhPPjkW6lRXWCo8Z3U8FsR9XAJb5z
6VAF/C6nrisG5VIaMYVSK3NNFbKWNCN6S/6+rnC7iGiIvzDsgHLaz6Otngx3/72v41aGzPXXIJDi
xq8VNcTXFJXAommFy9l4Ae5dhlG1OGfY4+OWZjF1Z3nN/XFy87AW1M8I/NtQ53X1sm/QATXRj9jO
vDjxDHfBpfMJ6YbLGQr2xH3BEcczXfyLnauBsXawPkRYOmhifI5jgMQQDRvcIzCTBrj4ABIVsE/j
gzJ/OI0SdboqdYGMUybX/Q+eSwfQ4OsAPImZHMVnOUTGOCU020qx4CGkWtP+0fnBhKMOIjW8L7Qt
souq8Vx6Dgm+qM36eiEe0ulv6GORlSr9XBSGzvOoQ3aLZpFeb4QspOex6vmBhpmHsk5q7N+Tq0BK
kg3O1pE2NuI1lBuPvKOZg0TRxYex31iE0ROkhmdygF/+jL2Ridqq6ZSD4H6i58HcgpMIqGaV82AH
Xdqc38JfcXf5K/w8V+Ne+kXtNoBcOTFD+11DA3HrORhRluGLTYNKBqE5jagyu2uHIFWBhNEHk/KC
73D1cRsJ7vz0BWFMRh4IBfnQ0IZtpY7F+8NhaSg+fE/87EyDdgZk3QiJUGIDAV7Jk+lXxTVFX/gE
SyIj+LeBdAvk0/CRpdlmdg+MXQDeCsUoe5Ui98TVms3s4Osot0vVPGLpbU1+kafww+4LaI+bHk9Q
r8ZRbQbuOYCDias+pFjxCllVFCD/XDlpL0hp0CUwn6wyOWjVf7jwYiSgbylkqd6JTkA1U0VMIV8y
PL5zltO0AX5CrmLxCbsXKIPPLjZ5vkA9OqK7Oz5ydwWqqMNaEAjQl4m0RIOQahVSlkjI76tzQQEY
3LWtM+UqOtctBCYgPcpQNEaVFj7rWBuABZY3lJ0iWiC33LFv/i1pF0lI8DhBcuZ7H1bvDmrNRC9w
0m+lFHPUqB8wOX/oGsnMnvVK0RPuebMxjGqJr7qjjiKWkIRIvIzQL/V/Esqbi2i1uTLvkIZD8WeJ
t5P5PJlFeGh36YZQekD1R3DkUjyvgZdYKSBONEiIpiDjq0HUGl9ovt6T9ApyXOp0h8yLgBU9RK3B
JWmHti0VyKUl/fQeZuW1XqRl0xUP6BLCztnf1aLZXZZcnGEveXEhSKeL0Bgdb8fH+BmDA63B56Qe
Ja4QDydJ4ykZiY8y0dwGMRkTIVYx3TO2O6Z3ZVBEA05VgD5RpyTWM0uw5MSEVn0dHupzsEghT8W1
K9SeGT8JpDUaswtMSHx4M60YFXl44IBGELDQ0yycC2uqqnG+Xt0NYfXplcoT40S+bBUjArzzf9AV
ln8ZOIgJwNTXfMZstb8rziPDcUh9pF2VcFFwQWaI1FvZ6XNRKYIQzEw6qSN98nWG7KcCYWx0rwkb
NhdmdDTOFr3jFugEqKzZs7yqActV3/nSMG0g2MVvFUZrEirrmrmpOBWH8eNSPTt7NKHAKrUDVHqL
7OhZVroPRGYAN7Y/KOUVtEiPjyYU+GXeZnN9kCF/Bgm+n+LkOaNywaBIocWpsoxj4LN22t9ETPPt
mZ6XNXRUim62WFqa6Xe7jZgygs/RBbV6mTQEFlXx3mOiXpsMbBxziLiPj9TcJPywupaicynhxaFU
yZRyyciVa/dgiff0WroSagJIUqlDe04/8rs9VQhypeSNe9fOSxRCvppzz7jXNr5dwx6oKqGaKz/P
4M1VsOORmJK0wXwaG6VzCqlIdwojgCcdSsin8OF9irAR9RKsnFtB8za/wLmyg8bnNeTKvJNJ2HXR
hr6aqbSfWa77gLmdYT+/Owo5u+sGgSnl7J/JxkUV4kFFnQZyjH3OhKz6o+LCE/Lj6oemOrQfHPcp
OeZ/+S0mzGxpoUX4pHy3DiCHtj6JB93SMVNz/ge7jTQdIFhqiJxLJTYVQTuiLZFeMT9IzV9gWhrV
IVa7D7nPh/ZJ9ORa5E83irFzZFg/IkuThO7HE+iFpbnlfLLDbnRWqccF/tE+F0Dv6wkVUVI1Ie7r
FujHbY4ZAaVAJ6DrgL+2bl4qzP0drSZHhc2zukppqBwIH1KnueejF7vEyoBC0t9IlqZlGuwHyF9Q
Npa4dnGx/qgfbIArwkoThEuqqgxqyGOt0KPpisZfjHS8zR4lQPKDLZZY7jWXf8zkogW2LdSGqSBT
vjJoeUvMeyAPR4/atjrjeVUSJayMYgtSVZRif3tVNZVh2j3wLoz5IEf5s3moBjd2XLpRQ5zt8oh7
6JhQk3Rk19sedo4rk8WmQCA1zii1NG9QsPyJkyCiKgEwYmYV8hbyye4sYynqBmPRHr2WG7Vic46Y
pJ9lvpAG5FHFtH3cDqnl2ppHwb5WkpQK/iJ2opbOFvXqG/72SU7Xytu0SHTmgYAs10Y6Bzkw3TIw
2zkGDDXi3XoQAmKXy5yVPKDn4AtOM75HbMxpDBepy7eWBTd/zGZBIpJJH+KhS7sglvTSZKIssieN
CZfmd874FcOJzX+f02TB1DrkTH0u8QXdC+JE0Zjlg9RlcLACB1n+wFfQTHhwKt3St1DKIltwxmN3
/SbF8hh38i6kIHF/cgVl9ei9kSv8IkU6tEBrarROwxZJcXe6pbdn0rSjK+504MPmz2Z3MeJGwu/H
5yMCn1xDlpLUWTcIrkzm46C1culL7cUuxnMtErT8PHWtcFDSPiIevYaTqbMXr3GKTViIiROomjHj
+GP0l2x9FRTbolHxR2TBDdTKq26M5xD7PZe+HjihVyGx3eRa00V8GlAY6dCg+PzQLpTPMw7XAR54
7vfYFrtDT+DoELk0250WocCRrGcu6psn5Mwn3ZB6hRXReXpsAifUvW9PzkVPPUYRh3dQSpOvrknW
9zFr9Ryu4hM2TngF0HATOPb9J0hBJoKk4J9O7tCZD8Zf3nYlwzHC7AAWhR1u3Q5bKo3+kHIq2QN+
Q+nYdLq11FuPn6NwIFGkTQjbWsR7TlLipiPQp1C1bniT7cFglG0fMQpkxqwz9SuvHoJ2giXZ9Prs
B+oLI+2ivaHcgJ6x4hvjgnKbU8j8LQUqA84NBsN+WCGaPj6GlKiMbMdyvJjcJKReFvxF99ni6oQb
yCYIhzMbfPnGKissxsrTTbqQxT4zbMVX+bQNCW0SGNz0xrNxsryo55jpwkJsCtadQRW1D2LRtc2k
nS7XuEq4ZwVpUfAX+AYHnZAnNhxZoaQsa7Zc6nkD5y4O
`protect end_protected
