`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FEFZZu1l9hQJOxxhbXmhK7veuQ71uiR7AxCVsUcjBubc65cAgGNIST9Pc02kjcd6JCXO/hjV/bvq
2Qzv5hQYhw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QgkOLsTRByjOZLS5U/dfI4ro8ogV3dovLulFZWO7MI/krEKJykjyv6LgN2BTssbryEGwy88HHqTH
lJ1vEPNUCP5sOgIdzdMiWvX5HQtPicwOARpoqhpD1ve5zikITYsz4jkiRpNV7u/YcbkvWGgjs6sj
lXTHJiCNkuXAeVNDu6E=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zf9OIqlUlPTypL99ArButPLHVDmKWmnOaCmh5SibIqvbBZA9hlwB5rEFaJ/WM368kbSJqTKuum4O
rbZlAMmkHcecTDCIxqsXs+S6wFjDkC6df67kwQfrlfQ7wvuDPFZDLrPSFwrc8Zi/6wwDPYkZ2gZ4
fiZ0t5oEGChlN6BK7G+Vid3UiKdcyqYp19K5UU7mjHmmE6kvXEbh7KPKO4vlZjoF2j6l/kCFfvRn
hApIEG5GbOCWMra+7en2rQyJP9OdyS9U3RAhkAJTUgHPg5M55r9saO5HkScEFNnf9mfKnDXXaJul
9i8+Wi5S8mvdHwXM/OPjM0Cg/+M5FVT2ZdTNEQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m1oy5VJY/mNNfhbXF/nUfZAJcWZD/dn93lPunAzF0yvFzCd3FFAQdsLaWO+BM3PbxzzeWZYYJWZS
vn0Il58zUmzKXklOt8sOLZw6NDn/+WPAqOKHoAymSFvh+nRXiG/5zt5iCylPmNBqWfRhMOmwa+pL
c2Y6/3yYNOx4gYMBcHn9c03ioT65UnL5Oa66rp9VDFrCZiac7e9+CeRvAJSj3yWhhVrrR3w7d05I
CN5UK+CIaJBxeW+754v+vnAlU8VitN2knGXRstNKB4vWD3hRM9WdcRWZMmztKybCsP0LCOrp80io
NiagQwKPpWOHuudoL+3vDk/FJE7iCtrpjFVXuA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o2KxWpeWWGlUSYSzbhVpCcP7bH9I3jMMPxq6/eHo/pjmBsyawQ+0PoKRKvCty6l09dl3WM+gGNqv
BtUz/Jl/pdqFJs0w/J6izzNsvcdH2jP55IvGDTfZhITATTIU7JvKn7hiOLEH9TzxT1+g1uKFfx5c
He0MzZ9ND9InmGr04JLOFY6KyzGDjEqWhbLxHFB5utTtVkpKosViwHqUMwY+xPA5ntMWJ7GPHDww
IBFV4Huy3Pe1KyU4XGt1+DzQhnIUhcMwtxGjg9qXL/MVVGQLioDcIBJGbE1qYaNgSkZEUtrTWceu
FwmnZS27XaLAkOBolIqNj09TLXvnL/p6ijAnCA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dljmA7zCJEWM+olxJ8hx0uuuQBQD50jBXNUibL6K3+/DLpvZSGgohDoQiq/FSyH0pPf5t817jzOS
RYKQthofgANW9nenpuoag9MwBqX7xUGra2O1Od+UchZ7GZYNS0CumESrD8yXs98Oi9I7lkU8HRFa
FlI3VSOHyJJUmCU+r24=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AozEnr0AoDCXiAMaxz/34GbUb1U3G5cQ80ozTxzPgU7/tqGWYwonNM8ad5vxmIURSHe2SLcW/XIL
8mAPg9jQk121PnCZoz6atktuuzqDAeuQRfBB5hgzh+u7sFP7030nUTi1CKfAKsnxNE/Yeh8jYQwt
pWDToCdq0Ma4nNzUAotPYcXuU1vAoCB0sqHhmPsVCe7/m4MUUA+Auzl7eSJcK+pxRYjXSPoFYeL0
PXkiCNc8vjvSnXuHLCFYjTZiY9s5YpfoFP6OqH3iS3nG6K4+XEonpKMJwjmJBp5H+vxuMxlblM+G
7Ac4wjB2kNtA/hGcZT5hNsMZwcGQLHOGEcKmCA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432720)
`protect data_block
V+LNoOY5GRzYBUrgkqj5af0FtYcbGfRk282USXcD+sjuoQWtuMYWU88Jk71RhNJamFZ57eAbmgfY
wJIKTdmnVeNuBKIyWNi2QyOHfpRs6BAHT5VYsAvQcCL1TA+X+AP1nZ3tKoMtOT9aZV0rXlm61BCt
9czyqQx79W/7Nc+HY7eES7W7Dp3OD4dEWKpc9Dbd4gzSR95FOBY6T8qK74efu9y78i4scNJMgcer
81ib0y1KTrtScIX37w6D0kcqhlmlPUQXyVXeJfYOxrQeXt7pkDzs/zAN2cXw3IW4qd1VKc/G+bEI
KSvy2mPbWiytNzFErtKPEDLJZlzsrp8Q/hNjLMPaSs3G91Lxp56acyyUBVpUZSL/kQ8D6qApPHf6
0SKDRuQT573fga293uQl7hFS93B0oPuK9yPoivEwX9o4uw5H6KxypUcsbiwEyfBB+cTUwuXAiENL
YP/Eim94inTolEuUaH4YkgHkl7TeAt1dHY5TFln4fC6Rp89cXBQAxANXvP1IT0cqvKbOm4xyONlV
1foeR5rzYH2GDf4oopd8iW2DWmbPV2kBS0uCpg1tryimAZrcpZVPuzK11B8isE9WrGvHd/97pcJk
UtfewQHVXbl6z6pfPcfTv1qidDINkclUyToiYP/nCnlGlZp6mpXamF5bx2mxJ2mgz6CE9ID1RiG8
bW/5ItJSRQ8Y8sJXWg0rZXNey/c47ZB0/hkr4vzGxGI8MH9y1I5nwbK5w/3xYBtbG+88WEBKINR5
CIsbSYK1KuRd6iGWrpphQ2wsYUk5iDTRJ27f6z/hlOccTEsplHrswO1NYYqr0W9YmhKXuOQTg8mO
ruoY4HD5PE4J6BiF6U6UBppXYqXm3NxNVhaMto8hla9RKDO/25cMDtYWqIeGesJeliAL8bEIZmJO
RAthXfS+1ID4WI8/ZTrsDXXfGp8cbt4ny3sefIvrZaEIz0GdEPKEwP1yTM3p3jhiZbOZKroakewT
/9hyIFhP10Bpb4pNLvupu1CO54Awpst/OgLvq/D+EOqOEdGlsHcgiy9FQWFeFW5/6dgjkFSLuQw0
aumpUpIbOE39N+9fG6qWDroqcUY6buiGkENeuC16KDFegs0xyP2QsXxbSXhFLbBiHuXlXF6rQqsq
2kgVzHcsj+EhoC4CZDvLTYsE9tlHTmplJ+F6KT8wKZ6CapJfQH+Ys0DGw4Q3YkDN9KAzpg0W+3HZ
NT1QebhhVY76AF4aHFPhiTNlffnIbnfPwZz/gPaUQLX5+TyHt9eSWGgqINoNPLOZc3y/xa/hq6A+
RG5NNMFtvQKM4+WYxy86PsE92Q2Bkn9vFtgKtAl1qoUVaZh5lHKVrrS35LuVBYzipeEaox+QBLqq
5v3xOXZkeckfWu/s8wTbNzhI1QSrZW1ZFH7XveX5xPY+Ymrqdcvs8BFdWvmR7d6jyJ0IEVe7jniB
DBgQNhfm1ghhSWpB9rX+coWLNRiIr0IW7f1x+wYEG/Ac2uueyjVccZZgUsjQpicLb/wp8UvhPreE
ddyCsYYSg+XU5b6pTE98aReLtxcSwMex6VbcqroOCfWce6mnkyIxitFIgV1QyUxI96fH4lD+M/Kt
ddnkPoWVx9vvQ8HwQoQL7glGKiKr5oMvb2D9P9F1k6adI5Dz4dJ6FIqL4I57NE5Yg/+Du5eP6e//
twgGM/gyiWnXqcO56GgGGNedTwcLpv/TfA43RoAyuOnMYGdjXx53K/ecfTgWEMl3b1u5k7JL30Ic
lb59guiIscGw0GIem0hVo6M3dCNChVJmq0/+aasZFNK7Zf1CRA8j5Ji7mBRI7ohhIaE+oKwYp6hG
KvTkXg/414VJciB0ANjfF6wMInomt5pW9i/AsIX6UUexwvxZymEYz3iu4OBnEyK3WkUCY1oOG/KC
XD524MQeIC7sDjT7zENq/MrzQHL1e5Md7w7TuZWYdrKvj56CU0IxyGyZISKUVg2E+HwT7o9EJhPe
o4U0QYRsznDeBbtMDViYZQuYagNZF5V/XirbS7PANpnVWgQHXb8Ukwlaq8M94T/8HOmE9j3uVr2x
rjmuJyH6sNVrNoBwZhZcV/I+dDZpg/taib/huqB4X2PSK0MUX626hyHrl0vBXE98Q8zx15X5VQIA
W3vBZwbzq+k6CzVkmz2qLoL0lTsRdXFNjiZPMFl0lX7RJ+gjomJd+3/HzQs56W+Y80N44yls0kM5
It1g+lNQJ8NwFhyTNKTaQUctDcswGu8/HuWKWzU8uKtTy7k7dsxWl35V/m/meCUNB0D8yOv2h+Nz
GYs42+mEiPvMeaTQVGyMrpToDUmWbfxU1p47mF8Sg2wsrVJGrxJXEFbW/9MQcvXeXr7zbUZItuv0
MDoVLPd/+LDMHE1y8FkYb7lodWld9Cx02aKSCfnnh+7HFkdAZKnjvRHzlUkAWaTCNuzK4tFX19mh
+uo5oea/YoxaGPAxoCap4eWqqsTiFzb+NiwVFT+wWFnm/h3+ia4fFmoRy9d6YGrCgj2S+qvo2Htl
kiWTQJki6fenTunigE1Llj4Z+vkLITmzW18OGI+iPMot3Pm5cVtYutXl/V3tAXhDsi3T1wBk2jZF
a+FFfcP8P26P//BaXzQ2d9Nr7CcYTB6jd8IBD4m7DyWSyrDvDnBkdZMLrarUfnZJdcLXNllWoK1Z
aT9oicZodEt9WmbffmnM169uScmhs2Bb3xvW/E8v3giZjvflFkqWWs5GEzT/29tJ1HPyaL+pcCLc
0k8euvaVpIGTZeXoBn/59jgNJrxlN05QyZH66/Ja+O4UodxOSByaMXfCOYPvvLyIYwSCNZrPUz+Y
wkqf5nWpjCV1NUm72dWqVueQC587GWuuplZDy2HB8+Gg8QZygJZ2WiZqUZxfLViKD9wBbkJOCeKs
7itscq028baJcwLxkAMyDLPbMrAuC0FYKq5hD1StsGmdxDlucE96OG3/H3vKj2E/RDZSJ+7Zz/aR
gEGSP5592p+I6ZdViNE/CDGoDkYHGVERawF4jwPpHe5Q5NtUZyB3CTswT468LrhWKzXMHVuJTe8e
QuF4rnMia4cA/LuYpt22jSFp+dxXU7nuBhOdfFbeiIyugBxufewNv+QUGNkp73YrqWM+0hbKcg85
ZBOJYeF/fZxhUYgH4eKHlwAr96bmshqb8m6jWVH8pbLJZjBOfWXwDgGw9JUgVlgv1EyI0S8Y4tuA
5J4FkIv+NXEEH2J+s7Twme5oJZESVTZUgEe0HORXc69ERk+A1ay++6ngkuu4c+vdVUH8I0tnL5D6
riK5O6hO2AREiqj6X3SLU8585nJ+XurshMnrdqqTZr3m7a6wxLIGIJpPVZfTkKVYyaRnv2X8H2C+
Om7k64WTK/lSuOZeBNNiWp58m5krRFf7FHVkSdElAsVksNI8MMMq6MKFRZ9sJHDrg2JZWXYPtQJg
13/jiGYuvqQjq1Y2W2RdAJ4HnNA8/Gf8AMvTwySL7R8mwyd/c+gfjjsdty7KXtvI9FRIyitA+n+j
Fdo5gnAKpxeRc/mswSgln9PdlgmMtYJC/22UOm9QOIkUw8U1A2jt65FwausVgIN8Ys2IENAS6JfJ
Un9/9vyvBGjmADbdBZNgsrAWYyLaykQTSW632uE6Ray9rn4CuKGRlKcI1yAWJ6it2QCrBe8oFVcc
HceEfVUwESs0opjXgPL3kZ+373Yrta6sw3hUXEvmQ/1kJG8v8gA5vpkEo2uXyjGWIQzHD8U10YZe
Lu9Rj33fjVZ47Nc1tJxOL//lP95zBSLiDYuFpBTFSwJLgCLz6idUgINBROkKWDgpehswdY9rmE91
1GfjIFbw90pTxRUtRf9CD7zkrubz8GGMkRvgPlgnC2wD4N+h2YilCU/9zjrqJ/DEoOXuTqzq5CVM
QcycaAeDZFm9l3TSGbG6WL7mrPbfa9Ad8212BaH9OUau3Y2bnjleDq1o1q6cbFg9l9OTsm0Z4oAM
bCh6qJ/1ogVd9N9dTTskiHUzPHMEN0O7TxO8OlhByWW2RMlrrUhuSXWG/lDE64/7JFo9V26fHM0h
UpLcENwXXMwvOFR1cnsIXP+G8kji1Lu4BTrGkQRcbZchEAajzYGcJ6QXTy56RWMux17ZJcyJY9XN
X4vlpCjjs0vOQglJ/2cGlA8o8lLxTgLGl0J8zzze5F+08VgvUQVmHuLZTfXExQtVq+OzywOMZutt
E9uT05FgdiK3pMmtYQTVuG8inb8ESWQPp+CZ3IqfKMZ4FEU5LcAYJ2iyF8TnUJk0x0vJOggY0Tdn
xN8WYfP4kNlWp1PRnu6msH+FoJTleKIKNGNmBIG2mIsY9tTgljcYC7pcaNsY9k/1rLoGPdic+MKL
EOEIzGZum1WQVxw31xzZxKpKJwe4qB5HIsfx598BFdFyWHvearHFPsjL8PRk1iNCf8sLb3Y+kc3Q
2vC5T5tMSvyKPQKo/xzlibwQvPhMOkJ7bQ3x3pAoX7gSm1GNRnjNm8I2loCCbw6g8oGtYeyY05Mr
5zhB+CLVdlGfh3yGaGgv58944Fz0SCAHnZ/FriR4LxzjgsEqDUqAvo9g9LcODbw5uGPOfPygEbFQ
tv3oJWEjNz8ouUTbtmDZ1CrBENLg3qh9q4+/SOUK+fVmeO03iJda+0/ULTj1HETZGxDNFLnBFCSe
P4cjeXxEvyduceKPQBQNGBWTT4zq35TmIe3iT1ctFYcHytnuMO+9sgVLrE170tV5BS42C70cEl9v
ZPJvJRvbKFJ9VDfB3vd/VyEYQ9VSnKtrD3XUTinxPq+jsFCXzGPgqbBePk66lx2EkWjZb8+DXiAF
w9V2JZbgvjt64VgkjYJJ70/LNW5UU80eprBpP/lcATE95y/Ow4cg8o1IJgifolSYQKlh5iFsVjlt
0+QVdF83bpPItlbPcr8GEgXU06vQSc4KNhW7TxmNb5NzZ9Q3wT+KR6zqKdgz3tKxaju+zhHTzkbN
TK7qNehk2CLjxxzS/LMfF04KN9vIx0Z0ihN4bNjQJ0Gt6kOAzZHUiDkoVZf1BM6dxs+ECm/+UdBn
SxTRPT/rCHJ8fw0CRikzUS6FC9duFkOFWQJxf5NftIkxuzHdHOhIxbQLbgzS1U9jxp+YboYExyKv
t7tzB2BWxiHp/G2td5SOplcukLuRq6dDktz0FcrVAKZEY+dkSJCKbZNcmrKkigyQUzlEONe383EZ
NSNEFm0xmy3Y6MxNib+QAcsOHDPxeTdOnQPA+mCGRmJAcRAXU7vJS9Do6Wi05owyltLDJ18xUeGs
k3UZnn5aOGKDHtMGv+QRvDTY+p6wBjElEbJSWgqwuKY4qa5xt/kRy5UObBeyPz+t48KQWM6kMKsF
mLriqINcUHTJT/v2CyoEQEsM/VDvcm3IO19CVgDJTAcNGt/BQcP1lXISC2upnqiaKuU0nKwhFcg/
+F3ozo8SQyGojFdws/019vSP145IJ29OCGehVCldUvXMJbxgCrH4GQsuiSHVBlEozfr6xdg5umCH
Ym9852rrWrKllTUzw6UDewi014zJFLxciXEK/JS2ioFH1PlFRQvfdAjMUCkGIg8nsrxrGpTbrQEb
reIK4fiHm3CPnqtTftkRxFWpQuPJRVPrNfcPkrdT2Cq/+gBQ6OPlTvBp5DVMHLEPWTvdyt/YXSCV
MrZ4H+YtF4rioS+osfNPYXYlLYCkeuICgkgUwiDFj8a0uM3BWdEyjpkIwTUG/QommdRiYipCGNxk
DRo/Hl9sdEDHkypqtztBv8rUKJo0GJeFbTq5ayOAAH1BSEPiwCdow28POay6ewROQxXy1r00TnBf
Hsl5OLw3xHDwLESdmBcjNDZYrgpmcyF1g8minF0xCaYK3WTPeh4GT33XxDj2+Es9vB+Lp7N/DCYq
TTb0crVX3wEltYFzsYtliVnWcrKQmcxwTztM5NheSsi+H2uQNSFdZn/5vYAcv2z8V0h87pSXWpYU
gRRKEY+HMuslHYKnvNEBnYlCewJPSpxc+hPi+denbTG4Fbt57BZrS/OweqOSnC5NLxqgKHmo/tco
z3jEytp6DcsNsnZ4nK/e/TK+12zflWl2k04IwNXwjCXELJztNRWB4c3qvh0MqxFOD6yPw2hvFPZC
nRv/Kkx9OcGp2/+FJprJpx5fw9D2Kdx2EN3Y14eP7wL5j9f9EhIDRotnYxHobvb9Kui9oqMuYNTY
u5WbgMrvniEGEnMsT0JFn5AVuUTz94V5A3+kXzyhuntJqF1Yfy4g9yNt9AEkMdsqGTaYHsL1F/cM
NzKs5sezQkNll63k+J8CsYsWDiybBrCxo3Ibhd4C4ymmVSBIp+pxCZDnLo9VaQkAoGhb1Xzz+bNV
f2nyTOJ+1sMLqKtwqi9N04yJ/gnSnMNIrDs5dKZaEtSfnlPEdRYCJ7uNG4M0dHUIsbsQXNVPtyH+
btnaaQRIDAntipKr206qAJQSOhKpFwAxFseJ/YkJSdxQLz6Pl62zbZCucvhNx2F/ScG2Ic7WZIwC
royQwPPywc5ZFT/gz7JDMaJtf8t5tk4FH34bMlhCFBVJKUQE9X7BT53fBRhGWFEbOaKzR7xuDE/2
/+0NIKvoHUDiSCvMjCf/bdzBNawK2bbSTHDm2CRs+VwmarXodG8IcApC47TcjLqHkTlVvQtKIDG+
2v1cM8enVJZCoTVO6T612dic+IYS+yHm4wLCfYcktldv0DaGQPc0284pdEHJctmZxwvGd009sG36
iHHjk6kXJuQiwbUs0CQI9ohh7WzRCl4lk7U9sGYNAWFPcBnc8WAd850f0lvunkWu4d3jArHPzy59
thCEWDRCjG0r92H2tUX0Dl3CExV62+sYrk6R6ZHlblZ2+zyQ7FFEhuRqT5s8bdffOwe/+7Sz1rKv
HlpluSKJU1e/gU5yfroSuHa/IWNYBrbXr1ECBU9h6VrwWtI+8lHS44QbevrW2F+ckyecMSXFZ8g1
pxBzut7MY2L4duOIZQCW4jPw8Har02maSznETkXiBNk/Ze2/1v2nV+iLEwgdT2SprqOW3LJN/hqX
gew3RfowUy0sJmERUe0x9+24lVQlzFXGxGbVW9oYzdwWCfRoG3g0cpjntE1+t/l6c/KLdmSYfFtM
gtbaFkql6IPR39o36VuY5BMSUcSQ70Zvx4Obx8FzBktT3T2yjt54SX2ZeWrkH2UCEjSIpuiRrNPw
giILaXw0/2zB/sYbXPRDk8ukF7eOR3RRc+Tpr4TNzREvy5m+EbCnO0pzIf4FEw80KZXYvUbe+Li0
rv9p8M4fD9QQgkWW3+3pA5q2JCd5PejFx3RrVLxh3Q0S663mTMNR/g5WWGrxxBdbf7qd43UbluBy
acj/Cwpu3ZYe/h9NT1H3DP5xaB7JztGnvM8p26b78t4We1WuX+5iOfGKmm88Ym2Qm6AIPJq6f4Vr
rpvLKPAfBD3XqbyYs4oklOu7kk8CHgZIch+kz7H7Fp5TjXPxIJ2JGKOMbRSQbHbkYm2GYZmgxy5b
WOa3H1mS8fknt+U/7GcXE+E90t7yVRlhLs+wRDNLK4rxmArJBm/N5RLrL3GKaSFgCbHM4W/bSr0k
jCDXp6QgOSbuqsQ5+Aw5JeGR/sb2FOS5D2Tvs3vSOCphNLa+cOkWG0Ie6sa8EDoXgHvfkBjE96Cd
vefcxFi+Erx8UqpkGjVH4nAGJCw68MPBNkaZbwU0v656KcT4jXEgx0nJt2gckSaOIKWeYRn0R/R0
ywCYSAUlFv7b5XKz87bFR5SRV76w89aNS8/ntbCq89nfc7EqCgwhnhp+tYljJlS1gHRo9l4TlQqk
G5PO9zGr3YU5uqAa1JW+z7LHq+2OoYhYpuwPUUoHwrSSH3FBZoszAfh9NAO8PzulsvBgs8jQqCTl
QGXlhk9xy3ZIT5hGHtXsYdAvtv8leqftOXCz/q8iTAzBRuXxVxUr71/DmvbvTtb0QH0+eoxEwgiA
F1XbdFbM7afguUq5F9sJ9siXbey2P0Z01xWwdWe5YBMxTUwu4TPTB0Omz5z4VGYSz5nDciOJHrPx
5aaSztI5ahiEd5v5kGrgxMV47/61pKu/pwpDRNbIy4ctMdrMojGckxcPQMeA+kUK+yNuY05tP3sV
+VGWWmORmVhL8AM+JmE6hoeJzdOv/QvV30s5stT3Srx3LDBuUScBu59OcOwlOFmgACLBNLrkhhYs
+yjwGzf61hnGlMesSEXmC02RxYWtRPVEKzrz9UVakmbIzTf1PqwZ1GTXv1xRSze1iP4DQldJu8Et
mRezE18F4Bt4PMEpOABn6MJcsdsmlSfw9HLx3O/5LhmbVELIDNe4IR442HCNpkJ21LBr2JQWbZYJ
j2D6xU7xGaQx+DM2BfwECmjnG4w7kbnu+8ayaQJ5X3CTWCojKVzRBWPDJFrJfGc1tGiqnEzfH7df
+E9k2l+W3bu0bUJxPvkDaSTn6RkjflkvJ7LHY+rtYE8dvKymvxgrCriloNOVirnwohkrylwlHEQU
7sqM1fZ6GsF9jGZVaq68na0spk2nGldidSA4jHjjk/DZ57QECiGkHpm0htwfCxxaNTDjt1i+HkyL
7fQndsOftSxSeJP3ceXgy9oqVYJVGo+omCeOQ5ECkLTBSWkAbVddhw4lNqf4pgzRlWRC1uXCsBT0
BlyFpyF95hS4Ea1WXLb7GRtnBreS+uHsfsEh5oLAf6PQf9bcTqutL2QrumhqEz1DM3xNbOjmVORm
Sdu2kKbfuY4f7iih0Mr0kmSauVxudy6IewrX7aV54YVuLe3sGlyduZ3t0vvNXTxWclyJjyYE++C/
aXmKIVEfF6BxYSS7mapt/XChYuIw2P5Ocwl/Efr5ZI9NvJdRYp/TFZv8jqKgDvzn6Gfqfwg96Cgg
x6gud+EtHSIhm9IUnjEH3RwPSF4TSybqsSialvHGQgWNwEi1ZSDMJidf7GZQOKtZJ4Vqi6mGAbRi
ywommNxxwsOsoMBpU1Cy+ucFp5tU8JFtgyNHNRmeCH2E4Dr5wSWpSJuFRtbHQDrTcAwYqL6pXV2d
T0eohEXLEwWquCCTCF2rnDDisQ9X3gXq/1X4K8Lk/MjnNk5aPoMmD4T2O6exrXmqFdr9szKS7HR5
B3NBbmiCyH/i6296mlpeDIP2rOi/D2QFd574H3aMPQJ0e30dRF8PkpRF0t6FE0CzV74MauAXYkaR
d9Cg3LYrmnNWnS3OLgnn35RV7/rkFH1KJK0VwjQsqjE3CdcKDtZv6xN6oodJucLKaSsLUxTgFcID
sqOIRWTNA8diEi/B9ClDLdT1RRK0cGXYraGfnMbH6tbox9DyPIkeEaBavR4SRaWwdmAARkalG9hF
Tvr6Ovr1GSV5CZLD32quc93yDF9h3c62HKRv+XfuwvYN2Y/5h/I2qf1sp+lpXke5ktBCwp8Lexsq
a+JnKN8QCHo3aA2xLlMSxFtc3Eemx5QWtp+cBLnxP7EM7uyL7ZNyDqhwFWsDa+X8TuasQvfJeZId
pUf3CbzpVwNmmVQsGw5H1P/sC9uh4frGE4nQ1bVJqZ/soG/o911EfxWTJo8mw21hlb3TiYGur8aj
hD2Nxk5UGKuKioLcMJe50Rm99chH3pZZLiF+K/UWgLwAV/AzmPKdwpHwpNN7tdidOqljtEykH+J4
yT2LCzx5Adwp8kiwW6xdIAiwC41eOpjyq/lJvSxubdII79Upwc8E9WY8XfiFvZDQAEyV/k4s8Kn2
a9ooAZg8rLM7aOUQAYRxe4UhqaJqBvz40HTxmF2LpigxV1VeBzItHS/heNKtkLvl9odJ/jBeKSsh
apsMZbmNYRt/bXlninC+qnGmXfox3MYFPQKCyKr4k87WMU3vLx6e/kP9+Q/xe+o/2cy9FawCDDtz
lfFtxaqyGU4kbBBEfPKdELbCNidyGplgqxn5gWlmHROQNxs3oiyv4Sq2qMHrLpFVuYMrZSuR6Y0p
nXCuCZaBw1vzfHXixMEn2VjFpdvI/0zAR5D4eT5PrebeQyayv4Lk8hOjbWjbAN+PVPrvBs6acRU/
aJkIMMh90bEr9gosV+tfOnUTONyj+HK3DT03a5Z9AoYT1Fi4pFUNQJMPjZPJRttc8ZA1JnCcZtfc
CHDfS0/ohJtEPa9x0wTE9hBDAUN4Sy+uR33iUM2SNBM8UPc/55ST4m6nlcXMCIZ1NG87AhvyjMz4
IuE1T/2bQ9LhCmWQ6Hp9XbBsxBZGbU5fajngMEchIf90Vaf8zB30vrsRIJ6yBMxNWaNFAJ7cI0pk
dgudjej6ZqvvxwHAkpMkH2wOYYexPxXwURZtpV6y00IjKKQBkMBgrYwpVBOG824WBsSAXW1tjLtM
voYd7s1cfjxfG7QkXTffk1PnS+Uy+E0WhcYOz9Z0INIbuD5HamW788ebenfCA0uAdfuh6UuF7Nxw
irWp5c2vEwwwDGDeHUqvbx6Bx3MgGoTRwaD8DRLQJB0yxfSq44O+28fAVX/QyG1jnaNNdbaJ2Ah5
CoaKpzI+FqRqbzo85Dhc/ua2c/pPgJC8omvZ5WucuK+xdmoNuFmT1prwc70IRSNf6L/P/Vi4fMIs
iKS4FeGaX0swUhxN1OAnLTNpMdCmvhzX7xJl5ewYv+37M7aSK1jBNJeOBW532kSyE5E8T6/DWvtZ
hjJA9vyDNxwS6muoqRtOGYYEIHuBxgrNjbXM60EKYm2XPRwytz6zBJeUMF8+XETpQiI2hSkSDeNs
zKKg6B1TP0SfsFukOcPHmudR9I7xFnI3W/hNz832xdHsHo0E/NA7TA+m/b1vIFP3msdPz9Yv9ODf
khUc+xz8+gjzauujI21S9uoGZ/H1tSYRoq210sHZ6lsq72pwpVYxBp4Ng6fQDiiMfR16hmtVTdI1
Xg8V1iLsLJ72dyHgX2rlMZP+759XpeIOJVPd2dYq4DVVWUGJpTJxkueCbSOr1f4lvUos3mdbbg59
L+KqUM1/yqE2wrb6xMpb0rqMgiSWiTomuFyp+MUe0joYYa+03fQcvL8nc1zXcqoaZQ1vLfZ25HMU
JQNWBiAV1q+vktRKbvoTEFo8/qAFmWslwVKAZO4tZuMDb775/y37UImx0zNH0z6AvNgYVZItflVS
moJyHQ7WNEkiXigpNR3FEQVKZrc0EAJU4gJjA8QOsPRiYZCzLzRvw18L9HvBrs/S6+dujvUtRzK+
Sj59+2KYsU8dnRJqIg8JUB/AUl+KichPqg8zjEOAiKlEKp7Gg0S2AEt2uIAp+YIpglcKmIdF9avC
gwM08LYkmafe3qUIJyEAY6QzSlkbG0nKnpfGpaVBC8qrNGxYz3RGhaYdykbhllpsxQHuqLFOQFLO
9BxbYWNY4G2htWuLNxH+B1VGee7Qbe1JlQFNw8WhjCAQPgGR5ERX9R6YC7E3amwv9tXD0/RtyZ2m
tS4t5fxjXs+Imjf9SbIQ2oSm7RSpGlGwMwwAoAxhVrAYouaMuJ6AmN3gaFvsX9Ul4AzwmRPRbp8X
Rzs2nufzjpAOFj87n4s+wPFEKP5qP37rKEmUy7JirtWSeyKmk7bRTI8FTNJYwO1SNybh1e4yUpae
tauACcy1M13XJCnVXVDUVoga8wxupErzhHIDuB/vYQiAaWWIb8gaMkMDtgcGIf26qQedYpcFMmfg
SLWvF9/67D5WqexQhg5f1cBZZJcmQZOsDcFwZsTY6RwnxDyY6ABiLIAj6JpQqhZBcZK+j97tmNkG
HaWyozovp+TR5zSDAseXjeB+FC2VLjyO1dd4aB9tYAWCXF1Wy8OxP+UyFxrBIRHiU1AJCSPa+9XT
E1E5ieY9yQTlMt0s0LDI5lxyz/nkhupbuhvin/SjQDr8G56ejQt6gjTH1MBQAejClkRGg/BAnKfk
lfcT9vfVhc0aOpZdPRP72A9YkXkG+V9gDg06BKsQ8AUU+Q6sGcO4+2eIGxNAJuRfG+Zerx6mw7gR
hWSiEg+IkEz1cKD0e7PZOJeqC5q9im5H9aLJOK6Bgijijd9si+1JtxyRed275zZPeoQpVZVe2Ejm
pp8BGoTZDjABXOH+cYyyF7TVlPvavmC1CxYZCGFPQRheYVZQW1Hkr+Hx1vsuS8ie9bXcxTk19J4z
YglkOkqOHxDSInp+6lKFia+RIamIk9VuXvhSfHdi6xWA4KxUR7bRYEuQDKcX8uFPfb3Tl+GskGjs
YDqsZSICEdQbulqvKEFbyp0nI1pfiyTgZuHzwNU24UD2Y7Fc6Al9knngjli8xkady6yEa0dLfR74
mLInTjqGO85dDv8kRvMOyKdc85swLRqUzBKId43vpqGT8v2PjPniUwatu7+a/0tA5XDLb3Chl2CJ
SLW+Cn7P3582Yw3SszpVviYori71LBSApc2CefhyWBYwQqFMKBloJmpYPly8hW/X4b6I1HeqQZw4
uXMIb8U5gx2OlepIU2MArqDXJh8i5y6jDMANDBTQV30wn0y4G1ovsBFfkPxUx52Euiro84qgSftJ
rJfM1+rMPbAyAdDBz5ToAF/1bi7ZXUaqiRogHnJvV1CO8tUzUi0pcTMmT/HmrbwOk31Pk0IHgTXC
Qg0fUIfcSl49cpuhb25pfmGRxPbrm+Z3TMRWV1UvN0swsGi1PYEyVp9R3fjd2vEK1KGoQvsR5QBV
WBXdyr9cTdu47+z8CbxAHfeqVi1pQvEmXHTuvQzr80AT2Vnfxs4o49smufbhdq9efMYFczmET9os
v00ER1mO+oWT8fOIVTJjfIX8vpt/RVl7UpWFFlCSzSlSKaDcqQq8N5qKcegscf+7xZAg30wx/DKb
qJUcRtM8WmICv270hOli4rgdlhKnbNsHSuVfP6JLE8I59V4DlOhXE78XQ/nuMXe0bo+VIRBifKko
rIKK3x5UpyppPFwbUCyXVNdyn4BtPbWoyuBmTXDDLF9oXhm+g8xjxQxWkRCJ7x+XWuICQheiLNch
omVr3wDkvuVXA1TMZMC9biJFFjqeX0ssR5cM38HFgbZl7LWT0yTYTZLb4p2e8YJYSegPhbTn2E/v
f3VTK/vquiIkIoxnABe27Jw1V480biRUwb3q8lXnjgFVz/UzMSnEcvidp0P3/xiS97Egtvu08AO7
GRCuO17qAZslwM0Zl1tDGN78iMysCZUnual2de+EFYzXHTrILP1Svjb9f3bqHARLWHMYOO+7aBKe
t5F6EVUnZpGzbcKpsnfUwAAlpOwXccSlmHyUVcmGgSUWrGY9tSFQ6eAXuhKmU/WssFbavBkitEBt
7EqXaP04nP6yfwpOFpCuDSOFpL7m/YUFjKNrP/pUewrt7OuHNN4DYG9nSS+rVc7Yeg+Cvo22JdF+
FhbH128qf+g4R0U5GnzbQ/xLsMM+DaU3n+mevkFZG2H7Z1rPEuybMRog6TESyx+8YNGQr6yPKCZq
pH0NK8DOl5NfNKjszPatr9WY9EusZisVSh0U6VtvLORzkWMc+9IrbYkv9GoMy5W9xZ+mxvjiFKOb
W2PDph/3kgr+bTo5ijfqu/PO/1dCqqPC+/iZOIBy/Z1pHJWixkEauqrbAr1CHUVRPRcTk7O7oGcP
eDAx+jn48EhNw/wVY51Ux09xAtiM/FRNrt32nddM9Mrby8uDlwr3+T4jPwMU5uMUs/Oazi2kNUIB
Em4WVJI+vb1YdE/n7Yiw0KMgx8MvvasUIo+JZry9Zr5pj/epluxR4BAZguDVlxOv5tQgGBmsqIy4
pGETZeVMOw2U6ZFZ6szo37BR2EZ5KW64o53RiqrzXFEZgdfn25DQWT+IkDTUaD5SjhAtpKafca7/
XfpF86AamXK9tfhilbKfQBaa9mCcCuDbRQ6IcXm97MQTg3YK98PAYhn3MzXyQgqS+XBbfSZfTvxB
mPGVa5HpZHU+1F7ek3vpG2lxYCTW5XcPjqHFExPS9Q/YJ0bpDwbcdllQwMNoZI4iAS1Ezd/3W8X3
k6wsIoJwUKk/zmPx7c6EviqnR1m99Opo81Uumr3e4Wn0Pj22XQgPGwXL+n+0z+3mVVnNwQUh0IQ8
52mT34fCPxJxjGnJdCOrwHZrD4gwz6/paPb/bIUXZJkUUvUCVNJR+8z9zUDRwjAsCrNN6W92KJGy
nhQBlB/P2/tYwT4CLZQvKSoMcAG0JhpOUhcmCNl6o6PMwEOIVd2Kl4xAiLF8UsPFCSCmuctiOg7j
FTklOXfdA31NTbuU69xHnfRf+Zuu0qLGylKZ+UexW2vQUnXTLhHyu2/1gQehjowV2AXrYgswZ/wm
lplxPRh6+2i4jharh4z8NnrJM74ayTvx4B08qrfYRZ6tr2lFOXLYkzpJnLgfc9TrdZxvy0hmjtAg
+VE5+B9SmxGliioLMXOlOhsXHc1fnn6SG/fevGtlZpfUFKKnsFcwIigOM17zFgt4p2j87lbAKZ2X
fhIEUv4SBkhVCWI7xKSWVrRE8hVVfOKyvq0KFkRPbDbjeeOa78b79PF21SL+acXFTyE1hwvVfkY9
n6rXmcMqCVs61aR0dDGCjjGFoJzPTuJqIBAm76nUMi7b2HmVa3m2pU2S3jB6zo63I+AJHXGc/Daj
W6j1jWxHAQE6gu9rqvQRZcgvuosASXRPRjSb2s48fUlOkImCP3h6EJla1XNmaopgGU2m7ETHOXOi
M8ty13wuOVP7MmMmuQOa7FgDpAHi8h1nSyfP2iKB5AeRsXK5PFwX+APBjBsqIXfXV/Fug/HdtdhZ
rdfmuYJLWkQdmXTzoemPDyyswebygfdbWSyoeUNxiYVD6GaSmStmSPWB7qzULbYUpAnpbefzTK06
vHE3NTvYUlbJZnO7p1NmNjAxmoL6c9Peno7BqI+80BpPOGNI/ad/iuMS9y5ugSo+65m8wPQWkOld
SmdOjeD7Dj85LpHm8e08iYBY26oy3udkwudl45Al0bIsl6Tx05G5s9NxWnA6n9iL7RDvfKmnEDpq
RBVU9bvJ/qI5SlKw02q6ZfBbGjR+v4oTFNi2j9OUFLpFWagmpwCvjNu/z5vFg2KqtdlMJhlwq8dI
rds+IrTDBEMI0cn7C+W/iQ6vvxhMzl/PyJg+aM/R0OqiUqLJjzAWmJTNkHkQovdavnCaxYzJKSOi
/OkTgW5P9AesCGi6WITTlmp+AtxcCZ3RhbU2MdtXoCLsjQFridQoI2mobdyiSjit5u6jk/Z4RKJP
w4U05Zbt8MYpgNN7JYVxtFn8mjVBCzg3UU/nWFafgDPOIRgy3dwsowTZ+6TCSJedywHYE3pEg7jB
ty2FhrmkcfUu688XI76g5D0gmJLLepuFXsJTeOBOJwDmcUeh98XaCH4FGrZuxNKYBHNAvMMg2WxQ
6LWqxWQsY/VM8IOsZBGGskLM6+hdqx9X2RRchGk51nUvsnCVH5bd66Bg4RICMIX3nPDGJ6VyS/4m
AWygM2+hSQ2e616f2/mKev4yTKAh+uGlsj3+wnj2jRtcQZkzepSCl+AylLSV2y6dGiCXCUnJ7L/E
5xHSOCNEeZi9mKj//ik2DKr1bm683KLjBHyNLke6ngZ9R0RBsEi41bbzrEpE+XRbRhY/dH9YvCrM
AvlfMiYEI9ccgE1eiUOACH3HKJqUwAPzVW3JMa1VD73OHMv/7bH5Za0S51txqovbTT+QMxZMGtdn
NGwapwgeCgNr6RZ5qAgHkgjrO6eC22WQDrnvt+lPLOJfsyUbJGrVshCvX5Veprswp+k5Q9g+FM4+
mZFzpFlpn/4NYQNjXz1RMwLzbhw1gb2xkPFCwkg9bv0HbTJW1QsZoHkuvEURbaC2Jrf5YgWqhwFh
8wHJR2IGX9iei2UFV1OI1fcDJMmKPXs3JmO/MPxC8Yp1shQIKqYXOLvLs8Q7fHG/fDnr3W5KhqpL
eRdI2xY76DHfvgULRUxaj2fDMBL8RktsLC63x0/VWIUPM3RgOa+YctR55n2tEWZv62xS7p4dwmT6
W7RBWIz01nL/BPEdg/ytw/Y4ANHYGSeeXNNhbFk5LROObPgyyebJz2LTUzgTIhbt5SKiE/ub8KI2
3nWx9ugmrteG6Li7HZQ+/ig33DWUOMKC7bf2jHjxEjuIzR2xrtM8Ff+rwB6rogBZ3UMCEmgI5ClZ
7hm6l18XiiD1RrvICWCx5p4D6O4koiUpXW3A1vNGHpPOPrywC/dwYNRRiZrieOV/MTAJOZIfjZAo
lRQv3Q3cjmMYkF6ok1ovObLycgInt1ZH3MB1uJsrNKVhYXWh4LSRAMjzhMJgAX8KYs7Aue5HKPQ0
dXCr0Fh/nJQcHwPPndgbxPz4YrjoCWxAY+DYCBUnAinYAm2xAuQvMz9EWs76JZT2kvme6Rt0hg0w
w4WK1PRUg3QBb9X3hHWcVCTrwbhPl0+reMKYTBlE+PWRnrYw0A8F652zEIgOxUDcIBwLwErGH7v3
dwNrZf04uQmxeiCGrqzFy9e9DIKUBNLtnUXfAhgF2xh5mxX80wx6G4M8q3Eb8s2c2KRjyaJySpQ9
g8zkJfViaTCauXYQv1lk/XDsME0PJVPlgGsEjjC2ewkDzLlt6VFByN07WEidspRW4+1kDTek+FIZ
jgEIAHEKtTRSnOGkHZ/b/9qybOgO30e2A9e+2Btz+12ZKvKaPImIOBeIg6oWa4MhU0xaq9aR6d9K
d+34bigCNr6KZSuXSlK69zDiUCab0dfrzzjhaf4Q9ExYAO/ppAF2KPFLrg4vCA68obVQQGTjdmZB
go8YNvRHOW8vkhDt6cPyDqsoQ3hBSboAlBvorasxYwqK9SIa4BUOlbDfmKW9T0TFBKJG30KopxhW
1vmJzkee2xeGnZKn1k41u4l/suzRu6ajj+MMnTlSPXznmrSxn6SAHhbJBoiGbBqvnJ3G0pWM6OUi
fHRzMaUapqCL80avzKnHyaifUz6BqeaK4hq3FPZlshYGgN5JsQiNaWBTXj/uMksdFQlNuaI3u1xq
wLWbxfVjsAsl/ZgCY2199icnH6m4bEyVzU0eLMV4rpwP0E7+EaEiPlm0Zk5HNa+KWUJ1i/z5gpl+
qfo4knAl4ijH9upIGTXHorU4NOqc3ly/lr1jnRiNp/bBbUmetNn8zoKbnO+O27kpPwWulOWCrn/F
8U9aQkrZImKteEdKFRH8p76xHH62CApvKNOXLVhSAvJRT0765HhWyjVbeDXHk8J3kjFLrKKT9mBX
ebn3ePCuO7NIHXZinYg3ybTMj1vuvd7MQe77WNsRGL1avIKnrv5Is4NwHQ4jhfunYlnCJ1Tnia8I
ODjfaVnuk56DXyh+ZZMhd0H5slAjVtJJKNfhXaHlSlFUvtu4Xb/vjWmlbfw9qCT8UZ/2pnVMYKEw
Cjt/mC6yt5TWpFHj7nK0dw8ts+hnjArQ6IvKBl/yvt6uDB3N6IDHiJQaj5lIM1XrFCfw/szyydVc
QhmoxtrR/KsfrxGNAA7wFmqsR1AMW7po2S3wHWZq2c8aiB0n5uAz2tCva61b4VKzaL4vFvfJ+aFp
Row+3J01Dt81Q+rQtyELIlW2MLIyEmza2B6ez2kqzM3uKqQ6d/ZreFiiGAHvmtaH+OdwE15LiN34
hwa4Yg5h0XT7Q9eoRCdMmf45BKC1w1HJpnUqxsn1CzBoHfD02q9ccj+uLQWm6FZKMKFjd5T2AbUd
nMGTvFu/6GDREBl2PISNFE6qBVPQ+BNHZYGYEAuJ9dy9BNA7gDSAEr0I9pO8gHGiFOwK1PUhhOOc
QQfLow6LoJ8LHfxkvH3iZ5UOSvEyAJjgty/E/6er2J5CNs37rsuhzaNjyD5eH1D6yeEakDnLlPy6
PiA6hY8GAnrnb9x3aTc7w4FNkT5BO1l3AalRyaWlBYvv9H7Bs2xuRtaIos0wMPlGimRsEpr+48z/
awPaGGOjuleILTFw//PxUCDLHByOnfPwUtkxgKphLiBRUWF1pcaJaMoyVyqzWOdRUjbBwZrrugI9
gnBqwoWRpdHD92e3ZUBkEoXgABK/7Fg2uMDx7opq5hsptYDUCiI3ELPM7kUnOvFMb7HABKVhYokR
b9/VFejBHkvhpRrpEOwlmq6QwuM5gLfzW/37Xf5HT3rx8cWJYT7fN8wA1kfyKaW+nrKWDh96evSp
SKFrhm4xwZm+IZTinS0IO7a1LfQyAEtbqHFrLdUaxwNE2/sNSS2ZkwBa7D3LwzeEzD2qkCJBE/HI
IVs9hFnOLZpqQ283uPkI/Mt0TB/ebtXOaOntzG735O+XVV018Fw+XwnpdgQk3chtV2VgItv3MAU5
NqXM/R5lOV25OKd2jDfSjNv9lU0J/WaEtoJGZxGF+sDtPacN9E/c7aP4SC33PvIePWQM5cENiJg8
HCk1cL8t7Ctw5qZPso2MIOm/oTqsv7MfY5IVG2vAl5ug8trI7/7xuCSF1d/dqDTt6w7kdVPsMjXK
wUwhO1v0Ww08G6TCOLLvvIj6lOfPskUiWR5UuXRYIkZ1lkpSn/QYEWysAGzrH7IWZkUYgsDBqmel
hXVXC9ttEss1YaeZy2S23j0QHjiUuBlYYPML7s+b+Mi6H/5LDG1WwUsV7iys52D/eH0f9qKyLjkA
ADtB1HuBgLKd9769HlCZ/20yMLPzUv5Gtzxpjxs2+JfxF9c9rsxQbxf5vpj/ltSNRJtcmlxqn+q2
rPc7ZIVjObEnZQz9o19KISfm5t8FbDCbXpH+BOz8zz7E8zkWK2es/4/xMBCY3ZNH81ugkESZK6Yn
6iMKLKh/1pNQb7Cai/XMZioCLcqqIn9ABkKVfK8YalRw5/Z5Zeu397dhrdyWQwU30lpPiRNUA3+2
FECdAzX8dcriTHoKtiJWCs3zi0T2qgcj4hoMVQ9o1kDi/gjM/aAqXnHESXeT7noROgONarOZ3VdG
f0zn+7WrBRvryvdKjiQ87ozJVzOi1bA7ciD1hEGNYdpIeENtlMXIlQAM/+4eEC0DxJAV6wew1bsQ
IOc8TfyAjkeXvke2eqJPdKIO0QFx8pjtSg0sVkM0H8hdlSn5tTHAKZlT04QgPjE1Apjg0KJOl6ea
8uygFI9AKRG7oIlFad/DKtSYCrpdjiBXiyEaMbD18CsR2Pvy25Nhp+wxZhWyTuc5s0AxKJCjguKm
+WLc1BXqzdzaPj4aHh2+dsqsNwXqoYD62FfbcoC3QD4zxJQliemzqWwTrL+E1WOt+JuJKi+ttv+R
9UOnbTIXFdsZjsxJFXp7iVYhBb6uvwPRCTpHB4BueSSNtddxPtYOw4QrIm5VRecroP1zPh7V2KDI
anDaAKOiO39ELhxejH4b5xzQLnNh5vxI1MyGYmEzSndrP/ndF3aSCyohNvtR8R/9RvkG6nOkChF/
Gb9fpkPoFOsIOSnbJ4+TC816/MRQtkFaQR3Ok28XEAQwWVFyH7cd1l3az2o82mNacnb8ZiiUDegp
n8IOEO+wpthf/sdzcJfbVt6XkU3YAokfggG2s0cBKjmS3OCdIQ49nmfjntacoYnyxu2+cBwpzC6F
Dn3AjUJWCDc0SeHnf9NG2ga1N7OhvX/qDlEREkbkX/WYr3d5oCPw+iPDKvGwpughDCxljXVtd2UB
kIm9OqM5jnkx2yog5PeSbOIPThzimCr70w7/kbKI8IOBYYgsD4UtT5Ssqup00NPyTpcIZ4TK+ZAf
3GusvR+smdcUDGvXfntQxi+7nQ+gvhjyqFxGSITWhnZ0AvfubCDoFzRchBqb6grbQS4CKjzfEOB/
elH0Lx36seoCP3tge9OwGHr5gkCTmfz2/KoXmKdvvrliv/+bkHv/bTruVsZ4u5C/UPwWTGHQW60V
Ao9m7WqZLlF25mhgyCl8YrOdYLKb7QyIsAOmLE8cHn6SEYrUh3Obhq7q22Kz768dTdbQ39Tjq8Xr
qNoTwAaO4yd0iYVbXvD9yZhNmdiNun3zGNu8xqKZvq5u0Z2EWy8TGU0g525erou/WpFuvXOUDHzK
Fv7Z+fN5MjPkHyFNg8w8PbQiNQf/nZBv6lILKqLZ52Dk2WiUCP+gcgePHB730+deLzghERUFfBJF
MdCaizz5N2jvBLmyylK4OQshArpyQePx15+F4HXAisook3TKzKx5Wijmcl9X5O/kt/cxAxi+m1Mx
b56JS3r9orIVNOyPMDpJDHzvcbsINsPG/plKuFljsXb+gijDrF70J2zbPSpR5P1r7wYEL3J2j9kj
bhZcBW5n9YM1/Yzu70ckPETf+9jlvFYe0x/re5git8QxhzTMIBV44+c5H6zKH+r1fDpBvCVEYg+a
b7hEc2urc27/bAokKlGvg8RLaYRTTapXW2TQ8Ru2CRW3wlYWcbd5bNFrrL6YwH1CXkIpCzSCbfzq
7zZn9Sq5e0eQaitjWBj5oMth94dgwrxXELkxd4k3A7jpkNxTy/6LyFjVlfhae44aQWF6gK0zH26V
57EWPIfuzvB+pybGVJagOGcQbT5eC4100Tgh3cqWCIr8X7lQeps28GudrPdDOuKtuY3KCy/OMQj3
UoXNh3XRh3TmVTYnFeYSuRfSMPjFYA1++pd9tP+WGBS7gzFALRncaRNBrGGa43LC20K5yv1E5BAi
38zGOIC+CCnlkVBQ/+Ajj4Rrp/PVhza48IT+zY6I0CiTns3iA82DfJn0OP1LEE3TSAdmLMXoxX54
WBxc/kia/SmkITmcicd9/5Zl3IOIKnwiujiS2KRy08yK3yXpxf9J98XqW6QAlT+htvQPJnx2gulH
NCFrsY3g1kiAFK9aCvjgtxJpfUVEJvqkopSNZ8XTthyz6GL+c6m7p62LHUz5bIVClIG04ETFpyjC
iJZTZ5J57tz7f9kEkSLsIN24jBMl8WbHHMX2YOYtHqamCRh0VmONtijTSR4ChHatKeYX7hcQRZEg
5DJs3KO7CAO2x9NK0dwy7Oak4EoeT32qSexeK9IYTIIhj8bV2sQH1KK08mURscJa6cBD2anaFM5D
hWmxLtXj88W6EQaE+VmqvkcwhwgIWusUS8lmIIY5E2V/N3G/AzKu9cwaosoosFFaG8BCOFy7Ho0S
PtWpwqUevPZwVmT9czbyw+Vpvl2LSqy+4RtqDyU/MuN37l9PpyW/ZDv0ZZGWioMpTjfiXHup7O3B
cDNNe8z9ap3Yqklh4PXpI7qohqsN8KErm/US4VCM/efz1g3wmdMimVjZftAEXraoYH9aGHFVhJJS
RHdZZEijdXs9XKF1YpEijQdkO2MoM9mO6RrTqbDRTXgxk3g27zOOXZK38V1q6+cnsZ8NsJ/8nXyk
/BMx2NFDcUvCMMiPNUF90QorEeCkAjfVmIQ9GiQJiXiJo7xFpBP24U1EwaSzA3CT59BWxeJXjy/h
GzAUynWJdKskURn56rDH4AK5BjpYYzBTbRlgcWS5//bsGhj2NXtLGvj7sx/6kiGMI8JiPN/fzYvz
lS7RJzI1B0G8jZOtcl72yVhyuHWAl4d/u3sSHfGY3lS+Cxu5wmI17+Sz4788WSn+ppnfDau0FHij
0woUtu3m6OyNT0V4AI82VlWgbkStMG79yigYifKJkhl/z9exsfs4GFGbcmrt8w1aqEKOEjmcfcb7
JuEUX3OtvDug1ZkqqJAqlxk44kdl0pqktAAZZrBOoYaqA+bOrJ5JJW00vfBgqcxXG0WTQCFwgvu5
bZfmQdi7xBh8HIqoA7TO8LYROK98Ghgjz4Q4/52ftuHSutWnBceHQA2QQBb6OY8AptxaxvXqEnq7
dyObTwRO4VshREttsqmowNNWirnZug2AKhcFeYhY9vOSYrvjt9AMmpbtXRsPtcgZCVPqCPup/gC1
6DJcR5pfCV/e86ycFbKfJTrPkfvzUQ6Latg1ovrN7fGk0gFi4BJtbNzY9l8DUeK31sk9XCOB7y9/
Eys3ZHionyNtG0y/VucxVH0lcW8Nu07hD+Qrz47f9e2pHKTeo21ghVuzVek0DAXgDBDV11Da+pdi
+DDJFK5gMIAUsgE9IP5G4hgUqjpSgG+JWUlMQVKlleG1X/vtaRhlu2jWgfS3HA/CANZY+7xAMBOw
uG2ijTNIcIs7uYn6uMvM25U8dr49/FHp9crSAdZ2UG6rAbwlTdUPlLJAqXs8EX9IWk+jReQ0P9pl
0+aPuKMU8EF0csSgokZl3FN6rLOTboMQkFgrfKdFkzDW5aBiveY8uhfitBgNZ2r6PiGXBk2qrL+k
Ihpsqwe+aSZWU6GnK8x57Xm94/VxnsW+zyitxCGfkVLdeFPaJoo9afXywVPd+nrJAQ8bLqRRbcYs
YnW9v6bxWpix0mp/wRA11A1EcfxI5rItlN1NPyX6nbs+bAaCoSg/XDJXMJlCYs/6nSS6FzCBKF/3
dOASQH5VsUP/LTcoG8Hak7RUjWkKN+l1F8H/RISZGS9Vcxd0zZLStVEOHzEZ7UtA8UeKsaR/gcqO
s3l9NmVJo4bS2Omb6nWN9unSN+ibXZn+fmQBxHsA95fjLMdJYPigf8TsVp61xGP2DqipVhCJS61G
0AGHtX5tS6fP4MTGuhrcYU2Rfh7XZNYnqIJcJA5Vzc4qxUHMd71BdKzlSSPcqJKXFzbe18C1nNDG
vwAht6sVyFur0PmM3MrbnyXBJIPhkDOrzIq21oAsxu9pm66RAUOLtGQQaRAe7UknHbSl2BidONqn
ZTwpt1+4c1T5TYACV2zdI6VeRyc4FvkW/CaZcckAPubvvxc9M+8IdeI+KSuzs0dr3ewpnbQJi8Lf
/KRqnObUDvtdDLXgokcCWeuXgvw/6agkqJsRJiT0WIZcZ5q++EjRz1wN+XwyOhCnvh7T9unINRQB
EC+sinhIJYbWH5f0uTggsvVvokPrUvfwC2bD9kv1+YhO0DEE47Z3lpqYklXqGSBUqKM94kMlPL9R
tNgx51gm4/Oe1bTqoBmBaI15x1GUhFPv8wev6d3Q0fvEIFgSRCEoOpfxwlOPmuydW86Cx2LkFpNb
Ilk3OR72EEfCEw0LnHyXnN49Jn6b93ZdRjsjpHzHCgUgNFrnqj/Qrbjzq7RHdP/3RyKc+uDieZRx
3ghmCbPDJ8Am3qvA95ai4B7q6gGUZmoRCNBNGtWCxFGG1JPMH/aVED7R4Y96MonXv8VbS5Ltfw2a
ku5YoOXfrXDNebD1DSk5j/a82GgYD9eup7Xg0Wy5XpJKsFxH3cJqJc2K6eeeYng/m52f9/zj7M6N
M+dqO/5yph5hwKCeiYtiw26dSw2ny0B7iS4FvZGcGUhj0p6rC04KG4i38SZYgZfyig6Xrls95NkR
kwH1Ampv19CA9YJu6IxMFbSMjQJ937vJ82UBi2XWgQRt/vN9ZpElu1q0BDzKS2XyWN3tTnHihXjg
NScxds3OBg0ZYdTCzk53ufSlGBmovGv1XMr2aufEUhYbmty+q6r7FYYO3LW8T03iPfwRwDTG/8Bl
WUBMCE6DHari3wzTzZDqZOXfgdt7cZSwxUR9m0IBDauc/Dk/bX5R0NUXv6jX2ZVOU5KyTAsgZFRq
ym7s1hpISVIcM5DBFdNRjzr2U5TEc5T7Ez81RGTdf2RWy5dOMcJzyH/SeDQTLEJn+Lp5lMlqtx0M
nGo0BBGdmtNAzMJsiigRx6CO7b1I8oicfXKCgUDMC8OAz1geuWgI2+Bc0XIY4orG1a7TYC2SLZdc
aK/ePp4/Cstx59ux2rrhluz2nJNpmnQC9zf6D+CTyHQxlorOvdN86i6mJmmjCNSKsWwZ6SVVNopt
zTj5vcYqBFXCcphbFLTWyGfICs9GJn4BTgS53/U+O4puPgYS05dRZuLyBhyFK4fScfQ2yzwwzFEz
6bXQrcGBePctnYtlKgwFc39PVtWoZ7Iip0a/vNdgTTRbdzXqlnKy0EAv2spliRXZTxpby+GDSIwT
XPWxP3KkM51zdqv6VYzDyc1BNNM0FLKrdW+mHmsNMbRnncXpYTM4jl/GbaM9zLou/57moinYBByW
4dynJWiyIPd0Vwe2htG6vnv69FrTYcEAfgHsKNcnrsVT+/81tEt1JdPnocl6kSmRsR2bA4qjpWeW
u1kkZszOppGmZnDh2Wm7YB45wCBBC3OaPM99pRMNxMAtY9U6rrTv/viTWtCQWTnCbreGT7xfOU5M
fqkdR46SrTXgd84EXromf3UTVx3GLcKfMPUuZTeQLBbosFsVOaoIPaI6WCLzSrRZfjPzdJsBeSQx
6DD0IHcjoygbqxRyvwNyKXKX0tFZ083Db2M2IdMJ6tzBcuWVd8j0233q+dgAG4dl/Q73vXT1S4W8
/lFedHkwSOob4q/6jgZ+dW+rjOX8cFqqkJKskQA8Lzikn5jkmmO7I/z8aRzwHNPStHVnfCXFxhH4
M0kQzhC5XHT12MvbGelK5ytFavJqWJP7r66YTCzxG5QwejjOCx5t87rga41dhzjtQ7Jjigewp76o
ZC5SwQa795tfOb50/NCItEWiEs4gYhkSCYB857uLIdbE8STva5YQhk4DnV3xyx1neoG5g877yzHW
wv7J3Y+Id2Glw92fOAufnELDokGGydQr+Bjv6t6hdoItmKaBFdsIo8og5PHiNUt4h0QPAS5N68O+
iSDWvyzmCFPi4GY014fz4WklE0cKw+KrrDP40iso0vNcF72zp555UgHqT8OtkvW0D5KKmFMgPu57
6fisNvTlncewXnenHNPzMaB88cYTV1IlEwnhzwURvweS+q747qQRjFQ3Pej/JRZjPtAQfQU6ExBd
873Pz1erx6YMzqRqH6PqVGt1Y7I02kO4/lXXxlwxId3aJgOY78v3dOsDAlE+3mWPt4YpL7dvFp3w
oy+6KGdirsPvZU6uOMO6tdv6skRKFhixY3LF99MdRCOoUvT9YejyMnXCLuwhAwQ4LOotkPOaxNKG
kM4cXlRmvFTwdrWejD2N7+Gjzvja1VvB9sZfHtcILEw6g8L92TNOQ5tfPXjyvYtlq8XWmSB5sdLg
7Ueesf/HdvYJnuloO45gzrUCmch++gLMtwYxfTHd2HqwKmromZjtMEEFctX1SgadTkjxw456VaX6
ITmhvaoGZrjutAsXkGQA+nscpzruobTTQaMZlgvwmPhdqrWVMVN0luI5JAqQ2t9JXaOs5CBwvwx4
q6HUxzrPAuct16QYRWRYlGI+mnatZyIDZ7p4S2Nedaau8vXzghZKCmECiqqhzqQ/kofnd1YlZDjd
zbsj9yGRm8doMt1oqaixw0plxbpsfj5jZYnV/iiPvpwP+ky3igyOGqtLxrw2cKDRY+Rg92PtLjd1
Xon7UePUVt+pCHEpA4gl5GTee+XQjybCuL5yloGugjssYwHe6qU/vTg4Heco4sTFyOxjb6PYtbfd
4IzqOWX6aHFvu/E4qvGBub5rvZHtr1oyL7asx//qFEyTueUrPTTcrKx+IqveVs51IAU326bIgOjT
eXQAQka3R66rwBhDJfwy0/gvDfhr1krX7tqGgWGNxwDZBIfa9Z9cAaxB9/KSbGJHUjLU0KJNlzjw
kM5a9mWTbyBVjMclS9fPzn9dDSDvz8gIIWBekuz1rXomZqQ+i/wllj0BiRXnS5GQLDQx/NzGowEY
Zmfsr/aLkLXiObaDHzq3lgg84+ZPwrT7XZv88UbP/GkarHeCPgCGjh7quLqOYOWEEmJDgBieujtl
gjxEZLm8GaM1A1VFrQ+sSzHwlYFwT9Y6qD55XUra2DmZZI7y4sF0id6p/g/OSQCNgTmgSeJIWTU8
jHBA9PUN/k0/6Ft1OUuczASOts6nB7cAELkKYAGXI+JEw6QkZb2iak6PnhGAFAIbVrvehHkaidfg
jj2zss3lAjWCXH+HLtycX0eSUDlyRDlCD/iE50YWnlP514asRSXtRGWAw/wr4qjjAbCmd5edSwmU
+1Km+G11pOniaXmiPf8qkL7XN+GeD6LVJ58F6MZ4QSysMWHcSXnZaFFEPeK3NWq+LU8oTGm60/I2
A/m81uhUYnB1ogD1wxomQuTJVCPJueRdzaLaWdKWkJmHbr/B3YwqLIkpERTZwmY6NBIjBrE1xrJn
AzW85qPni9MAr55LPkhv1nStQTqOI+SySfHykkAAK7vcOQXLlpoyyQjSa+LCnCddCv3aSFH5wP43
2YiBWYDY31IWUh2B18VDD319FIuT3uXz8IDK5j5NCLicv8oFf7BS+0E+Zilpqj0Fi1cpru2ALM6R
+OqRs5EFkUVJwIQEgdStDg4YeoTwCPIG9DHzdNl2KcMcfLRCaxH+2uJLAMk0BwLCwt8Id4es7Fss
mehYizDrQFbBLOL6Gcwvnkb9Uuf0Puqg6EP4MhEAzXvadaj+69j7vafQsMbNYS0Ccoj1lT8ypJO0
tLpGW4B+xOQ9e9rotg4S2MmeIfs0tfgFghIWkx6OUjDXsIVzAeAxb2tWiV8DHKUMo1mvf07Acnub
sAjoDen1BtK3TjMz2NSx6IxdFiyY17eFeRb7/OBLVV00vnAOsvAVv81mjEUzEKjRngduUw0gtwKp
ZUz9OEFbPfPwgUYhYd8hixamBCyPeHEA0Hc9IObu1GjKV6T3fXeWOpDR6IW/JEwH4yAzcsE7w0rG
/RtEcl/6id6tETF6Vm5iyo4VYLpDgKSsQzSnbbA7kaawn5bE0i1v8SnsAkCB6EmSwbhy84WoQqWa
EUr8sWyLWhjdCRBMsH3LI4Lh9QUIPUTL94rkBBIGa4gb5a+U3pyQ+vqwGntVHizAgFYul2uj+aI3
5GaVOmugjVe+3ENXCo+WIv8rLPt1fvCTNPBKdDAQ+ZP7V4xR/1iEKuc6lVJkwzoInUU5eWAF1fdh
scAY+LWEpvwUKjz6fsb7rlDA9NGyxm8LOZ5/DlcLxh34DYv7zkrhnN6LxM04jKJr/Uvkl+9MZ5rh
mw9olx9vP0ZVbzriqcB+gtdJwIz0kKzDagNrNte/mNqlgQo+TbHeE5ZgbOZZz5xBMdKJrZ5ioOtb
lnDtFa5GfdaFK8lG3lUb0fcn6KsaVPN9989Ik7a2m4Yctn6nOtyHntPqskY2SV7nwBF/gh99wAJf
RClyVMcq+GmoD9j+WtNymgzg9xMspG15WPm27nmrP559FTdDcpTGALZzwo4Vav1BsfEDXfZl1+HA
MEokS3dyO/4/hi+JlCiS9TK0lFWkjqfrPKFLYJOr0iZZVd6aLWsEe4pqjcj2u+/kn+WjXF4e4Jid
Zpoxbq9aads6AO4VKtH/lnDw2DaYtl3+EXVrpa9mVygT92907apd6SKq+hBO4apKVk9k+G7x7hiG
ZGT0B+tX2Sn5Rt9Ql0YkCFFkyKZ0Q7YJabS4wJR2HMFkhvHrnsbTNST77+G5MaodxAsRTQKLqJwG
0fW+gv/X+dWxboJxOoT7Sy/jsnswGYDvgyHgekN0bEovXyxTGzBZPZZ31B2IBbDHmPdKrBT+22bM
VnI7Ch0SyRErBPFk5cuYJIRm4SrAjsRcOXJxZo/hC8Sfthff6kEmtr9mDJGWEDyNn0aa47hhynLc
H9IHueDzyAE98006csTQXaRqYx7E7+jJ6YujH+Q28XJ4ytNYuNz9Sk5tiigkS9e5kKMOhYwhMb7H
YT4mfKIEQIrEMetWCC+pHj2ktA+wsGhdIyCiE0L+Lo0qDG1e4Xk9RzYi4uJ8HBtLqgY+qkTJoJay
+23ijuJa85ZKfPYVFC3nV4dU6/L3ZhFnC5TFHuy7uInjzwudnwQpmq/LsAZ/uypSy1SpizSfucYA
ookd7vfSFkMkYKfrSOGM7xFtN+I4e3SOWysnNv3wL+3CN5+YnBwhOx1mf4wqe/1o5GlBuo7hWyFD
EE4JSReL0Z6MzckNxb59acoD8qre+KzRuISdX52V5Y76mbmmUEUVBy3bFP97Aeyhbwm4bNH7E5ry
HBpOq2M4do8d566t9sMWqP+YTbclmjEGEioduqAIVReVbfAbgjLp4UHHeRy/PQPk9AnxudAdAaKz
bA+yyV4TFotj9fUWwzELWXDIZmEIvlqw1IeUA5CyAownhbUA81bS1eewbT4e1KEF43hdbhw6Z5gz
BmYz7GvF6xMiaviRnP4lvBT4tcvf+vULXdV2o6UFa7SmvNa/qZnqGEBmWNRc0OZdLBUuP+JnOUa5
G0PxzCqtCK5hR6bTT2Lrwigk+mYXQiT7TRsqvBhq1g9XKHbjEWdvO4CrjJszxdRhE/ghG8NmVQZq
zi96lI7ajuRNu8FYp09MJqLVmiYmmOg7ABov5jd5G/vlNy6T10sO5/S2JDOkuLntlnKVgHwmEng3
WxI+NOB0Po2ZTfPntcqsrhpumn+EV+F6bYeWUOKz5yqT4tCVg61q8wBhUsGIG81LBlbWMT2aCtJ6
2atqAILFQpavqGPTzgbKUtukUA6UAAns6wnyN2M0GKEAE5vsEq5eF4GxvDq/S3Gc9u1fRB9bP6sr
3/5qK5U3RLHhcRIvpmE2PUusRzD6KZ2fzIYb023DnHxAWRNeZ5sFKm1LQmmfDLVX+L+xBdzhf1v9
mgIaxj6Dw/TnU4xdfpK3sc6kVp+s1cje+EGK3nApb0hWxSDQ/1yY7d9L2ArUaJbVQyoO6bjjPtai
VNxuALY90BTYZ1dfkXDRONmr99YOJbZxEElSMdM7Pjjw3LRcJ14gTLcEdAiH21uTb8TdWYYDv6CO
dClolc+NERZi/JrDuNaBOiGBdkmp+wq8U8iF0edcuKj97gtyZTJDLPYKZkGDfJEYL0BG2HrvqISn
yVw46KQDDVgk2o4py1ES99qNi1bbqhNqD6WzML4h/C4D2KS1bjpCol46poZGF/KBb5cY06R3+S3F
jzJiv2kJlftTzVkfDQpHiH9JOXfMlB92zHz1CqNqEOWneaJlHoq3Ok0rzVfNJ0Tm60wrfloqLRmp
SlrUWAVO4Kgjw08tR8wog9wN8d6QCKXx5SzoqtzbnCF2WRcrl/QpNfyETqrHaboeYuwzox8mTrwJ
tVpLh/lgKAjHPbw8eQKYJi/eV3P1AKyhOIHIhGb7iWZxLiwDBU0VHe2QslYCgTUlTYyYiIVgpnWD
1IU+RQ9ogVgy4ebHZ0ET5bPcHIJwZnKu2sJXfMrZzBZd3AJODo5V6IDblfUyP4Q+Ni9DzD7K2W3g
ZpSdDd9pxm6Uf1v529q2QNukCLFUK7JdkLS/9NbntCTvTMPjXPAlrJVyEnONR+8VhXl7/gu5CZ0n
XSKqn4G/SB2MnyTrZBSH16vXSiFDBhKHVlDB/pQq0ROTWSNdnOyVOjryPcCaTlrHGk3vo0V10Azr
DQSaHgHnJhvF9cojw0XzTu6rN0FFhAwkmVowXbcLfzMEvi/bmTcJm9rhDhBsvfljr+9fCjTbar/D
WjUq+wpJTiXi+dmIu4wywerB2e9bAOG805c1ir+03QR1wyX5iL0CQqGZK2EA1dmdk0toS7bXzd2G
KrTpRxvdxTtMNtFyRsdZ7ANMe0zBuEQcUJuESBP7599efTH9gtrUjTPWHenYY87GofOx9GWxreLt
86HOO12UD1v65xK7BaIAqtAxLL2ptuVambGzb9LRzPTfhycJiPH/nT984XN+lXs/13FLAoiLvLNN
3spZFVOoNrPSKpQBposp8RF/X3wxUM3zDkfLtzPliX1Ypu/eGpBTC7cAOQBmh813oDuI7lUNs+bH
ETv6CWb6FZOtydifEt7AXNeJZ8Q1Dv/8iW2MDhJujuUXBVn+zyf9JdHJkQSgo543mFCBTseAGUxX
77UOoEE777UQKhV6gA4C/QiO5cZgEBDBqmCF1uHxG3BTrFn4Ckz9mjLS9ER67rgUDoRML+2E5GWz
gY4O3XppvA0+enNk93eMSrztDUl0FeQ/eiWrmz47ZgAfkqUSqXfmtX6TIFOh4VGgd5v6YnukUxRq
pdiwhXVaOjS9BzJihpDSryFWZDFlR9HI9NA0HyrC/2/IPc3mmFzIv8TmeOpUQHy/G5R5mal2TIvH
hYooqZZHlB/bWW+Tq5AZ34JwfRiF4pxaWGaypGLncS3kMaHjWUSxrjm0zTkr+ojzQOvJBwqfGRh3
siJK+bbD85gBQLP++m79RqFusrWn6yraU71SsImdIhoH4yTK+Ehpb/8HTM/ZWvy/CCRw1mVa2mH6
2uL403DMKSYZz375unHezE42/2+a04p6rEQFYyZKdaKDfSNmHXcfF2QsWWxjc2v8RsPPmyqW+VSv
HvXvtTZprlppHJcIx1u25fX8oTcIQJQQ5xR8j1iYJreXj3v/B+MH7prySkdo1rgMXadK8zij4LpU
ysaLweY8qUvjoWqDy2r2Zc7cM4KNB+n/sh5XBLwbXkM5cjKqD3s+sEboZucY3KGv+a5TKXJfVW/U
NJBignLQBMS1HrOW+LToijqEpPx/cBFWLrDQInLZU+3Js/jNo7ngIF5zmRPqPAKZCpu9rC0NAz2t
gK2QEk7y6VnFwxu70AzRtBJKoqRi7N9NdpeYygWNuWEP8dts5HiBvPxrgXcmpeTsIYsHWE8VvaLk
Dd38K6xfdZ4CoFebYswrpg8XZsYynMo5R4sZSI2P+MbML5O3b+EW7rGuBsM6mJOfmDU73PIBcn36
pXhRa52sDOme9IQhFD7WDBymhtGCY2rzs4yVHAi+AGDCTKGdu4dJFZpNHD9uiO+dLWjV0HWcweH8
lTCT0XkotILiWAlQNHJCF5Ii6dMqrri7zl7t2dhgDU7myjZYRfXp6BR09ySTkIemJsiL/q1Ap37f
DrXYyWtIFWXR2Nb/z1OzCH7myUXfRAQ1FYMsQ4Ke0uHbhfSJdPlTENpb/JIO4U+O8KrwwPQZ9NVg
QPuskx845jo57G4gl1XVvol/i4b2NO4+/mGwjg3Br77sRLG/sbvo2KDNy4tA2W00zc/dFX2oLROZ
zqWN4QWC+sAhrG2D6ON7Dkap3Gm3cU6p1enfr2bkMlBXg+Vfru2aJ9uYlU6Flw6qbVmkUgDnw/kn
AjeYEn/09d3Qpu0hTOxP0dmN5n7P7F9DSkyouQybFIQTnmts8yWsHGv38PoLM13zJLz82NDUM4w3
MdDa4OI2UQ0jO+u2IAkwku4LcuYrHR+oWaiZDtVV8rcwu36tybuEDVYzILjqrjdOQtZlWfLAteWi
dBScHWbDhrvLsX5kGW4k6dGADbTQ/nZ+zMM4RKpOdnTqssFGOviT9/0RlRxbQQbK55uxYrcbzrrB
0cQAf5pIm3V43BgRAmsK2QcGe+LNhwgbLOMjvyxZ04H+vfOrLB7F11xeOp/YY7ytZF0U/y5yr6i/
5f7U7u0KqpukWkOVDzZgnanRqhtPsFvWpxmGAC8DN2+XrQWQSs+xMRmLZy+LnBN0BHIEdUXKCp60
f1/6IbIIr+h+vSlj0V6TW/DhiYN6FK6Igh35w4eljO8S80dkEumi/7bujVk+BOZcn68rDrdsCpoj
vPibouJKoNzQsdnVV4ZPhkKX8s4ZlSbdpx21Xgbdt8zHnv5kECCTgL07E3MQ5Z8JehO4sh0FCVOs
28PigP7F4va0w3s62doHF/n0TSLtBBC0F70OE6X88hL7do3cTI8KFq5QWWi4QVj+AUC7FOFqyeik
WWqDGVhUPMQGtMOK956NEi+vHWY4igAPYNvFb8A7TgntrjiOwyztBvWD4mORaImsJHRv2xBm/xO0
6YflhO8IKmyfDx0IBQuMA2u7M2y7t9DfAl159IN8TGskRFUi9n84qEk8sc8pRZEZyXNB/xod7RTn
8BqFk7fqv7tBmTvLNgGP+h8e25JjMDR1OpC/SaMycR9t+APKOSsisKIX/M02WCFFO7Pb5lHV14pn
g9q89C4XdsuiERyArGLg5qnsxFQEupwz0pskByhcLCkJAG2fzb0e1sKmXHV3I5YpMXF5ayU0xNmP
Sx32qppK2CLWA97sE1R+wswgWr2+f+GpLT/9/ROjhrqsBJ/6rf0I8rnncklhqu9GSxEKXaS4AmOT
TPHs10NpkhP26cZMWDDb4yR1Kyifb0KIZoOYxvyMUFHRO/riRTt3F+zRdn+43pn7atA0GpTmEDn1
0TTQ5jtHpHCEhDUqQTVwvVPqa+mwJFqo+yDkkDhiAJ10Pio1z3nPEMBT3IFIT2dG2+K1TrLQ1ahQ
fviaS3qfVIyMjR3gjljLjAJDCZY7HWNHl089df4aMXMQItDbapdB9pGavRlvx4emRCtjMNMcAmmM
CxoYyOGXfQ0YBoaEfjHV/KboJHuYD5nwK+KtMKrzre9IHmfednVpU2X5ACuT0av/QqEU1d0Y3imW
je4s9IO+ov2XJLzpj7BiWkiLEl9UwKkFAOHfFfd9Vx16V3K1tlT2pcKbvc5YuT3iZwrYB4stLsrc
w5TXRXvEbJ7wC74oFvYvUFywwPyuypl/Z077dO50j36xxyU2rhMHo47v6HT7YaimQuXXxTsQF/xU
SmUBqDAWDhChMqLdr8bteK8YitzN0ukCe3xm7FK+McF+Ho6ahc22rNUOlr+kGnrcA+0WDnWdXrjC
Vw0OsW3zX/GAjB/ikB7OuIwW0HL6JVsSMbsaPoUwh3tzM9tI7Ls44hQaRVVfZZRMeP3hCU7YF+1n
ALfjUtc5P6Lzc8buu0Y6hC/OG13HxhSmMMTB/SpYpZdHYsmRuNBdJSLhN5vvpG8JTbpMZWwXMe/S
l8UvGueTdGFBIbVhBpHy4EhGKU5upwt3yR5kZBTlwTBeUARd8jgbxVYNba1p1xgvuwPkQxu3bwzF
NIIbNz1WJhkdhHqLtMnBWkj4wAuX/RC/v+GFh+NKeafbSaYXUigdqzk0cFdslYE9fOtHSJ6AyMH5
27DODmxvlqXKdvzYWRJ08W6azNVKEjxXMaxN3ZgFGCDiVWEjjnNQXPKiYHzZ6Asva3CWB2lJB8FP
f0qdGrhgwMkiPyn5nnczUIsZxzUU2e7DinUElRrbkjkxMjZDOTTDDR9HT2961Ep3N1t9d2Rus/3a
sLOXxbGGQZ+ALsSHR2aqNYPp+FbHg1td6p76TRFK0/o1PZdCFFbUBLxbTzs2O3B2HTHp+cdcCZfD
sH3b5XGzHGQtQwPKJhuG2gWj0mkclNpaWx32RnhB3vcccDV2+bGFP1CZ925ihS7bLIIcPac48Zpj
431usAWCokR6PVBzCJJH6sti8Agj58Kt5hb9WsEbsVxEtMRY++G9vnyUHfkmgXhCpLlbIi4sDqD+
1vDp3zXdqUd7no86Af3ie2cvpOFfZ3iLedFpTmJBJPUg57d58o5rkyVe+MHYYstMYCrWCECSQq4z
bIcIMCKkrA9MTuj54iAfU8p4kR0tYYhBKhIITALVi9bkXbF6mBmctMn+8nHkXpnSPjAOOgvI6DZ/
1qYBq1xIxTJcAUNRURhT2n2TzQoDPxau1Y/m5lyiNJg7A9yr0dkcnYVJ8FDFk3pY8WihUrrUKDwM
fRnzZ/d4l5LoSOURmnxRR4oOTHsamAa53BcLbpS9wXfZvuruKc/kvKqaGEF/hZ2bcw+vEnIOhGbm
djZ6rWFauAI40sAyUP3ZHR2JKrHNfuNuQL6YM4vNJOPl9cU6bKipGmfNAzmIjLIPXCVmj7TxgdXf
NdyuN4HfFSlMo7Mfm/B/3gArhYWztatnB+y4nmOfE+O1dSHEirf4c8dPW3lKvIXafv3loQPlvIOq
0RST8b0TBkr4DRuEZxSswsUSDxtC+uVMgNrqMjcMbCt98IAeTOzHN4M5PU6W24ILNunSDDZcDHCR
TJFas+5+Uhx8BxRh2iwprVwG/l8mXfpY5R1CyqA4T+8r14METEA8G+U+s3WRiBD+YjYd8Q14p/2k
o++5dKIJIffMowtugFjsscaTgFiitVw4XGLsxv4Hvareld0B5BvHOG+KD1Pw9nFN4qVidrwQKtot
Ys3J6GJ/bNBW6NyPu13IMkzXK+oBv1PCfW4OakRLX/uwO/APJYwIp2BKT3zUT9RePB+JPlvCGSaq
AStUVQeppdZUIH9Ak518nO8hhwbFWJKyr6aADGM7AK7eYcEEh8yBkSavjYpAFgI4E9KCbfFIMvfN
WGXpWjaWg7ybinkNVhAxOM/8+VRfhERrgJx5S2vhs/BmDMQYfBBYBvV+1tqe+0xJc98xOoMyO35s
S8JD6IysC4KhCgaIeHf2j6yAiv9nylriTpAjkz2KvBcn7s5gITR9tXTujk6EZlmf5+HOtxMfNEBY
2o1g+LC7Bn0LzDk0fDZYBxe05xDnignFxoMq+F+7eoFk24tzLB2+oL+LkBNaTLwl7LvJPvGpNTh6
2cDS5WNoRJzU0o7iDjnTahPl9T5+P7p1sjrAiG0anvKhd22/8SyMKNBFmdAAF/8QBUWIoGeuY09W
xVY9NIi3d7QLcBPlPSI5mFIGhxaPhCk3m7vXv8gtkhg6UkG7h5hETV6w4/CzN0ilIDZNm/FpHxLP
HYPIO8iYB5CBsywxvhXU0rUeQ9+EdcyM0pDPP4GPTF1yCq9C+orbFmlmAXR7bSVz+YBwwV3m0U4t
0hJXi84/y/PZ0AEHvZ46zQozeFkM8adxO02R2OKWz9nEDzF/LO4PSE2Id8e/GFIFdViV9EVmWMXX
ge6vpouFLeaLohRsydwLvnxMVnKKaqBwjZeHVNrG+EYoffkF0G4KW7iFMpDW96oZPxQqwgGxIigg
HSmH32uA7Ycq+p4CDbCibgEkUkQNCgW5XZtVV92jrzgrK8OM4W5XDH9y33lBoQtG5vOe7gSU6joj
3dNXpK1Uj92YVb7pPLzVGWHpiF5AQnjcLZfkNj2oZwcN0J4IifRNmHXNtljaWFbp2fWJLlVO6FII
cAltuHSwyPag22om06QjUbqTaAl8XDmH/hE8q4xYlrOLj045H/54dbOWbXBqHgXgmO/DJ4qCb+Ao
vbeRzMuhIv4MFfHaqRd0FOyrc3Lv0wXuUiVSWHizGdtu3CpjNGj09caT24cQ5FEjdJgctfMGtxSU
rrUuGdSIgPgFMMfe75fpIB7B+Qo+Yx7vHOhu8BP/aje2WZ2+kwuRCn+TzgXGmJ3y4rGFu0+6EED0
WHWoJ5NaIl7nAEYohjtQfzW1+wuevlgydtZg/aYCyYI8lHUB2Zjwn5NUN+uU74YniLiLy/JT/P7e
x5UsxmeINGm0/xogZGS1Rj2/77mmc5vuJbykOCbzFNu6jQ+aCCG/RyPQMEadP5pnVDNSDzm8rpN6
XksLwhxxiEd2taq3vRdQ1OMC3Sqd8vWdOqCRDTM5bTXJc8xp2z1WBiUa1A2dvC6csfGDpJD0dL/V
EZOC2w81P4C5arsQgWop5I3G9bicWYWdCH6NIlnMgoH5e3zy6e6pmfOF+sHCaf0/rVk26LEuU9FB
dnc2B1+PVkotYvzH5yck0ZumCiuwWY3QNi8rf8UCQb1gHcyjaheRAfs84tst42/Swk1/G8hp2FEX
IwOLBY83jaKvyvK1a0939J2WCMUB8B0bL35TCX6mc5FAgXomFs/N6PbvXo74CyOVXmvQC0Wej2X5
qq78GA8IavwVdvX7ToN5893WyKnIWepEqtzpDsXePv7hi6r8nQ6BcLa73wRLc8dMCUuFl/AtRIL4
otTzHJKXo1vHGJtr+qU19Zs2bkNKDJLm//wS2Vdvsn6M7m+ZnrKPCEYjAPIi8dwQEHLj4EIJ4IDz
E+/oPbU/JOKLkj4D3wcTCXhiEuG091nCJDkouRtR4kPqLS+iaLEqvKyRQu1xXi+Qw4i7HK8A/9Yv
hEewBEGDZBu/QiaCHeOvURXURF888qQTBg7Z7LBcRFkZ+u++n6DmGG0/qMkLdo4LjUIE1/ksI9qR
UihX4hS1vIkOqV8uN7Y3c1ZRhsWrZj2S5PKFS3oPl72Zelb5qWUP17mwQyld7jrjKwKu6bhtQ7p0
n4CM3Q2bkvGxvnnXJ+raTT1WcmA/3YLWhU+xto6SvHukrKwxSP2cwLQLLl7sSrQw5EdQFumrn+jG
pYL4oBivECRxUTTa39wOyFd7CL0za8k/uQv0BLasSnOBLB4l3Xs+5mWlRRi7r/zm8F9kpIk1QVxw
C9Tp8YoMhhVVIz4uMt8N83WMxvFdatCLtmbXKjYMUfsWg2unY6qBaBGoOF9DIYpQNB71ZnDHlSjv
1h5SyHSPjTBkRQmP8xR15bH3rOaozL7mW3h3ArfyXbxw4pzmcOvLUyc8DZ5tGwZGcLlu5oPs77o5
HMWCfqaZE+zgvcYi9smEEuO3LZIBEWvVCw6o5LnL2jkGD73ezBmCulesSrnXNsFVzxYZwJs4cuRx
5PVK9LwonEbtI/0+0NxWXoEbbZK/XOhDoX0rnw+U9wp4QGOtCrd19XHWvTPvqjeSRkyHZul3Nk92
8gL2XA8ih2SqbrtRkQspnTnE8DawHAZ7qp2by9Cz3tIADxMjLhhB0B7URDwJU/XYVe8WJ9lNNNlP
0uZ2zWGQvqDb+vl+TyxQMGp+t+2hoNZDCEHGHaaZ8NZkJxryBhWM+3OGZ/k2ebngPeDM2086RZwr
kdt/lwWBYz8nfb4Z6MQ7a4MgLD9jzZzvi0QUI00wA89/tpofuX0CKn+5543DA9bphYuN8Xlkb7If
xLGl5qnqWKPuqTvWn5CP0ZOOvJxTxHNNx984LP84CpTuMIr61D8QRBnIAR3mAbgQbi2Q3PY16aK6
5XMMXZ4w7bzydIsfNgAnch6zgIEzgGmwlBmXid7AxrbaSoWYZAckRqR9ujXF/rp5c9XhWk8dzf7J
u/yvhnrs1wdFGyCFTAUXGGbIrUJSKo+8Y36HOykW27L8i4QxQDd6XTOPk0V/oXMn+mO5dsFGMUQk
ApPCuTjQkSc1/AcRecPg3KaJwWK2eMu/Fe2lPsWX8uHCsSu91AdVF/EshmcZHcbbAC85fK6YLIC6
0ukxUPA2aTNE7FudPnrKjqCubts0tMgrm2KlDbJwfw7dr231dGRFvYo6MDBxm6PGkmfosatqi3J3
KCSR4hbkViK+7gZwKTEPKCxn9zA0fSBUgFuM1Nk4fCUQYZ4qVkgIUVOzu7abBoJ7ehppud8VjYZ6
OCl5nnlKLD21j9WRspUtdp+tnf9S41rcJ8i/DZ8syQdlYENH/al+r577Cm0wdCDYKKP2ug0I5Fp1
vUDvdpQx2SCZMYIkOJDzAwKpycsHBlWOv3cKb33GSs6pPbpmKiHOp6E85EwBzuDqsfNOX0VLxVeg
sGfpMWYxG5CcRXM5nUVrLV2I1rPzepq+IOTpAZEKiA8FSBYkk93rIEwQC1zWLGkEnuV25Hkdu8gR
9Y+Y9tYmbt6O/A/qDy35TBrOnECECKpYKz5noMdTGLO5uZMMRIpfcMY+ZSAiPl/UGT7J9PDo7YRT
O+WsgbnURBwamtUlIKHBYD3LIMoD51Few2RdS+qlJGQ/kykkuuLNJ5SqXEcvLHL94PGxeNEE+Avc
8sEOesPIQWeoEGXk6UUY4/3q2E889bH5t7ODWPFwHZwed2y6uaZ7iNA8ICvXvQ8A6w/nRemRDACf
SJzx0jkw/zLxoecWFOipwTbMzKZS7KSm8BKwtxvN91pYbpPOJFdigWRHYQq3QS9b9N/pe1+IIHa5
FIWCmY1k93ss91UeYJdyb8He7nEjAABf7mIhkig0tTLkiHOfScVlHfV360izNQFKhuWcM5JPb7J0
I/KBcVIkckVGv4XAv8wWPqRvLnyNnQKDnKJde1bmg0Oxm2m4rKpTlpPB7QJ5r4ohZTjShA02jdcC
R4/sbF1lZSJO7DdIgjKiFTRJWsF3z1pfAy6V/h5825oboDBkIYathbap2xSdv71gDqYRFmkWzW+H
A44bU5DGYVUW4zlifLET96H+ZL6Tc565ySfeuaJFGnAm3BxcOmjOpstMZ0X4KIeHQQnmCxLeRZx3
uBpOQ4Ii+KrJ9NuQ7oqYsStnoxLAZF5aHhJH9jGK3jaRsEkYgvdAsCgaw+fB6IGh0sN5tWpADjC8
TQWVkf2WLl7f9sjB4IQ/kwmP9ti1KR3mKobKktGmUsXeuvuBa5wa46B4hD7nvHO/kmI3M43KMnU8
p/hV6JA8vamryaKRnWUdDbwCHOjdT9JdwDwc2dB1BGliwRhgnziGAPR6YDuNZtN+LctELn0BHOam
+WmlX/LRweLoJ/z2QoeGHdPwhTjnIMArzSRdQDMoI9w/fPbUQ/ysVjU3Qvg2YslPMKFmkHB0keCt
G09hfj2EeScZSgc7xueoBSwlUueOC6XMrMWx9NeohGObeVHdXtu6cCMN2pk6egwZyvOYVCNbmB1q
a1BkQY5Of2qcM2nytt/wefJN9MPwsekSqqsOP7xCpajPQJKGTaqTET9lcREb9sW8fcBRwBQy3iu+
y/yjjCHT7kwfCruvFzk2YUjPJlGiBM0Nk5kmrMrKtutFH6DD07P6Uu9BoDg2rPCt/RcNlpBRE9do
L0UNnXIckB9lHLqvhgzE46PA7y//r/X+0qHD0R1F1+LnijTOq2433/w4TALIC9TRqUpy8NjIa65E
ZHy/EEETXHkCHiUx10lWNAnKoIpBBw5G7OolxJDmJqg59s8jreHoN9SYrm9zVSsHXuaReLU6n6E7
CPp57V+APGdJfEe6qujV+yJTyXOLI7pncRgY/dWnWdRKojFv4BJMgrmYl95DENYmemCd+q3dLxST
epXDkIVALU7gt0HBrTdf7Yx2K3FJzrLiQOD2irmX8KZey+WorQBgGcgeuUbzVLX/A2UdaslSIaiJ
f0B1dKJ56dRvF2XzjsitXeoWOFwd3s7xfvCtEtqytEekhHr2a/f4cDyJHnJ6wz/bvbRJ8tuJV8Cl
zBKP0n+loug8cuAXrN5LqSlGpH47ixCUyXL1twyRe5ZMLU0dCOFkZFAou1z6Ugsd2uGwSsHRM8hZ
hgopZHYJKAlJectQ3k7JnoTJDVQ79s1jtZ+MoIPdghNsgFLJl0hFTeuzC3a3+xsXiukhktJCeX5u
5Um9BMtLJcYpxqxYhs2W4VTJZM1tDtR8o3Pro//rFTJCY+Mb3drZRr0jOGramc6AemCL4zjnCnIX
RcCPDnkx9RSdQclmupN/9QorgXQx9hkOsTJyr/D9V/eNx9KHfNAZqa1bjjWXUWgRkbp6sZu2yRxo
n6MvmORZxCP6nrdjaa168LFoScjdYFpCW/uGGfYfDK+ZwCiAqVT4HDgvNu/bhewr6kpOl2K+MKG9
R+wE0B4IvNqiR4h1IpvhBS1sqUZVvS2GXPkvp7CxCxKY0LHVWPaOmE+IZ4ObrsK8s+UCzk6/NhAk
xzlviHxUMPB9Og0TuDyHX0xTLcG7B1g8KFqbN8zuWIXsbPwTJyuazxZ/cBY7zUsbeFPeY2bDYbk6
ELP+StsniSsN0J6GguNkUuUFhV6m+g1jFeoI88ZuYFdTHjqKZ4hw7OWsAybzqogP7TM+0OtW8YSk
kDaEGwBp2yum6ExrqBnMlVQvQAFxmHejIstq97cT2zPeI25AjBuUuAKmFnyKDy/jJn5mf2itgyuz
NnuB6ne0oiJ7KVef0GGn2IA6zneOGYvzlJoVQyQpcip+2SKo2GDcHd48SvmlI6ZZSwK3EQJ4TxUl
+hIMtGOnsE+sC/9lCA2ddhHv5QrwxpeyD/tyf+DjlAE2PIIlI88rgS7PleRT4CQgQX2tor+obSvx
gQSduL6sa6CgTIX+joMlAGnePK0vX3onaBdbbZ/mgu8dkiOKQvQhnz9I9t5TKLCdruFxINnChgBR
r0E44ASaaarbEj9S4wjg5oChSnrXx9huH8J/I3nDDg8dMD7CWqcJA2UK6cQ/q0MGzkYYmCRxsNVs
eJFoQ8gtk5PhD0Cb9nM/XVUTOiCCpF8PsfGY0WQk0M8fBDELvg0ziOEo8WtAdi7ZuQj+41q3xQ43
+adqt0LOCOpGkNq4gZNpfT9gALlPL62toSzDDdoF1BRXQ8YvC9zWOgOQ5JhCzFzrWVwLQH+ic4SA
6u2tu/cb/etHEPaHIqcS54o4EelvADKbZyw0etIedTJ4gkqHz5u2fWrYQHmfGvhWXzSw/Bj657CB
8yDO3QYcpOEAwRbtcJyA0txrCELsrY4UKFcyQikKoniVazjP7EcgoaIgsUJfoXEPmJnnNSeOYhVT
IyL02JrBO9IcEZA5JTbv9yxm89+AMEfuMR3oham7gZIR8zxTlhz7Tb4mmmxMF2TmqBTyHVMSO1P3
QE/oYAEPlPd88gEwROSmuNn6TP+jKIZ9by5v2TAOhHjyQgJk45V/NdX99GKvtVZyS/NmonHP12Yd
qBmphX1205f6zsOLyMl644uqiHNsmd9F5Ov4szZDQx4tm5V6d7PDRdxxUEsBO7HD0nPuqcO6ydLq
ONWew8P+WR3eUDCqSd0EZJ7kFMxSLrpYtdurEvdaE/YsoHUqhLh4ZZj2BIW5+8o/pdXNp/4ilR/q
kHWrHSeNAKipAVKG46+NjaBv51uJxjfzx15/+zuKXmTwIwt1mGOKBc6atHxD0lEjrNyAp/L+QV/+
SmcKPdgxfmWX++qAGFxA8NrLqLNnMcw8Olu8+sO6hjdOgeB0HMh9NqzI+u2ELtIVUOG+4x0C67s1
vRo9kZNQ9JuBVCi6DbRg38J+Ev8BE04xW+g7ERscUQWlCTXQKhsddfCe5k2fvZpb2ctcoI/pdS5H
of8La5frt5Icuf9x8IplbGmaWOqIpmb4oKmS92ykRWavowN7GHmp8l5ejO/9TtqVhZBqaR+XRzoV
LCcRHRX6Q3UARyh1gNyDgC+RYMhtlhU5Q9n/X8JvNLRULNNOhEluSVG1KZyh0upRT6NVLDFjANwF
1zbYfgCHb77kq8t+p98HSB24j+1qgHONEmjZIgbZ1jtUOgQVvada+o2dJW9NQaU754+HRWHvNcm3
DNy6SDKjCLCO+Gq2g9XEHImlcvtzw8ny5CLATthSbcbn5qu3sOucMQHg3/gf0jowOak1goCbjy4N
HA6Lt8SWpbUMxjQSsmHPcFfzq74yQlsyqmKWIS5eBhLde8x5I/KyZfwTLBUDH4B5gWiypI+t2854
BGlg4BCirSXaVbsVv53PXmLW9dM+5vcjNOy137p0BxGi26PFjh3aoSiJmJOEyEt38lZFVmQr/gDS
3TxR6+UfMN1Vg7qQDf+JVKNzSRUmxew2CsB6FrTtzljNaZwugYW5ec1epPM+Ex2g1YyqXDmWxfLp
4V4RK371TVx+sG5y0MH+EryCSZVGJyhHACACj2pFpZCTcrBq1TTQNivpMm3p10uz/fNHEOulCmeB
sGJO6mO5bGHoPRzPAvgZ0akZXwQ1HmkHCNBCs+jaaincLCxP59tT/bRmcrUPHf6ZHYHsTcpn/XI4
L8GLTQAtn12UEW1BG3owPMoIE6CpKyVYDWkJTB7qxspW2dod5l1B9uIx69J6lQJtr17GtOyfilMO
39XrTJQQetAGMihrTsU2RlmBIx4DFjFE22GG/4VoAIg82gZo+tSkcGGmhhyRFLK7K7q7TujuX/h7
WNs0pDtSeLl9ugDOC+s0MTNGtkQI0S7gBPMmkLnFaV2QkLwvLZaCXd9dN5Oj28K0hIBESCsM4vlx
z1JINTsZaEJtz8nll/eCW5bJ7gelntlcmCT1OaBNrKJwcl9mL3X8P9zQQ90X4C7MDCJDQzRAiTrY
75WBqT8EMWFAZBgNf3FobTXv7Vwz82Sp08lKoqKquCbng3Gu5E0x97lN3iWuu6bchxATg/yxJWrK
DLp6M/vrs/XqL0C1fdi/nEk7TwDxZnhu0fGPj2N8aPX2KtIf9U6uhM0ZETMk3yrsoL+dCwlkQ+dn
7bSTpYhH5++FcbU0KoLdZtotPN9gmoXZTceLQgX1jBZihdDUVSuedvzW4sb7X4a6IGHQfVSTIDCJ
4Z32I15udjlEeFHAkEZnEKCAfiHrbozQ3qo1QY9856YXn1gDk9iUjbgXDmkhFXuFSZ/3PmA3Z4hp
OiSLMbpWvJg69XHzB4OVLZnC5KeEh+ZAWefPUQKG/VqPhoVX/PZrAiMAgq+CQpxub3jYQrxch9zJ
Luaqkv6QxvpRvVM1YD5hK6Ca8zvxX0UzqxJqoxtiOjM5zotWOzOvVjU/iJiVJeCqVt4PaB8SQR21
inYidDjj4KJxbgePuTi3bFvZ46Scz8IYCe4uhyNHBoqg8AzQlhXOuCjauCfbpqi2dZGEejdjWhMY
rDxFzMfXYXaCUUxwLWlNaIN4W5m2IGuIwojP+70FS3xzDdDDkaWELQtpFeCG0R1tmag68WR4NLpR
kQfzjd0mbYdXM7YlKtXLIEX9opuWGCbU0QBVqlGIafzKjJq0c4JPMCwVEaZDqoi9U7x0NSWjFuTp
wBQvOJtBAPIm9wjGJ1wh7QyMyP6k9bg0AFonyJMyyjWuIOHKtOp+CCsEU3Mz7I6QiJmsgmrWOrY7
aNh4UJ+1jku9+XYb6IaI0GYwfnoWu6UquOD8ImEVG4SYHUlD2PcHuFU7i3K42VCv1ndE4EL7g7Je
yWnqz9X6R0Tw0QpG4CNL4ThdKUZFbhM++KR27e+jn4h5dV9PjH3fmlAFXC7E9pOTu7Gbrg+wZG3c
8dqJi9hjxCh3HNBJoAStCAZ8eorG1hcOJw5P4uQfVwePx+ZyGQ7CqLluu5a3uPmZWoFLqZXxLIXi
qn6CqjQIiEppcMVSdjmVIjJeEWeup5PcHUWCd2AX2h0js30u0Lwl1hHRt0CX9Z16kIbUcupzsJ63
fHKRgXwlQeYywbS4rcY2TpBgrdeNUoCQATgcwhz+ad3uucD+7C9YsHw0zck3SBL+Rcfcf5jXpTZS
T4Vb7i0PyN0S4TA/a6Og6MkPVvPc53Froq+zg6IyrdO3qLO63/4y0vP3xTMk6ICYiX1it2mHBJY2
Ex475t7PYGU2MYxeB8QNMSBTLkZHMHCl477PO4GAFX7mBdNkcSxw8oKQsMOIRY2H+0cYXCon5tXZ
fLHRcB54H85y8UHqJcWXQRt9ZsMPQciMou5snHHEYkiF8gTOTpy/68zWkVyg8GX1yg3tBYnWXO7w
lK6jfmSHYhNSjv7wmdFpcM7cRZZ5piPKc1PTvmopwUDxWVPaI+Lur1vF7Yyifd4G9XpGx3TQbfVK
/4ZC0li/ZYOo/2GyAU040KZSUu0JFcP+IGKfLj/ATmIWQQ5krIpApyxnpOaphhWEZCm2i4RLBz3l
jeIq8IwEJHgEprPKkRSTVD8vwb6fatE6Jq/L5VpYnptZXpi1pLCh2Rtzkj00i2CPURVjwztZejiJ
PK8YsfJkvtJfYa3GEoTL4B9S1S4UeM+oJYQzKhJlPqgltXSR+QEBH0xrcUok8lIEx6p4k8g7jb/4
+H6TBqAPJI8OaQmCneUJ4RMsM1OTgkHYJGBT6PrpJg8C629ehJpLSsr606PlrfisEEkgNQmkALGS
9NvoQDyP5lwDU34pVmhJUofg8l5Y3BnoHF8LManE1UqFz5z+RVQUo17Ht8svvItNQ5euyr6UL2c5
aZ33HpNwtTa3ZFRvBTnbiZuEs3EDFBHs64RRCMP6na9mmT8MG0b+ILPMnFDC4AshFHao2y6TfymC
mApZ44P2nKqPVpnVOnl6w4y9OxyT3BwRQWfmfNS9as9AtYROqzvQtssWROKDuwJO/sJ8a2eAS3le
9THbVasLye/IHESxEMb26wtiMqwqWPuqD/Ag9iWMxXUWCgFyZ9qI3866WWgqH994920vNvfbJblF
JvUi8Mo4eFpjQf2+G/tFWkik1G8DIEvo/UdBqZkI1h5eoeJHHY8cDCKMGB2HQIBCudCRUXSc6zJq
Y3i3R+8KC99tiHaA2mC0aIXvMbTg0EV6xWWauoKkUs3N0yWqLA5WyNasqkGhRk2xeaooP7jOa8Me
7MzcML3x/B8Eu/vqHk+kbqKmVou2gerK+moUFRNHdBaWpIYNWgDoAxDgHOjLgUsCSrnyxrGCsDff
wPrJxy5Zc4wpeoc+NGGQJbecdRFR/9VIVc8j5TWRTecgD9NB9TFYMXQCspAOBvTLoCQQ9QWGaxL0
+fhBkSzask9HIGzr0cTNCc0P4G4gx2N/y40/tCwB+3S+mZK0sEa6XFeLdkch3tsBKBMDmmsvxb4X
bVux8KUTE3BGr6fF/dkuNlimyKW4sghl41c0R78PxvyAdsLz3BEDxSak/i1ByYHkjIXFvsy13vGZ
3Yv+YdYW9U+P7eROJRe6aMPr+RNqHYPObckPUmoQg3RjnTPjO0lDV0bxe/yxyAR5Ho72qw04fWcV
On/WDWJ2Xc6cCkRiuwW9xpR7JEjB5E1OKsFwdgSy5AVSpv1RTnpf8TdWqmvoygRNRos/ippXb0j8
IpLAUzrq7hvBpub+Lf32nTmeq3roZN8L7nftyKV5O1eD1S2BJKkw/sEI6xK3ilsNGTLKFRkvdJkT
BmX+JOawDCRYNH6Nhcj6XZF9aFTbKHObwclTFB00lna8nZHbMh/pPob/Um5cG2VrXLAzm+ALjmH+
hy+jAwy1yKJuXndf+a+EE9EkACSVrjUX4IOgWcPs30Hlw9PrcWVF80yMTz/UraYyNAv6rY+Mf7RF
kAjrIJ26PntfXE2FDZkTvTbMpMVWEN5pteLVk568EYE8CGJ2t27z3JDX9jTxeM09hV0E3LgvORwR
w4EfnGdiTxYiOQAcQ9fw+TqiCLGgjLO+AiYz3SNGxnAIognTKF8ihnDnQZmxCtQawlAER9SQmV56
s5AJ5iINHY444PBcd7mUDH4HUqoMvI4dvEZcdljuFcwgyuV9Mx+8tOV+So4UIynn5/4DMe4zi4rq
nxpB/tBwg2BtQQTIxCR5e3x1rRbdWvZZAkhVxOMggoL/rNeyNcDhee2+rvOkWyFQyTXnUcY+WKt4
9a3ERIqKzW8aE/p4rJmgWyuf8REbJpO3i5gPmdRugMXxNqwr3ug6nW1+D0A8NUFd0c2cOydfHo9/
KlS+p1LBAGCPcyGd7MVey3Q5M43oRyBqPV9hFQCs6bTEJgmgy/SH7sa1lS7dkojhqD5hfwlvn2aJ
aLqt6n6BoZAuOhuovqA+D1MA1+HtIMlSh/B5/96xIF0oTYvLrUhDk2QleNCDGrksRdOhgbIyBp6b
I0RAboVUOBX4cmOq/9Tw/7/EeDbMYy8Wz2YJJ8YdXR0kBS+SfLuSLmhJND8FrWrTWppf1Jhhvkc/
7kCWM99Dtv6a4YvOyjxxWRKUm56i0SHYiuCadvh0hHuEW8uNubjNuB/2VG4W+QRYF31ai+CktcEr
sLawo8cXgS59eyp3BnOditWiMjt8fose284mUJPCa+0aNV5taKQLn+0Wm1zefZ/1gEm+mxMXYPCm
8+u4VyAV+BkxLmX4bLoqTyu27as3SwJpmwZ/JRQeGhqh+33qrjUjzgaTn/AMcRyOE0nMXRd/Csl5
6daerdtFbqA9MNz2M1Si09Q2uibnyyzKQDRmFprTs2ESYqyes4GDTBIov/kqhYZOO+lQ79c9+foV
TMLXh7Dnwpl071EVWwpa6nHL6SDdGXpEvc7Bvb6lNsj0HELG9MgnQ5ybKhE6XbTO/r9LNh5onobx
O+q5hM11zS+xbbPEMdWynfXUp4tbJ8qG3jeU3cscWPXvSHTPTZ+dKjOXNPpsgloosphen2QyoUuc
IYd7B60LYiDaBFtxEXdXVpZFliUCUFi311hRVObV0NnlmMDMghOltEpgTmj9JSRdK31QaPVg8COF
4Rgx3UJ1QrIGTpXSdLWR0Dt4j0frOxC594ibAflnWUEmmGfSE9lkHgHJ+Ueob06pISqQIjgng85e
RLP9bCeiem3wvmaldiizNQxYfz9tbCuqf3oYGj5zlSOeDmp2pLwoTaNfKQXR7s2TQF2+sev5ADoi
ucpN2anNiufTzf0ul4V0I3QsY5lR/2im9C77064YAw9BWoOaUrwNWugRXL+OrMgfjCHZ0YVkpryH
3VNW5k6XzWBf1H0ZmLiWM6jOoW0Sc8Jxsixdes2xpcspwuFWTIZ2YsnP88A382sPx/h4W2VSGsQ0
t67vLel7aTigXbffkG8rA9klbzZ2x1kcM78Wbkd7O9WVjyUjwv+byGRJYN9n5i0//I+3625D2wiu
wd7vc8B49KpSbId4ZctRe8Cps+ulrXvLGbJpRZGBq8QGdkV9b+/2b1V/qHjRc/4DD66l9hLjIlhP
rkOCtvvWXVd2hrVwR0FWaTaqdFt0BuQQVYLKPzagMLOB/jjppAAl1JZ01zuNaqCGjr/bT7rJQ1ix
WWOndyuUceYYM33gn2FSXymN1ToX1C6XT4R5rXCP70rdJwWDO3SEtke2U6IpR+Vsu0n8zrrXfPBf
DDrjyITpLsd7mJus8nZJlsZh1UORp/8vAp5x1AABmziGpmONAE7VpnCQEohLuWmgkAB4rhGXqcfK
5ozi8NkysTF2EtxA/DVROOq3ra6W6DP5VJMi5Jmzl6vPzJsBLyDdAuspVloOH01QLxvwpNJoYaIa
pHUBlyWxVUY4uGZ98B+4aCCiR7pwE3cXfq3OvTmYEaKJ74oHq9+SY2MVr59d/osQkxLQgdk8Gdta
luD7s09Zgcioe3/LxlHd4wMjjrF2Ea+01P5m3mhgch9yXh4/OMOVUG+8KEwWo5Eu/+qgaMSmS9Tc
3o7/yqyscyC/PSjCWkoP2Cw567Htq0R+zQzr2RAWsHSSUiGXmfxPPsG4zEzHEkslFy7MmSe+crbs
on1NeSoNwK+7qN1ZpK4+1Z2sr/22Vcyhx3EidPGd5qkZAPE3OzsSVPnkEc20tYhAAa7EWPgUi67h
FA7CMSTGZJt+61DlEf0DgUb3SMTpdiZ8O7y3fuxNbwRlwPzQRKHsLoeGxOCQp8B2WUPrE5X66qzi
lP/27BvXsXdBfCjkIUTPNNFOY7cuDyM7p2gkvzQGUh6n/UeiZpmlATSyCfwJPnZJDc205IFRnMWr
Nofc7zvTVfVzhg5wawFoczbO58dAjqrcjAGhaDUdOb5kAe+h9mZI+fB9iCJWQqvI8TcSuXEmdO7J
fB+ux/Y8PpmDpJP+CfHY1huoQ/gPENETE7wXHJ2dKrmNjjHbIOdWtYYC5WLlF/QyevERRZ8IfiD3
8hgwNubSo04iXwAHR3ksJmL7JeCfhk+MmQgeAZa/otFVOrsWMm1QKNXK0ruMAMRG7SLjnBZ3lUuj
n9kO06kGNgzZL7XgpoYTMjUi9eJ/bZ0LVxltzG3XvR+KQMlyK+jA4hHbIpQ41s0ow9bBLBz5HgpI
eNK5bI8RYXdGpMqupRPmfJbZJ42UueWYNUOkGaNz/F/x05fQjY1/Jvcc8Bvt1GAPiQpXgf0ZIia/
OSVLV8czzo5XTvpn1Vvl/armFrhvKwg768+LQT54H8tqaoaxe2P6cuA1f0+PLdlSXg+djWMFdnoT
4zrlai5Ov8Pk1w80K/Wa/tGpg42ifnKdWloFJsmshLe+FytQhI+OXlRRdqzhu5KJJGzVH0555vu2
oifSCiqtychgRUO5+4h6YLkfOeAx0aOcCS6iQiktmQGb8AjZVHWbfitD/Vv1Gjl0kmdVbKfGjY19
mWrcKKSfFVvSTuA7ORSQGW4qU1Ge0vUO0YrgV+Q/hu7dGb0pRoXW/sxdpV/Q89wRzMJtdBJAtpmk
8ULMbWI82+RQvhqgNHvSzqOfoVMqkE4ZY1n+EIkCRSoFvqLyDGLBioyKNy8yfcV1zq87emi3iyL6
MkVUNCghLaIFUk/89U1G0eonREbYrHxQYxDr2Gnrcfm+3BAy5xat8YSZu28AONC1crDc3Qk0rexy
vO/73O0SXsH6rpgY/DNi2QOxCLBNxxz+ItXUXAJFrt1BnsOLlEhZEid03VRl4J8P484IIUSeTodi
KF5yrsOkEtXG86jreRtPIAb7tapHh49D6BATPfyp0EZrSWURYVM1gMCtr8SC/AM35rTRB+wKEnXe
L7fjw1V/j43prsxgCHIss4RmwS/3uGCkbUYzF+uQzaDjVlvXx/TrSP2BgiNGO0yMBGl3WWtzzUgO
QShe/p9CFGgncI32ea/qGHQkSotEnGyn389I+6dDaFg6DZYUYd4lIQgt6L5K13wLbrhK0Nfptjh8
cHcp8VfsFvBkg8yDpI8OnbkCl6ZHdR86nHVtZPbQoGfYQvIQWzR3vsjW9pDQpalBg2z8NhN2r38m
BiNHPDzefZmVkuwzWgSXC9bwOtWxTYLcChQzfeKq4Wr/gVnfszeq0YHLx4lOaoeZxksFmBCkwLmh
CMU+VbbAG3XQszBqZhk/4JegH4c0B14rJeys/DrT94e6KIMatYQPsiG4UlUeeiLSqY17iGg0uWoF
k37ozzNkQ4O2cAjibw3gEOEgw0mHDFYdu8nWMWIKXT0SXnciy/gTYXCT1jP8E+tInxok+crgWhpB
bN+jl7TV6CndUdtn7WcM17PYU5KMtmT5z6L3QKISPgirQiwritGR4OR0KLnKQda1c1RVl4hfcsDv
kNr8dLhBzO/1+Jc4oCHVY0u8hUlgTuBRQr21m1vq/WIv1Z51Fy+FYuJ1cY1ANcoWZ9UDEohj9fhC
+6xmUvE6pWEd24BsoQRCpBqdJhP0aaCdp6+uKKzkx/ppeLMjAUZQngMA2yHbSSt0OrlXijBApbzw
CdBWueMvgVPhpBJ5g79vmtmK/D6zeK77a54T7NNLRMbnDVNCqkIlwXvPDkt3JADqpEBIOHNxg9qI
rdvbmrVaLBiWXBNlREdWR1OnXXwoWIlU1MoqAcxy9cXyV5UR45NnutACMmSky+UdrF7MTKkWqlfS
UqEJQnWzP+L2UyQSAwjoHqrJIjSNS00Z4vQfDZ3ucZMWJs/cy/ncckkYSpP6KQdHmcpQ1d6oQ0Yo
+T2emHnI8Gn1+zF9BENZG1x7FVopwxoB7eoQe7ntj0nNpJBWy4ROUJgpNJW5LTG/cynaUNetGGge
RgnKZmb0V8T048s5tDw0boJ7sGuRaJpxdkDLC2rOmTvp2EXbCNauoBKfxKrVLglMlErUHm3/5DnK
XhISbZdjhxaD7Y4byLsErTE3syFL4bx3ReXoIGMSy6l2H5x+t13BsvMoX2NhWD8LtkDG82mSC9lk
PBG5wldrM02Svfd5cdEK/5gNhik90ir+rVIhEaOxmdU6d/EKhUFhDRNYruitPc+B2/C2CLFW33Ql
3QbCxXLNs5ewgcJvhMjbmmF3SrUZzyuHCVPnFKLgBwbfUXW9DzHREP7z6qRH5l3+d3V69uu96ZMB
83zn4M44UTE5PUtYRKDAWojbi57ctUw4eGpnRYVw2T90g/Jj9RfC4UfAmQaj1/DxJhy/guOi/58B
U2o2gFqNmsWfnAtccNjpNQu5fgLNWWCFOfWtzWkJ9vWQjXfydaRzLsKusMxVEC0ksFCXhUd9LpVE
ab260JGd91nok6GlAf4f1Tkn0TmPKTDuwJFjIwmtNn8Z6hKxMZ38gEZsiKHhjCnYXbztKt/FmRUn
wasx/5Q+wHaZvN61tCy6cU4rldNOoOwyQx+pcCiRFd+kBj+u/xlZG+wxwF6kHrqQD1Wmp45jKz4W
VDIDdXJUZrqD9cmJabxRarG1sSQBLmqwQSCNwbunOvPsSKKOfoESGxpdA4Mzra/5xQF19S3Pog3I
Xua3StY+pa4Qztq56xEbYAk/kaJNDWwH6P87E+3p9ge68djwnzQdzWmD2wWOUIb4igXum3VV8QxM
DfTtclLP9vyHscRARbPBt8KfYgNCu7/3xVsQhRYrr6vpHXcqmE0XSSSsDV6okZwmxBAJxZK+DoVR
uhyQj/InvpKSqeaQOjGXELHSYIBd1+Bl8j+4rsP7VTDY7j8srkk1VTUR+a0YuKii+ihxpJCP32iz
gsp3zle1N9bHT6js3EG2QLb6tFG0XryvYfvsFmayBkJXRZxfuMeMylzJz3lv7g+CMOka9RRc2zAa
8NyGy5/+G5rsUKCyYxMUG91V9bJ7LJIQJh93XtZspTyEypGAycVOyONZLFiZ9UmfZtNuXNYDW6tY
FaUlqEubkZG4d/Mae7OkFpVjxnSqSfA8gG5touDV+KN1xwah959iarjvtNj+tQDQKZlyWJtN52Kg
T2EKiNQzNegBaKUo3rPO5ZpvXb0dgs5cq1GXVwUpp6WRAd5/L6NUj5OHXGFN0SOrUAHx8pfnloxl
VmdrNRe0k2T3orykPpAG4zmx8pkGhrp1vnSDorxnNFipIRI9n5KK4FvqYtLVJvHRDHwJ+cU5QqFY
GPVdgjVguHy3zX/L1HqKzMH65IRM1CJnU6oXn9kj1nYokT9F7YIiukeInjmTZr0uYRgLS/PcBkQO
eNJdpwUTJaldoXh0raGoxRfwjVtnHRRkv3ldLPaqJKY2hlTZTwOOmv89naYMNGWaQqHsa9mgRe/9
sKEzWn2FQnH1TlqGG8bLC0bTXswPuwKtmjZydOM5uMUzmjvyt6QJYSXWFMptqDpJa2UzndVO+Nhe
RMiwfE1seAgmovqO6BPwUnfoiXylHo2WLOSxg7cVDxxsVjJ9yzcw98MYdz/G9CzfX0nTuKi/iltt
A5CzHFL8ohOUFR81MOawywStiYaSwb2+VqmRkycOLRMcxi+NEJi9V2RDSk72Ii2lQeV09jZ/ND1Z
CKw7m+IZ+kiWrQ9OuXPIFWRn3ZQmV8+FtySlFLc9S8ooWbwSi36Hc/6bgb8Z23tcZ7XxZM4ZouFV
myinb/Q376GR6jIDsdJIcWTdZslpdRfw/WKZ8H7TmS0rUTep66uu/Y0m8QYuh7k2cfGNkU2Ehs1Q
1GEI2bLyLPdNYFBMTKT3LDtAUapw14F8md47KS88hmOBvY+WsLJ5ITnQUiR8iFnIMGrf5XHO/UnG
iDFw65MjcjKtJzylZkNMEfeRhafTLKhunqe+wpSIViC6VP9zNCclIbWMMlltkHwzxw1Pe4BIMQk/
cQBKVyQK+T0alkUIi+1SL3FDbrOYozzs/KOdw9B07D/2Q/PHBscAwdPJ0T6RVFDRRyDvFVqxzjrV
B2FNF8Arb8N+E+m57nGJe2u4eCgvREgqY6I2eNX3M2uVWrbWSExM6rW1uXZhxif+abEEdpdvI/nr
8YXHt2U0wpIUodNGaQSEd58sc2rCHD4lxgGWCmb9qx1l3fzyt3liq18HSiV7vTxK+rMfCl+JBWUt
RWjiOBkI8VI3CU/Aj4RCjnz0KOMIVmBpHHh4cl1G7TF7vb7mHEJuLPFq+iw47wzVH2zO0lJrdFAo
YAX9V3hkZ+yR++M527BmkoIHfr4Al5MJ4YFcuWxJgWSbCP/SK6bBWz0bhBgMAJDbRd+QbtVBLanM
lfLxTC1Bk91rdFfx3DzldU5I+aODLf3ZJkpAlrhqWyp41JiBIKLxSdkLwqhWpm13IvcUNMdg1UmO
wBJltweWi5GsWYUBzSHBjGmxUhIsBYEtcgmSx8TZZ3Kev0vab6XPPTvLTkJMyggN6UiYBbKQlgEg
FJVzWN+YIc58xde0bOuajCSk527nngcTdYaSo0vcwAnOnEdJrFoNj3pHb04rSXksNaE5WdFSuDBv
ozi2DA21AiF608ron0Vs1CoMA8/5KuEwHLxRyUO89jGEmkVq6lijT6V9HZrTlg4c6qBlDtBLzcrG
UqqxIylE95kkisWp+QpXQa4fJoR0LpgNIMaLsN7DCZ5r+NRrsa810nRxffnGGItU8Pw55RNWHaig
72pXFV37WzFRDDir4qz1vcE17eBjSmnOmD/8y06untCtYl+ZiHm+b5OVUF0bsgThmgyXVbd4mSwq
d04yzXMNlmbcIlQTUNsPZpopAmfEuUWJp9+P9o2YxBAUQlngfE0JI5GVY9ViGeUJMFl8jP7lhYe3
UUcjU64Zao9rAFWuryCtDdtuaIgYnBbBDWeOrqm9N26HZ2weG7SdeO0kocJLQV55F9oeseW6J1su
sQAm9IICiOF2WUkAulU+RVqgsJo9a7tYjevnMW6xXPOE7MsqspuXpRXSNC2+JfCXMg1UR19AB8cd
0vUnaIfwgO+P2YAABZ4vVEo8VGt+bVG17+9a4tpIwf70OrO1NQmchv2+hgHdH6WkO1ATIiqOh9mb
1bMjjwZetFeWPuiXtO3L4qnvHiszmN+bkqSKprNqhMNdpWXMkUflIIKhOAep8XkCB5uneyQ7kemk
Bbzo5y5RfUfxwKYhmIjwEclx1n+3uzFTataHTcGM1O6IEbecpNclFDrKB2hsRmeRlbr5keCeScAm
zq5V6yQ960Z+6JMVJtxEUzVyzwuya5BfIR4dBTplVbtZ7VoSJ29bM1QizL2PQaF4wrutHoHFYS/r
9OqIHocZPsTjGzEMKcSSYOiOvUfWJ7L4A5N9G4pOKCPN0MBMRC4nGADGwip62jKyycLmHc/TK3Vg
USv3OZHUbGMufxoDAGSpfK1xkS/zwSG224arirNl31X2D+hgp7w1r80zSEYCYV+igr21IDvX4GHx
EgCaJReerjaB0O1G+j/3G8Zae2Q/0KBZVYJF0QF/HVJkEaPn7naOuIiOaWCskrFas0DDcckiODZO
fLEf8pqAxyAh6YKjXiRxtDJOdcPaSsWxqfW66tSj57bnQ1sV6ktPuThO0BaXb2mTZoNTtG7csm87
iQGTejgvyFvPDT/M3xA/xekj+Qvi3BGQgjBq01yiz6n3T7X8CaGUoQhj+Wi1oQLA2f7Ppq4warhX
VbxX4ztRgeYcnNSQTsg3NFwVIs0ymdExiZRHmesxN139+odADflLl5leFfkZ8JA2eLysZ9lZtiW4
QDEQEIVTPETG+ECrRocxvJSRafob33mDU5nac3sg5nqOzGyTzhtvQY1CkTvliWW+4RF1zR4YsoHi
D6/8mQ0V33r3NqxNQS4aQGB/JbU+9FFl4So3c/cT+FTHahYGCNtSZl1Nb6j1lIc50bg07X4/hrJX
HTB7ILYNTc+aMQjK9+3nsZkjoAf25OlbatwaQr9B4zvfZuipjMEbhD3MYsk/fPJ+GDMzKBFWTXcL
Lv6vT5LQE5jcQPMtLUtnT8pAe2MNvBNnIZgyoOPoGt6LE8pqFBfErsyGyrcmC2dN9U3eSnekuRp7
3sNDVGGQEjSG8U1RZiq4p41ddHOJcbigb0hw6sBjtGIfc9FQMzirEDbikpORteu43X2NQABF4OLI
JlEPgHCaG7BW/bSfIi9zuaZe8G5/JDs+/KPYCCp8JuepQGrXiqFh2My96d0hYtoJj1m0KK3kj6NT
lmd7thJ20OlmSGAWhPAaUrMHjd4LdNY0XmYuhFOL3BKKe+JzZYeGh5hXJUPtZ3+EpLiBHVfif+5h
ariJ2TjlnyvpcevifkOmiq0zMwNvmxRGvm/Q0YmO4FxywoeoYrvilyBK42+XAtpJFQvmQ3Qfa0aj
9494RGhq4mPaTTWNazB+t8mZmGOHeUxEBmqo9y5vH6BTl7WMTw7n+zjfLGnkse58pjmpMmfwZqwN
HaUpghUzLv7Q2ehdvmg6UjNwh20nTszGjZZJpz17SDCpidCR1XQMFtQkpO6A3NHBsVo3vbEeMuJu
Bs3B1rAt5vJX+M+yHWUDAalpaS7gkFAQiSfMIcT/bwFWSmFjzVEd3SWHKHOTt1BGGSXeRc2VUPIN
15eVVLfd/+lCg0AWtgOXlCMvBZPqmrW7BlIXfhMwt9gFZePg/B3gbDr164dmezLC+wUMW1aLIRaz
WHlp6HO2aEzz+CZlqNM3L5BVnUycproaXWxvuNW/dDbIJrTwa6dAbeBCKqRrpfBCQVFQHrl9pAm1
/dFHyX+TenlRciZ0Og5nRNB3tQDm2zfbXhX3a2gDygDc2KQsn7L3IAo856lol6RdO42XWWWvCLUk
2yimeAlYIULw3+wX6L8GjgeIDhTsEB6A7lcyYPiHFYNbiUYGlXVgkJEGmHhahFBfqIlzIMLBbxf5
iUoCpK2A0Zhs0M+Z3Brnw9eFXo0uthOvJRARFI2frLq2QJKn+eJWpNdCsjJ7ISe5gyzvl4H/xWKM
RtwxiPOC3kNo3D/ZHuV09cB3G7CyvqSSiZFUd2AdCM9BWB4pgoX1xb+IfJyqWW7IFsnKumMKsBjm
HfKu5XwMEdK0BLsm5UfVaPujNMaJQNS2GjC/6aQTWayBySs+KQSIImXMl2oUvZiyjPYLmPvGclKb
i21xLSGdd4fM5lnLwYmWPINWvfBDovQUh8SuP+S9od4zSWBJuvsgKx6MmBaen2+jB7VDnP9A+kuw
cICABmYLHqCeDouXdDTfZ3kmm+1SbcLUmPg0C+WActyUNM6LMUSQSsGVjHrncGhmnzFVm9piqvP2
O8ln3wL1hvUxQoxJNvW3WwB8YgfFUAYeOiOG/CQluRhYsckFgEKi/by+ViP8DvEERDqizzI75c2A
PpYBa4MLdU6iisMqxuU6Z10WFguilekrVkDWQcmUoiaV4lm2HTdFAnroRInkPAx6eHGHgXqqSySs
x+u0qKyDJuMsX0VDJJU2+wsZ7Xx2bYhpBqAwKDtLG/H+r2WNyzMIEx3MQWUyUeMh1o4AEoyKLe3W
iemOLDkbzvCDun8lfsmXCKC1Q0sY3x4gEpMFGuqZa8zIgyAE07c+1tgQTfXoejmBeIUCc71x9s2o
RVvTiiQSqkh1aj3Y2rojP3FqTGIK0NlilkIGTjtdRIJNuv14zOnL6CSSyvx+bE2UPHFm4Lt3G4xV
tlV6NnlvmKdFtP93R7as4NlGYZTpEteHVnAkJ4TNu1QKpZLY0P93xdWh9N+5SiOt9BrppcZ23tLT
oM0RmtvJekrIIAnyHcbuGiYSEQJ4KvHsAAfn68he5XGjj/d07FbvFm5muvi6Ll8pzFrMQF/4xH3r
Nv80ffcL/ooQUwckFyojR2JomxccPQb6VDPguZ5d4UV/V10I6XeDWDCOVCLPWgKEkX9fHSNQZV9j
TY6+5yNcBL/eqmneedZUFOM8eqVzzFbfPd/7SnorhzSI7Id2BIJanNuo6dTdy0yVltjhlbswFw/S
TdhV2ASFIlOaHUJAP9gmPTXwZfXQRYh1NphE9EY0owiAriEikEvoc8V4995G9GyoGyGUBbEN4Kgu
RlxpEFQMiuhSaG0Gxbq77UGkQw2Mno9merO3hKd+NBINGIUkTNEXk/uPhQlgYLBTqatN83wEXOEd
GDplgYjYJaNJ9cs28OWE1mUuk+BT2aRGPRxp5yvwMzSjznOzIfwZwnNYvtIVvUDN1iGSbEqSNlAa
SssUUdPRDaYrtvOeMatkT611GqFUVfkz+acq9mPRtk3ZrwcDQgsEViJXyVw34L3pXqhuDkAIEXOT
ENCuZzPhTMoR+HMI+IgfSaCNR0UoFh7bWdrF4iaf8QVhp2qyeW7p+tElyQQXRv19po4IGJZNA/yv
zh7LG/3uR0TUdk6KQ4g4h4VwxOsVjFUoxp44BuYq/3xqc0Ms6JiZYCSQSR4Tqa8Jf8s3GFALqqiK
xOJktZ9Intc39V9zNO66meaY/C5kCGn+R2YGLAUPzh/Hw9a3uyjpsU+361qbulxVAGoEXfJD/4wl
71VBplYHbYf3MJ9PwjKIRVLWs16ZCP7yC3xYGv8SSjGjDLRnaoclcTb2miUorbZRWvpiue/iRqp4
SuY/PxuCv+yb/vzx9xe2/eK1x/KkOELjispoDpGjjpdEzYTIZZcRnBsPu85KQkxvu9c8a5UTx3YM
1UYgLeBRG5XlW15d5+xy5w/9xsqUKVfUb+GpR7MuaU3Akn1th82aI8ljGDDA94SDxqExT2/BuT6H
zIBTUZ7HNs792K8PETyVXSht2JiovAPBxvvEMsjkI0/ADa602TEckND5iLmGLg3jSSBCTfdoJM2X
7mdrUu7PuuDPGMSkf5fMt0qw0M0M9muf7f2VUHB5n2B5XNqOinkK3Cm/SO2nuBTIGLrN4An05eFu
hOyqGWNF4cBc2ImLEcQLojwdrSdDihg3ITwBqSjUaumh4rN5s8R45J7zYxouLMlyA6guGGwSqR/u
wGmbLtzAiHa8aIPyqs48yC5KyfnzQAagc5uPNDFX9cotW6vj3Mb+qzgZT4ardv9h0WRNgTIa2vHN
5NA4/W+PS1/KeDHb2JnIlcBQO/Gulb53DGkmO4zNCf9H79CDGX7Pt0F3EkhJQ20erMmkcPKLgVlk
1VnxRm8poTh3xQAkHKLjed/ykkcL9C5jQVXFfr2beChoq6cKVEUKVhQaoOsjtlyOm7gwuOr7kBik
4cvWH0VPjg2K9pJvFkBEirKEi6z9Rd/zHa2IN7l5eHJ6FVmYHiVdjjaoUl8Q+SuSqOndPECdF/h1
LnCcLng3woh8537gpBiIVU+yxPA29vHk37wmWWOzc8J7d43PbhDdaywErF2+r0/QMoFDblq9Wul3
wrc7hiXo26r8ubCJF2QcjcoBSqMTo3HPAW1AOMFbgEsmvNb7YjMPfCJ6/ZX/MT1bSKtHRXrY0JgR
2AB/hbSMZGdCJXOEDuntLQbsrvAEn/Ecd7k3+4h5uPy+BTXfRyR7jFRXUG8cT//SycfRiyJpCnOM
+pIJm315FsGO9kpbtDpX4cwiGuxWgpwJTRXCw5MHo69r2BfQ7AIiM9RUVCkC8MPn/jsbIaMbYQex
vMhUbGaE9omes5fedcfzBsDOqT1MZU41iwIo79/e3rT2poCv4ztJLzzjVNJALDmCVXILmhffVeAM
mNvV4aB6xfs6EeAtGGk+kJpOoyI0vF2uFVEdZy82gsTM10MytXvjJNmy7XGDQXaSsD4ua6fQjsUC
m4TpvfAze/5rbMFN1u8L7E92pvIoeRqqPTK9GTqdXL+Y9iHklsr+Puf1f815IMnlNV5aJfXvgTd1
1avbysHOA0zmxwTQmQASfYheZG3ZqAgwTI747hsvY3cKQJCm6oWu1IR/OM76mg1TKAdMbnd+khJ8
FnzvCpwgU2vy4SFfJZVq+LO27nnfzxaoOqB1ug7SCoE8JZLoBwZbJmWbs/T1F83kie5okH11gQn4
CLS+ZLJQpvOt4mHqyR8KId00O3F8JD+rGiPaXoIY2GKgpWbPi0La1p4VcAJRvR1jG0L8jegRACGM
qLsQicxg940XfrXeQg58/sLsbgwhlXzQv45u9VonUMOfRGyCwq/8WU3eEpca1kjV9KpE67exk/Nk
/Xmc4qcca/VJgME5OoS6ei1w6vUpcVpqBxdUzQRIHrLfgEEQ4f9mpZKahptSMOZ0jraKG7m7TxGF
RBDC4e6vwuAhnHUhwgB33eUq3DIZgTVvhCavEw9G2924isafRkkJA+qGF427QDdg0yvNNjEVuCnB
iQ19It19KH0O9x6cRyXfDS7w9xhbyzoLRxjXjBVNlMTPljNlTZw6L3GhOtj4O6V4jAhcjjway/GQ
BFLsqI9oTM+N4pcnlQh5Q4SNUSvNQjyqI4/Bog6ugcwq+PpGPwI2xVHphs8NuWMcVqLSnpI6GiJS
cbT+8oMAnUgOYReeWAYGaUkgOGrRSc9Vmk3RBULuZLaeCOXHvwcvYK8jPZ61NH9pe/nXpImv/F7x
gi0nCn0mo1GNbBzZ5mQJ20MlPNbnCdGAKg1jCA6f18wuvxb0ENz3txhODf2KTWhwpb7R8yImtw9l
euOnzSZYlFLGbV/uNpA/jnWCaCdT2syM1X8nW1YV30qBpmKaXgL/A+KqF3z2F+xK+EtN7mUNv/YX
fzq6TEHgi5jARuX4u3PxAp9dwNNsdzIr00qgj7ACTjRQQQLnWVItxEulXQY3yOlY93VhrOAFYlVj
Jp09aS7YkjPTGbhq2kq0WTcCTyXEBQHYLRge39KFvP+qbiEAnHTHw4KfEYADUS4iOVTgj11gvilX
ax8hjUdwolZ9M2ZdtR6zn41/CqkI3JYfGfopqS536QtwvVBqQ0Z64kcyhHfZXF7pnWfWmxTQunkm
Az5hFAtQmKlXrd2sBLcLwlga7ILK1mavMqyG08qlPEwx1xWkjYSRu1s7ddMtCj21uM38u42riBeb
GMdBC2+muRl+4TxEl947ydTrDvMl4PEKQTVIEdz9y0JYmi+LvQYGXf8xInID1RoarB20ek+3d2Ke
GL2cnyhqK8zPtZh/ewz37/bbZLC0410kwakiT2AiOocfeFF0zbrUg7hqVBqPXWJom0wVFZ5reR35
4R9Qp0Bi91GbQnfOpqGpqZcfrU2cezwdP8oyFFmsrjrr5/6xcQ9Y/nl3N+Q+CHAcUZoj9LgxpFiP
6I+fH6FktkptwxZNjgf7JFUFAhdjvabXOqDwH0jYznbVzolvqpcCr5rjC1mwgz4kgr23QE4XJ7Mx
e/8P0ipOvVKDT53l+ngeMBJAZMVw5fmmcTXzYkWPS9jCExlefX67YIbr2Jkr9ysFvJUhGCdMYn6k
hwRcC8lwTHnS8GzPAKwekqQ0Umjzie7afo8pyOtieyxkCyf+Yl31BdIu8BUdZ5XLGNSQV38q5IOz
vUlIxp26osP0E2udzX8kzeWyPsrs/lhUua7o4PCq5SLqdB3Bp4Ygq0CukjP/ugK9Jq119LdWMK1b
QyDARsav0lHGtzox7HMWHDXmgwN4cFUWKO0qSLL387wisXz4+WdAV68IJ7Awe3VQvdmCHKVUaH/L
h82IQ7s2DKozhEyoooqR8XgcU4r/5XLVt3pyBeSUwuwgxkVYalAGDqyea9glt0UUAEgZkLSVRAU5
OpBHm4sBW+LnY8A93yzkjhXKMLSQnAvcIJeRMN8nmBkf//R+A3hILKXuplnAe6bZYp6hNyN8sTvy
hihB6DtpnIMHW2mn/3SKcQDTVTbyQ3ByNeHl297zO5Gc5jBEc2MDF/FXXylRn0aXlU1jbyTKMBd+
P56MXJSnRcGPSGGFUvkQa3xIwLdAWDYVKIF/sXAbg+7lqvqwAV/zn2x5RC31CVwllEGY4txZv01g
ZnAYTWRMDib7QYLUcEXU8tATxvElOhQWplO8v4LrP74qNtKuWMGqeYGXBmcdcuVDyj/rdLtCMFum
YLV3DpPCZjrQHBm0AfJyEACHectE19siV66u32XrEKJwMTOpMmj45vxHL98um4V2wVx94Ny0ENdu
1SSDimxxKhui00bEUMhHzNQWWiYO6jrw2Z45D7U+18CBjlE63X/x54JfasrKjS4J8cp8pUXNB/hT
981l74z3dxxQEhYo0sy3PWj8x0smNH3IzAptx770UlPveASQaIlsNb6CLnaQmJKNZFsI4GznXVYV
NJ/5/WVjAyRKVbBjwX9dl01DJFTj1ylmR2IyeD0bU7EK0Se+C/Kmv36iHy8yoFKiUnHIkib/aJIs
qTs5oor/8xuCgYBvEdXAITkR7GdZE2Ze6HATeLnWZb0U9jVSoxn+KEaCLEPubv9tOXUKmX2ehDGm
t71PknZ5E/TFxU+g9vpyZDDfz9lwcI4yW/v1jhYhKscYa+h/wTdX6DIvx7lPY/7pHW3Gv9kNHrwE
XYMMrIToqcXFzdvkMX5wXb/3tJz8SX4TgPf94PTgdI9mFl3kWqJ4LmjL26KuFhFrhoeySfGw+3r6
sSJa80cKq+Ufcc4Ti/BSwdPO9F8nuhCGfVU7Jo2+n+L59DeG/ujxmd8u989nRo/N28QXW5dsBRxv
/VVoAnvtmkP0m/ZQ6p6AWMathwPfjb0eYPe1dlwl97YKlVQ2xrYVl2D3ZqtAUtd42yspjL/czua7
tJZCoxr6a4Y7saItIlpo5n8k/9aN6qc8DD9OS/Ufdx2wojwcDU7gH3IGDYcxl3k7zGnftHJ8UegG
75UoNGZnf6a5Gs3DjaULeCzH6CGakaMhxE63P5TLeBE10iTfH4gGK1Z4P91sxFXlT73yHF4J9ZaX
DX8BmgsO3yj+Iu1pTvm/QbHEgNZq9mK5L91PYT92Sz9JcS2w6j5P1zj6xaeyprIsEiJ2eLXr/hPh
g/e/Afq+JuoHWuTvtcoMVjn4obFQD5OSNpyS0b5cH264tSJE37u/IWvg16FsuPN7DHFOCGQLIhhj
si1ylEVdX2JcGKEiF3cRE7yVTMM7N4YpZ1msHqmpgS8bb291NvYwEwye+YWKqmvgd5YWxQroXzeG
c5DOFwgYiIiNPDqDXm2vIg6T4AqqrNgY8VgIwWvQr3+p77zyk02Qmqe/qvoPNaRl4h0fheRGgzzo
Q2kJkdETJAHUBvkd0WlnmcN2tQQvMpk8lkJKdf2OxqzCBASFrlK8dBMSVYHnJgZFWS9X+5y2eL34
IqHosxxI//d5ZlC5oGKPW4gOeUiN6OaHtcG0ynwZm0vpOByv1GPyhEXPfqG4ARhF5fDS/9NyZ9Cj
qzbEDHz8dUv5RgfGuvhmz0ucK+sniCasfzQcP6/g15qyqXDXMGmQ8x1X3jha2d0Rbe3cldozTChF
6rq/ngM7DqlH60BaomV9jGPmcB2qbtEKcg/2aHPUSxkXbeqyMciXsL80cdfu64WXaLFy5bYbxJJ1
ScE7g80kvQtghEPovEDyeBZePGqoIf0IGYgRPpoaEvgbTklU/5rR8/0nj1prLg2rY0xSf9nGYT4S
wb2Mvr1yWZz2cqR4FnBJ3GToT2aFjQCRxYiw6QPOhf0Hhekqp6zdHQhnbC5SAUyYnSvgAzxm0Etf
qEuQt3pjQiHjtv+BeFzmyPI61f0E4sj73QYyzq0H8TXY0gZshJOtSaC0W/e6xb03XCkvUWLwsnqs
ydeURgIWMAcLqzZefnFxOKTwRfwH5E7Rb0Ct6rKeH9gCX+SvkYEauYc0jeGrtru30lWSEXWjk+VD
/BhWW5QmYUEjREZI6SWgg6s8QwUKARSuY6sVLdUKY3Gr3L0zyEpnQK7HUufMu8zgwWI4LRdrFNcT
X3QqIiVLfJZQQSWhjEmWJNOZJT0tc/+Xhd0gAHkiPQZuNEXBEBl4dL+gEpu4K8k9B0LNTUTOYMe+
XvsRsByFdcMxKSF6mwmT9RJ/Bsjm7/gZyr3hPat6p/YICYjbquunwmnNZBQxA/2mZ5Z45s0IRpRi
N/Y3eIz11mCCKi6TXER9Keajq13TeN/tpRpBpAnOa/SASsgYZMP0VbwYFV9D9p/hB8eagOxreBds
/H1Oc+mTlrqhcmhUPKe7kB//IuxS8MOyOJRtpHaf2EeP5YUj/J/DReCjRncHkoA6ZxYs7ojIwcDC
mthg0YWuHijMqc6jNbsEvBU810l1/VWCIBKA5AFMIw+AVG2b/RQ36pvSVnCvwFVxrlzp6HNdtv86
2wVQX2WoZeV5FKxNiUOgmPM0/wTK8N3HXzW12XxvKE7tJqtgay+3bYqVTf+cncimWiIBa2vIVmya
lVur/xNJoTqqe25tPbBTzpLDS4i8JV/ZJ8y++6c10a3pT6vd8iaGoq+ZDhXIKd2BAWIZySgu7R+t
1fJv8JWv2gauhjmATgSjjobLoHCcd9N8277AukTextIxnXYUJxWJ90NxuW6cWsY4MT2ekaaGl8t0
mf2nlNxfsZX7Fk9XsL4mTR/A909G6bmnHSK4mdJUApUVNxhYWg59pwhNoTtUnYOyXYWTwQwl2XV1
jyoS/BZoeLOeR0CLY4CIhqtvuZb6oNQ+SREK+2SfB8uSkkdJk3CFVbkyAssH2pN+fIR2IaTaBA/O
2oynp7C40di2pufHMxwgI6JPdaHdfsc+bH/vmC1FzF0smtqt4iYMN3biPn4W0ZZBzYCss5s8jaew
T0BBWWXormZ83m7lDRAyVhOjRyzBDh0DMsZODDd1vu4k6+5v55z1o/SrbWrkrHOMG6KmbqVaM46n
/ru9qFziGmyhI4sohJ3ymUpIZF/tCTQjCdpH4GpBc3unbnj/IfxVN1ljvzJ88rI2C+HDjX2xZOM1
n7QmhMGg8SgsOp3D9dqckvt1UDKsVoqLHe/jxP73kKfu60kZbrrEXBAUJDSjr+9Z57r6q+09X1PM
vfu0I3YlgGg2z90HH8tsrkyCrZWda5LN6FZWq9g4yc1typquq4FqCK2DTn+uOZGkR+E1XWJjhmt+
SEhAIgjB8EeSsrO41/THEHR53Z+Hc4qI6L5uTV8RPSHhlMScK6OEhQZyMAEdsD3yItxkN1z0yJ+j
GOCp+nAwg8iIC/6rKncS/KVoA/nzCUpb0VvLWgF9kOjdx5SN8Kit1t72ZAhkoM+loa/uPr3kCV3Z
NRzmWl73Tj+4db8za5gqOZRSuwOWmZU3KuFxRaH7UvOsnuB9hYZlmcQnnEEkiLf0y/D2Lo4PNawH
/CIV9+kNNRUuf0+FTNFUW7pQPyFTZuizaO0PTE7ljU7B0RZI8nvrcNBT4ytOrAkmem16ax3iX1en
zW8svT0B8qWYj90YBDe2O0h3AHTZCAElX0qbSyrqZS/PTdFQhjg9tLgC+6q+obeN/Cj5DFY0U1rw
Cuuw7uGX6gmjxcJuRDEmKCh5R4eoM4s2na4fa+rKTdWn+HHn3emit9HYVe8kF2nc8paq/lklpuzw
FPbXluv9jl+n8Fuc38PkZdMlr1NdTLugXCNo4VUdW/dC/Ue1xgzwpGss6KQquCeXVyAU+Kvc9Pwt
1vNi45QcXMe2/S3RJHpg+6VJyBuzafeHTr7jLsA4lt7LHs33ul+G1TGmEAgs8wgO2bXYYqiYFZch
kT9nuFTX/UW5rMv/R7m2wxHAIJh1f1sD1dRZ1Dpa2kUrdwSGgsonUUOQOQ72d+HfdxjI5U0Xg5ks
8M/pnUq+9hHs3dNhqG6F2S/HFC1OYKnaZi1q1LKJWK1+8jEDI0+DT7TFckU2J7CuTcPqWrM/7ffE
33PwS6xbrddy9tcRJSCkFYupXWqZMXbRSvxq7TsJQIfWJaRTORC3Q5EABezeN26N5/KwDps8kI5b
IJoPcRqm4wtmhxJtqCEoFWFzC4tdg/vkSMVi8O5vZNJx5rUPY/cFzM7ClzGlNNWRIrbWsnukJZGY
AEmqExKV60wZmxSVK0jvDFtUTDRaRJPmtov1ZrGHUHUikV4xzOiRU2YDgYbiae6W9HvBHJ/p6aef
A+AyARHOnGx7ZN4SbH7y5/8W4SmAAK5tsb6xKsXEqIBKVng1CMDsHHHl7gSJv4LXtINtNnwMDD5T
Oxd+xTPaOTKxve0gKgwgoQYL/F/St5cX+HCzluoW2GN/x6IzLa9NFtepkLUlJkNUCnu00KTqIria
5zD7QWmFwmgBYqVbPzxhxBRs0wHFwAj4+B7Pqu4xjETVqRRKDlHnklLwufRtqQnQylGHB7/IKTwA
TcKLQFcPGvxjgUvNbYinaHOFqEJ/MZgphW6QpogTtpAhmHBhO10m/WX9/UzU2+PdSZKRSqDtOQ1i
I8tUFfj0+vpKya2TTySLnQhIeOBTnaPW2Pf/e13lH6TnaKZvncBNtw6uj3OP1MjB7zkCKfPGG+MQ
nQ7+Sub9rmxikhfhpe3QxDPp8YPorx+m0QoWlPbzWz1Ufrzxhdr/tO5Eore6rk7pXEg5GwRbnCXi
/+GXpNnH0RcoEq0j9DynGfPH75daTxaCMiIoTaH+nwO6CDjtTvIOvHFGK5UyJWPKrA+Fabf2/nIN
obCDG/7C58y/CVTwabGSuTBso17WANLFdoZEBgeSDBwvytuyP5cMPcwsCwarcAPO7cE9SOAnmges
NlpZyP/VdOCWKQQcoXgseiyZf84emU+4eDmH1msw57W2qBKrXBDfzB67Hc2wja4ktvFvByjXV8yP
u4aE9iILdDkE3c3jXp0X7Gj//lzCJ/X+ot4j4QFs/Aek9aJeFIXB3vtsC7i6TPwc4zu1rxGBTAjz
Qo/gI4CShIuXy3t4BItIGAiESq2O+mb2mCRYqceCQsRjSfh/3W9M9EiWEY6in5a1Bffho3d0oPii
+5VfP6lGxDq9Yc//spkJsYIqP8wAo91ZJKypF0KFejosP9XMqAqDDRFtf6qxyfejnZwywizPwBrT
Ka19Yfl+/uo5IhT+yydqmcLx71YoAMmyQzYbPfgu0Z6e1DyUbGFBSjuEwYrbFmKuqPKqM64b9bk9
1CW52JZ5D46qXTkJ3By0RkiYhLh+pkORksfgzEMd2+ym+uOyBsaEoc2cgc0NIfyr6cAczmvvBJhi
q/mHM9nyqiuFeJtKT3EbtrJGwxbeSggMN5ilTitp7xT34D4BC3/8R0Y4ejT7fRB2t2V+5oXPbcqh
VNHU1WGHx+4i9ZWRSEOVtp1WwbrGpWPfGRIeTBExCqdU/XYGiS6EcvfN5OH5fsPZvgGJw81jW8QQ
4ClKqCudJy39AJIA4jTAuxZU7/kXzP+QthkYW1ftsvJnN3/i/mK8s00EIldb62vTNJDGsw1i+h3g
o+h1NvCBcQ8toFPWRS5XDveaggEPor0u9WQ97aOgYGxhwZuNbKfPX+0y9n78tW7SfRgVDJOrlAhE
+CzS/BgjfEx+NJfQTmdXVjUtUD3ukxjtkhpclTYAsIq3xQ5g8KAgMAab43PCmueD5QrcW3brsx9U
7AliClft4cpCHuu35J0WoiFROQf82cZ0/J1cWpfdNXDFeCu3fQuVn9a45Jpw30RQqn9crzT6NDpX
0fmmSuUuwy6ao072GrdLSsoV6FjGUICqN36nsY5Hk5bC50dmrC2kyEp3YQdrZxiDy2ctiSW0wWwG
PkYP84KsbOx0SAXVlb6TFjmw7gE6SULX5L6NzOSnn2UpMLt85995986ucGhAiyBfWyvJiAVhwiJ0
BnAkuTfDRTe9bkQ2Si+3KdRv4RyiD5vmPQOKWYu1DbFTCgdiIZ2NLOO1oZJ0a2ZQR6KoevwJRo2U
enA4n1DZKFgFwSOKwytVQY6h8Bi07XF4+jRTonCRvEL+BfCkbXTeo52dPAQipNA7lzrvh9NVGD50
/tjhZYB4MKfmfskXI5koItea9AJY/cgNH9Fj14sSvi+OSqPBpnjSKL0d5y/wy1YgyNFE3tTJRBbT
N0AK8vAEUoWRsamH6/74LRnlSd0v6WF7XvCbCzdqfbYpBlwUwsFMjWmR0bfhYMVnI8xbOaeHW/GQ
LvDPHR9566YOu5tH8M4KYX8yp8nNidN7vsxuuBVPhVXEauSCJG00fx2DlHhXOy8nvY8YkHqjUpF9
3Y2tJBX3WSFQuwwHJNVWkXjY7uSBdqJbMVtYczu5TPX00rnMWfs91SE1ZhVfQbdoyvr0r0UUN2sg
g73LrfWnTLfRe0qTwLbnJKBUqHVa1JboXYnDS9ZPuMh8M/i4rC8ZMFZ5vfrZfEUK8zSCST0kUe+u
TUo2snYhvVPcSNHeH1aQS6jbn2a/iSuHQdLXwJzpIq3v8yVIcRX5K7mwsKxzdsLsFkrt4sHGaDji
lM0TBWQzwl5apHQwYAlfy8JU/XFjORN8m3jdcrvMK+ruq42X8B/f7DFAyeU8GG1yYJxjbZWJCJL2
ABTT+K1Dy5pb9q72nvKSKWRvgKwe4dgWe1CF/IFqEgUSUy8CMy4BgNlxYOBzzM1zdi2Mx6meYdhk
20GCXgCo8ybS/NpRujHNwCecOq78jVRg0RmZQHTZqjooZEdeCLQBf8EbzvD1O4NkWNue1lhJDTjy
CDInfFX9O5EykfVdJDh+RHx5xjr4iHYmD/imAZFTmsr8SWS+/83fGpnMRuj2QGI7eU7s8keM9w1V
dukZqZ92X13tOtk0ze5kCqtIkZkTEnvMfOTPi8tS7OM4jZ+RHlQqIJbx9vZ4fC5UqFERNWp7QpP0
herbAqO6m5O3k1KsjGgnv3uX1sdyXEjp5y10vH7jr791dFll1CXNODac+a486Y/i38GWxElEGXma
A0J83DlNrqBe6Sf9/FMYjvZBancLGGIju2lLVDk3YDP+5HKS+Qg5mlmNOg7HjcyEXQ8U3kNo5fGh
KYYlYYcfyZaLNuMXyH0KHRsSPFWQqU4mQJnMt78UtCJZGrTSDgMvknbWWjmDb9UegfCuFJ0OoS/0
Agb8fOxM8ERrddTGJfDFSRQcEaUWuzdB7klodXiQlTCspLD0pmeSdrDvQpqNKMX/dw+KdbX3kf3e
MK+BB/SzkR+g0WoN4APBnHX2oDJppNHXmv0uygF331aeaff4vGuclUduZ4reIyXaCve7Gi/vwYo9
rS4RaFEeWjJSh8/CTCi5Bb/tIye8HXdr4JRF4AbW8n8PZj0WFJorHlt5NvspLAk7+V6UccGuxnFJ
Q3f7lZWQCqjYC3+txv6UYv2MaQk9WPlStIbff9p6yXvYbMGUDeCebBIw7NMtFQO/x6acUhGWRqDH
wkaZZRotGs7FzJAqtGrT8iXFiMfpBWBZgMbNjS0JURAn1Oh7jTah6YyF6+o5leZbi6NvQ+ARA4zR
PGBOzEAP7ctduoqsJdqs3hlylL9lPPkY5TSw8Z+eaDiwmFqIzDxkPMEYQTM8yTfZr6ecIdQT/pvd
dtUuCcONw7X+ijP6yDuKZ/XagOgMCkCO9PWpdVJ8qcAdeWKxEf3HxBK1/n25q3WWN0Qg4Yxny3PG
Cos+XiN7UwfrHEmWypfkV3tS+xfEKGAKQzKNth5YGJsHoQiNMkdMY4QgY7NxIt42cj/rzvp55h0y
U/SMQehnbZnZgm1G+TZzyvAgOmG7/wfNdxyxbEw4tRgZcgtZLZyrdMis9BD502bq2cEyfwOgawzW
Y2Z6JCk1KWhqyMTjEgZqudLZfZ4ckcpGKrmQSTDs9dZbnk5HW8vd9wr6J0ccc2JWSqw/OTWjK6AB
ReiRHU3ZPj0SLJabyDfl8Rjqk/wNF0ONc5iLBGy7+oPlfrMPq8VFqDJ5h+bHAAI9U0stkNCxKEYh
R/aTo/3dVIeOA/EqmPifZ8uDDqQzOpSxOGerxCcK3NLIbRULQvKXKYjLuLp7XhPSCDX3FObOUt0c
xhseuldyXaz3PvXxI85GIkqrpyaut75WH0/B6vLglyd+1a4RcVHmRhGG3Bo7q5yR9np7UQ4olSJR
0Et/dV8sd+irDrPq4XKrkx30ZsUH6y1ft2dWwVWyEeYD5Fsj11EUBMcRzrjT8po7rKbp7i6+ssac
UyXXa1cA0cw6srvviZlEEjLwn4mbK8rlfS7vjOGT0Zd99qFojJrRFcATqAtMOgKyUSY55lwFKBVM
PGTiZHB3k4qAJ6YvG6am/SFu/dGapCidSFE3DtqCRXL0fIsYQ7sHQd6EE76Z9rg7XHj1tcMm86Vo
cG6Rf5nkO0/gMyrXWOz7JWRuxw6/4+94vfvSVSkqZ1XgJtPVg9KZ5atI8NGnc2HJqysbNUqlbcgs
x/PNWXZnUKnbNOimA75uhVntAolpNXeXHxCIexRcCw//1LzPG8nMU7FV2ATZXC5MP/Lh8oPQjbIZ
iKORq4O0jG7EPgGLZabspzBZqrDeIdC8zVcDT4UTY7Xo/nMkVK43ojhgKBQ/Jtna4oik6x6SnUIp
Zx2+9ZlduVmBB1/1TrV0S9sp4IEBo85TDrUEb3Nvud4eIeHVSZkEgnoJg6phnXIUI52AnVGTtuCW
gXxwElCQN2+gfNMIE4Y28SzPMVs6Raw53gxdBxytFkaCTLGE+jrAsj8Do4sZUo87f7hZU/pnXGKt
lwsUwMckJvG5fV9Q4yAE3M4LNY7kNFjTWJIx8IATYuc7vC3aaaE+d/VuzhHNB/H8g5OWsRd0ohbA
wDMZqTXmhiVDBEP7V9ODVDTenSoQgACu24azXWjqo1S4wDJr/7ywIvV0s+mGVkESRKgrMOIB4qIp
f+8IIp4AUEN9Cuc4DEbeSFzaeRSH/u4pSeh3t6t9SOaqlrm/6g7Uohyr/Tz07unLTb7oX/mm4Oio
9FalHbPNBeiPGmlJDAAvgzzPf6F1BQrTpM931DdzwwDokNUdIrWSmUHxQvzankJjVx3tc8UOwlHU
JONarnT0P0cEEoFUmwpYonvkSTDHeRP4oxvpiZKqsi/m8JRzpyOGkB4oqpuoLstqvSFwZj+jITLB
LmHJjbFvf5aLWFVZxr/bY65+Eyb0ndqknibRqeFKCd5OOEWshX+lAPm3DEzM1jCIJ+Or8+C5W2HP
eZLeHIlg0iu9euIHxDKEypdyr8NXcbnF+fXdMorS3ZKwsYUWN3JiqrYcQHG2tt2GRYkQ4t4W6rx4
P8JSQDVuRhyW+Smh01+p0scCuHWHE7QCVS5BuVkzT5BTA5J0qmA/4JecSnDeDJ4MVP9MfgCPZXCB
fSh2FIsgXSpYciIn6TT9H5Zh2xguuWWCdVsuXXtLIPtTzD9310LpOGEWn21W45x51qUt5dI3fm08
lCJQIcxOtJ4i9AwesHiR+6XWmVgYhWFFt+yYG1i0xmNoND+krnfcr+vicu7KRT6T/3c/8olFFT4U
aS34m6eZ/jNhsqi1+qoLGltH9VrRRaScXs5Cdmr5FZvkn7azmpUMrC8Moko6hp3huIyOK8HAtUBH
BNW500pDRq509nYmqIdaUZcL76s12btJVeiMPTts0JwJfxb3Zt63/whMfBaetOlHFaCbB/iiwcXD
qIYL3KGptK+ony9Fniz97MD/jAF3GsVYprY8ueMqAEuCc0VQ/kxtrLLqr0SeI1MG5TOhLNvJ8Xd6
JChQvrBSYZvWuxXPnnt27urp1hHFVlQFL/brTESW24s1YkhmAlMolrLgKiEGj8XZpz4oGJXT44p8
eof7qYzZweWgJqiyTpiLTt1CZO0m0xcZJ2fkXznLWOA9KtbULGneb/WOEdvs4tU6ME3E5WeOne4H
BNeyA4SMMXMZFbr6NztV8In37VG9YWRAS9AR5tEk+hG+umroL/eI8DGU4BQxboVpJcQNw7vv+EO/
9TbKULmZpKcu17AS6DDzFeZBPElEihbRp9i+cdJ039GuMMqthADOn6XXwwYA7Yubcj4rRiXWH7Yj
Y8mwPUQWC0IWGrI52S+gEbOHYVoVTMHDwDhrgAlZjl4P9bCS4I8/cvZHnHis5HXA9ibl8+UoFmPO
CID5kmtBv3NOLuu8R1RlsNBvuDe3aKlTFRqD7g56InYdzaH7mb7oFEPbIZjT5SIu7ZzRknsDvZjX
pGQnIHkkh0UhWdf2Z2BzBSUSxZyIprCP2GIGdX/OK7FgJMM2NVTI/VAMJSv7CKpKZv6nsNj0ELxQ
T7rEoHm2LWbGG4vhz5TYM1TSsVeGKJgOqKyvXvzMnnurfC9dksMj6FhfmPhxvyOl1gklJT6ZVlzG
u0o9Nd5j55qB6/wcWb9L5UfpckWhkM8RCGyjMsCme4RXG6Gp9kkqlrz+RMkfUnSyPz1ODStFKF6n
R5cQcnGiQzaWFQmOWBs0p9If2rCRBGn+XeDpKuA7iZ4kF7uKhFCYyICsStHSp6v6bUkuwmn0lLu6
iLrMFSRL9R/GOVTZBxA9aSO5wMeyLxSfwvvUvtYzahLwcgajwHs/ygJ3IFR39nY9qDHuW4bbj/MN
X25jjQsKxjuwpg4R9ZLB5NxD6ZWj7zB3wSTxoMH4u6ZZC2nJ62HjZWsm9xi1KVjLjMkCRfhBrfVT
lCV6dCQ6aWsyKPAqDM5sN611KHNBYU02BTqap2r40DJ0YQ35NMx8d0vCQbxj2MOlFJ3PJhmJkwV2
TOHEF/ucUjcM+8W+VdkNndvTiOOTmofLIJhO4Xk9cybVfb8xu7bLymWnU+WW6iK1/EEUaNmQ4+ZY
ekNhtrqFik4/SfeZ16/kTFGCUugz916TMtFpFgSkp6J9g4XWgs++E5fsiq4/zrjMQysnzV0rcYk6
pOkbcJTMQKksdkKvxXPBx+WjCEXAVqCPJVEng10sBpH5zqBkhfbnUkOqgl4kgQn/VK5p9TqRpTGO
8Le9+UDSjY7+BXjkzU/SLWWJQvXOhL2t65eHyY3AeG/tNFLYsV6SujmB4oi6BzpgFClILkh28u5V
mjz0XsAx7iEE7hHYZuS7r43/Em4wRTZj+RTsyfAZZbv/Yt0s+JkHujY2HQg+rUI8xjlTcTeTCN7d
x6J82qbGdRFftb9Ko/zI4pH/WdHz0/gt8Nn7f6JcVK/MW+IZRjI8LdtzYwuMYXyIT2dUN7UKvbqm
bJAy/ccSceeWMb8ZEHo5pZ5lfhzSEluK/zV3Gbm/duevcP7OHozmiyDSh7t88B0y0iS4itawwOLC
pbAnTGpopgRG/oXCMnkLIA7J5MjS9SaZDPY7XT9mjlIN0MwEX5JLCp2HwMelphMHa8RJsjdf3Zrm
HMw+I7Vo0OjfbYg1bhm9XePvqUrkUE2UUDYC4oe7XMTA7fNxqPfIBSRHqnrpew7Kl6hhh9D31g9Q
bhrQy/bPDHTnwALZAaku7z8GifVBwvt0Q58nyy4Z3re9fflSWh4qKf3WFqR16FqeMxcVrF8PY1Zj
5YIV6/1YAhvFev4JhK7Miqs9AxG7JZlXlBvTrGNV2eBwogYrCXZt0TL6osZiieij7OBfRyFqtiBi
YKbvhNM7+czUW1Jb7+qVVj7b0ibJUXjRhI8Pv8QzOo4iwBmjT8+ZpVJ6/4WNRMErSqV0NV7KOTQU
HWiYOaelIFFJzNiOyVnUa3u4O5E4UrBFq/sTjNA58OtLI8ykAo/JG6h28agHk93PgAvJtbfFlgEi
y7WATQXvQIsZ0miLXPcPTkv3Ujq9YmX/vNiGw2Hd9JXQ7NQmxYkrz8VkUn9Nj1E35e5PkLxDu4dI
p2835A/HZME7QdyJy1wEr0kl1tJsTVC5T2LQiN6amBzwMAFEUnIg1ElF1eFLVQinrW/9885Atuaa
EdEnoDovqF4203+NBwj2zqS2PptiE85Nw4kd6H/xJpgVtTB0wGrqqfYOzBUfQ5p75WNilVOtQlkV
QvTnRedEcT3EkL7oxNFlDku0GcLBetctZmI3E3kp5KSDOmHyuBFwknXz69cRHO14pqi92rJBW419
x4T8D+3Ra/zzJ+BH5W4nDEnlPExOE72gN6IFw73hGL/i5tpycRFVYDlWAajPTeZbDqCCLlOJ12BL
xqKd+BGak8NoAJXJRUHfsF3XaZP2FZDFi2iLr3eMhs7WYz/D1o08TLOHudbuIPaoSZCeMo0ksINa
/TWmg5R7jOICsMTa21uxlEBsPpfvkiai4xpG+RlGuRZuZlkzW/jXPITj1EnkYXcY0raBYHw/hGDi
vjSx/mgHqcsob1VLLYoNhs2AvbQDHIRfzskwSVPt7pRiFY3SRQv6rjv6slClIYxXMCkt81uGwV4h
pDqpkckyDPQcAAZcL/bNlCcOzi+U1jVbqQVTwx7xs6IR5fKVfeKLfyub+GWVRejtQGUCDZbcB82K
GegwKNl5FgqEPzUxBJKzOrqdsfu7JqxN4r7MTBvSbaoZYNdjy/a0BiO68IIspRYHlydYDlQ5eCg6
KkMNL9pz6Y74gmMXO7DuOrlHy5yEPkfmqIW3EWtIpQoOW0g/cQKTCIl1uuUohQ7jYHml28nsEZnY
Nugy4VuEkXX2rPVkzhIrhNA+Oq5tvg7BULvbwzvSzl1EPHyKyDLW5fITGmIYEJ70Tp7YzAKG1VB/
yfIQjh2Tb9unKXQIe7Im19IJYzDY2MLER3wlba4QD4UM7Skplj3GoQkdj0sv6YjiW/J2QuPtgUQe
szeLrfBKnPvXASTd6ZfyFUlayBU68v6P7EaWJxwYFn3JW+1N1O1J6DbdnzI7EkAtRutVncAkEkmn
aS0oAE8oiuqongciXvvpzT3IrZelYCXOZSTkXUhNPtTNs19y6y87AlmDe7mJnKEYq08fJbcLGh0S
PcLbp9u4ey6oho4RuAlaLKkU769XJoCiDdT154wYb6h/uOsn5PrCloUryKUG1oBBO9e8DCA3SNAw
pgZ79RMh3K/83nFuajXRQeV2RxKougqzC2WYExtivBs8Lju+Qd4dq/1ny9FIlliVwzH2oMaWshmu
lOngN/4ik1f66wT9EbaF/peUSbiqVfj/+bJctJsQ0kR0sNeSAwBEdbGGe3XdkpfWah767AqSFf9V
m/qnvNzWN5SRj0xQxWeDvbu8F7AtdekdzSmyLZbWI8UhLk8bQuMkHLoJ4OJPT/uM73blVFw7zpko
4ptRGM1xopUEBbBhIY+8ZUitt1DYiRP/cWN9Yjyn+QnV0yhLnJTNSnhfhlsNektSmJ+41xmTdm7a
u2RF43xd///RxqlktF49capvQAM5XqwvLwlurFO5mYlGsZrLMCztT+KKoOKtzGvwGmj9US9lZJ40
Nn5J/8XF/Fz95/PHYQJ8W0kHS63BoW/Y4CDxXKxAUTSgVpZ4/BDNLxP2rTQUcX5Zb/PCjl1iKnJZ
dcKN97LrNtEqN8J/Sqy8cew/WzfLbCttoismPIsvA3KWxa2IDqQXA+nDJ0LeE42Rqq/PJW60Bod8
unC4L820O+6QoadNVLh1lEV6mjLbbvf5g6HAAlA6Zh6AjFTtutpr1BtPG6gTNhFX70UiUbj9BGY7
tGcjitGFBK+BDumSlU3AosjFLSE2mH6fT0osFBsLhuI0SmWgaZ9yh5keN6fuxGVlBbme3ArN2mtG
12gFZUZITp5Cjh71t8OLc/e/YAHclu5HLm8N66Dpc8o7jWmGOd1Ur/qXsBhEc9BLlY77HbVQtrFJ
ZJLTy0i1dFIw2GknXCqiiKQR/cd3kRkEi+tQjFM53UI3/sD6nsy4NrU6yuUsxCvUYopuW0aQ5xX0
y/Z1yebe0rvG1HPrXmdWeEp9jjBEOLR9A1P14oBykS821S4VBdI+uaVqFZic0MmdeHvqAQ+H3RO2
7Y7EJ0TyA7MsAsMSkVsljqK8nJw4AbTscl7i6SIi8U//cso2Ju6DDtUdma6M1jBkbZWqcRpZnGF0
O/JKSfqW7DwHKLtNE/nnqFK9QIed4aUezSZlL1rGzTn+CWpRjQREbUci9Fz+ZDltjrRCzF1goMdJ
ch2/eyXAcdT5c3pVJzCddZ2HF1IQkERTPlPuupr4TmGfL+STA9cNoJXaqe/1upKWGcJeUODdzJrq
EKBJA8fBCFox34joqeHyEVJM4tnPXg9KTZFzIHleLqf30tyKAFE+o8VF5k+qGC4ty6COvqdFi0sQ
c+bfykReutrXoUGy1Pxlxzyb/XTv6/9Kj5KRJTLGOpotH98bmP+O0IjMDB2j6OQYpu+h174dsplH
eqku4bQPssdT5JXctd5um3JEZYuwD2Ha7behyXAqZOQzrooptQ+EFDzXys3T8BYcwjIkqxTzQVAf
p+l5GSXokXR3tm9CrKK/TLDttVCZfaaaar5PObbd/qSfpYkNMbBLMaXmG6tOgnhJQVq8Qd+mMyOw
x6GRHETdF/M6aF0m65BVSw1QS1K7nuj/ticSrIKPqaV2ORfKHttkKeRpXpQ+YEUDdC4kA2Hb070N
zNkxsICdGKOmCkekZegbDu8c0xFMbZicMSrnslxbO4X15hjw4VvdDfElJ34c1zbQa2aZsgsdObUP
KiiWTOGJtaU78dmQGur38kXAcy3iJcE3axKpUJUEbx6rjSWiOKlvFKCUrVle8qpf362Tf25hS8D8
G+t5XtaAL8Daha/YllFlVR+pmmjJwRlTdPs2YXeLugzkj+TQ40uS8873lxGke++crbPR+x1osFyv
IxyXHLZSY0+zK0N4WyDYeCEdtbq0VfSjhgVXsG0mg465X8VE6xP9Uzh33HO1yIspiXNYEFwCGKbD
FeNfVELeuE4O/o4JLK2pObQTBAEin6AYtiPaDaMo96KAawO0etWhA0sPAPmeBOK0CWmS8U28WQe8
qUFzNe6rJ2okkerf81Kft0alNTWSqh3/5hS/9N04lvOPOVO9fEz/1SGK2jKRn+v4IA8SID959doQ
OXhRmKqkZpBKnhrMBQB5ZzTjZppoMThtAAohXKTwMo7suvNuiGsqRR47e24tl6yT8ETfjZFSvms3
I6ocqD30jIwn7gxO2YzEMBA2sW8+CChb4tCaQwRovvYbm43FI92Y/xr8Amvd/EpRiFEZXwpsmyoS
qLTJk3TA/dcrgctaQlqjoCNVtFJHlTZLlq8EhKY3d9OJbEc6BJygPFBz+SgVQc0E+E0ejq9Vkn0L
/xah+w6sUWvQ/r4lPAtTH8wYfKx2jnNM4hXiNmbXgEwwlX11r6Lig6dBY4UXwyfRVc49xc6OA+ZS
LlGwDOkcYyIXE4Feef9lknVPBd1HxIkGaE6lYQ38gC+SvqBaXWZaUpM9+M1iHOYV/IHwOjMFZwXC
s96gSuFA6oEoF0cnZtPJyYMMmBKdBHdwBshpalqRiUuiui7EtEh+xLelkXWDkriC0a500cFcyEgv
bnVlBwp5VEiw0osobzGXg6/GM+jVBfJgtU6GaDXdQS073NbHQvUYiDjsUTR4bfzpjdHS3hK88k8k
OjspWp/y6ZXN17ZVAuo/mcHoCZIkQ1rWAIHKoRJRDL+c/Cg4SbU8NlE/UOfEzgXmoWkEgepcFYyq
bUn0kRUOuDeVmb1TMKZjcIH8Y5zuPMU/stq0rPswG/0ccUhFusgNIVR9xsVklqyqLv0tvxCJxeQZ
eitOT4J0FCLv9tB97/gqkomvK15IyQUNnXQjCoC5Ze3o21O24lm5dcm+ajWJFIamIhtP7VLPciog
J3hqsPwXR6CegVnHAmNa/stwmk47wfCJYDWpH4iZw5s+fl0wrSbTfX9hGLnikfW3PJ6f0kRphQ+Y
OzYN2Mgz8FH0PeKxYQWbx1HJzHzvU0Re4iQzeyj2rZlSyojtEf/ZdbwAMqpfx5j26/pECsGTKr6G
PpZwE9e+BHbIWSmfpplsNW6cOG3RGDJ3ExEMQwL46wKQqHw2Xfso42U8ZZTvIiO4fPeoNg4Rqo/f
QAecfSrPr1OIukztJsPHQGdfvF7VVCSCXaXe5cGK7gZSuYLH7nBcXHsv8g9fFr+7J551gLjqOjub
VDilFjY2O4v5dLF+0LUrL2kThG4LQD6Uoa9BtD3Q2eVWBy6ZOTpbpEqxW3ViF6xGIvnp55mjVc4F
cVmBomI93Ji2WVKCdoGhhloLZqqfH9KbmaWMmOwD2rWvvnKDHykPUiR/h6POG1KxSZH7XOz/BIIs
frOk7OKRP+kI6+IfXKK/wiFW4A8RaHuoWhoenR0lEWQmZqtfpIynczFLYaaIHDfkFiwHZ2lgH7PH
078a5UruBbxeQVZ1Z8Vh0si5t0UyF0DhHK6GdXfSQNQSWLc4+xj5lpLAVdcBFXMdpLWjew905Zfk
hOFhi5BmEty1RDpBavJtzcjNtFnZ8FHySoxs4x4wW/CGprrLRGT91Gc1D65C276nZPUWge8hH4fR
iFF/RbdE5E8hcgm0XtTwTYzHTovAqebUKjlifN3TFUHT3OX0QFRHPAUPda1QxSkToGqA73bIbF6Q
c0M9k+9xnm4uBvH1m2z5w9o8Tm9NdWB4SaSqq/l/ii+XEoWDg1cKt/8Xny7ulmX0g88bykMoo9Aj
WbA9sq9Sq46Xejzai81C6tfhFFC/IfLS2eypbYtuVNZuPJof3dcijn8KJ1Icj6jqK9VqGTFgzdFe
0tckb4r5bFBsE6PTjJBUufop92YCo1FF3eY57UUEWbScsCDJZNn1CV0rHPSOeKF20L8eb+iDLAlc
6/smAb2bqrfVmAJE4oSzJRjWXrUkNhVATAb8aiKm8RJQnYAouBpx1KQ+8ev9k453sNHu/LZL9jIq
KDYhtYZ6kJkDSaX9Xx1kDkplYF0x6h2WY092QTLSi2vc7QUqLYRHWfoz1V0m99zc0qmfqi1y20Ol
o+YwvEeIgEmpLaNdKrTkB8SUTrxzLOv+soVNttmU+ZwTOp/L/0NzlMbCljhANt2Wo1ZkoTYagU8W
xBuiG1WLasmQBAZhWkhNcZ+EANJ7x0nwfkOZS5nRB9zCKUzGVT7lRZurSrq5y38sso56klF/O73Y
MP8bd9X2s8E9MWAu2ezg2c9lF/P0yS9eeNP9xML5Sks0ToSgkmHYmO5UNWm2oJnRdLtraq6Uq5VR
S4ycbVJtucaahOWgQSYOnEiDkrLBuqCmeJFH4J2ajLRJp6dvV7K9Ngf6fjb9l0wvR1VIiLd4Cucf
+7PK+iERWjN7kXRf0OI0P9xryxhGCkhVPzzgsIzG/co7hFZW2CkrPW92vCA4gSgXmcCf+5j6nLe+
SWN+LMxq5ZY4l9uL6gE/N55hJjE/BNtKTdV/cSEW68cHyKUsZQnt4SGz3/rzCs2EiPauxAkMJSPW
PZ7wHnB6DI+qXQwZB4dEVPJoo9JxpVkXhiPwzxQPYTIW5fu6deVcEIUS8ZZfVosGPOA1K7szdBYN
cCvpiTu02x1pPoNh0lQpzUTkGbPZw5SHocBwN6KDFR+q3OqLmB32n1pREdJlVK2+kATKGiTDILZe
Bx/eyNUsww3BCxD4q+6BGGF+cweILQrTh0QzWomEXP/zsngCYhraV72niaX63bKLtZoTAB/kD0qG
LGDEktDBaQH6CS0MdHjSFwd3jwzaATxACYc/jhjTXTBRVWaaFGjRkQqdEkjKZA0VrRaGdocCU63d
FOredZEhtPrCTY28mB8pDDWfu5HpjE4++vzGx2SrliGs3T4RGgfHahB0jR1KxvJA31LTnMK5I49Z
4vx24HIcDA2TtEUzTlqd8y4S8pFct4jaiiDT/9x8foZFNaQCTBIQdR03gBafk9A+7ClRhHe5KGG/
8hv9xDBWAxt3cRuAXST+bAYvdMaBz3PB+d2UYZAM47ZXkpXgWjdvW80PjDaVO7Tj9t2jxCw6kbH4
OSitW/dGLacxjCHFWSz0cMKCHRU5ECvQ4LH8KRXV+XK4OZBtV4qN+R+hzzanYe5NE8TFQOEOQlAY
oeGSYeNAXbgzOAtAbKkTzFFAZSug0vLkbOiaYaaPi9YOgTmG8JN6Jfsh3NNdtc8s1hP44284Udw7
SFY444xhRgshkEmdDW+hCrplIA1geEcr99XvIinLz+yHmMnYMdoy9avmtogti+2892+UhkL77t5t
gnsYyQWPddgKWY08VS8lLbjUwEyMgguWRYsQPkD9szNqIq++wXTbGD70Cr52i12xjrhCWvLgUXF7
1Bpvll7NQwKAe2sx+I+yWEmsEcTzKge1/gZrUL7aNLe54okLVJQFHrzYV49sBPfk2V5wj/igvilC
CHJbT2g913xEbbGYJU82+BiG8LAHH+LZAgmoEx+0z9m2pODhrO4fKX8vmCTbfZloqD5cuJJigtie
ktZqJ1io9GihOPNfr1MFm3b75q18HQDozwH9pIZbD3V2Wk3hLERicvSq2npvl8BcTht1pO7xBk53
+r0t4fFuPBixYhiXfEeAFz2O1/fToEhMb30SxGtGGUOqmbQjdbPrwAnXJ/9jzl9zRf0xTmB7o7w/
d39dvFLEsp6M0Od9iklGKCGNkwo/R/VLM1YpNNWOfI18u3Gq0dyHkCUD+9HP2j0zxGdHvTqyQa4K
muDlm4bslKhiKxX7Q9o221mR+w4mjk6y/eh3dLOt2As0NFplHVbF08dyBaWz/w7qkwTQ44GKFRrt
pdViliD/KGA0j9xAyAwJmP6+29UR7ntf0ZFi9cd0+6iET17B9ZI2E+Ct//U+MH6/gfZ+NgLcSYWH
C8osKfxoKeECDw0mPyVX+TOv9QzezSdNMlhUv4YfvmhwHZ/T4ClF89TH5fuYRggmwsaIaT5WMx1f
PyGX8ZPgtcJ74f+PBvJ/YzmYtjLz9qIQqCu9Z8pYzo25omN4OiyVHe3yNECDJWERb5SmN1ALcXX2
N+4PX3Cs58vc6AH1VUK41D1BZHPf2FiqTH9dhnz0TghKaHpvvnUXBdx+ordqRj9w6hFyHVi9S4jT
2tWzDfNz++fyQj+znv0JhHEK7FvPaxHrNa/UFRuXJbm3HW2vxeRac1wG0JOZtfsHY0VJRRFbk3fS
QOY3lzODcA3mAgUMqfo07DOgIFWbTwzUBSYP12xLBNaYhFj5GDxIxcxswQGfCLzgsg612XPVMFPf
PCEOkll+ImuP/LHHvNpxkAtuTGPI/Q/M6Kh5PY1rGIhxgUqSbLH4s06HC0lTICIEXswKFUeIZKkx
kfDnWc3NnQhPBpqe/oyQTonhsdfDE3r1TaBjdnlMADMEBWanuP3Yp2KV/MN5HcKXDa8TRYVptm5J
dDRIoVhrYTeh1vIG6uBkDogHkrMrQlNAKBeHIFdkypd7f7JRB12PU7jDVJo9Zi0sYDMEXupRnc2M
J1LeLp1cD6MQuOLRawIsk0lQlH4QLe1izza8YoOfRpNWr+UQn9DVVLiyKcGWrl9B3SlSlQULw82s
ldMRLJhpr/tO2pDxRRhGZql4zoK7IdAZMd+mv8KHMHcajSKPJn+mhduHkAdDpaGbf1XQgWtRG11f
5sZrejqAanXK4FNt0J2Abu28fEV7APjIVIsBIXdfCw5gtrwqbAr8etD6VC85vpYeB+g7GNLF1J3z
Pn2/o9VQhGC2/Yf60ZPq00dwjm8SbYxUL8F4TZeZrO0CVIIFzrqI4OFoOpzLotSUSV70yGH3UH/S
mUr/fQahOB61QTacijqaI5rjL4hYA+TRtZsuqZhsLbEUVp6AweiEiRCEP5ouQeoBBurM40CmMSWr
i9D7bWESms7OLfhLeQgSGlQg6nlZeequcyauN8eNK81CL5Lq7fZuEtVBNgNOSzr/PE9sM+891uaz
YT1pjR4g7o5kxTOD5g6gNNe8z1u1EBGAWKbTZGbTysDuGs7aIt/v4wZXAMtJno0twYLgn8qQpYjj
ruVIYylJLcr4e8RZe7knk+h5vBJ7B6gX4PkFoCbr/35+bAL9kmxmBdcN/ksIWaqH00vF5cPDOHbT
Bu3nvJoGa8b33DKsthk4hN4UJNDs6MwIe0hTs55M+ZCosCdNbdAdDQ4sYlH/7U1pnvlahJRi3uQ6
Ng+Hu1drAbYtwzodT82Dn6JgBszxBUY9CLUCBUdsNtCbbG665ekHMsrsJE6ACONGmBpqlzMzYlNz
geOLX2VLDiAFiBXz6uYG9yH8WqrlbO1Unqlt6TC402clWsOMUp0NHXQuKvVqAYO23DCMNhqK6vqP
oCQvdCoCWQ/DXOCMk60w8vMFwRWMKQBnETRj6f8N5uWX2RCAKee1j9Mrd/ol0qnIIoz9Dq++9j84
h+wcBqduRJHN1sCk/LV3ADO4z0/FutIXdjWVUEL53A3BWRzGRnf+ooFvRtzcs0RYlv1qstBbf86v
8kyg6db9UeNLNi4soUcW5++yZmjHVfezOcrearV3RL8KzTfCORpBqEZ8JzWnRr5SYtrBSmFbB1bc
FZ/CRyuMjJddsmPNPJBuNjipZROU60bNJAooLrVLOxQAGjPJLu/aeLVPGPjmfhT/9/VCpT0TmaOo
iVMk+x4iACrr8Rp5c8oYau+a/dGqU1BSE/hrjEEABa09Y2A5Djui8sb3jWzARWuzXJ9Sm4cwdQUg
XRD4LKjHAsrnokWBRLw30taWMMTgTlBVnWi7oulWwkCzpmQwKpMGTLAm8UyrKgPDz7bPTX7kexH9
+eV2ZZDP0weZZkT+Rk6P6yhOVkUOGcKFbIecczceMdRXy7svd9UTj04EWSp6QeK/rcmsvPGbQeKq
PsynGklQxMw7beg+0DPLG4jTW5pGp45lPYAEKbl7q33I9uFpypdUrXWae8osyX5rQPzhlbHo/l8a
Cibuo+OS+lA3y3nUBvcefMsFfiQiPFWjHcdI0+Fd125j8fLzBKLDC7WxSpS3aPMOJgz7/800LkOW
e/08xcMaCavhMHm1vdsVe1kdp2o5FB6Ma0FBxN0P8w02864gpiHbKK7gNHul9yH412yiGPfNZ2Ya
k9nkTQHCYW+2ySBUGtfuPR0+jT5zHLfaa9r1Da4Qw9aPGhoA8gi3b8mifImbKDtA6+PXrcFiAopK
O2cOq498vUTLZbkZ9B5Aau7k8cLfy4xnA1zxPAx52aT2v7Z88CeCm6a146aJAm10CZobIIs8vCm9
MR0lAu08KRsjVFbGf/oAgDLboHnNlGQuIU4O6dWeFsuvXqnccB8oCYO9ABVbQ0ksVTWcQVFNsrkU
eMmsC7IWh6HmDwKlVwSjon1m2Q0AGNVIxOl6B2g3x5k0mPAOO3NDUuX34YwHmiaMOwgJTHHn5mLu
IzRHMsHNbOLf+2SwP8HEt9KEcoTUNDGDryynXCdtScGO9bkVMclAmCMmqIu8NoL5gmoK3B+6CZzt
zusBP01QD4qeAAy2dsP79ab1XS0anFuShu+hdp8fVAtaAU+5qIQMXxImCE9NBREvQX04IaEsbGUT
oY2rBLdg+tTyV1Pii+5xOIhsc0Bhx/PplKnWNkilfIGn7AWM3X2zUFZ4BpHHN/ZfpHhvR1nAQNZw
SSgrN3/V7Ne9zVTkzKfiLecbH2i9pPBO41BGC2x/6L19p4I1pmBOiztt+Pc9g8Ry88wdFec4+j3h
ZxUsg+6Ktyzch2zBiRM7Jl6xrGtfEqUSBFHdBEuNN9a2O1gJNbrBjUkPz6HKwBLnXoGzQ89XWT9G
V3bejtst43oeDOfKcXquwUb8GTG6HF6km5QHd1ZVrAcW5ELDTFsQ2B52XSuq96cjRFQocPC9PnA+
xFJAbPjyW+SxyCt/ar8DkjFFL8h1LNOymR2DQHfj7gqkD3apI/Y44BvM76i8x3ANhf+8nqVidLC1
+lE12pc7AavP8s4slN4fhVT4/K/3AT1vQWzPpvGuU1lIIPAZtqJGIoVWx1r86clfr3z1o9qqo5Za
SFANBXGaY075Iu6mkOGQ0BjNt/MraQKKDOBwnAfUNV2ckey8UcFM8TWpWDInGrtC1sRucy2QBzCW
8MI4ejf7gXK0APplQPWoKjsIhy2GzFjfdVWx3wpWGgz1zEniWC4rauLzBSS5tE7aJTIxR6r9URHS
0wOJ0dOGzHHdVEZHxI0q3cCF4hyfoFUDmcf79+EwPLqs3lHyN6r4cjn+csU7EnA+zzMGNNAlVyng
haNptJF79ydu5yL8oObXk6UpO9bwEr08s+TWl+WDb2Qa732l4WoBq9Z2GoyGB0Pzio5bCt/crXHe
TkXpOdjkOChRwExOLK6S4TPxBQAGBUiMfFApc1l8UCks8QYCtDHGGaGKvlBr+G4VbvwMiSd4l/nS
gDnNGriF12YXmjKZo3nLLEx2MdTw4rzlxpbM/4hanIFt9aYrScV51P2itr5cDQ5wtHqI4GS39xkj
wnd2deMAdzruuCpdnALfZsm0TIfv9BKi9ekfm8tTOjVjiI9VcDF/P11U4fjc+QDbqif0Wr0/shrB
y2upT/uchY23tI7gok+UEMrojiDKjKPmraOVlYB8x6oUQF8qjIPTYOQ4NI6c25rVomJ5oNiMfhnI
+THtQgNl0Sj5vmt26SEOGolXWNY9cna5bTGB10qn0fKsMBBzjalWrHefMW8mO9iDe0FC5mdBDjox
YsDvwITzVGHdi08Kd+h03NB7CFGbOrmKDJL2nMzieIMuTo55UVJa0bTgWvVIZsyceV0e51Zjdp8r
2345o/KBBHw40l1TcC2wSdZXppybf8Hw5d8xJApNEmCPLUqtHaH6aABj2qZ2T8r5ceY2AkX3neja
tJlUZf3UOsslkty9x5jCqg1QDXsxgEV7r5go+d2VFI0ZkFR/+Oza5yhZ/VL9VbuyLOTEt6jbBQ0c
dZW7R+e+I3Y3YYYYYhNWvm91BHs8tBL73TovEzH5fEFcMq6D/c9tSCBTcFf2JEpLdEH/6BpBBXxl
aWkUmaaHgXWfAzc+tRZUz6M0DolgNEdTsSYLfSbNmFOsebSQTarEK0SX3C1w/E6GQMk+/KTiyhak
tF/Dzax3s5/ZiDExCPP9SW+X0afc0Flo/bbaI1Qw1gKomFOTrh3oO3v7tVZubchdcW0uCIUn00ky
xZdNoxa79GimxaFZieTmLo4RaU/l7hJlI6rvq6HunYleYZ6+rN5w9UToBeT9fUUawaIkeSompRcH
w5PlL0EC2LnWAilucOyii1FjU3vTW08haCxOQPXFXPN/DC9xxA1qk+eBeQiwafuuuV9lEdOOwhWT
QUBIZnFnn8tsUI1ueRvJlTHlVKc43sGPtMchtXzrsQnKaWsriN9MM+GVijN3xFeyQifGTT/lMibY
+8yfc8WJVqJafzGNVcwKYQU59reMjp8h81EnhyvteP6F/4dvgN0ZQWdkzFR0gWKpCi+kPpaQpsLK
indDrAoVJ5vs5gpRxX6G8z8/R4epTwKyaNB7Czt1W8nTEiLZte9hBGBzCbc+G1Er8ZwncbmB09Ou
kr+DuCDQuCharMclYgAwnBFlrnrhFM9KMJLs6UCVa6iqhR3BW2DWl9JnFiSowzOx/uyDfDsImYVO
aFeenxrXu642h5PfbQXrYbAnsdddoZ6Qyn7UB1bm9d9033fNaBiBB0ttwFioKRrAlufnpc3BAK8T
e5fJ8J+2EAawEekhvY1oLu4eVLNJopya6zZchasmUSJglfO/szdzwKV1Y+Zo4KJPGLZ5/AdtNaWH
L/fNCeIYrFAzBTZvE0uHeKBZfcKBENuR7C/DjhNaJ14xWpzNAF0qMEW/PWP61Cho3xw4UZZdEPdN
8q+HOsqGa9/LObMJKubQRgHI75UYuGY4ihFQjjGZdqNcAIUWNBGY3aOzfMrLjIv3zT0Oh0k/gmsN
hdrhTOQ5REUmvpg39VhioVjM+xU8tZAUp2yJ7yOa6oJPKjIODEEKmf8WMczdEl1YP9XW3or+2ViA
Z5UjZZKRadG8h/aJ84GM/nkeaZ7ObNrG4rdUFSoJXxNkn19evnN7QPqQjE3qIqu8C2k3CGRl2im+
WxlaRzrlxegrDAFkKFFrO/PZ6xb9lLTBrnO1oHgRYQ9BaPwJywYJVVcQek6KGoPGlBra7CvQYVLu
huV8yvbRFgDzPkpTcmSfeNfFvP6eRW1ct0ua7SBATQMFRCsYpn2UiPk5YLfG1L2oYaXS0BbpLXKQ
AeJF6qaVaTF71JfOa2Sf+fSdCX1vaPFDQ088v4EESDHZ6nIsSNaufxPmfwX4I0QnC/DmA9yNcmni
gi2aOt0E9X5fFZhvhv2HYX+PKgOUKVLdIpFeEmQGvF7LX1Iv9R2yZwjBcJ8s8PJY8ho6xKpQp1NV
fHCbl9tmATokUDM/iNqY8QIT1GuXYjjbGmw5cf9rhGiZ6wjupDtAqAAcUJ5WCIjYR7hDO9czjnqf
9eIXksxHocwW3gk24PHssDnqqvNicYM/JkX8xHbtcp9oinmyfYZ9FEnPldOScBsuwjVRNz9OtvtK
ptdDuZSeP98JlJAXSPWmBDavgZAcNa35J2NNcECUHPQwRxsYBE8xKy1Jjl39h+WzxN2LbcjJpm2p
bvV7hkCqJ/z4lQVb3AIBvb+3CyOupToz7cPBC8BbJRB9bzmlCSeq/6RnLPwE8rBQyxIOv+65zt6W
xB144H5K1Crj2spfESipldNUiNYR3rrw81fAwUo5YGe+qQIYE3GKTB2h+NBQEGkZn9gY5Guk9Waf
d9GA5BvI2fIDuzUl/ActESumzPMy2dYWsRraNASdGEFY4McThuXD3LIQGA3IROgsyrV358LGF2Jq
T1ekVyYwr+ZyNBdT0KnAV1WW2d40peBgSChaX6kTmifbVVaLSvsf8nmc91YhyYaTAtYhOJhkTMm6
ekp0v6J4rjhbgj5wTTIygGqx/c/ITwdTsSM70ShxpQ2rYhk2FirxP70frWKOxFGcm2pJeIK7QNIP
a10lAu+q9RuzTBM6YYAzLIwi9GIphmlgRw0Tn09DeDJl6TQ8rVqVqA4VSyCeM3jlkHaTQmBakPF9
GG3iwGTx3cvUSi5MU12nutuuPisJveYxOdeJF1ZIzDWto6/fCopgCH/2ex871jq+KD2BSfF8DLwl
LUGG6vz8phGnHKowhtNMAWN7yqvXuD0ixq1203IKk0NNyFQYsX8Cxmw1XX0RmJz8DLAn5asWZ7mM
FDjYtR1VY5jr/iQHZuba2DY58kpB9PTryY7/JFJT1e9P6SI+DbE0DzVl6L0UwgdGbHH6P4ZXJwuS
4Yq3YtPHmSMTjP7c62tthktn1YxYfThO9HOEYffsqQXyVe5B2agteO+ntdjjvOOBguWPO+/Jac0i
2nKKu4FJmOfWPTbXU93QIkUqrFQOV8HpmF7XTircUqi42H68mCSHqKenkddRBBnEJPA76KCB3mjq
flkxCvQsyr/92R1ghM0cBUIXZvv8aZkZ7vlo0VEDkfRYWpTv+W6gV2NK9+QGi1yxLre1k0BNeAAO
RI1iImIKWnq7Uv2Dz8Rdl5FrLM6pe9SLjgh+utwPixXD+BJawq+CA99ADcOFJsdPjFvhSKK9YYri
mVNzGuiQVSdx62fmZfvQBGWu77wqKxqnE6yd7prw4d2P/6ohM4dfnKo002kFpe6p5Wn5FrdsrJ//
6/QGVrhMo28CPJ8r/NuzEZUm0x2qaILEt9TGG8HYnI3mqD5uLCtsORxnZpgBOHougfZDZpTAG2aX
g97dsk76sBnLxujbbYmSofU5cT3hH/j2eNEHnCCTOQS7keA8SJXwdI077Y0RxRb2hmUed+9GPb3u
r1VhYws4dNI9FFWr18Fz2lbDB2woMJcgmJ7uAUqCeZaPT9lLUngEpoCK2a1mccVL0Q9pWgquw+Yw
2bdA+QZnPEHyc57RmpLnlxvbY3X7KHWskvTDaipS+9G4z54lgsDuvoA4tgEsiLyWfDgLs1BaGRrK
XQp22EatqUWA4ieisaDf/kKqyisQnIXskUMU87Pl+LbABBwNAt6MOKz6DFczrQRTRj80r1d268lV
iBG+/IF4XmVMLqbJAnCsHN9EMCtliFIsFKSpE1+kr/ci86JuLO8yMjoWYnO8B4M9RGpT6t0adOpo
UVU3/1IvmJHxZD7CvvrAXEVRQeBHD+6E+IPVNWZZxKRUgWRFlnCXknPI1D8vOU5EsTbfprphaVlu
zaSUuqtb8Evpb9q7s/7CaFUCBIFMnjG2m9uF/X3pZyhhPuBYkZ+qIXitXaHfKJQxSAHOEdfCM32a
f3cJdh/r+n1NB4FZmZzqm5k2ZFavpj+sYJAKh7j33mMnbCY/7RG3gm4qcyBkrllZ8EGsZMzzaCxB
IuSY59jvS8G7zZl54clAb3BCypd5GkVNMTHv3RBhEJLSKyk+OxT2rTNDAEqTltg2G2rY0+a2UrsO
1UTR99FRLb0EhcRhrfGYvEnMAvD2Wwcwg2qmk+jOvdhA8z1vBcYPgE0b5zEHSI+6qhfz7dc+hhxi
imzj19jbTOGeCdowsjC7q++E3vWkHXqCoDMtsqouLr+8WnU0cW7kGFxCex1Z46+ZvF9E4vXcdfpo
6qmz4U9LBvprdXu6AgU3V6Z2vepXLbsvVza1GYJVszLoB5emjHduxa40FOs6+MFwHV7SL3ly2Bo2
6IBuRas1603YX7SPoMtQWthAxbVKCU7II8E41mhSdX6OZMU7/34a9yBIyA2Sn9Jubwnv79jSvij1
4C+FYxXNsP4Jt9qYEXSHssSGOuqMP3Ipw9HSNUI456egxj1UHe8uAuqogywkR2B2r8F6lXzOTIru
gW0R/IMv2UThk+SYsVai8l1YDU5mv/V8AyTwHW5xIqtzYsu90AYi2dMFJeav8Q6FtC1GgMEm6ADZ
kCsU4gPGlrTqgJmBsptmjp3COLz+VX6XTinh1GN5/9hmy1fobm5A2RaLi8Ml1b5eZpM/lAZvkU0y
1IC1IBv+Serg7gNVf37ymDRHhNXyRmd2sixUDsNoMpf8dlDW/Qe9SuPr3ZGq4zDCpRneEG24XDQA
m60MW0LbIEs0mjz+16YnVyKkCUbm3tHp5Nj+t+EDwRsTPOnpcXAANX/Z7s1+se6dXBA5JqYrRoNB
DNZeCrMWRUBNpwr/Ix41asQuHKFG/wy+A1gkNefkn1feSMUSTdtmEYf1nsqU+JGpzSthjW4ZgZ5h
IYTt1Nu6+aebPz/Cmp6Rf0nPldAnzkRvA5TRlT42Ey6/awOa4OrWOTTvR37yBBmTu+tKIhOZigzo
mpJgjXNpzJS+F2rfK84jE+c+rrvVty5iPIp7IXVDXzHFQ5mBx0PwM7jXfWXBOBYZjYPuMTnDCq8H
j/InTO5+U8n3+HR71J4wPPQBzGYuPe0gQZruyNdSgbMIq6DQHlB03qCWpT7tlagtMpEMiyd9zjYX
M5v2GcDoBztgqUXZBJs5tK5iVuo6p7OFbzEniJ3wGKzAJw5soH53vzlmvaBzC3YmIvQyc9v06jze
4/0QW3JHZ0KpI6iD08E3nOPzgh7vUngKW/muiO8ZAsVfcy9eA4pxenT/CRFf/PWPifU36UttZpLh
FzK+2LULbD7wjhuRTOoA3GBaCjcHX6hpwLXcNTFvDZ+zt0rsBxoFDd4VCJEjDJfzY5YounxYv/nf
deVjrQWgytZSCHb5aySVyh9/IyJH28Hdpp0t/8wHzECRAwUjf/tBeRMZKEg5+0ouaA5lEiJsNpnz
CrglDf6wnFwbNzPfeMkl8WrbEeHbkQnWCwLwHRwrOv8l471SlGIjrPcrghkHA1hxSRZQgQD/9CT5
gRsM1YiK+QZbq37qk9IdMdKhtRzy78+HPIL3yt2B8xgWPpr6yuduLhJDSGE6fUYzz+Hig/oQ1hFF
9DMvpRCsoF+BYsBcQtb58GMz1PrEhBxSQx08lABhHlXbUokCmOrMCadC5zSeujw3fJCH8ERzrtZe
8qoLv6NGwOw+3lmfAgOf9NKzbe+XZH0D+/DBw7oiOqp/EWuqp21YcShnX0mFqabdY+B4l98h+jK4
o3qkboh3apov0JVjdNEcuT91vx0oMi3IARCwu4opKNJLnBDo1aJdctPCuECyBHF4kOL93cq59UAk
jjzfySa6PA4IBxsRAIabE2gkp8uec3A3v+hvGYKeMq7AfMejQdh21j7+lZJNyF9lrkDcWTpZALd1
j1z4e1xO/lAq24V4iDenmL+ofAuWvEnd4y2rY1GCHda047/VyHRS2X1a0/eHC8l5DJZkqMya8shT
4uC5LC11T5kYOvO1+I2cItgkS3GszmSXa4dxVrbuonbSUIqRmT9zlmSbp3r/f8NYzA306UEYdL+9
XCRdkHGCJNiYTUw0R2L995gDfqpoGeBaQ5WbFcb8Jvh5R97LOuQmXfMonIWPpiIHMsyd6hPK+XID
HIs+0Z5Sn6oLAcicKbu4p7Hq/Gtnsew1jsRBFw27zb32XWI8ZZZqEEgKPNriPcFzG1kh0dqDuLuW
6hW2HS/Cnx87/PouUlXvFt1LDPzmFvl8ymI9nA2Kkp8WG6sZWdOi8XNNdUkke8nled4IiM7r4FYg
rcaYg2Q8O0Ogv5f8SzitXNiOHeg/VUg9gPOIhVSzizuAxgl1/QZeUzYpSyF++UNZeToICkDP+aDF
JUb152JI/jKEHTkf1B5bhLea6PZsQ7U+URiEH+YxTrTrvrTwzD3hShxMkua96xT6CCEA0Ukw/MR6
6Q+Jo3ilkw/VGuLV0LE/KPat7JcArVT7ziOseyto+sADUGQWmwOw8pll/ji+kj+7xLLy9RS40IpU
Yn6kQ+evOuJrGb3NrwUnuMv4PudwxsLj+apTSjkJVuTO9q7++OyutqtSp4OMQ+UZ/LKeFw0gckJ7
6Q5PWMFkpXLwWVMKBEC2U8cnO+jXeLoQy5RHogzejRV+G6hxtkUAybBIDTzTVbKZzHzdIrfteuYx
T6HcknbRYZRAd3eJtHW3RLEdZT5wXrmVNaHzV7XNvKaNwSuGa1gQx/d5Gg/GSC59lmr0rRUHo1On
b28To9+3DG21xPfjamBatC21AoeJjzs+g0QkmJtoBulWyuUF0a1fGyKcN4H0D+Ya81nDr4xbi7uf
UiJYhJxf/gyN7pJ+sY5onpFZpjlVOYoFZzvAEOXa36Hh+61v2sE7eqvZxqey3uZSzaV5smGYSAEr
VhjyuHMz+HO6l0qbqb4OimUg/OhPWFYPRXGCMQHaaOXxJ+GKsg5vdAyq93h8Yr6ld2RGC9GRh/8z
NTiGPOD+Gg3zXnnz68/6qB9odkFnxmU+zJqYA0i+zyg1m9whJcBiuDXLrOhIzQZYfaRVuyisxNO6
ENAEyAmdn5rrh7kW0uY/mhCydp2Y/XPDW1ugLypPG/fsggwngpQQ4Y985e0OjmynYopMJUBC5xVp
tsXnjJTPt+dblcezQIWASdFn8PRKT4xNwogAmS6lDc5t8iCXso4VGHEDdjsd4MBEbSEiqFXEXUEe
igA16+6P6AjZrhBzyPKffQSeP7rhaNGU4n7H+bOppNL5yur6ReDxYQ94FNmjWr+Kuy9XnufmDxEE
nJZvOJPpnmqO+g96VWHyH2+sf+YhvL/yydOEEbMbHszU2Mo/0+DMXrbQ++1djYH0+5SeNj+lRmeD
n2WkjpkkkVohliIW7SUVZlyGp8gBwTz2L36d42PSsaSOR4yir1U2G645ndCmTO+AKuqgX+aDKXay
yXoIYWGd0dp3kzYB+YypQNA6do+2ZgA52T5cmcN37xdopuCGtzJVY4QhKwyluV1oWydDjwKO8A2j
42WJBfvXvOUZyPHsTuMFo/hnVKlCKvxKcqrdKqQO5wDv+lwPjRbbpuFMy37dv9daAdMjVOk+1LzI
mZCTCDtY9m6myNLazpEdTrYe1flllmmp9iDEhbz//dZ9Z21vDf2wzaiTd0blLTRqNv8sfbCjrXbp
daF7y2ntvUAqJdYli7qftByOk0SBPfABQJjNKqYWC42wtZ7AG8okgRun58LptGPIKl3/yAzUXdB5
8rylWfolTaej8W+NjwwrL9e27u6fmWPuMcoJ7FHiKgMwrnTanMEkEFt5kKluz0JH33xuuaMno2jP
/9JU/HfeOder53ZPYN9tcGQr4yGeepu8emWJWFUl4Eais626iiSQUSmBR1vqZzgOk6kr59rIQQ2Z
fWu/wuHFKpOfb4iNOEwfmabhFV7WnCKBhEte8MWIRUqAK7/NkWxPlDoBRve6vxBf51vZv6sDxmEW
cm4WDB/l4nVdZFGEfaPtV7GXlfbmPjklnxVWzZyRpMY2kCUjoFULkJUVGn6B/3In7vi9THkNuOll
z8f29SUaq6isChYqj8Hxo+TTsEPm0n2M4/rpHQmvJHJUqgNdWIoWj4y2rw+CkQquX5rrDtuXebFh
bhLDC6+5vGQdtFPLTvqUv6AhPC38SgkzhIf4/4x2fUijYlyO+/TaPb/ouX+twogS6HnHlN0R0Yq2
TNysTSR5mp7K4CgL9r7YhidVAoYnyZ9JhKe4DnisE+TSxV2PItX9+K5WwaGmAgBLE91gxesZ5bPw
JGySxagTTRChs0uybv1NuaXdmPwS6HS6Y0cM3VNSPV1YeE1W4ZVe0+12zW2uC3agdDZjX40zxjMF
5tVKZuHyIHsPcBp6WyTS2eInyzGtrQwL+WT/EItMXImA9Giy5t24gY3eWJpCQGwLNw3KXpn1CXrF
GxGw7OqNyxX/53WYfu2iRCcooCBZ6HuAsCqIPsQ4xDkPNfTUBhj/s7Ys1z6JTQEtoHDzriQZRtpZ
DscV5O0a6eqjyO3DInn31CclvC03P1c6zPJTGIW1k9uAeD2VkQC7HX8Zfc801nBOvWJYWl4Z9vZs
SrCt9UD0iWNg4N5BVDLjPSMJh1rfsgVfROzPzcRL9IT1XpAbf/oIEUgoR6dykIhYrUkJmtVzHUMR
qTDSVLwfrxKjCHubacUQlwCLNUQ+fDlPyEfYq9rNsqgQSaKPkQEoOmS35VeqttSdIqNM6/twWmvb
snMwrHrZ8kOkz5jBLY5fPzEV+i+fc3IApnvPnBRetN+nFc5uc+VVRE0ABawS+66bgRWZk4wgdOZF
ckVdqRNX8Y1a5F9viUBlYqvNzDX935luQ5HghO3f+wK4s+pB9QYcXjv7wCLTcT5tVW4C1A4GkzCm
DTIOoiYQgqMi7H/AMiaXDs9SACZ4DOyT8hQkoXGx8LCA8Os6uT0nh+EvnuPBasZe6y9rVKXvbllZ
D7m23NiO8oE35Y+q0kpKJOk9P2vX6kwUtKkuZjcJrtQxZLXxArUrCUmSGUaoNTiRuBXzWiymHZWM
qPHZLO0iyVqmoOYuY2s6v5phVkuH9BUS0gT+zgwUOPw5fkZYn65g4ReRusUUC0gzgEn0NwfXWbCC
TR7mCVP+oEHXjpPMhGddhsnecLjpllXE/3HcxYoFDeUPSAi4UURFK4oC9l6Ups67v87YZbkgKppR
+3jlSREWYXHiWe7svjEUfwYm/+RmAyVxlVcMQ6bqABaXmMdvlG/gxVj1/4b436FMTOczLOUFU89c
tQABTw5Y74PEJHKtJyL3OoBaw1fyNTi0PNxpVxCN+CE3JPl3a1cnbrDTsw/TfOeaelgPSdh7WlRu
Mn/PEUdPWhkHEh0eK/g0fsxUzW9qTdBQK/kyB653g50Xnpz3uM0biNatiDc6n2QUSQ9TERVpYYZS
9W9942aHC0vWZGXRXcP2lLuHGAC3YGolrD8+bLI47nRBGFWQwSqVO1fLxgOUT0mFLwE1eCZFY0kd
OwDa62Dq1T+Ry//8jc3GbzKSBFvznZwUw96PduigWkllsP4bQJDKSChPe2XiUDd2NdnwR5v4swvu
sP4VcGbGb7cRaAzitvCAvdw8pjNmCtiwZZKvGxIl0EPqySP5EWuj+3XO9xYdCeRddqJLPuR4Hj1G
PCUe+UvMlEAw+kbfhpbwbIdpx1FlrktqTNgfImXOLX44bxXsEa3zJFbj28b1yqIntsusjx0SoaI3
aaIbTVay4q60+CqQG6LqOqEOJDAEEBH25Fbq6CIwXVmfAQBJg6uVdWNBTHO24D8C/19N+k7J5gyS
Qn+neWNHotECjab9W7jGYKLhTTlBXdAs4NHIfljMMyAb9YFEl3uHvL2GzQcqGrrQKo7vjdLyfFFn
tTvy5A+SYF4oiq+8XLOmLaH/DBgtgj5trXoqAKvpV+5ljZASMEM303+y/LSdPrUk233FKFZBYTH+
1QVsK1CKJJ11c7NKgg10IHeKomR+167A4CL7ec9xI0nlk2MWudH0x20360RvaOgi7xfCkDGjIbGQ
sOfCpJe2obVEhlOd7d/h2kS5JX7hdGan1VvHmsdnFbXR8jRUOrM0mTc/X9J/WCzxMZiZUwGCdHwD
htYHXmOV1bKTEeyKStPSqtpJs3SPaaYnurxQmcdcfp0V3yYDuSs7JvU2RLN3e05Xsr0Hmh9cLcsr
YvAw0fDBh5bsev7L5Bm+h0Sj/TjCyodjAmIDz237DfrzpiK0dFd85VbmACt5XlvBNA7tj82P1Duh
O9QOS9GSRL+fazgsCv03IWQciO9LSsfnc30PEKsWm6Qu1sfKpFpGeayzXeh6ZlMEP0vqHgzInejT
ulPfk1P97ytOl3u0AkcNbQQOAa2IB7hrNVABKFBbp7grAaWRQ8tSpuTzrUMsrjJ5bU2seok/z4aF
5AAvzPixc5LxK/E4lmiDktZIa2liWWC1AYSx83IYcWEsypdjPDwGtwYZDnbnNcRt4QKZvPeLQavr
I4SzxnZ38z+ZPAhlx26h8wEccLzdvlSgXdpVzfSJDTHDDdHDSgzoZP2rAizhMhUzHGjPf3LHmIB7
xDUhgFKxpSwLjgEsozhn3nGhBHoyC12wJumByO+4fphw1A0P+t8Cjv9XusbVzkd5LPQUemvOaB2j
KH9HWi7KfGRi4NlijcopKKZ57EZ58XZd0xG+e9YwhXIN1CB1Z/WgwrhTKMT7BivKoKEAp98yZ1Z7
GSpsmLXLIB8hMZ/pALrRAth+F6V+TyOly1zGqeTz3tU0+55knMP5ejGHb8D+t7m8yyVNoWMpL3th
oNUh4jtZLXLi/VaMlsuGVfg0LAuShBLM/7phuUghoUDbiguqTcwwI35MsyDy4QGjHiaPuUEik6JH
SIWdaZA/BR1J94YULWa9+J0odIy5pznw7tcKSOOHNr78KUEim64TXp4+oqea3A3vfsiX8zxwKuyB
cp+pKu4S1NfhIt3HHlUxBruf/9ftCCwTMFSGE9PGpAFI2zWrtPTZAmz6KLZYetFvs9Sogbb6dYrH
c13K+kl2IVkupdXxqExx1z70qAy6XUMacCmzK91jPD1vlrjgOYJCU0A4lxEZbLRS6rKjTRzrhK7e
5Z9pARPT5zoTSFW4ASrBaeT8i24/S7GkieLxmf5p+fNSDwJiitFHBePx1cGaVQen3fT3axkEbkOB
q7wYcfcdQF2cT5kMCy0brHhny1LCrWVYtnooMmOPa+Qui/YIXeAhYM/4lmDvGiHao5bdOiKiREM9
CUikWMAlTqYBJSafh3VqrC0Xduqqm6F1jHBU9v0r+RlfY8xMW5tQlVIPkHyydYJ8aWsmBmV8PR6r
TaHYX22HEqeH2pNxwapS23uFmwMyL2j0oSkDYYxFHNRorzo0xhm78nHDLj+G/wIujwPC2ZwXH4NX
a0wsAow3Up5rQu5wEsjz5Rp2RwFUCtHdOm+Oj6vawHV/qqJXybVaugziboMbx10WGcaASz3F+2ou
GQSpTEsn33BR8CESMRPpEJ0IoBN6tDhBQR7oEZdDjmNgZRi9HsWR0ulIlqtFTrCzJPL3TUhc0B5Z
uZaOEat8Kpsy1yWKk/Du1tMuEIwsAHQZOVMb2YfA6sN8BjhWtcFPwCLiWKxt8DqvbACoxY45rrtx
LCgtzeLn9dV1DAsXMXPOIzWUyEnCEDk3o7ukIzZ1nkFyJuFByDcHe0sOh8N0dI0sU/jM2ImAvTbu
v0oYh44ZWjoQxeVTJ2kJ+lJgl3o5sKnY/HTXD/6Y2oVeztjneRnLnP91DhJ/TRfsEokbnJ3IuJYP
sWwckMIDLs46RsEACSd9AJxxvNPnInGbDXT+ZwgOex+EVNowtQHZw3RFVFf7rP9dSvMhWiwbRuFM
oVNQCDhVJ52ihXNM+f8gKpO5RVQ+VNbDDiYrOun2kVHH6NlSls2IGAYlnUMzBmQeMo8W7FAfYgci
KgmyI9KmYkXa64+wfezHIE2/05VAVv+vBUfPRxsgBaY6Sl5eQOjWE4Q5F19Z6m2PV0WGQRNJaz8z
wi+GF6c1htkVj76GvN2E/2fTG0fQDIoAMH5xEvoAUDKI+WnLLQitZtEevuhYfiOnjZ52JkKmCYjt
gNyCufR72ez8PrO+C4DnUivSbjiwgQyRmsvO+H+FiIzKNVDi3pqMoJOypvws4HZh6yav9CF09lbf
JexdPwl2jQhiCcOuKgs+oTk/XbChEorOu69/Se1SYt50IJYfBcG7/FmqiMFs1YNmdTtvG5IZw2W3
mb2SL/6sdWTBS/dc2aPw89R4D9LtSrT1idVvElGKF0iXs7/VqN/hQM/WSjbRPwqBdsECDdG9MbpN
6bUCT3PIvHYVslnmUQryY4a/LRaLmvO5vvTUxuei1GhMNQU8iSKNQ1N2ldvYrXTEViZe7xabdWFQ
5Z0Ogxvmb+LMyIPwZA1SYTWeIVtHpKjSvt06C0oe5yiHmJPVRT5SgKJz3fGGpBhLSLNJIUTw5gjc
1H3rPoPvtLTxiFbDm+w/+ThYHoSTN+EBtuSgnJ5+ScSA+FazHeKxe6KId2+oq1yodTnax5QxlWaB
BqcOUW4bp3cT3IX7qwE3wWDCiCVEBbJ1N9ApCyMf2SuYHukDGI0/CKgZCjfwxF5l9iDlwoS0WL7y
lkqpglWO7AQM/TgTcAlIjM4IvGXplM5OS8tK1U2jM/IghqWbQPnH7JeiwhAfSBbZGSPwiGxu11D9
vTRT08WpEHxProYxNh/exMAjSrTaRyX8XoFnc1D0OzPD5xhKYVuLTTEUzrghefnGDrfwC0I4KHKC
sQeN/XT4CilnOvhmrhFcXBXgKzDAOQZTDa63yDb/I0mMji26z7kN6+/waZ6wbfkObJQ2ju1VJ1jT
2DQ8qA7yoWtvMI11JGzU+W9AtWz+i/+gVcRmrwVskS1phfBomkGkvMEoRRD0M14M3A3y8QhEoyzs
xugGea5l4yE9pi/Huhg2Rhp6hixgYce34r8AYPX6YRThle8i/YRXC3ta6ZwiL+OQQ8fdbVTG6QZR
8Tmbt4W7egURrfncD29rNnMZ8I1PAj/59GF2oKIVSggQ5VR87gLx09Rpm6pzSZLRHC1mggFJu5dc
ZQFmYw5Gdd4ULdHOypTl6pncSvFAe0iFeWMQsOGyK8IUUe6YdN2FUaMctZH0xLDk5JRUuazkFsWh
m8vvcUKgatADsAMuNB9TYjn0J3Mehj78Biwq9KfO5oaVle6ItCZ8CIE7aJu/S7v3PLyUS37nWCQr
HYjoshCjDEl1AMkluK+ALtUxnSCiEFFgRrZnOcfD2YdX3q118wBJGTzXyQJBiV9Hw6KyOgMrWa7u
bG1VX8fS+xWaNZJAQjS7c7cJ2lpiILki2c7to3yoPlfiuhNxVo1GKplg0ZZJpCZotlUT4J/eb0d1
nUa/WM9HpFQUIu0869TqExqIh1jqd09F3jrefd9Beg7UHjy211ZNf8z/AIUJiF3fHS1Xk/VDWR/i
2Z4cvzIc9sTiPe3laMC2qcSkB9ZpNcQ+g4Gr9FDsXKX0MtVlYl3ByKqGA8q0T2aD5q4UQvOs1q7s
OBfky5wxcyKxuTE1Dt0n2YNwQWxeaAMT00jTv577w6jvEnoeGXjPms54emvQhp+ErWD+Njo2zPmi
rRMGenhxQxcNF7+C+KnEr66RwrLk/Lj+5aaGLoUR3o00sBCoE+dXP4ZzwDua1dx/42/Z7D7M8R4/
z51ftTOJlgvLK+jr6CdBvTlHdJEQ0kFKFmm+k1tEvi3CW9oVnBdguL4x83RSzis9voyp14OkDoNl
LbxepslHf2OlZJWobQfs1Z0BnOeEkKOqKHcX8lpEzCND5ZiewJerVreM4qiyzbpcPm43Ur+eLVHf
AHZe2w8YodeAsKc1V7HsPQBZbKfFyd4UJ0slXKekRRURdq4v3pX0MgC0licZy0YOTyOnt73LfrwR
3WjrcUGsihFpURYsO7IVGbxtulcw81OR4MbXZCNHSkVejN1cJjjBid8uY0byLoy5F3YA7VVH7ROF
7DuMpnXAswPjqnv8s5mECROz9G1ZgKhwneDJPKgkWatTFvTaUcnmZzQAkoGOjc1768MwRMMgSQ92
3/JVMvHBFV84HyAjR5SRGrSvoSSYqlPTRlnMibGjCjwXzdxkmq10uTBXKPYaIoOhXB/i3TdBP3eb
BPz31IIeLZ/oWgfcaDcRwlwEGkNHdmnVA6raUy3vD8++K36LOwYfX5tyJJsiKb1wJFixzYZundoC
QdnHFElOZWbezja+cfnSJ61uiI9Bs8gVMmjdTi2uKA8Kr9JqDI/gXvDh7tHj4khsbDHb+fI9siSI
1KcgwXBrptEb9IGJZx0OPUj/gCrYk+DqgiWBPq1b3h0q6KBhk4jWrOcn+hfM1dAsckJHNYEg35jv
X+BEzL9Dit8tOnm/3Ooi2HrIM/tPInKN09Df7cIiPzSd0Inj+B9x3aEIoiE8T6uQhs/HK6k5TN9y
mLXqn6YjDtg9RqPMvfQp4D153S/PoIuJxH48g5rTLwriJRk86iW0tVrI70WV3lUbHU0kZrTRIhbR
tvKtMiPaTO818RbKowGUUP7f0TVlrYCjgRFdHwziNgQmNaTXrJXo1rc1QvYbL2u+BG9U0Ox+GTV1
jhLVUYR41tHXxClJ/aTvF/jj7mi6Ijg4rhshCo6x9mOTz5H7MmnSXybMJc4/P+TgXT9MoE2tezLo
TF4uUrK1CwzHnJKKQigVxVFdUWnfuOQO10HT9wLwdPbdVU0gfU+PLyPbm9AkVN+2lKsHWLVipKgB
50WbskN3c5IqFOCa99U7tXpYZROohPnz7h0UPxwVofd6tmfS8iGrL/lIo3qWTv/JjF1P/URnGIsT
VhBYq36qDuZfd0TU6v1t7PANt488D2+96nQ3oO5OY381WH21WpStpVcvItyEPmqg0h+ZLLBv5cNY
eu1qg96VFxGtd6Z5M8rRWFsSdoLFO8LIfcvOPHuZHyTbSDDdFbNhMyka2YExZydYcOnCpcbVgEYG
okWX1NYoTvACJIEClnRJTr/iI3WsUegv5FxV39GWXUjfu1qVOhOHxcPqIfNlQOMuWV9oDevGDGXn
zNyW2S3fzCkaotsxmgjuhcWyk4KnbKAYLwOHq704prJ/DyNmXUmFhZXnZ+D/0vreb75enmjryvOf
N3UfnApQqUEToSBE3fJ7LLcAA7zJRpunj2XeSHE+Ty1lobO0Bq2ek+d3icXIt/S9s9+jJyAbnyTB
v89JG4uEjjbNSklE7oMb3cawo++vZmfsayjiq235p5UCe6IQ6798u5QLUX/lke2dRMaHfXcqJz0P
uwfk0Ozp54Ow+hRuZSAl+kGZEv8sVF8Awv4UrHIXZyO09k2yeSUzT5WiDoiyjc84QgDaNLGZXh6b
0xMmzRkfeha4g0qx9JAEpm/CcW7We1cvyfq4eZacIueEo/KFU/RBCTddK4KEXBZmzmbSlo4MAD78
x34keSWAM94+I41JHdoM1dIAS9vJ86mrtXeG6Vpk5Epsdh5J39upGUBlj/M3pdHMT3WsOuy3P+u4
RBMPfbAi+Oa4Y9yZGZCp7veFZQJdyc5bIuMWy2G4Qg53MuazOBCSYcqnhR92G9N2QSkRT33Ud8zl
CUSoAhr4nF7C48a3Aj3VdA9WT64HFtgpsgYGaRkh3+yUExrklVi7CVrYpQwbNANYbKkGhgTY78Fm
H2nvZBkIwyQkWARLPfRSyFbQJcI97iqjt16/NEYdcqwNgijCQYiK7qTVLafD5Ti22+P/XS6pIw03
MxkzJTNHPyYSnrKclxNJZY9LLhIE5jw6nF6eOmCrX3MDXufiL6p8Le7AuHQjEZGz4KUS+LqADKGx
wEpqUZBwkOmv1ulGCPS9t0fbWc5NbVCCFAm48glvRvBOu0qg3p6mhemoZzJcMZdlST8GqppT9L6O
Sc1XjuGW0pNgrB+oJa4fxOPw6a7CsIkV06TdjAJXINiBRabM2r4tpzFtpvH2uwODZNEnbKYFjP6d
IyMqNXIYXeVW0M8RqcWhDmR1M/cZVTO9vlkZNrSB+LHLsXi5tB0iGDdnWsddz7ppPsanzazbFlPN
GUHnXJ8Nj3mApVp8W7ERzh7kjPsm+NDZ48tjL42YFkbssji+DvyUwxhQq/39XFqrUz9puQC/BeKf
b2hBsrj88oNGEm/u6Q3LSXtmtRZnUFuVlwkkBR0np3ah88SRRqduF3D9ElW5p0pa7iEJyRW18IGx
HGMDenrmcQRIFjFVIditiqf3DSm7Uk5//VcOV44X5/CyfHfiDQ5DhHIZh8x2Zm2dYLPuxrWREcUU
LLIZ0RpVWHPoEB2bberF7xC53n3aFSkpgQjknor2smFcQeOqCZAFg+1ms+IN/FZscrmtQn91eB3B
dsC/nRdVxncbQdZAEjn5zJoudajq/5bRTRjkfN7usx5aD2ZwGlcZRV2QEORHkwmhuuCFMgGOJnWc
atj1AUYCIbn2WU2yZVFM4XxJZKI0fDmgd4Gs6rIy2iZmyWsS2gwbN+Gzequ8idnO6wvWCM5WlhlU
V7e6cSh/IULdQrl2pS+6bG/iBD0Rs2f9eqzEZaC76CHGAOhewpi4xM6xqK/fkmiqNiViG93aModD
90LvX0Q9ALi+yZRLqyqeSqJnL0tKTS9lRYUEnpgnKwlbraHyIquCwrsak7IKFwLN+3fhWchzgd0c
xVGVTCqWHPvmz4sU+XW/ZwN2aZJjnIe8mX2NC9s2pMsWdM3sO8PDJrvGeuw5JhJFwQ5OFcSvCfyT
2BKZZIaibQOnnUV5oeRpXJw+dkBlpNwRb+LLZm9hWrUftyq9w6WFVnaoPWK7HDLLUgiMikd27Z+I
rdHjNhC2AGqj6lyrd+kikgQJy0MceE7+MJYReTihQg43eHZopbSmeL1ydXVgZiY8sp6dYhp5kgpY
z59mOxBzIlD0IPw0MdvAFLwIo4y1a7g4hBGYrG8UeN5KOVU7C1ft+MuWYi9v97lw4DUzWguwXDIS
7FlD5tBManpyI85PG8Tg4NzdbxzK98YUlZHIbyqxNFVbd6aVfXQHEFrSyBNkyKjWJSJnUsfobOkO
GCv2oAjxl87vm5S1uWWEKtQN1U6y580Bhm4yKG1PjOhgE6luVYBoKek35IPsz/SxHvvSJbGKfACq
CCe2A6cb6voJ7PnkfnjTvrZMdWfL8ylvfuv/U5ifArkXRzavCSJ0OAcXW4j2eq4C1+WIHFK8zeTP
TbLM0PU5Wt5Vx2+LmLWXFKlTxmgj0wC0h1ekFsJ67p491dgXs+XhOaJY9XLeyZLRkcymrzJQWDWm
xq1ZIEnO0fX2yZmdENVuVn/BzYvrNK2OlwO/DbT+tPL5bHCsBlQBjma5bJX+6MUeNWEjqPyhR/uT
fTPN2wmu/O3n/bcmU5DTUvIZwf+zWTGDLhI/sOsk+9nIJ9Up5IdhLHOjlPKxON6Z7GK6BkRJ5WU2
35CX5fYLwSEPvs8aZd1813shmZN1y0ZtPG72MaDFAm/KZ7Nzm6LXWiezosqwIVOl5HOTtUIZu50b
NIq2xIb7duz6O396ofORlixsxPYLNMJdTx0UcjU8gFfJr6SG4cJL84GPQjmaJhQMTJ+e3TJ4wBoU
wZ4DNPBjXbIJShseP+daRAj3kT5QNr+xXxyL53mZF146poPRyssL6f/unznKm9FDK9LerzkPLB9X
0s9DhaE3rQWBvwJ7IUAYDNO9xmbYgn9i0wpzgLjcfOsJ8s9O+X7cuHx5c42lJnji6YYVyoTDjE0T
/U8bgoIaUxQ8BxNwTtZaSHuebs6LEKEW1wwCibkJmDuLgaKfAKNedvUg7rIHSptQjk6P9XTSBhlt
L21pYbiiPgpyO3AxxmDi49nMVI9MNXMsCaaJOyC9sgVbdh1gDL8iFGr8piegM4JUyftUngULMEIj
FfZEfG932x/NheHUB5daFK8GucpAsaYcfn1aZDlXgz/kykK8fAmULzwYcOx297RaoIKervuDYMwA
KWtIRyPRhBTB8jgvdqWdZR/mdOW0T7MCv6UammvhostUccquKsehPQRvq5aEIuu9B8ylHgh0Wa7o
DZa6tIzPD1GmyexVe9o2QP0b6X0+9j5UI3GwRJ/puYr5t5jTVsWuhk6XJ6LFZz/PAxmQqGvGYcW9
Mp+BwOIthcANreo+Ca45BMHSbx/mXFk31O/IrDBPo+u9ikZYkLWMhkr1TE1bMRwLlG4cnb2+bhr9
3Nog+GZJVnHNNAAzZlMZczTjeRTh9JAWWuaq9gr92M+1xNb/wGXPCCQgg9aMOeyLKxUPBOsBaja5
/penzGTac0FFqAgdrMQVCgdGm0APUkMk0zoouNbBb3TD3QGjebIJ3TDFtX0NSp1CaSINBgXEnJ9T
KEbv0OBJBjqwyNTVnhD3FwA4B/jpIuaTeA1UomzYblosUjLnkU7khHgbmhOOWfxr7xWmgGLjySH+
VKdi/u13U4jNUmikEMAlb2tZma97X9H0ZovKo58mGw2kdyUBVz+wlVB940grS7dI4zZ5+ymc0uAN
AQL8PINg6Rd7nZ01stv8bFyAjfp74661LgCWH2oS1i/jgZh52We+DjVtlmZ029BiVzD62i2e3Q0A
9BUti62DvVgTHQrZk9lHeT6ubCWhWDJISScPWiW6pDAEBAsvAZMv5UqGONiDI4I9UzuYDtpBpedY
9IcmxTUkd+AG1rBJ9KVgQTu8CDMl58O5T+XejR8Zhbyj+uFwdRs4+YSyUfV78N+6X1N0WTA1xiSx
7oXewlDG0Mq0Y4J+i5QNTharvbRowlzA40QqZCLq+YhJU+5y/eqiWXNdf0hNRJ1DwXWofQuLJepP
9YF3tbIHa02Y7NIKEWaXDyiZi3OUREAJxY6x/zFFxeRnYdj7A+Znq0f6+15x3YAGpyR/DYAI0IAg
nOpsgtTLCkGJ/ji6gZViTJCBmFWb+e1V6FH00HZ7xdyMDb885HegH4YDerVDjDEyUzZVpJDFykDO
EDwO9U8xBBIcIhHNzi9ZEjuPwhu1+79+ZlOJ5RvkyBW9k4CoEl3RRnMpGZ7OR+ykCebv0Nd7MVr0
4j+itx5Y166a9oQeHWvoZGwub3MGyEpFrZ6xWTtZVIP3OCZfFYLzNyByI2PocB+vln1KbOjwQLxJ
q4/uMLiFEHcMeuCRpqdGw3cCdHVn9zGSzCgTz1R+MhAhty+vfSfgMrfoS5R8fFmGrdqsn3gN/pjE
NB283PJm91MXVpn/gklUKu+e9DJV8E7Wc6i9+apm2oTEcOrjI1gcDFU5twPrDv2TBI3rbjTetj9L
rnbIJRl3YzVxAp577IoON2RaMUpjfWgHuGdmoXHJLJGzb2rtEjTnE6buWVUoZXWpYK0/ZTb/c7q/
VMruLEjyxg0O8v6rJp1Am3EKajsCAGBrnXoWUEbhvIRhv609xFC3jh/VnYSEsywOFl2QMxHuKAMj
lD4i9UG/yj+xcmR27priYO8kEbMhPcYgfEjCkb/rRNOlkbxVdG5D9b323rNtnOurCPuX65bXaPDT
ssVpO1C+U6B+nRDtwFFHVzbdushvPsLfd4ZUzmCswj4yCgPJ12VuosfiHIfYw2u7ng/6Bu626Hnb
/qJWncXfNzNeJDrU2y1d7zrZHd6m0pnz/RiIYzVgNijrWopZll+/48W3ooi9//Rv6+mZCSLbz4cG
i+frIFqGSkMyKCkbdBddGvh+0o5+M/BDh0bVKOEbSZeTi8zOAoQXy9cDcT24fF6fh0Z8YXkAIeSr
L9eytoQi9I8IQxzmqjop4VmztnuS5HHSVnpJcbScGz6LhPjAvMyu45nh/iEIUBPR7G7f+zHhCktG
QDU70VwPcm8KRTyrP95nxF8lbwol6/3Q+fFyg1x9eYehqQB3yw9lZVJVU8j9Gahz6/doDfixXkCr
ooeWbo5WpQz34n3Ttb7DjvD9ZxVFNacODWppIWSvUlmIHUxRDTGCQJnUPBbZ8+wICmwsf5AbXQqu
8GU/1veFFel7oFq/hUIAib/3XFhTFFYTs0Ke4ZVseZ8KUf8xagOuGIlL3sYuJaXPwnNDhyuXgdxC
XYnljSkvUDcpyKikMFjTR6xHOTLHSA8rMf7WyT73wUTyFjdni7CsbtzrXnX2uxoBO8EWIpdzPk/4
T4uovUyJUtX3aIOJXx/nVd5Y1f8Gw9DoRHnspsU/T94rbc7+wELMLiAEbGOH2r9Uz9Er00bCR50s
KJ/LheXEVPPZQx84fFvGTLPhX3UDuuhioqjcXBRUEMerrVk26dEw+oms8VayiI4V7KpmP0+HF/ze
ZQe44h6fz4AuGkKRNTkNVvHnQxejjLwl+6dutAKp/F8mEOsGpgZaEaXvu/OnHoTo1q3drvt38pU0
g8Xm3oGqyp9tJieRPS/h/7yE3aleavF0Eyrb4GbDRYaKNeN2Jk64C6QnpcyM31veRoNba+FHJ1KT
e6h0lTkqM7+okwK14zecDoUYty7ve/zSPPdp6kKwzhIq67UhEYSp51Lw+bXmzj8CwsbqHGN2MHVJ
qFt2LPmjfO1ylr2nqm4SkrIkd90zqwvAxGX6tHR/4B293DgQYdE1GCqNYMb35SukbaQ+NlrQXq7U
IJ0lSMjipIvua5xAzJswWwRidWi+vSQJFrxtEBTG7dZPeSKGsDSrfaX2JoetiVPHjsuzigEq47yL
OrGAzku6Zj3c3XMPNmfZT0094GnTf+mXBPiELwvW3XbsccKaJAMcxKnOwVJrzyWLe0V7DeQLd9h6
FBctqks5rxPwWv74kFRPhB6oskZQfk9XhbDBKNt4p6QXJa0uKLw1knKI1P6NZzUvTmgSTHeMIisB
d2KlA7AhkkgH97jlf6jXPdAg71z2s2rfM4h8J+JrCVMKaieH1QgQoScQ3KXh0wNTAijdBNTaqAYg
BxV4AzjuTTQG7DGEuEjhIs8EoAh5T5R3vKBixV96Lacb2GaiRsXDsOI0QJ8peAqJcgx66s7I5052
zyX/dDY95YfEBYEfILVRbAFRo/iiIgmNbJJxmJOeQqxmQsN8QZj/ZpBn8FGiYpLmhDdg6gepiyHZ
1uTFxnwi7Yykq7GcSSI4ZasnzR+rp/Hgusm/f2aUdPkgcaq3hDEQYcOhRmxJFEuW66p8sJtY39fy
Ruw5jbSgS29rxLJ9f3stGlQsNQhCf1xW+849+8afv3q6LWa0kjvWLCo2Eydsj4yp8SNN9aztAY97
I+WUiR0/3RuVheN/K4GqlG85e0ZQsE+p4hYls3FMe30hLQiWytmXXBv2GA8HowFnqEEubHQ0Wn32
eS2sUS1Ux9R7l8nzE9dNJIpW5BYA8FQX5dSRqt1TUZryBsqPRBgBsLAX4xgTVWD51JSWMCB3JqNQ
HHSxq3+bWPNQVvWWUu06UGWayMSShMsnQuxfmk6l27nIor2mJnv7x62NLXh/C7KOP8n2qoox9uUh
Lm1SOjrxkwXO+/84PcsBE53zVP98m0P1d+I5OBl957pphcVrZNGHOoE9sNA0c8qJXCksLxpb+UxY
nbGI1/FdbVo8VSbtwakQePmckaDkBFagttanfPYwT4ZVMYUCKxIIqtbaKcMjNpY1GKWAsNK/zUhh
VLxDXR1L5YQLh0/Rs0L7n9FXlVvBqGIBJdQxQ9N16/mKn8IDpPE5wT+z3g3VPqFJTrGJn7uCvieD
Oq7RaPcuW3M6pLxoz2zK19pitvlToQ7AJsXYY86aj7MPmgyfbnL/6k9pTaNknuoILKkMkc6+sZDr
N+1PasTlX5jAK5Hzh4UfVaUsKV+mFvAFWnZuaX0OzmktQBqB8W3KgsD8EjxAVsPXtvTAYu09080Q
0zns3tIsvNFGDrRYy0uc5ut5d3yfIEdhIHpjl32ZzJcVNao+0+dOL4T8Wimqz1t0Y+RxFQX3KX1y
xmHIG7rXF3yMHVB5otBx2O8B6v0/j8IlapUv4TcFl1RkN208+FSipJg4hLEKJGzqdoPhtE+Z6sN/
M/CywcG9/qs63neok+8uMT+V8IgnTADZVD6bPd/rpUREWqkylejxm+ADRLkW07nHSnY6GgZy0VE9
edgUsyK+oc90n4DW1vG6SGEuGuKApXo1xR6LHVxAnG0L1Cg/CVNvxOS44F+9FX9aRWeXvx5ZsgJX
bI64J1mEfuXYiv8xGT/X0Bd+dTXnY5yCWhztC4u/xP0Ml6ScFgU7B6hYfdYKhvl9u9/UMB+ZF31f
e4H7za5T8tRrJuWWp/t4TtbGpDZ2tDuKCucluIF2feClRZxzIY9HYBFsd+GfMBUSwxiZ/fXOy1s7
lvgrdGFDxhD11sKidyvbr2Itidzxealvgop2Lhg8mtrbZq1FCp4PEEkR8+pQflR7NorkDnx+W1Zq
hB8D6rta/UDT1OzlS5BUXvlrDDz/6PjAOHuCprij+vKhnitOBgD3Tirph8QkBpFFSt1Cntoo30+k
9YpfOR0zYeRrJKnuoCMKDJPfC7SuppPygISl7Bpw7QwcueO/9ybUQWTbO/DV14fG/4RQVXXDCCsZ
zFdIl3cPBH7zfoEA+agH6S+vyTVQn8UO5D7fmpOBkfjgz/IJvty/EFpWEI7Zw797SpbAbDjSFjJO
xx1A16TSg7aVuMZP41EDV/KTAmEuBe6+E4Y9VOqOFS+o9cgDvXrfP8X306WGO+Zqu9Ii1gCQILBS
I9E4WhfSeiep2RYSVnFPF4PCrfjthe9kP8e6/yaGjgokQJoNmVuqUiKwmOBmQ+CRv3H4pNu2cZ5H
7L1PUkXT+GcIJTpOF50ygeSONw08gFKTldd55P6kxotSDwVJMGgv+RH4op+NqaMQQW9DU1dvwZqn
lPcmM4sE893SlMgxBVg9VAzxyo09SP4gjqVYEc7KoAA0e6BIpGTCM4PF/GhwqbFfrLp5aRbMgrLn
jPZ4YT43COzHywm+KAr6liCF/o5rHCQJfcH954kKq97otQ8e3/dJqo43wcmus5TYJtymZ6gm3WkV
5HDIP33G2EisN4xyv70skKpe5UV/PJ5QQKvTuMLaimnz1LvaTDPekxgR1Ixb3St09sKvy4KrM6e7
JxXykMHYZLv6gtjqbmWeSuph+BgtrWNUHk2Uh8dGzuFOzMC0KG9vkE0brDU+vRZEvQDzWCFJtQGE
OxuIo0nrO5tYOUvBx7bdFJEABOqAIllQVFFkpTbw5J650G3E2a9+IJ0ib/zNy2nteSJ/pUqb6r6B
MC5Z7ZLlW3cpWfyTsKU4cvSJu3YCT12hM8htrO7nb1BK0lTW50Cbsl800UIRDRHW9WqUIXS3mg84
dgDsvTkdVsk9R2TXcZJVhc6pgC+MrkkCODIUwidAgd3saE9u9kEdRQ9VTs0pFirQivcjrSn+9wpN
ez02DEpPDE+a4WsTf/J3mVLk6Ce64GZ6QKWkK8V9uwly77btdixWYVT3Zwm3W2mNUOLeNEgWR+Bh
AIgLxkS8fheNDug7wit43RYMyUFQiNMg3IG0128svAXYDsMepFFCyj00EBCQpqMse8gdOOfT4vR/
yMTp0sepgEzzC47OCoenQwgTpOoaoNqOFCnYBOnZ4E8WlT7bogb8bP0R1wW6IZmcGrOa2RCjA6I5
g5y/GG1zzbO4Z7ivRop+UyD5FNqHGpLK+kwCwmt0duTrhtblFDnIh5fMaih7VEDW/M+ZKXHvCmJL
B5fB1zYryumfzomfnHPX/UKHKczz787zIufZ3V/wNALSOCa8u70+jJWivME8toV7EccwOv5ubhWe
S100UFgte6OQDdVANmXkzjvn9Koql6OQ1BjoqaBlT+nPAVVEx9IOTzo3QWgCnGCIsk2w9dVyzpPj
6FtyDpMzwFFXdytNe+VOBhwkc1h7Hl1eSNkKbB+zk87BO6wFKwwx1KyS5fpadyHCZ/yce/Dzrdo5
3CZ0sVPXpOaoEYnO/Ke+HCvOlvHoIoCvuSmlaPHeZ+gMSZqAiEmSKTqZgUd+C6FdCQwg66s6bpJt
aqe4gpo/q8VQWo2VCSlL4l+myFeAzAykE9hu+abqjOSXg9ID1Qwbmm8B8GQKILaCndgG6hoWkCED
uTEbGmPlmZ54GDsZc07NAgqukyZfszAzDcuQMZpfbFoGJr8lpK0V/e3p91iILO1NjMYL9IW9gfpd
radjY8oSyfknBvrVuHEfxmxzdeJqDuNNUXgodfR1qtQyItL3SDiYeUqQsnOJ4a/MZggZdeZ4BRXI
Rw7IE6kJAJqQ9aM0q63q8lccqKm3QAnlP/odVrw8rJc64U752grLC7RD1q8Q4S5v4kV1y2HNgLJb
x36IpVpV4AJy0vN43QyuC8FuSIlbEc6seMxq3E7V6lRwwh/4Hkp8fYEtdzbJmZ8qzDIkycjAdBGg
0NxgTgSDMOe32M95L8KVGULRpgSb+YMLvzcv4keVQTZzBD5+gjZwgJQgSgZWPq0sj5gIx/Is4GCu
87eYQgoe77vldJ7AOz3oUir3i+ltbijSSHeoK4CTHQgLHgMSVwZCmHTHDf1Vt1wVrQX+k68WG/wF
thBidUMLjvB4UN/WKnKPrnNjW6KqSsYJOfj1XaGMbkXQe6vf0G2Kr+rvgqMDNQD6oJtR1GHt2HnM
5pe7DpMGs+u7J3VejMKNVooaMFoX7sW51aq+rbWxkdGO8+HJEdJ3aDoCEJSmk7IooRZ/zTBz9Qq0
/VljAZfbpIXDBUR8J05hd/2f91ine6ICqdYgv6KYOYyVagRSLrrjv8xwqS+gmxyEMXXmZ0dK2U09
Z2j/seimeXyBx6tHLTXfhPBDhS2fP/93gXc8mj9XhVXtlJJVc5oKuAthmeYt5SfCxkcstvAgaQx2
3HUrOWEJCiHiFnyKH5WYyjUpW6EW3ky2IEBivEeji91Xh//3e02wY4bGWo1PnuaamZp0t00aBlyA
CongvfeUPy/npl3/95eZZuJaYnsS+OwXfK0rc6gCBnIOwOUvAMI9Olc/ED4AUj7jnrnhuhX5kekw
L2A7Xr3+addSalVxL5O2Xl3JrmIZPrdaU3RnxaK4U7ufUlV2S5gwfZ7/EaNt8YmshbwHSKYrjo5N
ir3fN8gFhX8lyGKeYTz1zREWOVGon9knTvIZ2ZGHlkzBK7m997uDGIn8zRS3T3UM0H6epG1mmO9s
WcpCbgBMdHz/Q8RpNrRMW+Ft/x8AagpSV4Os6pyo05aq49U2p2tjlSPDBG7Bx0QoS47YvYRfmHIG
HHh4nLcQI6SfWZOBb2coOeNXNkVZqtj5QmMF9DJI/7p0q6ACfjN5d7s9FkKorc7g61Ae5NLaw8i1
W041n/5poyLU279AaEXLDZ78VdeCBygc37z11rc4GeLwZgB3uF7x2QKXv4Yh9CLeT/uhutq0k4ko
j1RlI1/NRdGLuN+ooxg3zkG621fTlKU/Sa5Uumjd3F/IL9aQOmrxCcFA5rfHIRGJU0LNMl9CIYbe
eQaxKHsiN0RUhOEG31Cy+jHHkGdT/fmgeEKWDJKntGw2nmGi6Li7rCDltGNEtjppLIPeJ5FXSNbj
wHZCsrNCaieot/ErIEWU5S70SsqsB6sN6S5PyaJihsA9cIP/WC54OhkOmqZp9E9XWmUh4Se15A+b
VZltKycHoa2rZhb898SNjTn76WC6VtgEu5KjUPu9KuLUZDlWfv8KcMCDEkCyTJdnbClu3xv89fR0
YoYlDRHJAS4+eSHaFdvT6GOdewM5cLbnKKuBjimiIXzSPghtH/E4VjM6T9tWrgh+PL5TaL6f6mOb
4bEF1B5zt6eIu8zMt9kTjLCqchpT6FASfflzNWMmX08Qb9zaPku8KVXr0tvU9VNRmhuNMnfkZqd9
Rr05wQOV5tr5xCr0JQbNrE77F+UEUAXbV0CX+l9CoEYKqwElcZu7iiib7jaWpKBq+yD0ePpicToJ
q9s3dyTKcUGUU+GKnusVagCWhrVgsSLvlCvhXJp5/wK8BbbFWopGS7JB2ceI3S+Kw4Xa/F7+zst6
YRbMVGqTNp1lTAdM8ieQsKxn3U5pGXFY8PV/Czj0o4a3BZiAJBQrGu6j/CQQJHVtiMxITD9t34qE
cIUZpga0PGPsW0BX/mkckKFpH/fbeAkOyL+QEaRgrcC6ydyq1QI/ZCSs1MXaqn7NQOgZv901kUZI
NrLEpRC/7odYnbFAbD+xaxqRA3G1WRmP5W3Lu/BqXEKgVuak/QMP9rp7BqehmpcyzGpzR5rLEe8G
2oh3MevML9J6xEGi9GjNDkIC/6Wy5qx+3NNpEy+Rff3t6yiDfs8nljDPN1WT5gKMDtA4z3PpFSUy
T3GTDfdE6VVnxB1srMv3H7VSR2teEXfyXrfupB4Ucn1PjcQH0O3f/Xw7LKGJcK4dVS9usOkKEOEm
pMINrQ3N1YlS4Jy2V1VLcHf8ab14F/P2zai2Q7YP/zxNUUhZnXyt76mVEBYNVz3KOCbyXMUy7DG0
suhgwNLf3V7ib9jrTtXLahsfkUa9INvC+sg8nXDnuu/Jxkr0aB7iHmZZsqC1zuK7f+r8zbh1cgrQ
SFnmIdIqdBjFZiwYUjT+1TzVlp/U47u67e5d+Oz16wG97UeX9wO4chMgCsklS9Uryzg09wc3xbsF
7AJ/GK7Omky3cwyLnMI+GCLuXo69btP39PtenBudYh19AZYFkCC2hGLcqq43yde13D23+HeXgpvr
qBFP7hcsOzEpN9q1ajF5FdlUT5p5XLq0uj4wiS+OVAiRMr5S44UBnrMOvZQVwdBomwQGpGz4651T
D+OrDUNlLjwc54kuFQ9AlgS7T1Rs73EZxngM5evq4Cnxr+zfX6GjOa4VAi7OlsRXZGnvYMtwldKd
iMF7EUzJQwo2gHBE6fhQP3xJgvRGNaqYMHbBOzkpMzbjQtD78QcR/oExOdkwkQ0LSMJagyvULlju
/W63RLhTqk8O67EQ806SO/UjTKfUKQKhp+Qqe5tu41oPTv7xZP9UwXA9m9SLd4dbzdtUkQPdAzbj
RaoWcGVw+wR2a9yZWQN+jL6cukEFrXN4RPsV2Buv5fo+NgH06x9HDCx+jV3bpYUGbZcU2kvpnhRq
Th3K/Lk1gUWDSQt/DrDahz/sfWv6e7kWJ/aiFRHQGuzhZdqhZsVh88QdCQgNePqsxug3l2v58idH
4UISaeKJVklLlb/gBlm8IC3jEvwkWZOrx2V0EkDKCCwqFRgNp4lE0BaAtN39Q2Suh4QrCN1ulW3X
XUEhS2VPvaZEVf3I4T5FQLzEf1ejjHgeLslVBYZgzFC51Yd97bFGOixK27yfPVNLMWLel/BcQCVK
4tzAHpDAZhjW8oWK2OURvY8KHTf+ZLDDVphS14ZfrWUz2Ivfplzoz0Tyef5TKnsrYeBGu2YD537y
qnvDYCpe64E8fjIK3/SsSvxQ9mi9dc1TaJCWqRVHqFq1xQPJdKvjxpeDW558TXmwuypDbtDPp0g9
fn0MX7zzRullBcw7C9ctL2ec3Vxbspn874rqNgCDpLsk1miYJOD2yzxPhIr3rtFVq4iKiPUm7ZcN
GJyOs7+dX6z/PFpsXK6UxgP052mhm8boMnyYjXbY3IYKVgFPyJGKm+hqbEZsgiOfT5uTQX6XoiR8
Zpn6/9LvyAhQZFiVUq/qmib4bPQEWz3oOOL4OIKNTttCc/AtQa7V+VRKK7jFPBTV3Moi/KORh6dB
1Qt4FC2LoxZ5CddKXFUcJPchXRSuNz8yoQYIaZx/YAC8loK/8KghndVHwg6QIHOUlPhzbwbXTAu7
MuK0y/z21c3sLg/T/4xhYw9PduHKpjP4zIl0tU8Ndj7zYWOh2nlgKA9JWSaHn6QXgC+yY0Xlklye
z8C1kkPzfFY/qmhziar1oCv6YHaulLu/pI/geB+2ECJzcvHg3fw5L6TcHZPK53gx6WdWaRL5Ln3I
IJv+KqGDcGPqIw6BwxJJzd1zYceEildyerKelzD5RaqS3Y4fNRlCt5SvS/6ccMlAdWaPDiqhdxOi
6mSLbjCRGu5Kvc+vfBTwc+jf84Lt8O7GTU3auG1jIKTyC9qPFSMQsPwvJKzfdFR2w7NKLO3RKWry
94y16TECz7SIaNrpt9iGLkkIZsb5usNez0zo+QlIxjbKbr4/UfYM+aZPH1bPDfVGHVkREW8hKFdS
kRUubVhRYBnl8WJXNqp+K0wUn3F/880iLehkBxkFh9ooESUPIdZZCGomCS5SevznMjNB3nW7FiON
B9D5x4n5NFGT9kqv9rnLaAmIg2P3u9UiSqU5HiFj7tJ6YBS5kPVkWOE556C+Ju2sanrGC8BbIYqi
LjdevgubfyFbJOe7NS5F3h97nBLoAqnEGFRUlPEPmJpvwwHdJC441G9FeLjaFj3geuWR+bahXekn
HuvCn9WCJbvdeGUUiRaMwH2IjT7WMvwXiO6gciBy7STHbbrK4wBChFRDJmN5UbOgK8Jzo9oychaJ
fPHjNNGChIhDLd5JVescqRqh3ViMtvvPLV47BP9Jj8q6YLJdTvSU3eV+VohQ5n4lywMlD3588U5V
/BY5lQAcDEFqxek+hlXHOaxGfPAVQLwFr0C9tEeZtEdyHUzx1CPpkzpw1wky6SopFPk/zPGrZjC4
WT3/M2KDx1N7BzcJXhYQUsYpsKIsLZVQlIarQ/Zfp1NXfMvdswewh+LbnDmS6h7kfqaYTlPrwHhW
6SoRI1gnhyun71ZRVeZn6lO92TCLTne9jUOk19JapkcB5R/ld49u74jzIPBFHZchdJcXiyV9PRil
wBl/9nQTvXCDBa8PH6p+qbee9ftFoGxhUlElLjrp94CD4YdLIR+u34cIcjwxXZEvjFKy42FAdV8b
IcEQ4PyhHFzRLuqlUtdDTfbP9FWhy7KMaPX3qbQbtdLIxmkhfIVKKlRrQ6TekQmwB2xAPSt67+rP
4Vla4E0DpcP89+zknaa1THPUZYIY86WUPoJBEkHUkiIFCAJpek+ncZcieATTkg7eOCTtCfUSqMpX
UwNS26Pu6V7dXKtQEENHJ1gU/syYAr6wYFlaq3yhBdSn+WeyfyBt/k5HFbUqlv/HDn7XFJdYzpcl
XFVzOAFGMB1BYn+FcKPGEDxC681oPOpFJJO/S3TwG5mtTnA2exvg4Wnnf9ZTX9BfRBaa/szLaeef
eQq9u2YsnrsqsCQXjsEl4DNXKyakqj3S5w6R7a9fLE76Om+ypf4DV1AMtc4xxHsR+KCWALH6bcQb
utPOlCXDCazC2AISkqOD9RPe75d+Un/rZibtUodqz/puDgLx4k+qbe5Ft3NFXcAf0WI3UPJ7stnX
/CUg084iEmXQVCMBlroR0BiZa/NJQPvmrAQ48cqMFV6i+Tbw3dFfv5gcaj9l2t3ER9K+YBwcTlms
ffCU9V9PUJTGNsJvqpk2EgdxKeutnGA04peClzQqc5f7OPL2Xo0kuCgeJtEL3Xg8MlXYNTFBkcGC
8x/h4S/k9ttFno4y9VptjBvz8JNXzzv755psWqYweW+HdAftafZKrWqMImwqQs8Zd5rRaygyy0vQ
BSG+ZsHJG9JgaoIxzfEZos8TarI937wiPINhCKeV34evJOZooDA+NM2roLspBB/jJPlfJOeqfp3F
7JFC05Wx7IDIhRKvyvn1uHMV+Ud0LB1KLX/+b92LtMl9fm1HzKPgwLWGdh5PSQetxCyLRWumy5qa
YSQzVomS+eOkewZYK7/vk6MmoBdOY6L/INqBlbpo7uD4we4HluJt7qNMk9XFLuKuogrznDqG8atf
CAFGg2Qg8rFhiS0A4I8kys3X67yFoOGOCojG+M9Tr+NP3vtundF4+c4ndfGnZRmoYLR9jxOtHNrt
G7VPFuFYT1aZUv28jKRE2wob60wcxuZqDknvLaOg6Rff9ElUVWKWNu++SmfhxD7PCrwPu7Je6r5/
x9UyUdNwkqS3igqMkCDYTr+el0fLDyGR3/eJ5kM6p25SHwqIHVKsFfO+afLeGOrMD7KZx+kAkaHA
nIY9vBJ+hydR9Q3XDqW0D6KJ6EgN3F+SJqszfFf/VrdJNPOK5UixTaSgzeG/45VwUx2LG9sf6fHC
cKlQ44wloSLW1qAqXBjDrKSVW2ZXjhjS66z9Yv90EK5AX0CzXxBBFHTxz1NBSDxJPgokSNSkmRRT
hrsCIceLzn9JSA0ELyE5qzGaiWwJkAAi5COidaJt4QD5c1pjOTpRLsDYT9YXsGlwRKR3EN0Xhwln
a1P/3l6Pa82rxqIr2nFcD8CHd+6QLeV/cxRUgYAMDC8unRTmTW0BEyvX9bVKGuyUTeUHs77KHmC7
mltdnYTYOH7cVVv+Q3RAoBsL0EUjoSkHSs4Jk1KE+05eqR/yylqTaLpxdJ7/Ytzv4IAY+eAt9GIC
elgjSj6agJ6GdPl36ZkyFu28+99poWPbLryqJDQOWSvAi/W0wh58S2cZ+LdkylWC4uYI24q5INXd
Spb9CdiGjtU+vfiuboOf/5Ira7bIK7apZVlVIj0YL/ThDc2nK7WajyeBcvxWsESyfIvYIYJVK+ML
wy6ar91CevMBYPUlFAG/WWp2iNMANz5h+/nO++g8hWspE4nrTp/qs4QC2PDDzFG8jLgEsQ0YGbeZ
7oNMYDRaDac6wTvgP+54q+uKqUteJNnvFXhyrDCHVAXJussIdD9eNAC2ezTsqQzZ4CXhZOZMT74H
SBoYwqn23vklBNDXBPIXHuBIkzjuMzIsJ/nFwOe1rfFOS/4zP0O2cmwVMrejO7R2LyhcWXC+k/UG
NxG1BINiZ+XAu2kVSA4BeCSWYIub9iBAQv5Vj9xe/O9iD/7vThDcQzFpEMBXW3hxV56JPgtiSdJJ
AT5AL54C0DR6gyNwmcq+x8/b1GNbzU50pEEhcJHSOU/U/iQfJgfF2QIWZnHfu4XcTh3QAj00TWyW
5r5JYve7OswA64lPKs36/wL5M6UM3wOwpUq7YKoQZcfMZdegofrCce4Lkocn8+veocJ7e6Q6k+ak
smWGcjkaVGqRl7siniMjl2mHF7d1oC6j7j6fyimQ/V+0j3za/2wpROB421emXS5/JZtrKkPfnOKV
OiLoHAlKpYsCYjZaepJ0VtLW5qtxvCkFavl2YyUM7kA+MRKrL7sUrig83PgMIAt6xJdRkugNOYNf
fmEeeST4Wz6HujXQSfIrENGlAaA04Qwiz6Ewm826jPoh0hgLHBxhxRDShMlo7VkcTj+cO8pRrB9R
706ook5whKgtdIG3fXZBCWCjjIpK/NTzPsOSHy4mQhUftARpt/n8R31b46b0JGBG3vdbow2fFNud
yCI56w+Lft4PPQgk2HniQIXwJ/fxaAbGaQafQDPr4NZlb/V8cV4Hw1M7923b8tEPfDKrb2h+eqmN
My7wj8KeDR4T995Ob/8Wt1MoOgiZXyssJmKv2pF9+PpQopbIaLcOsJdsl1NhZ7jhLsRpVAFbdORX
iSp8M2UHG2UP0zu3ITTnaDrv7Vv1r+9P/eRlaAhCXuhmkI3n3YuUhgsOjYWvt5noftmFbmKvTAot
YWaPnGslYEpGFsHJL4uhLN7RrB0x/R6V/BE8UmOxsNqQPWPcBv8+4JBmuHkVnReJ0KTLSWkh6zKC
bw1Sdl4yYllj4p9YXFVluv3MAfdXDmoy5WJBpwW05O2JBIb1COddP0/tKL1jS9NBFsigpOIkDHAU
gdEI0aD5DXR5ikPuAipAybckF2nwzltIc2bq7NU5D3TN4Y/WwMoYuR7ldD1m5pKNFsPc7vBY20tx
B7xmgmAwOVWspo5Oh3pHsMhpJ71CI1IYblT5AZCwda7cpIQy45+CU39ZqvHurK/4saT4dlj6kCEr
CRtC9P4QjU4w84i3BBQMf2+cB5TeklrErE031zt3N1U3Y6NVi9rINQXcZfgqrv5tk3oVahcycJBe
2azxVpaTmjfl6YVlnbgpHd1Eb7QFQ6ubOe1K4IkY0e85IkABcNZz2EGVb1yifjqBdKFQ8Gu0LsHh
lVCwc8QHd8ANW6P4Ki0cZDYiUWeedb19TVp/Yt9d91WSbasI1VWALd21ujogpLiAglowKUsG9/w3
NqmF/Xm3sdxYns5a3Axecysv/yrZGcBo0n4e2APEmJ+1SXucFf2HHNVgpC/QD9wyGBFX70t6lXTj
ciVEBGaSEwf2Kt+jEo3evxViFnXcp0U239A6YSoL7KKzEOOWQlP45K/z+nOFG2gPQ3w/yF+6Iq+P
oKW5aKLYDjIuFx1ml/5S1M6dnWbydK7hm/I/f4HDtYKY5LlFzdfequUZtX4fCRFSmNA4RXGps7n0
du05vN78C75id8qLgcLkgkCT0MGvSlRImPNoFK/6p9EfzcQdfN/g/Ej/j16zsHyeeykKoI7/7h2x
c55lYz7BiV53a77mhJVT7yGGvhQht74Qb6yrf8ie9K2owQ+9p54AEt2LTW2gzyC8ZxsS3dtAcw1o
3On1HLkOAYRYo1e6Pgh6ZWa6TBDive10v6Ih9FNFjSCCAAyLFCs7X3wa3zz4DuA16FSQUlUGVzNZ
WNLbd0QR5S7U3fm3+MlLXKw1Ybe+DzjletZtXkX96lfbbtvmAjTkqI8eOI1/wsvC5bkLw58qS5kN
yaTB3+JbSZMFz0oX3tTHP+ojZdFxxci5cSRIHyDiyR29vRgmRi1E2704qyY2kXJvSHXjLgh2cH8X
r0TQd7wRvRcEUvyrIHYxOytDbQRap1SA/3v+52qzhC/kxqPY3rb2H4IYzaAik9t0mMz62FymWlCZ
HAdL9A7oHbOzp/SLAHnbQXQ1vNA/qrxDRO5MpCvPgKeI7xgUtJzsEabWWgwo86BxJ7syozDZKkpf
v7UFLLnb4qKBQ192bDfmdvOzO4XEjEuNTvA4Fk7mUnVVzhcfnyTyZJfbzdIwHxxZRe65iZrRFAuc
z5hf6AVU3SYs3YYQSyTDavR6y922LTBQpH823eo6bA4vt1/NRwdTgFP2/xsnV6bs3cHZb+GCPPgO
Iuwsb4zK2sbaWVjQifLIJwULuaA9/GagzIgs4Idr54YK0V6SK8jkLMSHCZwRPQIcbAHFxiAdU0qR
YW8KP68Mo/LJYyiv7VouOm/mwu9Aav4woVlptDM5VlSRIMcnqWYg/payF7DUHHziZcSmMZ8i8vnv
1nlJCcxTNq6+ZzPBId9XRr/V1rfFVTsUcOcGm8R7GTQYwecn91UTJ/4NJTM+Kk4GYbfFu/1nFyd0
K4NTi0eqFp23FaT0o4HJB13ZLY4RGGD0rMJHn/DA/Ipb2/y1gPj9Ytj1le81svLb8bIThweXsvL8
DBQaEUo9t3DvXWGgVXpUVl8HTJwg5M0yGOU1GGB6hiYfFTAu2pX8uHnlTRa8cnXeEPVxwwhVJu53
o7tqiX8NxXdw+LgETJ/+ljtgGCoQZaP8pQoMRGg5C8n5A7hK5wumkNQ+DbPLmq2C5wxQks35BBdF
puS+SPcDawkI9JU94JN4VS3rnM0ASHkUoKm5cefk58DYl9xwklWyVbvv3RkInqABZkgHMOpQBYY9
QtcadRzH/YmTbLImlRtXZ4MP0DrMFqR4uNz9HsEx43m1o6gCvff0LxFfBIslNJFi686OX16aRPTl
rzLeTKrWmCyCjOvrDLQUIi19jgF2XaB9KHWsZGREIUWXu3W9+tCVQ48/rbSU3SoLs5XgJC1EhrFy
u5wPi1kKIEkEhIO91ykI6P9HqgQw3g398dwXqslG28eWHCr6RbnTQGR0SCyIZCFNCYpUg64xIpei
NR/B4fsg0T8Qg8PD8Yd/K8SewnZiTCY/DRih6zBm7N3snlh2Oy5kllqL5HXNT0IVLKgwvM49Ze+n
0tD/xxzouX/vmEjQMF7PDVIYWipt4lbCQ6SrHPiwzsP/HHqi8V/iJxgmaxTe+V3y2g2f0getkSD3
fJLrF2Sd4bzkVje14oTSJBCYryrzmAVaX33r+USt5RW6UUv2m89IeFJf1+4ScZZWDGH6NEtzzHN9
AKiQP7UGAu3wgG0rjVarncyJoZbd1k66szlcKdB4bh4SMAGNHvqCe4pWNIk36W6NbGaP+xyKNc7K
bGM0M1+e4lbZsOGlwkhRRk+tqF9OW8qo/EcAghfXq+QBZpeAqt+RIxD/T7XYgoJL+JHU7JcRLQCl
6iuVNFi5r3t/U68lYvQtqN92cudxURJ841lyVvEiP36EhKk7OP1B1vegm2ku+JUYwoM/gYW471G8
mlbUeAvIiK9Oo1qSSbE8ZKqk+WH+0dG8XO/fhlg+emjsAcweMVVP9+nOyG1cramsXFWkDcRKuQJR
w01B70pxa5j93DMlfOBr9+L3jCWYjTxCqhj9Z+ilBZnH23YGkLJp64ALxUDpRCdrO0ZIsGnRUYA3
WH3HtOs4AVKqwoT/N7AQIsXU/tF15WFrnbOwQEM9LHQAqOHGuibfN/wP6/wkAWABrG/LbdTixY0z
quPv4qTCyDmchQTKrbUyQVeoYh2RU0HPmT6L+45/BCCdrB7+MVntjsYxKOVLFS3GQwS4zYO853N/
KXQvE1/DYMsqxKmGQARu8N7J4IaiTVliZ7VtGfuMbGAyTY8ECOpGm1r7quMYcGphoYhdXBZz6bot
pXuw00LIbkkJsMsfyc0GDJM0XJVmdYmo5lqM8fmJ2Jyvjg+ZFF+KJhity0RsaUWRhRg9Buw/6jZR
tZa/Tg2xZnb/8nczS8kBWxjB5ww7EV6TsGP9H3AfO0VardG+KerIW7FRUoDsx9W2XCKfKJOmTMna
8BcevJRUScV9WgiXQbwNkDk2CMIEUNHAu1whI1KNMa3S/TNjUYVJbBEXp/8XYqMtd8q12lbHi4BB
yTfqj9xKh7wshkyXkfWTk0Er624y3cXXb9r31A4ICnZ10tH5f42ZCILIvn0lN4EklOSrq+cc9nOA
GZjC1vSKtQFy55JGF9mt0PmHuSa0vpLeQg5frRpsjOtEBAv3LE6RmCj2TKIOA1GzGlVTmW8OdNkM
sSjNixZL4ZY86cUxsJn5DLmoroEbroKEDLWdxGwZZ1wwuojbjOTK0HmecrHcazq4nqCta4Oaz1lC
o8LhCCJQEwfWZQq4iwGIqlrKShWJ+iE5QwF0hq/orOlGQMpy/jqLmYp0eL3pht3TId0GH3RFFGBS
tByedvwttD6LhSgY6DUNvvMuIgRkuTt5JP93U7ySz+xMeecGZgtFWjnifoI0kjP14ez28WSRsvzN
CTSnMYf+58w3xTbzC9iObwmrU0cmnOjdgPPzGlTInoL2ssjNBunUCg9P+aYK6tWZ4F8ODbtaMzOc
kYQ6eOLSmGeyYbdfDgFbNSL2OX25p3sz8oxuvEReZNkXwNneR5PTUCkmvruZXslwqsTZ5IxnPclB
5747r3ySe6y402OGUIyhR4SHo6f4e2yTOoWWy5G/m0JHJko1wXldZ6P6Qnus886epxc3YfhyVvjn
uJ2E5HeWDRtb8GGkvSihy4lsZvi37xBmz7Z8cg/+zdIUgDiVsYjZzIxERTwWBan19K9Oq9DsBK2g
N7wLPHhp5/b73+VuRkCHVrgCM3O/xwSNu3QMSjMEzR/OoYOhSWw1p3LYhWQtaaXMv3tPCeivoTtw
NdpxtZqda6Cr/1acMAjzoImrr4eUz/Pb+A/M/ESYXA7V7vrDzkm2XmUCCtlDLtb7X+oURmCNNaC6
sN6g7zVcK7QOO9SjW6BvtopUQ01vxgtcfB0XAanQUIePnBc9Yhnk9br5wleDOmd67RLTFQ8Z05/R
QA9//xSJAISw8eigEgOnPcZL3wiCZuEu1xu9H2qsN2rGhgwJrIDQflO27pKVmtvi5Oqiqp0cqxzs
FYpH4UUAVjoKqjgtrw2SyMzSfHBBP3W5AVYMK32ethSgF3DjU+4/YL/IXM1vCUtWw8ywGQfpfOpH
wo2z/Mbqw7rTCAl1oUEFatL+oYi1NhIJ1CHgIOQtstN6GxkiySHRVOyQ/jBCnOp7KMTwYvHMpazH
Onj/HSe/2undh+lL7LDEjgbCxDJHdqJ2N5b8l3sr/GEcC3P+TQnGdBWs/6OpCb2Ludu7A5jofpL3
CsaY9fWz8SWZgJ9olxXh1xgYi4aLIAhYT2FvLIPNDG3HouzqysYA/j6FCDAxaMRzR9GlZy0MUdaA
dILxCIHTnX/pdXksq/y/E3fiax/+0hYf44B5ux/G8eBOZtuCkeNOHvdGw7/GbXhUbR22u3jVJI5T
zhGdUgBOdqnmtqQHhkgk/+AvI/OK6t+9h7EBvA2/HD8bYgMcvztZO2HKOcQvidRylv/0FlD7U8GP
MSr2puWWvS0a+NXsTqQHU5GkBPVWycD/TfkytC11opDmmCrM9g1Ei5YdiKgvR8QuLN2ywQwUWf8V
eRJA5TZMn54CPfyLPRR/7H2eI1AmD+oWpMB/ZBzOhNTg1Q6tDpeE2FK2ZMu9jmMv+g3WjKJwMsFW
XlK4qrtkeSaL8RuwyT/ttkz4qEkr5YNHdXJUAUGXqIFdrAHpMmd6mAimGKssOYHzDLTx8pG5T9nf
CYIBc+V8o50jKE2ZoBMvZOUEBjxiBEKt9Y7yYwihP8ekqOzIqTDqyu7Lb0yBG9KElZchYnL+xwRl
KWBoLwiijHwmKid7AxcPf+F10hntg8O/Fgpti+jE/q73Y24YWLhJAOB5wJuGzDE+zSyJxzj62jdT
P4GEYsLwlLqjGWC2iyjNmKjD1BkPi1KpOMgq9VpIQib1eF/0ssOVSrPUyih8NPhYPIAJswygmlu8
FTruZH8g172C2K6j5iyKX7UcBkGG7KJmLjGx+DlkbFypWQbg5t/ywKEmBDa4pClcBxSIYVBDvl/9
e63wMfjooxwaXVgE7GBjB3DZ7DxDsLE2i+v9XVRk62NO5Y5ru0EaFTUeFIPGjbxRqDG3ie5fkfS9
GbN9fQCoku7rMuMWTcbZJ9/qmGzLnJVXTKbQki+ev22Hik5pHiGluluGtvpWyotqEnw8cFPwYwk0
j3+RjEgrEp+C/VtDTtMWHV8IIf2CS90Etb4y5j4SKuacbdY5uTZ0hrIg3c4jAXvCnnyOyK+dNHt+
1SI+Rd6HeykLyszxljlRwoCCaow0iFaCSi3sF92vPHwNFC5nqUvozP9Odb+wnoeAHq8/q2+mODr/
Y2DOI1tiPuk45B2Eeuyc8ZFhP0RqRaBxORMmBtFRhr78xJmTeb4RJZzm1qhvMCL+YEOh4cgm0l99
84FDsAT0aFj8glTOM49Ep8T/r5KR3Jct+E1A3YULXodl99kwKkMCHoP1PWZiVFWmPuwKQu5jMOgr
iK7eL+eBDyxd30RSnNEUuRmHIQqLo47QrBTkd3uA3uUKlT54e7Y0slwN5IRzHAbTmNC+Pc5XOmHb
Xo3cNzVs4lXVBUEalTU2K+XMsmdvotTnXrYiJcXniwxvvgZfCvUyPoxicUSeHszcBVSEy2g/Dh6J
XV6XXIKt6MXIXmG69+LaakNfglt0Gu6+W0Vb+BUWO2mpd8rL3HHlryxnV6S1THao3Ifn/Uls1Z10
klui8qsgybOVgNGLIMnINRbv5+e8+4ux1fdhFRVRpG3zXge/DIQpRjlBrV1ffgGc2NOPgBCfUPXg
gLKfISn3KzGTnBWFdJZJfAqGWW/aaD2iYQ3ntaez238d3eY1lvcBx6dOIS6jGZtarixMCPxvp4v7
bEW5vSv7VVtA6ZAkkDtCtVBH2DW4vVNJbqOdNd+wWYPjLJwAAggvpehWiLWZLZUhlC9HWhHVfYCY
RswI/33ip2IpPp1OcYOkKGNOmkvZtS5FVujCiVcNjyNrpVDUdoEBKVMlhz5OeMG/rFXMsGbC89S5
jvg0t/QVxRhBREE6ArF73PKslB1C3ss4IS63R9dxDQ6u63Bry78EHeQPyXYwWmVtHT44PmIZiiXK
nKYVJp9vTnqvAvihla35eFA+Qgu4qp95+jwmc+Aq9OteOMs/r/OE0EwgvzNzIFmVsOlKXg79tsoQ
rduWBs+WDgOIWfC7xzE5r8TI6p5HY0tah1VCFuYOKI4ghRfOV8IxumsRIjB88DpvKK4l8ACY2XXp
CwU6F4NW4a9iUlEMNe487Syt7VHKfnAe5VAD0zgucgtyGRHNxupdOBeXypECjECLMIlo2wyxmNDb
MWE/wTPMcF2PFbeRSPA7KMVoKThLaYl68H/pGLvqNhYP57HiWzvDgVIrAnT3f1nNwg9HDlXyW70y
XOLmZh+su/P01j9IJNWU0OWxnWoNj1btfLmEfFWqpHCXropfkQnhpEyR+AAVDddhCRcZYI/uErwD
I1i89++8FPnuy+Rtn304Sxa7KXmhWYnMJy11XF4muW6CvAv9RXJCz7puCsy8ob4vwgJmwF0eofxF
y9kLTOOBOk8g7CQJZI/crngGMQ0dciyck0uaZWSOph097neYuB94Oj6In1sOUMGzfN8kDjqx4OvY
nUqctxJUur76QhofLF4zaDYG2afe2cc7e7Mwm7q6dTGcvxLNNaR5MN+TB5vW7qd2ZCtdEeaL6dMI
c7x2GSPHvF++vjKWdLjonwsYSoTUxfAQe5MCWZFgLLiJ0ERiqI142z6SdI+oBcYvTtJKVQihdq8I
7Tiyma2s//qYf8HNoxKS0Y70pG7KVz9Uzuu+zyUjRcBavrmOUqXA/l7BCxZ6ElyIwLfi+y1RFiUj
KcYS4AKgy68s3KozaBG+uZxOG+GfDb/73Mwh05crh4exd3rsaLpaY8uGdzPAfF94qQ0H1utaz+E7
s3TpjHkWj5B0IHs86A2CzCUxOb3BFMb3jSUnFNRpzbiqov4dWebjQHcvPMw/TU70KJRHLg7qd/7N
M5UuYM7PEPUO78EUG/ShXTphfWkT++nos6UMRsF1BL4L2SE+RtHnJJRNLQASXIeHaxApAyWLDZpK
XA2l7/m3WxPW+VYmFpcBLvrODWpt8P0SBwc/b/pe9oAuW9x2XApIhwcWrpZZE5FXA6/3s+wPHcUX
NgjNuLrR+rX+Chqi+HunRVfB38sdmtgUCG6YX17cGyGIVKZmhUuW/wxdDlSENNbIVJS0wDDgOsmv
rqtvzi8w1WLI1DCZfKpdZcs82pU+7ubh0dHdMtFyxuoln9OUClOZHzKCA73LuXb5HrUYrBm3ZhXo
N+fKMdxRxJVDhuo3v4k1HpxUGTwFiftGpAab3anF59dotraLkjuew758wSLhnTeyjVSEvrq5sF45
UtA9AmrF8+uS4cKeZBAFAzXRNfiLHDPWwPZovvqZ82tvHNEAyQ8/QhgYLYk+kexLQnhzwgWGU5m7
Xns1KXnxbccUqLaiaITak7wGUV6R4usYxYI0QAsWBwOJHOIxMVy98YjoVTz98pTSa2HN85piH6w/
wMhhDiDf/oTzxGhD8XlG7rOKN7gcc60XfDsbIMKezvoHVQ7Fo1Da5I1/R+iIDC7zzTzwtsXGESXs
HtbkqXyR9BhEBqJJZVcUcHyXJXGqevSBM/lA0CO4Wpspxgf2sV+LP/oXu/Q8r4pmvUpco4oyXqDT
Sl/iAj+Bg+yKSpPp9QAQz01SSHfr+rLxELbx4dWBvE38Pa8ZdJwSLMX6K/hHZbqpErCss+xGjw5E
gsk1Kqt1Wvs22ISEZtObtLHeyDtS9wGIBvJmC9CLPeUAUXm0YwXployRTVOAie4Bqt7W2MszE2Yt
vkWSEaciMEeAdXGNNd9kKWBGKJmsa/n0wo4r8ZhWvKq3p2epvHQ+IcTdLrzDdf9UOsqai+glesWb
J7Vp5qRAcAQyA4W3hYujunM5bmwh62CJb4LW65sOgL8Mhg9gcA8RSLFzw2Yemk1UbE3FrLjSkbQC
aO5Q9zeRdIqEpLKcWVCeoyKh1PjhiohC0GnzqquGMaySySPpT7aYKCUUaLcjvDLSpswdN1br/TRk
fLbR9N67/qgCsiTzWObssHYtOrCyF9ZZ4JEJnmfnOTMq71k4ZUJEwljHvKQ4ac5P+k16/S53cXh4
PxaSMQqNiADpwP1TWO+Of9hj1ewdWsPiKcSlwyIbuBXi9WsVkuGzHp2W+aYQzsK6iWk2Oq468ekK
ao7LKCserfaHnoTByGPISEtnx2dIJ1XHbhJxIiTJ9ZwBgJaqIV/eqFFGxx1FULLsnhox8spCHEtf
QovEYre5KNy3YRi9gbKC+qFXTmhAEunirI6Zx2jAo1qwh+t6gXaqHbQYpKZaPwPbrXqKheq4DzDm
Gb6OhwhzQwPQR4rqRMoQmB/Mp705C8C2JKWZPV0i2uQHQnwU8EUi52rSphl02mx2MltmcclYu5xD
uxR+mRkPUpOpWYIsitbAO4JAqOeS6lXePU+HAtsbZ79Bp6Bw4LdERw/aPwDQxJ3MiEQek2Zu+Pal
9xGT0grXxkr1rp3pL8IueO+VwBS0Iu+jYZ2Pqgs3Yr9nFZ16YqDnKRUHesamAJR5XisetxJO/NPC
knZgPrrL1BIg34neBdNEaOxZ5iY0YjxgvfpaXhbTfmWYC9x4SlF/bpWO8VB6iELFHlKKUqKklvH6
cizJvym8CVmAMxXrMOxdZCIA7M89VZQOsi4E5952eVcDA1dRePdEf7ZGNASo0mYaEHroFXan6rF/
Tn8yP06pbWPsWjPQyt5xF9rtlxrDew4gFWYEdbB58jl60YumEKTkntaYNbsSEfXNxfoAF5YsBoqL
pmhqTIfKZcCrlAGhy9gmBMAnuBg61VXyHrlFgcUIwXgPFBwF++UQS7txWioRMLV9nZ81SpwlElMl
VNynwb32W3Nm2dzYEi/yCoIZ4QkZY+Q9ZICBuS0LaW4xa91RpiQxaw/LoTvfX9LK9ixISBpQrFRJ
gGi9hXnPCac3J7PZzzs4SXx73CZRvDzPt8/PBX/TChQckGD14GlvUmqj9x2OMwSW4Tjxtryg9XKT
4+kgdP72bXG72WzJwGZ4EvSysbKWwy6T19sqEaHwC01S7dBhls9Y2HR+bOG0FlfD9VdBKIVNnsJ/
4WQO9Kpk7S0b3PQ7TxDuHwZWCz7tdJEtwNIo/gQDt/oFVOJn+aV+hzqxry4z1oK01sxsG802HCJG
ufPfkiDAVFEiTIPW/lPGt/0hcvQIk4GrJ1Vi48u5FqS+FXxqDUXs6fJYagW7wabsBcxiMRERPVZT
WI/yI+F77Ub0U+WziE/I7ulX/nWqQMwwrkPUvbqDqHd+o1fYXYTSWT8yA70725AxypcIYjWx6ldq
RwQ3vFXasH/nOABX47diCQVUG3sQeuwtKAfpGIZY4W8xWo/zyVKtYHdxvirvytjlGf/WdjYda3Ge
1EgRaYswuUfq6LjmLRE/Syk5oiy2tCODzaPrQiIKgpVSlMQ6MppBuGS7gTvWKglbBaunQzFHn8ix
mY5WtCJe9g+FI40qJt8x5sEwr4vFK16BJgLX1gFdreEQ/IFNabnzwOIaznXTG3MwQNDJti10s2YD
GXPTngAIDytLXfGpdaDnr6gm4KpWcyjx3wl3+ka0KQpc7aJyOcL1TMqBf/YVlProOKf3w9TtE7aa
Px7p0IQujArhJNwgj6Jkk1LyhuURWTA9l6oQ4gZyjclnVyVTtujwYiVSZDjbnDaiYdz11xA8e7lF
635jk1X55SGDUc7C5rfiPvAZ9kGy6cI1BuGDTpB0XELDZaSoYAX/+mp7ZNVTidTvUw2MzI06Ep37
f6DBAn1yEfcGW96ClNMYVelm3U1FlPCL7ORz4G/apgzw7aGFwfc9BftYvGdj4Rlru5iL5xBvBviq
ybqBsp7MlnPf4lueorYFfOi0iDewjkifIGcww5jXGiR2e9IiRgPAe8tHZahlQvE6/chKqgwjX73O
k3GtWEKRQM9pOGroZFDLNziEx+Lavu5bK6Q1Iz/x4TqnZT27qL6Ue1zRXK423n36mMg905Ghf35V
NJSscFqRURgVY43xx20icla3gh1Je5U+cjImc390Lf24rk3+1UiVoKOjGuU0TELpEoc4poHgFI63
MoGtaAjcDEvUGSz8Js0UWFoAjjAmBHFRviVWVoEn+MZJ/TlV75x0z1sfCf8JT2HMBf5IejsCetvT
xOd9QMtJI/BzVsMRUjqw1YVyV2CrdNfsmV2xy2ywjIEABAvly1qPwW5cghUB4ex2FIhIXwWB5JEi
4+Wm5P6J+05lhh+gApftwnjDxy5PVn0kh/SiW7a6Cw4P+4J6x2KhbumMReQGbl3gJmo3lRhT6j8f
P2Qr6igA+bzsj1zWDkw6BivNjAht0Jac8OG27XIN5bJ5hG05QYgjgKWaBVzlK0Aaes/BXlDqFQ+E
aYWXPs7aJZ/1Qd9eFhFNS9i1BHpNpNWKdiDtENFXhs0LOXEJMH5ncvh57kXNoUcOK96KyCfLTAMk
lsV5yk1E46ab88qUbyEHfdjBx9ALS4H+X+KTjY73Y/c/0+MQcfvEX8jvWLl/RrR8Ob7N/E1buXQt
9PrnvUN09O4N9agumBpTTvZVoKwJZmJbqot6SAJPxgs3mR/FWqkZ2VROxqdOz6HoCWku7EntnS+4
qQmPfHBEfYoJP7R4ANLgTN1S46IomQV38vjWYyWTsuspwjyXVL1jDB5ujsxzQTxEU/qINFtSPaht
OzvfERG6vxJzPWyBM/ZylvpUoI9OQAcsHB51KLPm/P3Of3y8X/HIpy18ztG6zcxTb3F6GLhFbKHc
4bl9wyhkEydO1BMyjv+Yk4Icy4FrOly4zIAqsxeIBqaByZ/FMngt7NHgUHlZlZUb/V9i0hTdrx5l
C7I4cM1fyaoMBDSe18bYMzyD311lr8aVk/VPFdg2y4/QPBIuXb4qKHLVQHrp8cXkfSclcrE/Cl6U
t/ORcgAhfkXcXTVsvnWjFHZ4fEjyWYBCgl/96VcXE5yIOLHd4gYVSQv1MhxwUPAjTd63D1AWMPXm
tBHVR93+xCPvS8xBD5kNWBDlBQt2p2fqB6SOn976/70n+4yFQUTAobZK2epHAI+u9RfKARinK6MC
GbLxORxZflATGsVredTcmB0ar/TZGHoJpX1uQFZUw5lMuO+SWZCaHiwCdJ2E1CBzAkn/rAS5DeTh
VfWYem7P9Vn8Mo5aN+z9keMh2FQMiWqhQg9pUk0BmhZ8vXufAgAavUGHpCdtDcb8zqm6bgGCQ+FG
C2pnc49zytqRga06UN62OZ1ncHiAbTqJ9M8eejAMFv0SE6arTiPPydEBElMYzERH/ZaU7z6zurRZ
B6S2lWhoSBhbzbIY0Pt/QLn7HZWsvxwYQhxDHxTatlL/zna54vy8qKUAkO8AZM03h7ASUP0KXRCy
GtqErU7XJ0/IQbvLQugiaydGi58rmzrm4/fnCzPmajfsg3ojmtzOSJDOxumx0TKXq0ZMIIZlhx94
kzvM4ZusKfG2ZoJeAXqrAQVRdjjPYwOFO0U0Sd6W1nLdM0+CURZk4O8/uHh0YVkI/pqEDUmJGYKp
tN80hnrF+E0zP1+LrCSl+wZ4uHSs8fUDaKHmAifNiRCTLd5jNrg3nhXPK6SlIza+/RPx6/UipNWA
3jENZi/ZlfzTYEYX9xstdfTXlBwkTJXW8+g50goFmJHtb4cciMAaYVnHC/omi+ilBzEwAVgY/iGB
Ai+MLJa8N0dqM+5vRYOWI6a0cKtfP0snP5e/WOaq9hU6TTQjTwYmAyVZS0cHToyheqmY7ODhZRQ0
pUdtDue6d16AnMMrUzFKDNGqzG+IURs4Xaadxs1FWfvLALa/4hf7RxpixFLCHcUp6iewxi1uMZCx
gd9B9uR89P5bpFEtmjQu+hj5eaNABVgMIZmx1p1wMYEUOj+/K+P4B8Hx4sPs3TivlcVCx+e7Zqst
tASkknaAWivlbVBivGcj6KD8WdEjR9Jrl2peuqmH4hFyB7l8l3TydLL51lnZQXks7EbzmLLxceZT
CGtiYvZtjaUu5/swy+RQJTd/kdoVBlzf80l5QAlV6nRSG165pv0zwiSrtCUkyaT4ssljMMmcyXS2
3IkQtYX7s9OoBPRislLdzksBWMfpgzUV+nQT4lBL2OzWKrLIo2dJeSIjIsHhn886ChS+XrUQQgAU
O1Kmm7RUuEfn10S8lgCdN79D5PX8gpJbPkCTAh3kbcAGXDnNlwbuGqHRctgL6nwjSEvPxdofvuXw
OFzKA/Jnx45p2TOm3eBjNg6l+Dn0ir1UcYW8UGgk1P0/elBlO2gNHn9nkD4d1uBgUwUNS2AV7Bpb
5gUD9fTUZU1/Xp6FLmbLr6QW9eEkydl68vy7Rw6qHRXhoqx7S9riozHodoE5fCf5tTIWbfIXp7LY
0t6Sq98KbdSNoJ/CZbFQ2JDLQBM1nMX9u+8YaqzfmTcEnZuYUiUbR/9xOTJDLC1Uv8UsSY+xTzhQ
KNKE4cfe+mdIHHG9gDGMjG42Wa6e2bTNVRzFLaIJK35roVHKsE6LhOCtPKjLxpzXiTQFgtsA2ie0
GfT7YTXoFGcjD1ccljUJApsKBlSW22lukMKTzTaSVxotXM6zSZlEEk/KTmtgcyDeWHzZKeSbBftC
al1FiXafPnHskv2/EvSoI/uYEj+kmvoG/UsVgIEk/MAdU9diWjoL2005rpD/SXNcwveDx9WtCyv/
VdyIKfVa09cuZCBZegQs1SRijsbrdtzbcVhGt1s0vEoBJCMLIb6C1LUvhfWM+3WRByh36nKRfby8
45jUxSeD4H0RxxW8PdVbdUBxTOAMwXfiDzLbFMZ+ofXM6r/zH+EY3sWw/YgFvmtJt1+Cg+YUG00K
AyIhDEUN9R1I9IVdCbuS60V8vd1mViVD0GEak5mBdvOZs2P74FVhpl6foAQURv9bCjqPoBMMTcyf
G8+AsIKq17DTfvZ2m4jVY0RxbCpSBE2a9B8TKaC0qnICPOLtEx82I6Bn1KYLwUai9EeMSgSKpdD5
g86itCY0AJlqyE0vhpR8X0dwlP8SLxynFesTak7PiCjUIuAR8cPqucHvN6Uh3Hs8GhGeOBBdFFIm
YDbb5pH5PWYvtOCz1YDlK3RcrK2QVyof4J9vwKfkdg0lSODJxiBwH/Kj9gP+Ij2oZC0CsUERIvkS
7WlOIn0OWKnBQP/W4Lgb1Bu+cyfgI8zytrRDEwXQALLUwocOO2L+cfoDlpVoNh4v8e5eFSmDOTQx
ASGsRBTyOzQ7BMr6XPvux6TVCJYOaitCQo0ZDs7NwDqaJ3HfBVLcb2BsXLLbMYmbpXM5dLZBrUOd
0LqTzL24ednYvh1GjYpjpvAVFWwpQd6lxyAx7MwrpM8FKlFD6kn9TTueCqGpChzq+IL9NXTRYpYG
JTh5EfYVpkiE0tz+P4nF7RqxqJ8RMiw662r0tTV1dYHur7y0flkpSWiIGKADaXoJAWMdtLITHDRY
qMFfHJed8t8uy4t+NlW3LaHy/aD1yT85iTQGCUxU12kKSNpp5oPuYPkGwZUSrNSCyP0AtvS4UaiP
04FaBeuzXC8P36sJ4E8acQzXUu3hs2BKYKQ/O7gZTw+gOUXe87z9bCkeFgWTrVMXnn/TjdHHcOSL
J2XzG/JDDitpfgY0F4ViFOzLk/CAXO5vXdUUZ+Oq7IVPVDLXBXGKIky9X6+p43qf/iaaHAJt/ZSL
AAlj1Wa9lOrhY1jZOFjXuLvNcFSpCAYoYQM//4M27d3ICH/eqzYpqKrJwInfGQBTwQsGTIp6qmNs
SyLcuhCa4t1HmrZx+hlasZhza8bP+Q/8Q7Z+oQ+6QJyndUldUbzQCsnCNPua4VgDlt3ZjiG3QDh2
pxe0aZmsVJFmFInBQg2ZYYH6ckFzFZoaEvEX19yRnXrTCbaQft8mpczC1QxTm4hoL7nf/3q2RqhE
bEaajoWJ5VVu2d02E3i90vCqVx4S2sxvREZPQ7je6JGTR137EV1Ac441A4CW81NR1TaTssZF1EqJ
qZ0ncdFIh3tzYHyoElBqvahy/w565/RrVya2y9PCJAgYmsleTR6BqWzA3hx8zOUskDaF2z8HaQIj
6PGm9dAyFAknpzZI771SN8vgqw8QY3sah5ezUsETaBTi0P45fsheuwi5rlco8YtXx1PXUtQM0dFl
ig9HAhWWQd3IB/DRyCl4ogMUGQ+C5wChZdcWAX/mb+LC1B/Vb8IPMgXhrKOHRBQFJ+pA5WUaRuCB
gYKhx39Hr3zAXDzO2DtOoIvjfFhzuysoPipXcw1IxL/vfEV/6HbFGD/hrc3+UHAlzLBNwo3J7BSB
tJn0LNklUWXrIBrrsoE6K4N0az8xp4WA+hF9aA8SXChdxgLSd6Ioq0vCir3b3qib4HztSak40xhf
CMs5V7QKDmJlNA8PL4lVnUY+ShqSVGXDCVp4pFH/iXl+W8444OFF1bHeMRElXxpLS0Y4xF77jO3g
PgeLRdcnBLOwdbUWrtSGakfZvK5BppjG4DU+3VNxFGomufYwaCcDBgprF2Xft3HnlzWX8V4RMZIs
M/V/+IJyvd/TWefceWHCiOTkahpdjXjyNlfu5+hIIssbMifq3TTo7XUxHo6IBaz5GDeQP7iXvL8T
06rpuWJlMh4yJBFg+TScvGVzOkGY0zMGdNCvb9ofe9AEUY8Fpf2nD/hXI0/ST2KmMkcP37gmKfB1
A3oJ/cTHM1ciZtRQGcTHWIBXf8IVZlOojgQ50ucBl026tSg3XhDpm7qo7hVeTbdRFbwQRbHAJ307
oJH8kBtKqEwTfz6CTDkrBv3NqfVCyPfOVPx0clrNtW1fUios1HsjixMzl6k/pwrKBrRac2qn8bJF
wteqjdpKUMy7pnGOUpn1Zz4+BTFzz7Uj1hQApRCX2ATgx5swS1VSIDMPlXS6wSwQIulCygYwrrA+
tadHBaOIuBLqE116k68xLyc4s+jHJaprmG7cPbCm8xCnmjziXOHVSf9Szo3/us674B7pRB0vJ3ov
PComGjG2Xm/o5XjcQBCpNMsqzM9ZR6ut8/vR/t8XUNXtZBnyfw/5/DgZtwUUwtn+1VA+N0yKMfqw
TKgIhqZGbWhzHRGCgM72Bd/Rgz+8SnFj/NJYyA2RQ2Y6DuudAi1m62p8JIrEljYmSn2ipIaVliXz
gu/dNQosKrpogoy/Y8SmM4yNNFCapRTRF4fbAiZuETSBzdTeM5g49tH41R4E8F9RCXsma51UtMTd
vx6/apJuLZAW4SqhEuwbK0ZMLjegmE1MpBuaNjpN+C6tOfqba8x67NjflKV6QTrY4PNJRyMqwdTp
yRjAJ7dzRg0N7YRKczVLnuS/odDy1NIBNHCMKY7IJc5jGPpLrYDg883ngK28p5bg1sF/Yvqy71ti
3oKSbapUONQYUFag7k+WWqye26kwYsiPLdWcDEPYEeXXx4/xNwtIMKuTjYoSSbYGzGxQ2RgiyqLL
LZd1p9YcK/3bSSjsCQZkGTBiOaAlsPNGzre15D2iWqniRBL9WfnTJGmo0ZlBbw5jBjC0b/MzJ0AA
FlAL/yFeYNCDSZ26s27uFzKxcbk6iH3F++c3Yg923kWKu/a2hUoczJPsDPJpHmiDpnbzcOYvgd+K
cI7/TVTHUznyGALhfddVZRExKQpBlycxEAlZgHBxdBxwWk0sqK//DsyWdvDoPF+oj0MvknQ60Qa7
aFrAJYtMOXSlZr3iGs6h2xuPmOHuv2txAhR6E+B5YLU+CpSJ9F95ylidK+r3+3jZwszoiz2xRPes
KKSU093HE0Wr9SvIEujyr/nzHbj9vGR5EmQwkmg7OPluFJPGce0RzwPSDXYEEq+Jy6JmITFAZ0D4
/3WEKrFXNFF9rgzotWtZVHkzDM4mG5UBsR/1oEvmEbwgEOTMR88bRz2BU3wzCwoJBMo7tzNB2/YU
1FtKG/W4hxTtbgmD1R0nWmqVnU8DrfNVHF4u75BxM+ttXAy5YvoeQKd0hG8ghLZJQEkj3TLLNEIc
fCCKsZntaoaHmuyFKsUDY8bOcq2rh/2nsfkL4A0/UbSaMh+Zd3Ty80sjnecCt+MPyUhkgB8k1z/e
Lz2vAXhcaJF72UtQL/AMPc4/4ZO3+cEFueOkOniZWw0G8mvYnEhHYxq6NKm6JoX7LKXL1epMztLB
bP6Y/z9iOy0n8D1cjPJcizUg32ky5PehiXz31tdV+Vnzu68KWcmfIsgiTzMb3ZCpUfeXSMjmsTq/
OmAQJ/xpbKxmHEKAmlPr+UCU14tszcgfENDVq7zXgbwyyIfKwSBktB+adwyxnkstseryyAEqczK7
0DhURAo3vEff58abaGTN4teQs61Ze/nilx7j5NDmnbk5rv/z5STRjzRLTXrVv5AYyzSADdGTnmXn
fj9IrjsdTcyPsupDVepcaQ0+8XwmKW5q1XDy7UHO60LqtDU64PgeNpgauMXSnT5aGlb3uXQOdzVR
e3RY4+a7C3qPQfkAOqxyTy+HnZTRfICSj4Kj+sdXX8dIhgXRznD0tRNFjuBBvRHG6w6x9TtNcaFs
LsewaKhpD3G3lwxOD92mubcc2xSCfzlJ/g2VTRjczjvhrjv7OtzMw2H1aXthwQTleXYaLtlIXVWY
CsAmHorT0DS9crgRdgBU+shqo10cnGuQshIbra96SN8YFYSZuRLmtuAKmpUSK/ECjWMhFQtQZtGM
pbffx597IrusA4zxGQCSVL4/b4GOG5twRBpNE1fD2ARBvfpRYixj+0fNK8nIW7V6hd9sGUqlJDz+
uIVbOGOdJUCZrBRg5upM5tF+Pn1ZNOKT+efk++0pvUeqJxRnXJrfe4jzzkLgKOJIzKYA8nIswzzI
b9Dx7F9kTwPPx8b52PXdLEAf1PWSU2ZxUNukEJGA/KKaq35znS4+ei59qF5A6d829sLYEM/SjTD0
sxTQGCHQy+LB+2z3YHsdhWQlb3KNF38F4gx9wnS5MVslIufQccYh1A1J+xBUlN52OapYJGu1bsX8
6yUBUsTig5OoqW/sY4CnwELD5D3nGmMgeZFCjcQ05804H8QSfzhlSSeqMXvXS7cHmKU6kll+wq3w
k0yL3NGkSSww3LX0cEt9cXkC7nZVt1kH5WXG2UhFTrT6FE3mTHcxoEgcYULjmr9fbqBkaaqxsifa
bvRdlIC40jWW23ub/6tFEz1sBGQwMIvyW0pe1vF19T09xAYzyOU+TVIjuget8SZh8/XLUsOA2tK4
mzjf+zUNxxKXlgTy6GV8bd29z5O+BGLYbd/boN3vVKnkQMh1V0P3aoj8w6rKvQMui90Rzq5O6oV7
pOUGf8UxcyYgDMeCtr2jE+pEnQh/U0MCt/1vXVNscdD9OAggWZWDkN0JqAntqRltNJnbGE3cbQzP
5mmzarWwINSPIe/KObSKK0Ug6GXLrF95lpyPMFVQUmc5a3R8ehq2R9fjSiy9RM+KZwnMUaEW8CJe
B6D4ofTZoirJfYjI5DN2RLQr5ukNXyuCkP5QhYiDLIzIYKMBw/e5AxS3sdmM7iKq64zgGX0K5bCf
CV0A/53o0ywJpcp9vzSK2fGKr9/ZhkIsHHMNO2yMLZoxxw5w6TzeU6mb0SJdHDb1fQqYuE7DkbeM
uIYYvl3UUYNgiyEYZt8lh5YSrqyoqTfqHFM20uBrc16EO4Umhfx75KNDpN/ctvj/rqfoXVDS+lHJ
pKwwu/GSOIrgsNAnLVCH6x2R0+lodBIVub8j4Qhx+xO+6jfNlO1JyR/P0M5vuw/060fH2u8hy1BP
4zW5L5B5MZ9IMWHTD2xSQg93aryHQ6pf8dpLFbcVybscuy6+DWuILyTZG9kSFP+SdxtDKaibl8Cn
m0QOIrzEWAfkvFyEVnaWHezYmMr6s8Epg7AHDt+THiEDHs49uj7Zy6Un/uU0VxPrCDrpiyoccXWm
H4nvI1TzttUzFJWhzOixdO80IYt0ZTsPP9r2db7b6eYdU2A1OoM/o8xi5+vAwiSqel0NWxS8Y98O
IEqKdEPS8x9FOM6ueaUz/hH6mZKWTqoJjf7zVAAleq67FN+UpHiXO1AIF4TKA5CqCmHQlzkZXGft
eGF1VoLl4nQa4+VL1+hfkaW/UMbpKK8ZL0krLaQcLRSVRp3rJsz7ui5D7tCekyxtpe+RTYTY7Faq
g1h04Sk/S1QvBmFENBJwD+9SyIld2VdnB3RnkUWnJNX/7ecM8SWHRLLANgOuX+H+6pdqhCPBU/zl
CwQeyUNBHxkIKFChUr/xz+V0V3G1Zv/tZDEc2bj0L1k57QaM3Itrd82m2c1Mw8v+NcqgJ0TaGapF
Kgxw4FFvtrDZ8OuDPvexCr3jTH/ZPjY/+JCh0CSM+fAP7yDrZd1NtXVRFEPadxTSzHETqo3MGCwh
KRg+uRQ34hLDWU5BHDXulxfE+kuxUzJ7Pf6yRUEC3MQ1t52pY9COBAHfQiZ5IgOG3fUEpaWkabPI
UZdEMifKFEdPOSWJF71GUSUWu7vReCMVq+HKrQxmFU4K5x91MiitM3sUhla9QzBWFLmOMhq/Ps91
/+arcC0G9CFhFgx7bd9xJ3OZlGnXypMVpreDkU3yAOxX0s3ANN9375F5fXwfocH7NBN869xGZ5Ne
RvAPKMXwe7sMgs0gNTtZ0oWK6ZbAIjqmIhqmC/uCAyIzQjJ7C1O4nXVDQam7IuDVIF1bIF9F1EUb
DBRO7Fc1eMKYmQVo4mFK8RPXwqVggIkHevXCnkaoaq46PPzFcMwYkC5XO/mVXx0axgDGXkdFMHzO
prke9bX27MNFu/+6s81AZUcag8J7oXszsbK9seRN3FtuLsd4u+UuCsPWinPq6+95YOUO3y1lPRH2
U7Vwxp0PLqwyuCevp1LZ7dXAXeincB8c3NEd4rYpsiVHgxcU2FyuhuqTHErHywr2nbLvhhPhIUt/
SRsd8MzJAfeijIdLnVz+VtAsfqKVH9bS/UfknglLFM3cFUZqbMxw5+kVe8k2qKJneGyq6rZgxvfn
xFlxBJGuYE3GbyruZFkXMFulb72v8dSZEkgGBC/J5TcOhumWo9yb6SsOQWf1TeGEtW/PZ7OgcKw/
VtRWTQ0JZVmRjgO1+WnZQrQYreYZFELCG+LFCIjW+SXvbJ9cZcVp/x5RpNDyTFvF89ZCPD+cYDFO
znsF05OuFsp5dt8ZN0zVAUgMOHjHuE62DmTxF1G6vFJSsMXgUI91H9jM3rzdRBRsKkQUNKtiu1c/
r42mUtdZBPlYGC90VI2bn2PyeLKugUIpuv4eLB8bcR9pvjU3IKiam7VwnQlYK6e/QT3eghs63KFe
6SVPgN1lJi7EeU0V//92oXsz83BQ7OdrkpGwno3uK7Lc4j4cTcWI93iJXIQlS4GZZq3RnH8qElXa
yD2guMJSME0ZKsLM/Vuu0kJa7H1deBBIdtxGK4AnghEBVDAuJ/NxAZeEmzrzlTtD2ut/2isD5tVF
HZPr/tq4Y6g8vudOfLIZwNWQE9XTktXIlaMChfjcg8dWhuxD48q/0yNTodlDP5Z+OZIH4rQmC0tK
mnisGz/ZFsNsA1T6EbZjR370UY2fD3G85Rby6JtoWv7rx7xVJgmevqDRTXQQ4NxOXwo8uODbAHW3
Zfqte/Hnk7buXcpBsXytfMkOtNKF7vk94nbH0SrL095VWACW8BMM1lcF7PF1d1WaU68ZIOGUeSeP
3SEkydToXjokUP9e/J+ckde5RUvd2jJY1U7iqCicWUgCL5AT/DNAMKa2b0Y8B0X6A4nwOTN1zIAK
F/zfLQCh6MdkTPrhS9VL41sONn44EB91/rTFkunqIpskMDnSXiACv4gWho2a/qvcV+hUEnrvZpzI
1Gv1w61404j7x+RlYAgB3UD/AoD768yqoDboEi5yj2/4taLcW5jjqtuipxhUmGKhR6nOKTB0PyfD
8XobBkseTjgXJSBdJUDqNE+zQZ32D7OsPCn1iIZ/oACCfv8yzv5roX8fpm33BPWsYpNMD0M/2eMN
HgDuxbk1VAKthsXHnfV0RBfzQ8EI0NNoHXnkwTIv0TOsjtZ2DYY6oPRhEzm4Wd9otNzFyT5s+eF9
GpyJWsdoofOQGcJE9pdQSEatmNHGvsWP9PE1QQIB3B4eWuMkbtlh8KNs0BVjSWbtPEEjfuxVDM9j
NkfUSKPeCzNxfd4OkrrLVxE6yiLvV/2Qv6CwetOPZeLxVSU24Ybl9a2b4a9SgTC7hGGK6FfES3dz
qcZj2b2A3UcPmfgnN7vZNGweY0Dh4JQ1EmGPZjJvviXHxNmVyfh6nvw2uVOsvlLw4tZwihHD/qQn
FW9GGHCdWvgwDfIjsxfx7JZWfQOL+TfZzxXWlyZlT2bsrbvFvhi8WEcpxndUFPGHNIvTRUJJFPbb
l/DCnSYjg0KzR3YeJN8j4pdrRYnKOs2Exrgf3C2Y2cVE2VlAu3cfYWgo+5T5DMzT7BKdRfMDaz+y
VNCVmCzfgqv1bB3Chga5ObMd4eciMie5tpjXaQxBvSPwDfY2oRNUWkRwfou5uyzfCe6mcTwGCmAG
ql92R9dfK5hzowqK+Ko7mjiFPOcyl7FBIM/eBg4uw5ZiXHUqmsxDoxY2ktrdiDW2lsHBoShZu7u9
5sY7gZ1JAaONgJ79grMRRqBwwMRCjdyn8ZruHm+eyqbs981+XxUO1OaJU/+9bKfp0wQNOb1uidwh
1T21o53JLEpCGfBhdWdtEIlTbBFlVXAuFnYfnOWYAD+M4/f2B8TrhmVNJSw9RM58bFcn1FNFaPsz
DcbrdtFe6Ht2iMoWxYOBVeaf4kxh1y/qtQ0EJa2D/VJr2kl2QRAxRb1nPkHPp2dB5UlUqFCMqlpR
FMrg9IxEryqMDlH87bS7QQtYNxXGagQgy/4QkJv+r6oVDxdI6Pm8zgy5TIKZY3LOp6MhWRVUbdbp
eqOQvC3zZTufF9W097knHKA9oEHQu6hE4koZN7WkKlpWWw+G8Al53QLRzVAO0mDyffs122s/jS7s
ie29IXrofix2gYzyfHdUej8Z8IYJkLa/Hut+xO8buP1vfkWngC+nkd2lnjNbpw7TDEc5J74RN3rT
dddJXleSRPyKOvu6rb3ze02fuPorzWr+B+JuH/f6mvVvlPGUUXZLPmTZHlzO2nu8rRApIRFbTy6b
AYvNcA4ytPYnRZim8ZmHnIzrWk5BgzyAojGWVi5PSWLhh3nW9RlpQZopNw+rxeVTB1co7fC4fcqX
q17jPPnInILcVqvNXIvPnm6oQkeQRpR+Yb38zqY3GfHSlcMfmoFfv991noAwgCFJZ9WQhq7Jpg7s
2/P+DwpZ+hfTeBs1rjKH7BrKGI89s6n5DPWDexE3sx/1zLNGJDKPtakVtaHR76AhsjGD9PyrTqde
eaER0oV27He0QKoJ0oSx7n2MRidLkaWk6R5FJy1+d3T8O33KrYRL16/CxD88AZNebRD67N02HFTt
el37OBNvuDb7pnwFriH+nv625K0YLR+Yehd8+pWX+f0YTfhU3n20M4+O4ktpKSE8uVFQTYrk5mEc
DEUEubgYo+gustl/sZLMdPO8NZkriFNqe1YXl7syz+vZKO7b8eivNNc1AIwYkMvnmP4QT6BVu9Jz
gCa5Y2Mj0u9aCToZicw3TNbd01s9E8qCKgDRfiBwa5pTcWzJ0KIy6EMB/u+d/O/MWnPVCN7iAqAt
gemPuFJKms/utusbRPfvurKzJuYJIko4oab68n6R5katApk5HGmgSssT2gblzs02osHnAgyDsCC0
RRiII4lia6TNB4CMOXIXq6+FsntqOHaj3ICGuk/zV3qFgxJvA2DmL8bT8KbvL8IcvtGRe/mgDRjf
ZExngXXYJ8g6LI0XFMvypaLGS/y+Wb7sxpA/aSuPXQXZqSD/Vrp9w8bcnDuQvMY//aRzznYWR9rq
UxLhwuKOcxD0oJex+wAPOHUYZ7KD86kCu4lGea/Eqf1qaYd8cD+mikb4luJsaudsG+i1oJDOAmzs
hVqoEyPnL/OCyq6Vxq613GEwaZhVkVn2VDtuKnCv2EWL+R1XKPBalOfH4fFvppoAyR/hBu+M7ZQU
OX/g7cdiojEADM07dVmwCH6oQC3l0JPjm21GJjFA3asHo/ACbIdtnoKJkC33dAh3gVbFPnV1QnR/
xZLVWc54SkMSIksNO7f8E/jA3GcVPBUu/iKfZcZnBErfbAfdo71ukOgKx6+YRB32A4KcDESL+prn
ZcCdeGrCK/gWTFoUGJoOjG31d+J+hWQlzJFcIjYPAdAdlF7Q4WY7QbPmxuRvbMpR9o0jT4Rkj7uF
P3liqFYNpAXBHwXd8e5ihTqIoP0QguAXH24merfE6u0Cy/E5tSMBNHlhhuaZZcXbHQq6LknOoJ7f
LwTiLYbv3nV/n9GR6wrtDUth1cuvgf49T0kpcQlMDGKUXa7IKu0vnKLRnlcKdORtic3ue8qlVLQ6
P0hHgtTc1dcFFikNQ1EnIg7Kt0pSu3ocIxmCHdE7868r/PpEuUelCFjvscnILjxm5xe5gVsWkXRl
iolhNZT/QpOaxLVVWaOw4Jr+eEWrajwIQcU9cG76bYTtZ3m4vnRolC5Wwud8byTW+wfxIESopJKx
yCczJcZfNEVTl2WMGZiUGJ7eORd08yq84yJ2YB5uxfOgzB4dtTdklAY3h5B8iUIuEI5TXUkP43wP
/ooh4ZbUWjM6qF0qV6MH+q3U2up+Q7Yx5IT1DuWrKXT5F9sDfa/bC3UvxOzxOn1iC0ASs97y5Y1X
fgF3U0oOmUzgvVJ1rU6Xyblt1diyTddrDtU38iKz8pEdQJ+Y/c9bSSjaifjEWwuL2mwpEjeEDzyz
RmQRZbJzL++LyD7YitlZIgcO6U2gO+q4sBQuijLxvG8fSM1o+3kXfut2vztGubrlrZ+zuweZbz0Q
t71KZuHl2az7pNtksZ8fNS4/urdSYDqpDIrl73QDrDUEZ4ybTmCBdOjDNCubvjm9P/tscm6scJfm
43bDWAHgdjuye0Hgw9f6hvQ0+pN8mc/mCekBqqaksgcMMVRrXWx7yf1jXOyfOJu7FgVG5xJg1JK/
7Cyymm4FlMkd9EMlQW6qGn5IvDYnXqGQThC8drVmCkVCOy5pwQf58r8tC8kOI1R2WQqblZ0x0t+4
CFosBcuC2rGiJsWCultwhdnxrHXgoHo2tkYXzOurmEfDNFA6oznBrzdDhjGcRuLGLpVVL9rGig/f
57FGM1befpmymMAiqN8KYiZVnE3A/LC6ssT+OuSIPuHIsSpwRxL9G9Yri8maCxJknSWmxOYG7m5g
ridWG2iMwZ5CPdZA9jhsa7UnRZxzGXo83hEypZtMZcKIiPzfQUosZojYr4X5DrvA08wgjxNd9bj2
enHiEhgkRAK94j2YTTfXhM3CF00bzRo6Ljw7jQJg2L2K232L2GojQkcbyBmDxX1nBjJFp15L4l7M
ZPNU8N/MbNU2k8tI+VjBSrZ88azaj0o/NoWsQm0mD1Wfx3FBXwPtOW3hfHlVbYTat45SwZFUXc3V
XEHu2ukfapkS5+MmNSF8kGxuun1lckJzPlHT9L8Yhnphub4vbOHCu0Hpf0m+IA0aiLsZvSethi3w
odiEHRZkJp4dLN2gGctzVqGcYVlMwMVlbkJ4t3K/Edb7s062z969urWUyaI9Kscvs5Ri+khDXefB
N/th9Qk72vfnRv3lpuGFlTA/wblwIIptSciXgTkK5E73NjUR4JcMiM4uRRHrYIGHGjzcpcjukAnl
L1mDHUTmwGfGFm4fAImUJfcG6zz/kRSn8woTo4epEKpRv24iCnOnan/yIzhXdR4nptNZbe9E3do2
SKqoee1suYeyNYLSDp2pA0rOrEp1Si/tbMn8QXP9TlYbtvWRakdi1fzo3/fDGu2onnnw23i6RNid
xK+5uYmqYC8DGD4Lx+GzFIpyH7U+3W2wtvF8M7Sf8S+8WVzY7zWbYvl+g8e7l7IbmERJoWyPZJu1
BzhDYmLpTgrjFnhBhYD9h8A9ySSPWgqD8zX9fe/KxwfgovyAzwr7XL1X+faXmyl40Gj+TTUv8Yt/
sLbsyz6qK92O9/RlKJLdsnhZmJbUHAIWlCPJY8cJiEpg8v69i2D/KMn8eylRr5sKCcqWOD2p1Uyu
mnd4VfG/akkXOCvYDO158LKhSr7YFo0YegGcTlwNlqWylV+sk0tdX3caLXv5T1qSboMzuqez7c8G
iaJZactUxGDuxLH8kY0LawrItNGYG6o7EUjj/XvUKuUPu1wyLRVgiAhIdZB3ikG/Kx9Cryk8KoeC
Rap2jv2b9ywFPJch51xoV36wEIleUUkVVJ5sY1NJdiywN3fkJ1ZUH42vvAp3OkZWVswYimIDEqtg
M2WF8M2IKEeShSW73rI3zr/W2GZQLp9Lj2qbGEXPXpLoZNVop3h0Ooza3qic0eoiVwSb53GPXKZI
zMxXQQ9XC0J8QQOvu5z1kywojrjzomDCxzQTVmp66F5cmv4O6I6XmbUPt3TnshM7DUIyzkd80yvA
KZnbLt3UaS7FmAtiY5mRevND3ZfI2wB+f3BTKIdHyWSUrikG+Is2SoCMipfGicBAPOLjNSJT1EgF
ltArG7EV9ZW9iWvZ4EsuUOnFq2WE8CZqZgj6hPS5haChYnZ68DRf6XQpTXpM6cXfxvVP664+85eI
J1lJMZuPx16X0dsIdEuk3+L+BETDPUeibvIlVPPHMGHNwZbjNI7ftFcio3H/7p4/Z9O24iETEs08
DIXssmKFeE+RItx7MPoDGJZUiM3S3BxjvZe5jwULW6nJcAu6Ltq0vjDsb3qMt+9AB+7fxHN0RosI
ktHUy11SskDpFzMNcQ+BtfCOcgxadCmP+fUY0mLf2mmCsPP6lsxueSBgGjf3shIVuuv7uq32lHsD
iw2V2mDrd5Y2fHkloTljqwibhlglwj36GqGw2NLcca4ChRyzWPfaW2nSFwkv51DeTtWTywa6j47a
6uumHOYkFc6c9voDC0rlVpHfZ7imPVYrNxsE7frKtDA+aJYsmhO1RhOblYhdhLHSfLYQCDhsEgx1
KJOnQ3hc1ZEZ2vbHMczSTxdpowMvSBS6kO5YmY9ebwCdY9vCVtWAZgkaa74gG7zuSi7Hh6ndJarA
jYLu9u3S2TX+FSwmXzNpyApdCM9yxwuw3mLTqZSL7mwzBYoqeSGg4eJ8wpl/MKUpT7IHTEJVNxjm
yxvlP2pFKtHTQWU5yoUsTyleKumNon9Z7uMh2S8c0tvvecRykjMBmq9kb6nmQYS//093cyu6lEG1
noxlQ1DFBVeYscHDXngw/nIqSY8S2LuhCRJi/UGvp8QlJHLbOO9i662kSUmIyLLGJcTDaSYlGdBL
RSZRTqz8vQfm8Sb+BwGwwsXuE3Nj7eY1EGgpgGS5rfUAuRDvIXJJOxdtCv8HsMMS6VQk4Q2fQ+FI
ew1jSOzfG/4dcoAonC+FR8s+wrIwZveDCvCBBsANMBoHMl+958E9dRGV2fxhj4ottq14DLMQqEnT
peNPVeU7QgFqCe0h69/1WvmB2vzB2YYYVZ4diT+RVvzHEP/xA/LDoJevtr0X7z79I6HKAN2AivbQ
YiVGfXZkmPeNTKmlQvcYb9IM330bEe/BIRjoloGHpSPH4XMgH4j80eDz6cgdP/Fs8lBZVtXkV5wM
OOejDETS+ZVZu+mMz/Ispso/MWqr3PTEqCzC1DGByuGOaFY5kgBBZUJoWTs3nG8U630e+h6N3J0m
T2A7DgI7ZSbwr1ah1mtuhurO5MSq9JWEvTHHqxvVMLu2LmRKko1zFUREu6gPPN8rnSLL96o61A8b
opNLucrRYkIFa8gg0iqSo+cFGSqfm6vHCznPZsS8C/Ftmu1OIZq75qWZL5PF9JEvcymtpqxsuyo1
yH+KoVXeWgQd6pYtvM+0g96D3FCu7/KZAhDTSpcaVy1A2oAbMt8f88quhOkz1srDAhMXABElPMAU
O6RWDaK0Wss4YwjOQTAX11CS6jjsVqA1Z8GvBtmPe6hdL55AsRzMOhxnR4h8yemjnl4Hwyqd92//
rx6uZ1KRfzaj1USC08fQ1mFZN2eEAbwIqfm67y49wde8MzVEJLrVtF+ZR/gqOpFBrfuFfFr7d4hb
mmoNkF5r5HOb0cUlvVMa04aumKoMorDwbgNO0B6BGYOu7jbBbwCrWbBsWqd4USnlv6c5vED7UDjG
Bjqa0moo7XjNT9L3wDDRn6READrTkR+FOD/2AhPZJs5mnWZZV8SghMu0e1LW/7KSj1hhD/KLEVEn
0t6RhVhskHHvqDUhkoYgr9XvGlMb47AaCprWkBg7iM+Ss2ceTxrh1xBu8ZTWvLbNVV6HReAUG3bZ
kDOjtP9A/KOQs26ytoUy4JQnYaUiwzSHodN+iwnjPeK6t6YMqIemooVWwrTB2a61bXQsj2H9EGML
YFDW2l5979XVOrDP/D3pNGVwfBVvbPjK+SHKyjmO5bb9Zz5elelJEvuI+iomjlJVRwpFqTWznFE8
zfpLBdGubBoNU9oAsd35QL/FKERqw8DWWVD6QKf8U9ReJBaxtgw/ErdZcBVB3l2cQ10gRFiDW/11
KHBv32w2laidZ/uZhcUWNpPYlyRA+zAt3bZPYvDHqvArtSRqHmIMw4DeB1QkMuovKE+MFH/S3gH1
cIQtdA1UNcJMcnKd3c5pE9frm2xJvv3jhSbE/Aba644qUFMyu1ceh9p0WdBBFxgi6Mu+RiNz3AL9
QdOA277nc1Xhni8Lu5STyJYAf21TJOwBBi20og6jQQDL5mpcnm/1+kcAMowO8otK57ea1kF3NyMq
cSDEjcoJctr25bjFJ1CqvzD5VE9y6gTaDc1ilx0oMB6dFwFpQDVdql3IDM9RWXpyHnZtEyoqBzd2
5HDgvWsPbKjTzJyP9zomu5ATVcVlmdJljKtO7kqmzNw03GIUWYsQU9JjPiEf7Ql+V+akcJDPBr0o
Xpc8aM7Szo+GcuoZDUhK1RDWHPCHbB6sSUxSumxJWI4y9VzG8XqX4vbYmIyfWgZXCb9dPle4ueYG
LaSVqwwcTS5QkGSPJAYW5kLm0ByApmkG8dl6l30W0aFDf3KQRx9vvGygCwiJgFok1hLqra6rXHbj
yxS3I1KGL1vh+311thVfNm4mVkDxUjqzK3z+Ed6cJT3jnYpgAa0DeeIrh8kn8nnGn1NtE9PLh4mm
xNhzFhctYOTA2+mf+yZ+8zhIXxCOzJNBOHQwynnTiqar6SM5ubREZHQPglX74MCfBbnuGBddmjkb
L4Lu0DHDfNVCmL1+dhmal6LgaKbuFZbTyoCm+G2LCZ72x72L1kaus9gGCx/y71XFQoMWZ1ZEV4W3
ImbjLN1tWxOcxHlBQI6MIIYtod6F66EUBbeeJZQqBdw3r5Usc+VGEn2Unj7GtpWI3STyCrnQ5Wu1
7No0uSDdLg0j2piFll3ljyBQLTlNz0mKDfbnByN2FHrdETjk8cNSgebJE0VegyeN+x4mW/58ihfP
2RayUQp6QFAb/PcrOA1tPC7gBHnGKiYXDKvVxr5RSIwjCBWT2qNL5UY7+isINXJkoaBSEx+bK3DX
KZuvhuCGeGhbcfNz2/xjH/4DsLS/kg74vw7WAXKIZSuDGxNMy+sWIgNgTIFwI7L9TBcJsNJjUtuo
34QR7ljK91jb/0MtQTIeTe6U2DLy8U9m9YvMNmmD4b6Pqu+/0WwOHYhlG3uoNXTof7GxIeTrB9bX
T00k3lA2Fm16y1gKCwPe3CTJ4kv53RxLGu5hZHJ5JYswJACTZXPbnqtbvGByWvnrsbYHJj9aW7QC
1NxyidGurI4CvyVzwa4+gEl9rYLLhIw8XDwY3bACArebVtOdb05+pAcybmhwtU/bxNeBwDuOMgqy
+UkC7+jASzzTbpYprYQRjlwJhbBb7btp92im9niM53eCz009uh0j+FgKOH43PQh8zNrFwSDI0jcp
aTVgr4XOtXZBantoIafuVxZkCxHrIvvunSvl45QZz0gSSXPDt9EZ7/ZxziDsiazHl+hu4tz061Dj
0FXnF73KYyb/ZNrzNCr4khfZcKuO1cyPKfcvwHG4wuJ3SAJsv6YkBz10JQYgVkGfI1ItgCn0Y/Z3
PmTzwp0CuUuD1unakRr/M/19uRcbRU0c3Nm/GJpbwDH3Zq42ZHRskBfeaZmbO97yiUnMllg/tBiv
TMAZtyrW/+MEeDWs3NiP/D++Yml+2B3l0tbJz+qZVkFQJxCQHhiUWEk4oxBH2PmrvJUWrGROjDNW
QhiWRFUFTas8Nk8Ik0ElcrT/7rDd/2CRQaF67kSXSXRmKht6P9+rp+PO3uuTPQbL+56kmWlBSIGu
FVy+jcaJTNJWcs0sWO845LbP4j7e/qJPb9HFXs+/2lXJ5qKzjOH8fDYWRbdfxnO47mgoFHGB5V9d
/WCMmpe1OO5UiB+GSGG4pB1prH1A30qSDvtDb9ybSU0tQ5ruRY16wogXXbrcU8tLoV2WKbvaMBJy
DTK/+Xe5XGlFecVtlvLLAytbx05M2gw7vDI/47e3fwAU42O2RLRgMEamEoys8n44ecwtKQFo/n2G
1IjllEFNaMDDIUpuDJL94AeiyROpWaJ/PN/cE1Z7Bqgd8Ns3JJseFpCppVtMzIJ+qLDFIg+D2KGo
rHbCc8n92vAKP9u7cph66ZJoqTWO5EF/xDJhZxXdYYW4SbLYJtywaWsYT7IOWJZrXo2WsKio3T3R
grPsgOEHIhix0rRl35DRpYK6Z12I3hJDmeI2xGr8cGSH6IBFJFPjj3FQL2ji3F9CumO7DnGPNsuq
q2j7FjiG9iOr+sO+jxU4WD5JtuxVe0dazp8YovrRsgzxpsAUbCE1PcRRLbKHa8XLSE47khs7ufwO
IYZF71qSE2weeMTNSFsrWq/H7WtSWDCkrXJ0lBTGUQ6qbX5Q9oX4gSlxv7l/x0xF0Rmxa01/R6gq
+RPQt/ONmV+uiaoQqGxBV50kbMrv1cNZvgVPKCciMg66CrIRdYor23PDOV23yAWo56LodmAcVWln
zCr+Wuc8YoA3uSDUik1WpGToAtl+/eDe8Bq4hxRVXf2fbQMfO0LU2q44v2rsXDGOc/Qqli1T4pY6
Z4cHRzgA7o1/owtMZMgCNlxJgr5OystJEAn6Lkk2qh/jWbV+GWTaRR30hDTbRpd5G9snLvKQMSKi
TRktYpm7WM5FREyYcc1ljVPv1Z0+vX+qoAHOBAYyyKLwAQT6uK3VrLP9GIV8yZ3yHIe5dybSOiqu
OPy1HHau/P7Z7TCMdKIrvJSs9IYM0zaSAqV4UYQV+xxQOkcfj438mpqlj1B+BU288NjzL4aHXe+0
wSITFms8YAagv19YYdh0ZzLTtdfyYQKRcJ4lrgeUyOPuUQDgqW9fe84+JmsERNKkU16fpz6FPY9S
vDmTnWL4XyuF78BppATSmr16UQPkVgF0+Aab28XpR/aFjeYkQ6CEKHqtPiMrYtjzrtUtT+Wus0Fn
uI7+D/QDG1xLPx7tz3i/PhDBcOG1awgRn4VgI4e4ELfUqEg6Ni9NjhAMbbPaWfEHHc88hOGffBDi
jw5VrW53sYUWoV+iNPHKxaVL8iPidHWqcFLQQj5NHXY8wXEGU6iENGyvq1jW7F9W+eqI/muSw/9B
fUBN+PwshgaqeOYzC5MRb8XHGTLynjsKOClDDypFyc7okUPDYYwGSGi/hqsFMUi/xKqY41Fz4+X1
sTpuE3zWYyh6kAkhGELQfUS/9aKUw3lXajuQo79gxN9Yjmll/tDDcOStZh84/+eqLQKogWomDDmy
qymZFnjAl/HN8TrH+APhPDLsdWSG3rEHqenKQU4ommo4k6csefxLpZRs+oj80hHInAeJb2rlWp5Z
FWKKsBPlbHb8ZI8+1jOCJkAOWXOH1cbEy7NYckEeNDtcBs1H8zksjxpoG09+8BmJkWM7GoUmmoYM
1UPwwoTGljlAKtcD70pqf1lkPVv8SkYS/bdN2pAC+nbBY3PUxqmVQoTDJjW9Sv5zUUao/zqUFTNL
hQWUh6fgUfm/0+kuzV7I+xd4SwtJL5sLPYs8L0909usCkJURAfvUVMQ4ky+yIOylHZOQfomDbji1
dv8y2L/GWcN0X1dwt2pUAqm8IaYYtNu1uYrsWkoi4f9uuYNQjrkSAaoXwY1Cy/+Bq1bvXcXtZVwp
UQ/Zo6FawVBLFJ17gOBU5WxEyTvwgTqQjYZwktGejsuGcf9q7px6cdPy8wqfupmMTy+QhmM577PX
ajNc820agU8do3aQcaoXleHB54Wuvo2PwrJLHaV6Ktg6c0Qk5R42pCQXGY/TkdsMnFFcIR0FexHF
Yv4BsatGipsYAXYdiGObEcu18AFqZOuNMbNqFy2b37cFdxvVawjOZWeKci2T7Z+Auekr9xs/rVsn
mVuBBoZM6V5jGXXQvhUi6LOjztlmHJXO/NBLdqiJbheIvhjzu4qzTuBK3StMwTvd5tKXbzT6aYNv
yrlDnHz1OCLnoaub97oFsreOiVT9KMdua9JAlSAgYYK7Gi4DOTcnP9nl73AEkzYPQE79qGt6Trie
o/CB1QjV1uIih3Cn3zJ3RgAIjPwCBrqEUdiiWgvbF9SqNbP9XFG2nzoeO84UlNId6+0GR/+bft/h
qgOcGv4j1MHrtSD98fK7f/qvdI1Ymt8PygEuZ4wIsOjslvoipqOin2BGQl6TnPafdlnbeMaL6PSm
Ijcv4v4WLcB1042D2dHAJWhQZgObCD6KNKGzXZSbT/VypXU9qiOsgdxoIKFN10Eb0yZ3i0I81pSY
rIXsoqB6gS28bx1vI30c4dV6KX4AE+hyJGj7HAPhOczM39CuFYltqF288q1TEtrJAPZ+xZlBXvd/
iRvBtEmy0Cmq/8L0VGxVUVGuRFGolMaQdGY5CPmVaacoLELDJ240RCImMdCLcT1y9T9d090qJAnE
9Oc9Vwm61yWEVztUBz8s762lxtfLG4OYP6MFLW30jAZ0fYY+8Bx1FsTlwPyjkeNtxZntkvS1/FMF
kxt3LMdHP/cG/srrogC1uZfIylgvjDL0wajvum+D7kIL0TkADK1pISyP49BFNV8EG2A/TD7TkKBK
Gy24v+yxsFRd3pYwXsXsnnehdYAQmHeVIitRlM1Y7fq4CsgJx3lDPKDL1m3D9kdgZdAsxiKMXsQ0
O48vFp8FuDdofAacgCgv86CZH7DM81hZBQCANXa5v9mPWtF4Sm2O/YpIvdpEB6aU3V7pclGBayM/
E/CHdO/xDCX0SEaF7PJlkKroB17VHfLjE6vaKWsXR1wUgGxVbAfGANWVn/8z5EYPVMfxqBAiiwLW
bZUy6860/LSlfT6LuFZw0aum5mg4daas0ngfsaUVJmZHOlQaBlOISyot0WVUJ/lLeO+V1cSnfda0
QHLHuwV4dqvU+biySUh7s65fX3e6a9kwATMdr6pVjXTPm4SMKQnRthbRXZIs/VTVNKs4Zm0jWpF3
UHxCmAI+Hiyfa0QVVW90MDXaMskwzrNYW3QDSEzM0egRmYpOpiYvjy/CP0YhH3bMgsWPl4n54erP
FZ4G12rX78rBWw1F0tYJttjP1y2ieQzIYr78iMM8YlBy0zkrSoD89xT6iLCtNUYx31B3sSR/v+zB
sraLZEHaL/Wi+9tFrwzxl6rvQ/IIo2QtIJi0R7CFWm6/TXmg1PJjfv0fW2DRzGA3mJ0a/BVbxBZS
P5esgEoSNb3mKrO170FYyjb1wOyrYlbrA+ArxZtY9zsaUaD6lbMXtKMQ4LY8Qbql+Yp7aofdc0qP
TMtMYfIfg+NlaGXf6d+ccOQgVKwGOhsg7cFPRE/LXYug/JATxkm2cO3ClZAME1N1uHAm6sEreJCL
M8rc0qp+4w6n/3d1/c4C7cr1yyNrooJcr3OaHzzeasPqNYmsm8XofVVG0QXhsSvC6toVdPxiefZ7
xU38hHjZ6/6Y57bCoev8TK3JgF9EF1d3wZ7JaeLp7F5sEnn34jJMj/uugXlAbWmDoOpFAzVkNXMV
Lh4MFseBALVe2MhgWfNP35qsG9uZDRudIBhljpNThbmi9nNnoCatq4cd/eW8qh/dVJXpCVE2pu1d
lkzF94co61OZalZaWdP1+ZDlN/PORJnRzff6lVNByF84x4aTi1cmUcbVTG6zRoUvgfUSOUB7sAqt
1XLt/D6puTs9Jre0wQUSccgOiGA35SxNjuG2sQdoVzyzmRM9vNXiP5yUtbTfrk6myMRIp6mq1nfj
oLnia7E3Ml36ZQ+Irslj4mo1vVZMohX6yqjJV97f5TOnMCr2pY1/8j7UekF+qvWUpgdvO5lexdQ1
pxv+IX6nkcQg6s8zjXUuYqVRm9FRK1wZCPCbeDhb3XBu/34qivRPkNJONwE/mjG5Bija+H9Eg1zm
guQFWt42wA7EJe/dEr53xI5XPPWOPFaIXFNqkIoPSMcxoX8CgFvzcaO8tyqVcIXhlDYQDw1bMxsW
fGzYwKMBETWA9K46jqn7259NKCIe4spAvfA78ogXb731HUyHc21PREEN97U0Gduhirn5Hpfth/bB
HfB98Y7cJfxhaRw2Y8fulML9By3w+Ks9QOVCWzqNhtulDhMIUH7Q8dYVWT6o16hG+5FMQvJRL+Fl
trisDBx0u1Hqd705uhdoWDd+uonkwgli5YyLwO5CnUdiD6i76aamkbf7y+9ALYW4vIkL7yuJf89D
g0lZpkcB7UWiUTHLitswHRileKnLOWbQtM+cymmhL3T6ebRYbOgEqPW8MtPvzktE28xA5Jhb6xv4
Qv88T3JizVk3v58gIQAUnnxhd1zGRflU6RAc+FbxV5rRjeSVppWzKPCcVqgwYaED56ALsocyjL/q
qSeF372u0LckAJdfUKaeiwRUNE69do1+gRM0Q7+PPsCOcQnUo8u7r9vHdsPsH+hm6iMpIPG+7cCl
qgDfaDpFK75OgcYpD7IiVa9/2mhLXYx5wJDL1EocNrQwrL/MS8gPalJY6020b+697v0g36wZT3LS
yRN+SJuxVdjO9PbQN03x2zNv26sUY5loejaOZO8wCE09kMYY3sISwN1lYw+L6wfjdGrLM5fYzfcD
uodtoPhDJXOr0vh1vEBNklJfZc4Dbt62AWcA2T4IIxcD17T47Ae/woZ2j35UjKnAdRc2l5AVJ6SU
3LXWtd826XCb5Fyuj2j5oiSzP9KN2FspB/dPfWC1ZlTmO4gRQ+4lOB9i1EPxVfW+CGnCIF++FYes
JT7RakWn/FQykQEUnBMAApzEDGLrg+JwbNCtDxk6wswW0/4BucdrkyNQ7rqPZwRTacnSCm+klJ7t
HYC8eTceC20+htkIfeNKllZRysHs8za+n1Yef3Dlag4+4esr52lZUKDEyx/3+XQZjKJwsocfp0fL
+NZVbzs7P2h4hWqVSEhOiWSorhGGlFNHZuZhfcdeGwzgxbXElBiz2WTFWEHEVcI2SHmjdS8Aw9wf
SztdQTePJQelergO3Mmw2dld7wsToHDcyzFRZjs9N19uT0u2IfitniOJ0Zdo5pDvhr1HtrWlI4Rp
DULdoBqIeKfe97+5OfQsp/Y4FcsgiiurD2c4tfcFlmYakBniU1LZvgRvj1Tmlup159otAh4SvHjn
NRycIP/zOT/Y5iXyNa9aUWNdBwGXEISz9fyAhB4Q0aAs00Bm+p3CUjEyV9TyR1hWJTErsdSH54Cf
krFgSpr4Ql33C/SWHHsJ/WzU4awnpvY8SMbg1TnTVmSFMQCb3yGYpPwXUGDmpX/NspD+TEGX5Rcc
SLcFPVNJJjjtosXvW4+WoS5dfCOO1DXrTYyg8/LNDLtIHBSmIC6/0BO/wcFpGwWI34CRTeFYIclL
OaFNbjHiW7uZUBv8aRg+kkpkmKwFx5XPP+SIqBbt1JXr7t8YGuRaySUTnH7CzYpLgQd5OHZ50lzS
cHzayo5+XfW5KtZ0buoRalmzDSCSb7Tt5pL6dxwVbzgB0yL7V9WRqrgLbw74ezNr8crgMZk5ozTG
z4oKiAk0E2lSl+oSkd2BlwMz0djs9yZXQ4t0qJmJtXmhUGhLyuqcZ7Nx3N/117mnKW0rp+Ipvgq4
c4KA/0EsiEQWFFTU2pg5Xi/dhbKF5LCciowQGX0j7HMhh0wGNjEqljjIgvc0RZgGaeWXsDhPl+Hx
gJ5ZxqAXHy6xb8f39GdrSIt9gOtHPwJH+VyfogakT9Uk/PqXrmSA+F0AMYrXcs+dYCuMXR4ROq9m
JpaL2UVrk9gMMQ/OvcfDUpy59Tle5P00erqqgQR+kyz4Le/sFmhd/xdrSwH7nNFC/8KN7pbncBLW
H5fzLccKEJQnOotOaehlZrg1yuqDR6BNjiTu6zH/TbIkbB9XoC93igoGg4nfRFcEYcT9xkkuSqxt
lkbnU+JDdMWq37m5HirsTmBezwsC0yjDTLtvztXpiznpKk/hVSC70vPLYrgyAtxI9TfgomlVl0C1
vh1zZtPefx1F0cpQqkepcMvPF6fTRlISGCxzqR9IBHHqwJUxeQXmKqBgCMlmZfD7wEcFiYvBEbPr
3kKJAxrS0JLCTis8a9aca8P+9k9KvLMvzTFOJl36HcjMjHgw9LB4mB+UEUr5Y9gkPMo34orl6lab
nrAgdvWR1iBUrcCksO+gUcdHCl8vHyaimgzxPoGEqsLjN41H1xYJdBUT3w+HSwRBfTRsThEi/Jjt
h10x42AJQsN42tADK+cp7yM9vvkSYc2nYaynDvQMQ4S/15d2uJLDVFhPbnoJs4ndahv5/0EVwNpQ
0Jov++xdEu2wtst6Mu4pITeQTXjQahCovX9noFVQ8BdYTQ8lzH1iNG8vEjCML0w7K/fa+sTd9J6E
lIsowF9CSJJ8LJSexbnTlQ9CLt7E3vwUfm9Y/qOUsePE4bxNKOAdrJ0iT8GsBoVbarDpIFHdAv9M
DYGq5s++8Rp4ZxJOAxNU5ESTjlcQiF+sG9RzFmXll6z3yw/NLT7nxp2rxmRb1RpQATjTAEforbfg
5h7wyy6ARHh5aazYG6fj3QzFE/zNBeOL5j9O4v4pzHGPgeBp1yigM7dymukH1XDolBcnDXxjlhSi
g6DZA103fsma4ZCMPYMlueB1HkIvw6+j6YHywGxUKSsm0Fjp42XzlHSMBD3nctAUB1Fg3r5b2szM
HzsnfzcKpXtdWL4j5n8zgDflymkA5YbEQfuFzmOxpsvRhiAg0+xPmRaEKKopsSbpih4JnniKEGC3
amqbIY1yJJJvTDpoP2lQppsjjI3U2Na8OtVBZAr94awByT0n/CDEzlCNeDUHM/KA7GkOoS++dOJp
KfERJQmiLuCTqHMTY8ZXzv5H/GE460kJl9Ku3RmJcsDwIUsa1ULuxWctpmTfpsNCmr8MA1lZ1/Lo
gqb5RKssHPVb3+xOxI3TYg60bM484L3Ys0+yToGKAAEfhLWUSkYEdDPjYvcNl5iXUAZ1bubH14Fw
hDRHi/v/j2sn+0rkSlkzZPxx/WKM6NbT0rfpsvjtx7JL4dqxDTBIJZIGPoBgKS6wF/5cQUMmEs1e
aF9TpxB+P3UZjzec413CnoWaeuC8aKgEgCNaK8LnCg3tjTHPQ8RW+c2dVpbKKP8ok0vaBzQK58Ze
iiXg4iOSDNSlnyYMY+AkooonHEVAoWygaugoZE1mZijUIc0m/yWE8R7AN13/Xva805RB06NtjXBH
xYQ69/L/oUC2IbPGSw2ynWmtX66cem0a6zP7Hw5YkUD+4KcuL93qA0JgUd2WkiNXeFxwwG9xiJXE
VN5zDG7bScZeluPznxtTmHC8QKymRf0I0GYA5UzEjDYUU5AOStVbi54Y2N6jfI0fDUxV0SrM0TnK
TVSnnrB/OU63+yAnW67uTee+xn82IspD4wx+Ia0Qbz8psSgXsNZQe2OYM3S88m82tCAZOfvUm1dc
HdoVz7HYRoN5M8NRpLNrijmGgwCE+FksNUbsx+aKzwhzU4pHznaVJCOQJI40OUf4lWhG9c6kAFbe
VcktSWk+Frsurd9sVL1PSpokNb2Q9J2mg0otYbrA5QDWX2xXhECVmLJQ+Kh++RpTXImZXkElUJHx
3wBL2WgEDkc5VOFJKNb67AEtaIjwIalLUoAZ7ufQDSZV0u8Gvo63hbgFtSVtaSaH+yEwyyLyJhki
NDyfLfvk5PGvVCo2zBIN3giY016/pLfnYrMFcq5/f/HmhgzbTe6gZXL6kXpZXGKJJrgBFZtOrPk7
/D4PJWu4lknzFg4ANeooLRqjbDTh2MdY/u9UJxuoEJxjMYpaDxH9tXPDco7j/uX0u1s7veIgZbZw
9oT+/6aEP1SBMqkERYikm6bu7e9Arz57QOr3vNq24dyTnPNlLpkWj5lBNqOKScpHBxLFOx77RuxZ
kNNaKktdj6zdT7cceEa5BNlZrujc6xvaM3XfYmqddJvMJqXaiM4GqSTS4eA0HAtiJvpQnEhGWQcs
odadclK9sYEHyatoxFGDtQO1rm1IoXm4qJB/gahOrUTxZDwm6aULG/097MkR/qZym5oYD0WMhqQJ
MN35IHk4zrCzoeuJ1NKGvjVhRAqCtX7BkQgaoC92l1tHZhF9meL/xSWuaVbRI+QjaaAt4WgiWAW1
ngbOJ1ng4xrMvXrZy9U12k19NAXMYOr2Rjn+ZagII1TSI3MEDnmpjEXAfUtjQZnpxwSk0EwADird
DyO/QvgSc78wY6gI6rQ5ndZEaToh0xHfmXEJhsj/YN1HU6qIKdmpd9wrOYlEZZpYtm/35alS0MSM
0fUeT9W0tKz/9yCiA26O+2k+/E5G75uy2Q1l4TeFOQKg92ddLXgc3SmYGu55NYwyo4L4ekgwDUHg
8Qm21gzt3tvLIrzrRPHM0SpPCydwyXjdLSnd+/qgDNpqaBckkLkWnxkvfd/Uxb9OCIl4Yh2koAMD
sfij8Wo50zgjFPrGSFUO8IXzf7LEE+/VwJGkPeba56uphPVmGn4gg5WzC+5QZG9EpxE7h34zmuyG
np6N2deR+tZNUDL9CloPLU3K5GlPQAjD66DCVXzQY8LTGtEb49ENY4lVmYqkCTpOmWnK/bONoJ8F
mUD7OTg/hqoB3pBMmfWc5wKbjAoh0fNoqfK4VMvnn1KtLoyF/jNmsx42dSm/6BF6rVK3eLRP3Zm8
3yCIWRcRAlr3NTCqQgA0+07J1InZo2vkJSOdzuhwF+dEF8F60SEWDVIg6EpXf5DUQSJEzDMc+NR5
Wd76HYtVYww+BKMfehPT28pP09jwsDyY9Nduo0E8vXWYLgisaPYJc7FovubxnsYCMfA2HaYQ5RVX
Anza0/oipSPR57OLo3Yq38AvkHuQSKzwV7lX9HQKivY7ztdM6LVgolX5azFGECk+6bgmKNyDXL37
aqsh2Whvrm1+mNxCGf4muKU3QQbrG+k+DJY7/8vBoHhYcPGGtVmhWDbtRIyLrvM4BVoc7a/yNrRm
qBgAX3Gv8Hfzfy7I5KH8wbYrcx63SxfL0wf4SQwkHBorDWyvPQzQ2K0R+p8rtedgjCOtfV/20eMo
Ih5+YuujD/YaUvWtEHOq2ybCyhEvqDlRp8CZM9ZYefIjRm7IFrjqyO47LdMzkAME/EdleLl7mpGA
AfXkK8M007EgVy0/4hgOxyMkeQIJdeEmsmRI7SA3oCTt3Q4FgO9wk4SSv/QH5FNR3M9gZAWCdNwP
w0oAmRRzM1HewA6yzVdyw6daYUJs+o7TDwTizwrtzQhMvSLxHZXVIN8ZO7fZy8C08QFo0RTvNPeu
IctWboFdNECKgbXQ2ov0zqrORYA8whxwRCe2XtI8/snNFDTc5i78ha6MkSHr6SiRdXt1l7b4Kh8A
0jJtaWJ/3BHpZ20aUXxXjMfXgrvkDgITwGNa7WDQLX32BRcBp8JCmjqniJVBAG+rOkv5rASzvqc9
x3RcJa785a9Indu30qYEbJQTQ2V2nV2tnamta/tAKpaZ2xd9wJ0damjFLal+ripR3eoOHb+CDF2g
/2MJokwbtUmqnz0M0B+Rr68+nJMK7MH33SXRdTeO2/GrCpzmr4F8OJ1nOij4ApvXD9psBSHHJNg8
iUj5bxrObAMd/D0wG649qWuFp7vMs7jm8lme3ybRqC7gZGpVSDvhhjcWnJ6C9UFCsYJVKRdKkxwn
pi1IoedPp/9kOB88+ZQj2FphxNVU96CGqtDpE/NwzeHFuNAR2Y9XZ1I1sGLl3wpwasTk6Tj4q7/X
vqB12XM6M8XDQCjUPcZAAtAvmT4yoJyXBsaHb5jUA9pX0D44KF+KapuWvH0u6gLH+lTTpvrKQr/i
482VpALzMU8LdfBLlTUk+DCinZtA1/3A23KYYVJfpLpgmNUvRUV6dfE1BwyjbZJpJXhKtnqjpqdE
WfPG3NM92v/3zFv9s0yBlSPZWJicbOnTvC+ZtkhP4iS/SJApfH9nLDy4i9eY4rAq8PCkSsBkarB3
ubf+sVBcKob1IEqMMYHplMuSMddVy3SaPZB6dkVulo2dFPjFxof/znvE72zMR7qYkGwthZmp3KJd
3B9cGPioprAXd25C0vCYHoO0Vwg1b9NC+U+TCLPgpj6qtDWkPLWMTRtWReDHEj1gaJV/CrTFzPs5
mQtFXhwSNcIy8HlK8hOMB/LuqPIMvnOiG33hWApSUxam6V/Y2qFQZ8n2KA0YHPLKZWPh2VKlhe5O
7obw6Ul+GNSTTt3rQYrzDDjkl3tYBJJjfkYAEyZDA83QjipErdPwslgQy6/535qO5DQnonL8fimb
b1I+79vwLBgUEuHTv1lEAKcJA1B8iQWAAnJFGkrQ79hfSMpS2ax00f1cKtXRrNl2lUCK9+BWu4Wa
fazps7EbWQqh2AcrmmgPaZSxJF/o9hWtYpoG+gdBevZuj4NpzisPlzX4BHm8HwdtU1Iz2KNZ65sQ
GWGhThd15gsW4yovz1nxBuu8GWsnBCegL+UR4bHr/U/FKl3ogfBER8nQNM29AIsFp4CS2xliyQMX
mpiU72aA0rIFdXOGEn+NZnQmjOk3mRePu0LJckqsEqcDTmyH2R759GVYeedvEjVudhhq71p/vA/m
FeXObzrsxagZcJjVQ42oUP3o3snzH1g0k0rfgF+0IwbNdAUsqbjUuLECMxWHJluOfP/+7rBs+D9O
SxRUprIJMEmf0BSffmFqLU0gUkdwNRwZC23Y4eQ9Pew97WwrbaBZeo0OmWG8om5zJtoEWmXbMx8Y
mCW7bXpSjjrz4ac/ffO2I408g+ommg8+3yu8dCXmk0n9wI01jtCP4YzrDKmfBCS4buLWnp/VoFIh
9Uqj58w0EhKqEogl7Q0DE4Wa798W9/OhZRvC7NC6ZxwY8JuStKJvow3y8AeYIHKtKkWqjfAYOK+f
TMOdZfzLMJSzGGvHLFegGN0gnpIZIcD1KncjGVxfdJukowqk0IXJNFONRrkZ4EOat/PEcZxLhMRt
Qm0cbXk147Knj8f6cntOhWwKNjiHV7HMpqZ0DBEMqGxw61mSKFimrxOWpVRpH2vAfVL0doomdSMN
tUxuh0b1SCK49DzZmeHs5G90z/KUP3/Sa9qBmDNDS6loffgaewtM5hEoGzgoCHkHyoXa1Z8WxOnk
1LMygrP8d8OXNKvC33YDZPUtt8wdWDVbazoltkUl0PSTgrd0Mhovoc0Pecno0GfB3+Baf4Dq2xW/
jkEYg+mMvhILGZm93jxEWAP141tvyYRxYko6NVKp3SV+jjm41lh04LEPCLKdLWU7zNPne0GBCgno
5oPUm53ajOIGiPEqVeKMY5EOcPk2ZiEwnn1mkzV0gNB+QqY7w/59UxDA/wCcOu5AbNgTRQN/IP92
tmTuaHDkEbHeTXQwIpAiDKZaQeo+5gqmxurigINKTE0dGQg7R4C4p5F3ZQb51KdMRdIY/nLqm6+O
83hBaEDuMnLkkIuQZuTgCq4933xgy0O7La4Vbcqefs7f4mfh3kI5v11/3YT61krFXI1SPPJ/JQnA
WwOlhJBKXNysB9rD8fgoWpCkjMgUyMJkjPqyr8/0mr4xnVhxQfBaxliQRqGOnAQMxlwbQ0r9nugo
T95XBDYSRZFelDAbOoOyEadPi11lIrWxUM+JHnJabK2Z+C52QZZE1RgZKAsn4LqE+Fy+5fRPFE+u
sPpBqehumug0a2sCk/DHcFv4u8lZEAZIKSk/5pmf+5K0oIc3ZkgVKUcwHfVkF4nRI6zsNRNyQM81
YihlmXo+A4xS9qasngKmWjtas98UMO+HIPU1mIj4iG8v7qgmO58vv+r1giIhKgxlz1hkMTaJjBg3
EJ4lP3XGGuurb/5FePpOq1pqPnSFK+RCTznNxSQVuo/frwjYYkcI3+Ba4pXyus1VgTzFslnFzHan
1Fh5dPLgas0qyffASZgr06MfcHHnxddkQS8sDYeyBWDMlt3P+PKUBxzCj5ou2/CnOF2WecNBOMEv
bNRy0tyqk7RuArk0Ppt6MaTGepV3EmPy73c2XgRbo3anlcTu6zwnW3s1Vv02MdFCAIuvHAMxUD2N
KrIZr/oyzgiwgf9gYGWleDmguyc6ALRjlWmigOXRn/nDUk1LRyX8ySGRLtTyHBHzT7dzbRGkMjCO
r2LQAc9nnRdQzfG960WjT04Dm6FZEqwjo1qujYsISPpzHNHBMsUx0HX7UpN8QnqjoALGLaMdwrar
oI12neuH+CwKy78IwR3qsDGeNy+ls21LRqjJC78vhk+l2eOUvutArCeZDGR6pG0wqJxysW/GWZG7
C7X6qtpyQ+rleAfVhtDf5ynpOx1xsJK7o/VX2joXH70PqcBqbbPVU51yb3qWQqbCA3aCP6US8G29
2kNo66/E7rhTAxE9weHP/xuFOwrQ0PNHX1yaijq1mUJOuidUXomM9mB3En/iZC+SCBp4VXU8Vn/Z
chBLShXppXK+5hHjalSlwwa94HQ1e6y7W7NxGUcrFsQmukeCbCI4Ib2i5whgFW6R85NMt9pnXdpN
08Xg3xH2zpJgYZbRSi69n/IEKOMiW7CSK3j7yhV9h0eh/V7NCeds5Qsqv4LYKg382XYirtwG3E2P
WDZlL7vxlN8abKoQiwaWorEkVdHC1Ion1eWBedJczMP4sfDpkLhnQzcNvue/qm6p6TwcRyCB98FX
P9GR1eJZfh/gwNv6D7+sUwzwe7dnUdhDwYF+WD6+lkkHWl8w+BYved+LtXZy2oHnzcOORCHbvp3h
oQRJSTfgPGHzPCNGyvW2k85/cDkLD2fV54sZevDRT3rfcV069iDmONiEey9EqG6kHT7XlZuCwwJj
i73UPcLmrd5DzDkVto3867Z+G1zs8BllNz5YGkxCnzaYdUbZKVyAC59/LK0OTQ2kUpJrjL+yBglD
dRsmLMuCvR00ZaF6VEJa0BPQg/QxUqlTLGd12moFLS+4pcGe8HAV64F6x8uCJhrQbh/pPZjrouCi
XffeLfKf6r5XMYyO0YOvGiAs14oci3JW4MSvl92PFVfM4JrT3JQFSpi1CzusuRo/VA6Qxg9FQKZS
EOm6m6e9E0RYi8xNfOJv7Q2hkxo+miNtkChDOhZpge97FjxwWGTx+ciEOv+mSR732xdnfyYawA1m
n2jz23ccIXHxzBvRnxkfN5cbKV8FNSHbi3Fo6EHaGcfOZUId68UVHw3XKJ5MTgbgoT52mddCm/sX
OxcDToHlFRSrB8rvYP/CnYY9zvOOH6A3DyTcHRxXrHx3GaECWzpMPI3/XYed7hvev9/oKDdgBZl+
j7XG+Vl35+rttj03nO6dh6Jkzcp9Elv0wVBCpgfTYWCqMjAOUhurH90dABv0csPGI6Q7QOUHAGrB
23KPk/xUkQuSV6ZWbOyxp69T+WNAocZNpyf5Fiz+0eZ5D1AHxd3hutnAgAT/G8ddl4fxFiapfgXV
c9mzr140GRywV+fDSZFgAODGaegsr39ySV7LXQbYWlejuc7fuPsSvyHZCMxBBU0cvIdE1/v4I8fI
VhvHGqPjMisbYOPbscTi4H9+/T620CgktvM7DjGq7pcnNvQP5aBpL7hr3Zr4bfikA0/FB2XhOsFj
ugKYngFzc8KXMEC59k3rILrHdeaVK56zgDDcPzv0zmhB4rLMiTYYCqe4GUsuHB1pBo8I9QyvvwPs
aqTULSLuK53BymIQ43zzoszzEIGPzKvrHwTmOv93l54aPNPBgA3olw8CFqlmPPWDUibclTrEUmsk
HtuixdBTkbbyZnwAq7HUWLR7Z63cCWA05cC9/u2I86Ab08KyPBYXq5LY1wjStDQcUbrj/UsL76Zf
nTqcnN30voKCRufOLLDq4uNTXXqG3e55OouGKMRrJWYsaiWkqCUGWvN5G0n7vuBBwhKeSoyWYa2R
vHtYC5Ogw0mJn4x1kXWKBwYUnHKvs5QiUjfgmEkWt8MQ98pDlC2g3lz5yOzGqKFyn42utoI+9O9i
vXyB/RThnWnfXZd0Dvj8lRFMR8jmSFJMnnzbd5H9dzBdF4+iz4U1sJVDmKS5ZPrDAmE3zravLCHD
cR/BbqHEsKprcFbmEU6xcMCwfei7dB/O/Mgr5ffeYoZT1x5+ta/7kHYp5mzAcuw9dDtzffgp9IDj
goZAgOd5U4tehdrAyCQj1/iofEdSfsRU9wlwSv/+YlAz2wyM2Yr6w6aTpNxZQtlS/WTHQXXBjMcV
Cjwjim70a/DKsoD1EWkyHdVLoXx1smlx8Afh4FeROFozYZHGHC00uiW2WiatFMaPKHFUAwjxXuL+
lWNtP8tbxDbG7iSK7Ro0EH2R87rKOQg1poF3sMRVvpFsOwxyn883+hcsd4m0rXd81YAC5kibzW8t
mO71CoC8+alD5PT9Sld3RRMNAJ2QZghFPJ5VOLCCRPG573COMJZnWticCJAuFm/j9uOwloR+qa9+
LXFup+FSmeBTN/NjRxMjGy0ATdc3dHcuUJZACT02phsGg1/0Nh02y8R/5KQU818gGZGN0vs6umaz
JhzfgLGBQt+L6Yat0mzw1jmAEwK7obUjGuVdZiwiNimyiwOrFXzVprmS71Iet+TZqpc8n4im2RPO
4CjMSxul2nSzVSXAgkPNovRvgE4+AtcFnUkGCXpxNxVeHAOE6jRQPFNB+Dj0yolDNbrH3Rijzj/b
/qdigRX46RZM8qgWqcbACvjOengY5DX1jbAiP3OZbVcnW0Km//jEju3ggN1x/kGJcYatc1US37I+
7mS6dLNtT9BOklbQxfnUOK8i4dPalUYjub+NYIWZTFVkTPBGnUUMQ5Z3p1XXa5Ep8fOrx+gk60hD
nfJKfLDMkZDUYMxtuy/ilvdvc+PBt+1T2dDiHo80/ODtvpsd5Z4khf2tpN7HsG5N9nojmLpTBPYC
2c6Ldu3GcqTr2J4U5TG7QiTSyyk6U0vfXpliAZcoM2OYDY130zROU0kOgpTxq+gWO3K5iP8kH7Es
+s4aHdBkL0MZqEkmD69Y1Z7aw9gldLUoD0UCt/H5AHcEzuR28iMZ86x4Jc4IfZK36hP2a9KcC/sq
PlCpCf5CEENLrNhftnH641C2ztnlRSJoWmRJ2mtTIdPy3vWY2aIED7uRitAuIn3niIdwGO0b47tU
O1i9L/6pRFCkU+h/ue1BCkP1hrB6gIpzFckrL6NGFpEkeOzGD/Vm/MbRZOX25270/7MWep3D/XDa
qHTVSkMIX9uC4CRtuOON0mACvUl+VN1JFXPinzg6ilFEEJJNN1Fnp+RcsedcATAi8r4Imhhiy23b
9hWC5Bt8QckycGIkzUDfGjuqh6t02SouUdte1XijX61crgPeS/doGWaKKdRkATgNzqe7/Nl8be+x
2T5jmLwH1P4CwZ+92ESlh/MEGmGP9BMXG5iVHFxwKUl96Po/yi8EUXwbCkGPvEecHPLJSETEdQEY
lgBkYfVHyseBZ/kef2fXRQ4RlDJKmch54QKcki7GibKoDEz+lkpqOCyEE4nsWvFDQ9gOiuHjoGsz
+H8gVwqJXTK12JvBYdBpojkhBvjVGgFnm3r8EX5DRLpeK15JdQjaffcM+HBmJpfsqsHTwqcK5KfG
49gUEWMDoIf/m6nE5a+kcnx5gxMhHOeJs2QgZOggaQb4s3Xz3Mcf+37056Al+zQDfu6s3VmduldL
/8O2/lZ12uE1MrV5bf2xdXsWHwZmxT96izkDRJMLNJek4R3Q7Y4eqehvqSMP2qG3uptcAdW8Aiu2
hezs5BBgQxN7PV5fRGsUhELRqVAClD3XOCVHCHAykZCSrjLZ4YudBh26eYNLKzOvkhm/hZCRPXPL
VVv6IZbCyX3jY0w0jAZ2LaPLupKpM0r0KRhOolifZInORPXx2COmL4lTcynvQfZUhVzE0zPDjkFL
jRNXOaGwizW7x937DxjeNUBhPl7A8BKIHbrIvD4kzDzGPr/FsEu9wQhHohP8neiQXAxQHAsWZpi/
G8aAL8zrUn0A5Hg3XY9irqq4CWzDeQN6MeLVR5PzSQmvBtnGU5w4rgBa39XxVbmHd+Jp239Bvnpj
Cf1ezymrYTDqh4pK5myAgNZ6MBwS+O/TZutsA/SWWoah/kH/1n1lt+53eYy+0FbOJe31lEWWmuV0
54GolAGsjGt7FJhROLlJvdXgDwDWozgfXA1caAt9eZ9Y89gryuQXOtZmjEnzbMB5cEgPE+6A9AgN
s1pQDOrshRZE6dPn1r6V0+AJe+4oBDAkTB9FHkHZ3N9NqlB9dBSzuEn/LC2muCodcoX9cyXC9KiJ
rLIcjzm9ISoU/huuSdPDsaeWkIi+QGLOWYiARL/96W9aUOUi/G4jo6OlciPwYuDl7aV8bLrs4Cbl
hUzs+Bcdw/Yluz/rFbvK7pqIrBuThsa5B76XsYdOk5JUMur70S88DE3vdWTOym4IYE7RXA3NKxS2
+WIM2f0kLXwGUwVrfkvOdZCb9rMEPE09PWttKgyXWHU4zfyB00mgKTLfeDnP+W+Llj91WAuafLkZ
yMIR9j56RavSvAXlV0GAVbwfN8NWDxB79fdzQ2tPfvUvwsstizgxMzbmsjEh6jd1CSbeFa2QZhMK
cO6lpF5iJ2cJzL8BupVcH3QXI8+OiGhDcKGiZm35ujZ9GNgZ/pXXW2ZA1s44VrO05kaA9AbbCil1
E5vsmVZaBFJtPz+iJDGiJ7RU3cbvdzz1BaWLv+JhCQuW2lMufGQjUdqPGQhJ03GtW08+sjOr4DHT
6SLNoFrr09EnDykHqIUIlusw0TLR1B8824pg9Jc6mHorKvwGkRhNi/MC9MPSZqL3q1BtxLF9kIIf
vOAl68FnMfUlmRCyG6F3MbJMuVfwSbB0Y7rizwLJ1yp9FmWMNqAmPDWXT30OpkY+qkQiV4Gqbj/F
/4IhSgiWBw/D6I8kZiE4Pdc5NijdrBmRmf7ST0AEoTHfLaskM9+AQOofRcEUx4xk56p0QGJw8A8v
vurbmKhOy2XwN9pHl/2K+6J7vK1Ts5M5UwUXQDobvfa9SfL0LdNNpndXRvA0mcyvTp9SEIRXllNp
JW2GIVxXgFfFbQfWZAQGftQ7p7HLk335AC5PT9c+WwwxiG718jX+7GewdiVrRpJCL1OxnQLRDX6c
pRH7RchTh/8mMiVJRgFtGFXAg4Kl8rpOcN5iEBfyRoaSiPV3auvPh35rnsDnlA7AdZd1tsLqGvSZ
tRpU2I25RI5JB0y4qKY+av1G6aKz219TOPqzunE5MZ39GyXdN+/HuPjcgyIb91PVN2qLWPzGTP4X
pS89fcNVNo5XPr56gaP8pFxr3ejMUwBXRlh4ptldcQrZ/z1tegAAm7EXFQ+nAo/6JQmxR7sxO65l
PjyTaH2rH6CeyuEj9H5gRHseLGNud1ORx+hG4LUTfziR5KrVuaDZNiDYQaPGbQIoZaWQUS3r1OR1
G1FGKlTt9sqrKl1vJz0d6j7FAsjg9x1vw4skSb32Ii91bwS3olio+frlsuffo/fEng6vjgZ5xX5V
pRMb3qRc7trZ7tSkW0X1jm4bC+g8hrxiERQ5ET2bJx+QKUg1R3QNZpLxtyC1/TEYowl8kQxq3GRh
2zgvJnhmIPIvawYBnhhpBHRSGLcAq2cUpBV68IVHAZLdFWHrOfZsLH5Z0hcbI7TPp5vrkYlAzZy7
tfmz3TgCuRMviL5wRnrBU/Wz2RXEu5qePU6ha9RYQ0yrSUEqEKjNAMuAbL8BjIp42PcfA7A/Zjp/
kUuLowmwZHKgWNErLM2dLs7rFLzSNKuuZjYsS3Aa+38iq5uFkNHCL9jaeSwCYMR35GE3pyN4+b+M
F+SAJzb9Iodj/5bWcmKf1KBylcnhzOetf21MytOIkumaGbhkRvs/YWg8yNy+OXroirFuf41b+75+
PEcWz/Pt+jukSLIXPpeNRB9lbpHKMkjpz5GTo8a+94707xEoWUWBk4GQXKXvpBmDTb+MNCnBmq23
Yo7fyZxfm6RvoUcY6mfIunMYH9tsMc+sQiFA+GZZHwSlWYdsD9j9wuijwllAKIyAj28ynVAbx6cI
esii9Kc0XaUhdloeaK0ueCqfgBXZnzsiCQeIRuPqiLtt2jR9YV7iBBUHOP3Wc0phJovn5saS6O/h
iXU4NhF2ON2lFZdzlg4vAOjBZeJ8BhXTa7rOG+HsXfgaBgJ4qsSZvqdJYwnSpiwbv3wfHe/S8k5V
gDvS5V006wXGwJx7FjHza2i6D6Yy5X+4MaQdp7PE8RxTPaX01H5mJ2lloIZNiEfFnexMSDUeIwcO
CZlWInUptdZHJIzfcHYM7HA/uHQfTWNxsp9qOwz3zwF5vTRDjqj+ZfNU9+3PiU/08KLQfozec0td
9S2WRLra16Umv1A89NAusdb7qodFlE8vFjqHQadkJ79m0BQziFlGqzukddgnVFAilR1wwoZ1Jkay
FbZYlAZH3+183SRxmxsh1paUftPCCgp180fwv3lxtx0pkcxqV1bG5e7ESP+VRlRqmzU3ofLx9RpN
zFLj3mpSJGYeXIi5apnvN7oEL3FGQ9vUmQVra4+ce9/Ef0wfq6gpRwXLrPuW7VaRJqBzar2gcUKI
JMVtmNkgGRHcbLwSNQGZTjvEdl7zSuvVJUsc4wJHqUw/ZIjBmLj+rHPe2PAOdS5EAk8FqW7dePU0
zFi8IdOCCTCCErw2wcogkkzjuo9vMeXHwx3KPhFo9GcGjjAfsN3iIybMbVhOHacCEuYoJZYKXGz0
Cx/n4AVBLccUTdYXyDJUxXMRpYmX39avlGglinjFT3dDiEqg00Hp+CzMMcFL2VxsoIKKIGv561nQ
vz1Ca7OY1qiINewV0kXU48H+s3ysMf2wL4ycKAd4DYTAmsh81pekp5ntYngUJ8IKgX9z431BszWv
rSp1dZZ9Rh0sAdsq1OUl12X4LAYAfjo5438zBYo+eozk90WRZHKE8fP4fp/NvvBZAkaQdrLkVQkK
xP7ktcE15nV4l32qfRdvrKmmDwWuMAKPHrW5mnp2PNg24AiyR+cuFv+Vwj/Qpy55Idn9N2i4nzkD
ulRqdefA46vF8RspZt9pWpk7VNJMADZx0eErdEYMqKTGgxEearGKEgxbnxMn/gzurqZv5iQiadX6
2QedxCBUusUsW0KUoBO9HE6bLRDt/GwsPd+rUwUxy5Q61ES/y5l15oeSPYuN2CF9s93VieqxqE2k
YD99CG4zHMWsW1T5i/06nAeXVoS7vC/CgT/YoX2L4rmO7lBmBFbYMRcTqXzIOj8WtS7z8tlpQIK8
Gf1WJlaA+tFiyTAjhXXfDrbg8h6Ydg8OQuo8N9E/YtaeW7/b+6Yg9Tax33XhAfqZBM5yRKcZ6S99
wCmJJuRDwSInOHPEWnIu8Kj1UpecU/xsYHO6lnTR9E9yjXfkGCr8i0e+sp0q5oiJoX7A3UAGoMCq
czu4CxBzOabVX8FF+jtbopNzOvoMzrlYgVMqt4ZJ6tx+/de2cG/z2r28YlbCFGxEEKx1s6rHr/9t
evwv2xkIq4rpu9Pmk71XYdVg2DQi9IY8F4lBHafIsM2wrWvydhU+yFunRkR+JF7APPf0NGcidQnQ
hhypvOkP/DEeza7gq3nURdErXXwvdkilCIZ+/4WGIT6EQDTiFIVGDldw48LLfsGlEE6o1P7aRY4O
S/N9M/h021dtW6a3v5Pd30q1RvVkqdh2g9q4wGtvO8likPl16RSwOGIHPOx7HoyKB7GTd6iTobpv
GF3jOc76Ezd1aN8pSEWlcaRUtnjYTHbORK4oAEewEwGn1tXKBAU76VWatF/LtKSKBhtrBaxqEGut
McGm8OgrxWjKiad4+5WSmtWwYQoEl6bzfLaNhXAo5D8/xPMx6PPCFUHudIcS1tojXXHrqzfmuHgg
GV0+TgVmsCpn/uNz784p6OYBeZKbbzY1YqC+xkr1u36nFhHvu9Z4p1bWE+tuRLJiY86GY4hZg8ex
zk1irNfxZ3HtO1OP6xf5E3Wokb0He5GlCK87l97Emv9+wVEJgJLtC1owtbsc3HWmV67kTL2OgXzY
P8saa0I9Qe/aiX+mF/UAoVkyJHvFX30J2MaGWdCUwvHC150wUJlh11vhz3VnYgcrVD5V/8VcjN3l
Gbnhq+HNaPG5UZpPi2KxdGFpnwsiR3/9x9OAEawlU91cuAX7N9YATQ037z6t1wN5JOW8Fv9BJShp
mrIQyJPBI01ik076wpFKgI2gDgT6MomGgnX9St4uiH3Nkasl+JFuJ35Ikos6ovYdfX0tUhiwDWuu
pLSQk2mQjqC4mn/YaNnlgxgxLulHWQOwCvA4Zz0UhCKRkUEIey+dqrCiJLGK9t+ONQf8fGzZS/Q6
B0mcz1UcgdP0zDICk6CSLEPz/ElKbLypRhn8q+UFp1M9YszvUfJDa28NeFyK+fhtEKrZEiz5071R
KkaIQ8q7VDZG0xvsut3lGVTBznAd6TYrYkBrxJXrXTURzc0u/w83PWmFr3yOXNYRItkTy2/GGI2E
ik0+DkHtrYdG8AyK+sxHJUx81HUBsFNeF4dpvX32Ub01H1Zy7fqKol2r0PwnUQggvxD95+Ra8WCU
/OzBCpQBkHEsYKYpBq4LFHO7ZK8Ljt8czFj4989rpXPghJpwpOH+jYje0CAwD5ycuf6CIxiU0rKj
HdidARImPeLl0QVIOnr3MAVFYLqeJATwzHiDosoBwF15xgD57sUMSlpXBUHxKRJHVL8yHfiCBGtB
vFFa4tih4l5+Fy1xTg85jgfp5iADa0LuUIxMJoXh5H57DwvWe+mUia/Tn7iW7+cxaqj4pJPUKNEx
F7cVcFWlabU7xIXxWVEnH//KP02zqwver6Zo47gjhGv4kcZdr+qy5tskOfShR2Nl8F6vH+j8lQwl
AN2f9ok64wBce/Gm8bPvlOoRajgeYsn03kLgI5SNAeb6Cc3GTdu0J+zivGFPpuMw2lkX9H0AXVTN
JW2ARYdf9isngpQhF78D2tgXHis5N+WRR6H9P73AZwJYk8PzqH7kg7Lp38j4Fw4rZtX3/fvd4ZPo
JUb9vu909Dc/WG87TtnMO7mqPZfou6ZzarBbkC1bxSb9XLqjml7JOU6y15yXQf3ZflGSWIlUhwrj
XJle7Wu+dwSvyRWJQegRrjS9o2CL9F6HNbTsZCY33eU/nSFW0sNsNWXFJYzQUKsqzvC7y2+EyXK3
gysV1jNngobQx4cK6/3UW4eOlxvffkU9R+wVaVbTaLdbB5x6UraPe3CBxKBODVUzukjQfaDHw9St
A3TnOLflVCcGRw4BRyDJmLO7glw0CihriB6Pd87uJ+Wss/gVtlw73Wezy3vSw1rq7F+Zc783u7Sn
Zou3wViimMnbpCslIJYbaY2gbGcVRXZ7b1kBHL4AXBglH5GG+P0i0QXj5erUXFrNGaKRBRoi+jjx
g6oU4UXfjnxb3wvYrEHVTfT+FOZwmG5hsKggnzlvvulUNSyOqeh+FW7052KYermdYFMqs5wea4HG
jtzKlViNq0xtDBWJn0xzlCyzIaxQQL/BEqKU4cIvm8dSH4DpsjUxSQoFqiLm7AlAIczgmTVck5ii
iI0COv8lH8tCcOKFp9SbZSqRq1DiW2xFVV3Mv4+xrGG/gWEKbqKlW9UtgHQIgG0hQUsoeQbBUrbx
Mi8RO6vQTh+bWgtQspKqjAc7XYcWGAIeEFKuwrZXqK/l4gF2hBcky5mGkIKfXwJZz29Q3HfUVUfb
h+bVO7EndggCZXjcyNpOPHmDEZmeppDy3ps5Dl8DHoQICCkmzTJEuiudW2m5gvvEVVvYw9ILjU7V
IoiTj3HfQ9caVvwRgys8phN0yEuZSWhh9YzaAsWqiqIp6tYJgNF2oVyJ6epb1xKcw++5SZmvLOLL
Z2HEvIcBz/Qdeep8RR5BJP5kMTZVeC1vR4ixHhq5gAxJ2l8cXxVvpO6QpDpK9+pzLJlslaf+5iz8
Z04+UPlAk98NlA5X5wBVGe2opXrZ/auFL/7OrOmBh4O9wGQgSTmfmmPNYorY3mwgT7Br2A5ddQkd
fjNh8F8DjJUzfqdp23OEuMIFFFBWFImODN67RVX4D85Z/iJaRby3ia+nqAFDhEb8Xq54dl/aAQnP
QuFff2bcq+AqdGRmXFe5YU/sMnjIrnwy311oExOJESG+V3NmP8H34Zz/sxd17oQVy2iQnnhzbE04
mO/yruMyju366gaLjbkX1bxIxeCSjPGek6vA3ISY2bi37nNheIxIzGQzrWZWrQWM/0ZxpQ3zrsby
3fgsHeQtuSNt3zjYBy5CZA3ulox+am1hCYAYFjZcFFLit3mEy+dqIkDxwDbgCJOjur56b0PnWN9N
p9x/TXlbSKXBp500xZqdLMkIUkfWNxlKg29iECOrl15Ixik6UxZFJB7TYxbIhKSSZNtQmn1AM4S1
/dBhH22RMOf+Fo42Uybe5LJp/HU9vXZkhirZBXeYxxNcPFaSwzvAYkXgyF9ySxgNRBNdKT4M5sqH
lbPsU4pLrT/NBXjCfp7AUjwSQasJP4Zn3WlWYSfQZEIpLEpxV/ys8vB91GGwdwT8Recn3o4wcwbE
2irgfvMe8uwQCj3A7SQg05w636DG8eIepdKFPZaWga7A8Yumq3sov/ehg52q5SCOjWOe1H4vkZKu
F92u24tJRHmLRdx5pBNWTRFpJpvQu47wCZG3p1r/BsDcigKLUd1tTjSeI9n4aVMNg+YMns5/XY9x
ksvjBYSC+bKrFDHdvxX0HV6Hy4VASVCgN8jP1Y2LP/jTD3dJTMJ0bCDJtMmD/5OTl/NGcbiYvXIc
60aG5Eha9KnJS1IVCzsPNRyc7j+OjzKvD6mAbQ8w/w7r2EGQPZExbUwdmFfEBsz81SPnI+5bPhn8
w3tByImzt2pFlUOdcg2IblXYKtT5++GWFVsStdiwZJ6WyJtBq2vyyeTY+Va8gQq+EuqONeB45ex5
cHMU+2t56saLJAAfjC5aZpXsVW2IEQNsAljU6FO+7wJLzZK1PXfT3vL94OdfdOFnI1zmqNdo0LSe
N5Ia4s+N5++5ttCq3/wuzwmFMZSYvZL+54A/wKBgjIaZD0gMDGA6XlwSzlKlpfAqGFRDyW+hbIcU
Sk6dcfrHjV5djYOxuzhTupIYKTDOFATzAd968hZLngEdHAVXjKwy09OjuZwO9EIH23kxzGTAAe6r
xUSEXhQRCWJ5OTh/9RDtwDlKWWQXRwX2oEVlOcfZsOrBtYfSCvrWyOH/+KPIuyjNAacooGdxZUP3
7Er7QfaniiK4RgcoS1jiL3VzVQ7CYbuTwQsYD6gr2YE3Ky3kel6HMVGMaQF12mbzaygo4iIhWCTX
xuq/5bQVdaj+14o01l/YqsL6gTNxli/35tUzewH61NHlT7M7wD+HHEc0XDKm1d50lF6a3F9peyI/
fJrnBgHg618WQ6o91PdZ75NoOFWQaELykuIgyRSpjUvweue2ZBApywzQ6Y1k8Bd1S+U5A9cybf/g
hzycIkYjj5dIutjby1Y3h97O/R+0RU2KkCC3P7MhFOykuo9xYuJemAadHbE+YIjZRjMPbjRudMRU
0JiXm8g5OW0Qxum5cYCES+d9SfZYyLoasNuk6ghPrpL8bjBgZJhWxmcK6zM4fEkzfKfXCoCGHHtm
q/XRwFwVy/Ck59hJYoJ4uPKz4oQrECcYn3BV/AEqiZaIrqObXXmzKC/bBmtzwCjmkhGmID8A+sEk
KiSjAJcpDREG6exDsIF2ck/TdWxhOG0NMHlFQrQ6FdGivt2hD5S49T7QsrjK00AvhIDmxqf+5kmg
bdxSHATPiZG/sL2Zhd9hUEDF4HfYSmlAeO6y0FoYjchiql/E83Z00OiFMwgce2Vl7NU5WQj+ikR4
WD1xUF2ffP4nMmvrsOSMTbbzSY82bXCOOPPXnrrCra8GBK7+wM54WaSvZzqYJXSQXs3SYyz/lwFe
KAEKCjuWzqXP9s1zq+KkJNNYoSC9oyYnU/LjtWUJIQPA6NwIwlM9z94UNxyOlZS8HouWjyyD77US
9vpkvYw/EIXY4SpI6fGP3tgbeHSQN0C6q1rggA72xpkw/r6JkO0YhN6RfcpJImbRBCCiQVdZF6jC
mllueOnv4royESrDv1iRYtedaJsPaukIX9LIodJUoO7z/uyTnxOEsubFghD0wvzduWhjuB7wiB76
xbi11gOoTFuiTPSvk6UXQbDLozMNLZY9Y1D3F45qbCeXd4KWR4pt8cJ7+yFL7R/A3fhgsAAsVlsp
fFwd9MJNNZKBgWVGes6PEKjGQOC/5BdNWkvE2TIbSAnoul0fRtnGhYanAxq96/xo7OwfYji8jO2d
tXJZZ3NrxpsbGTyceOSE1jqoLG6Bw6xADAUFMVXhRjoA0O4HdoRJe9Ric9O29w5eUDyX6v/SWyyK
oNMVShWLW7ZrmPBuusH1f4Ob7YyAPD/I6eC2xLoXJT2/UZ9SJc7DP+b7IIhU2CyieFijm2aPs2iO
NtJR3fDdrEvhJtDfc1PgY+nIxBphrR8rZ86Z0DPhzVH5XBvAKeOPt3aKqi9xk0Ls/Ep5nQt6i7Ra
9+J1hBWj4eHHcme9IhN/nHp/OT06NMVWSrLtxrugnQI4B7pkPob8/qAsaJFgz547Ng0yCWb+1KgZ
v5wPqL1iQgh9QJQQKpzmJ1hJjpM96gZhOsH6ar+YLoCSTsOLa/wru2IGT/ed3d02FbcAfLyIHXkU
Q8zrxsCyLsHITE6NqcTbYgBW6QHU541TiRrgovQc+MmZDB6OinFMy4Ny68VM0vHhZVeMq6eTuRpb
ip6Bq2oeeLFx5AQd75Z2lZ/RfAVdKtz1sMEPjXS0aXVSOYIisS5GKlpFncduZpa+Eqo5hQp+GqrK
Wb7bLq8n1cNikhc3cno4+cJJnPUnZ8m1PUv9xpQn34uHZXpD+om09trdcQQ4QFO0OVo7iqM2D0D6
fZH7aIXzMduUzLWHAUn0oQ0ccm0HZBh09klVyEKJ3ZgcNJ4N4WmxGdgN6t3TeSG5rB6hawKj3MbE
BYnqES36jpXQelYBvxeA/y4LzMTqYi2Aw7kW8W/vX9yUlmFXnNrq6eziDwkq5lPNePe6dWLfwWZ8
2lqZJVWTdVnL9oAYKG7wVeRLkETB8yJS/NiPWPFIxBozYMWHGFuMp7eUeqPGNc3Qq9bMoboodHvM
Tz69VagPLb6kxJnrLWVTAnPdKttjjl4lhYp7i/mghhWYkZwo1W8Rz6Xmml8oZAo+AodFtRA3s8NA
2XUpcUiyffkjppiH9u2E/iwTQBKRcdAAjSO2lgphmqS6Bmn6ub2mweQ2eSQE1hXE3Nn0tYdmoqpf
esa3nQkdAnTQk53CKmrpDqKDA6choc3iO0ZidpBL+r7tomtTa3cojkNhFltqSkvXHat8q/dCOFl1
jgCHwxrdHIhk1TG5ctowB4b0i+f+v1EoXIOcDYEoT28gYk7zkoH0MHDgq9cJF1NMR7JcqAEGKXf7
goNU0+48fCQQGaIruFTwPK8p+vCAiDaVAj+lgHx28gMh0m7OQ8Kd1yehwPpRjgwbGdn6i9EWP/wf
e32g/GTChEAceblmOMuq53OBG1HaZe3+Cf2af/0gz05fJqt8acgtg3V2ickW4JBqAYGVM+nUIvIj
cX0a+OeTFxM5n0s85l9GNY+MiwMk6m+oBmDJ3lp+A6nMwZMtXKtEUo3QECL9JO4iePmfsjZwxDmH
givqgxR/Ln6bCi3Zn0arRzre5ACv5ZkP0Xl31udMusJvQAQU0UP0fhi1dBq6vjaA3e1M3DtEcUJL
tT4x2xcV+8Kwp8BbmyZ4DWoFSt9kYKQTezQ/h9tMS+IEw2XVAU6Ith7MWG+W/XW8s1YlrC7bPSlw
MftbjGNaBjzwCIZ+JksObUm8+mEXzU93HXR4QQt6IX5z9LhJ5AgE1YXJ/XvCtsYPDGze41hLNTIs
/dqn6HpZFa7+1TSusg089o7TPNUW+nZvYSX8RWylYBgXfkLsQ0jv9XdY8wJ8QRWg3PyOggFM0TrJ
5YlRYhN0dZV8S3aywVEk/ETQprUu97jFtNtN/dnvUbGcA2E5jiiCMGglHlBCcN9rAD4FVJWgWtxS
5rZe0pj4uNLHgeMmU+DG5gpqDulh653qr523X8b9XzOSGITywCQU7cMkdIv6Mrn92jtTxD2b+z73
Syl+NsYUxSojkrSJuVsrPFiOtEeT/9VNzjntxTRhiL3c0NeRn6sR9KdjVfcrSOjgNeCWl7lOVjN7
bmgtWJ5c42CZC+Z4OruVhJiSQjaV/bJtF0LvDt024ooV2rMww5MUwGZjuJDsp1cxhCJWpF9DetxG
9uPiN2nSzWRplolUYkP2P5H9O+Ub56NLPPQrwwWR3Y528x9trUBizZU6g2Ag1AaQVTNDRbSX5Rjx
kRW+s52kY35p/z5PnXwgWSGTRGiLOx18eaCCcEmJvwvNilKrQZNtK+uezPl+qlx4ptusKWVgYNgT
eTrmYPbj1LGAUTUuL0TEP9Atkv6mQbxMYeea4SLIHYl86FzeIi95X/m7GmHB6XKfkv41/jluu8rQ
4g45awrR4UO+NK7d6wvQrm8r46ekUZ6oj1nJiUgOWVeWQU6Z/NGeryBTFzaoEkSlkj/rXoxHpAtO
5jpOCgJFrGIaTxRmilED0sg1w8hNy+D7mdj4VP4uFuVKbrXp4y5UbCqol1252guBOxRReki7niWV
blDfMbEl9riUaUd2oVOW2Fj9gCi45HJtbmamCvWmW42pHd8Q5hJf4MFwEEtlmUH19hvFXrRLLHTe
ElRIRXPo2YA02fpFBa/AeACS+NdP/BmltYHXvXPwyRk6wKUJkINCbMJ9N1/xg5Yp0iURgHNJ0isl
dDvm/VNfZgpBj0dL4XBFgE2DhdcLgeZjAjcwfErQ3xpTeEXh4M3axayH2jTZbxQMBiJBa6zpEYJY
nrvifjFEkddrj0v86c3D2qaIcpVogs/3q7E1wzTzptYbUkxhGUPkF2exxtFSLX0uBEiDg8vqOpiY
h8cB6Z7kq3uN8eZBgt+3j6HlVj5XrEgnCaIlPYw9oth3ogNQYQLOTQB9DrYEGkk2gLihzCbKgUNz
+Gyq/gQfFPzm40b2p/667Px8jczCeLMSxKcr1tJE/ZrKlNehD+YTbLENIdmftdO5Tm51xFFn6iZK
/LIZxy9Kfi7xsG4TZw3ze2Jo2gfiu9ilQZXzZsz8M3P0gymhIHP0nG9OEH3oz4nF/3YT3GgqLxxL
BrPVyxxuxApo1cYV9f9hYwTBX5WvsVhtxgT21+NnsdG5z5lYLgY6pIro8tWd/NWZxOtxU0LMMtyB
eWQOhynteNmhTc5akRA6D8aGLuAne+spr0D4mOFhcofgEdKuv3Zuk6bqE/PX3dC18T36X9JRO5+u
IU5GRA5xzOkM7jdb1OaUBoUfSDs+xXC9UanH/gBSm4VrklT118/bt9+0Ui/Y1/ZjCv8tUQZamlQc
duPb3QIeUYxsbRMnDUQD4Qey0ozpQFBVhihMMYyQq9x7Z/XdcOg+rkucA5peGrmAdwoTN2dMpMI6
UU374ZLX5DwW9jCqFSA3ux3GGN/HEl2YeWyC8V8hqR7pgi8cE64hZq48McAWElAPYMBnP133VgOn
l8J8z5Dpi/NlNTK6PSObXMyOsq8Z7Va2j6uvQPzppNiHQSZYrp5pmJznMdYXZwz0QXutrErqw/E1
owV7im+EFhtuPSI6ZAiF+oaXkQEoh+zDM96327zIpUjrGSY0fvFf7W9RsoF3tef4PLx3vQfw9p1X
asrWIDRKmq7zl/epVA6bD00fT9PfBtfpJbozUjbQ2lDNiCpSL1ZndylzTbkOzYRfHQ43mnKKF0kt
YEHBLQ5Oa1ay55gb/PacPoVC0ChGpVGYKNCe+GzuELa6igKq/vOPDx6bs03eP4/K3CoWmicVSSh1
opboLneUPiYa8N2gutfDNwjP1szrpMU6C1Y3+Y8cIoH7WecdIa3yu59dQyHTzvwKYlqC1tO9F3Mh
VRqbvRtgwCuAvBmHjOcr2yBjedsS69uXUm3VLLGKMUknT4R2apamXxOuKNJ+jbFPHtgj9mD1Nghy
pCjUQOv3cM8rDNBnYLJZJNa1bLlvZ7NTfGOki8ZEbh5TILGNy1EePzNIdoK6djj6+an19Mu2FO4o
xXQi0C7KWs5Tg1j9G5J29hncNR0VgaTH7rHBNwNY3HtccdgsL35yYrL6PFGxeg8WMuQ8Gnx9fY8k
/pAy9oQB1x1AKaEJT56+Apz5a5RcOwDeSI+qmCwECa7zxkG+8KaEL3JQ6b+kGf3nmMcfywhbIkbi
xFH3MY6jSY+0DHkui7NKIzSt8UJ29Rj9L5O/RGU0Ozg1ANkkxHXgT86wJWImIqI8/SgV4FJrNiOY
eNeiOb89SK8dQ0OQnXuTDYY3M5t4sq9DrEQJCxx/xYHVgroVTVB9XlEalNPHu8Z4Pd2STSOqqaio
gnjPF/GmZcjHg5xSgHSBdar6cDRsfP9QfJkLQu3y9AU0qmAw0VVHTFbLHEt50Ea8tzAtwCbedLR1
8dbVVfukF/Mmh3u88uFKI10dMHNUOoAIX0OrNpRlfehXaby9Lx6ezUrheSMvxMLJCPB5MqIq5DIz
RmYajModqsDGuCSPvQDLlrU3XEBQJnPO6ooGrEhm0Ag6eXPAbjcW90hLznp1fGJ/zHOcLnbs8NFr
JRAdCZ9XLrW+1WA6E8cTXxjdu3uLq2vfVgupuAcG+Pw/Ws4i6p2DbAR3QPpAjRDX3Uj1CHd0bK8s
DXF3y/2MQ4timbLUBjUB2vzG8ed85XHDadv+g+Qvn/iVtxZLtzDbJB8Vm6dXYh/tZpQyfW6bh2SL
8SsaYJ9pvnz/i7B80Nj81UKZ7yyH2ehUtlireDzhhHoLYeENlJWF4yu7SJJLDuC9Uae73T2dRgc/
gbZ3xcE+8KmV27bkiqX6ccTpEKkZ4DtRI9f4OnOkmUfVLrVCZUy2f+wQJZjubFDsGzgs4dbZzwVh
AGxmjzWAfsDOGUtBvrG+whSMz7AzC8ANZJSjpTZhG4DWOHKwfAQyoP7Rx8bHtSTpaKft6sonAwyg
5k2dGoNEPgHMuKYD6C38nvNaEcL6zNpA4g691bViDs2t9mgTu27lzfd4oY+hEzIOmc3aRj0952HA
9eWqTGml4clJzzryDcSVAlOA5TJa0ENCl2gwkAJYp4O2bRjvrncplH91yc6Auua/AfbQWz7z7uak
nfbn9U3uM4OvJ9pCkMg3e9qhRA3tLXrmmEmIirGamT9C1BOodsh5IQSqqqOvXCLhOzYzxK97HgLS
dSDflYCrxX1YhxTfRJVf71SOBo1IKojy7B094A0SEtzNtLu00PiTRexN2MkBDmSKCrC9Ov1Jwx64
dnCO1qJF3lH+C3cQAn3DmQyBoBtQcigY2S3v8dYQA1iuiJVA/LmNOFvIyrv380AJJavplvIbtemn
smZN/K9zAihH24i1bHRoG1A6rnW+QM0fxEtFG1mGH+jrL6EcbCu1/1I0A1opt2yjA1iip+7Os9un
odUe+3fIYVhoYgd3m2loWe+7yKD6TeI3AYXm3PYoZBF8hhpDzZdeRdpe1gcm+o1NZlb84U6Pl1RT
557KjsH18cciVxiELvLWPekTWTuFXyb6sKdjZSew8uIAF3c+4BAWQ98slzt5sBYwGlHigPzmLg7N
GdTmo/N+O5RnfIWyVCXIZkBh+2IgiovKkgb7TZYwedc2Wf8cOAZlW/+Mlviy/p1H+mHYXgYQc4QA
kuK6CN+KofhmRc0+/hcLwuE0WSw8kx4agEgwKQVXL1Sj0hdofM84hb65tJqgHlVhkVTuBqRTxw6p
q6Fn5TEiF+yAsuDXdpMKYEqsqw59pr7g4ErWmxd26E5f2kZRZ1IvcQO7UBtKm63veaAJYulPgYRR
cbe9Kp675gWBTAkUytozOdODBBwhYwxl38g4g10OcLRvIyh8HyZXDrGXT6g6mFKBywb3fBcjsYRo
3pfGRzL3zAFN7I0Jm6QRPOrCLcImYIa6RUIuWoTchkQeqM+aDVgopN5NeNxltlpCDzkXkJMKn6Yt
adJmMDHANCyPXYzZACrIVv9heZhkZUKMm0zaQcP56+/EtQ/tALHqpLDnrEi329btJDR0Jca8yqci
BVOk2poRjSDLD6Aue+pubZ4GjVNoSY9yOwEFgRs7kY/yYDvn5jmWxAPK57WViQSg+WdRT2iztN9i
oYtA+OtdPwKqXf9egH3PgfefpQaSyC6yOWbPheK0vVoTyTbB/9NIk4rrCi3l/nVNfh9+irfhgKn7
Y7aM12sOTy1UKcdx5/6bVzSjr/BaqkxRo7XYHKQMw7KxLyyX2t5tNGu67uNtAvREQ4kSsP4wEJgz
6rUy9yaya3IgyrmeA80wQ1NPDkvEHhVemM7VA0+F+Kc1nZGoEe72wlO6+eHXG+UGUtCQef/fQeZD
DRYD4V9Ul/YZO/ieg/ieccsLAfpR2pYXeaHWiJyK6c4oGYAO/9uQZM9i8JvAHCIisYxcDOZYMpSy
jG1CT4J4h6RxAC7mM95Jl/Wf+daO3yWoovi2xI4E+gO6oOxAiUQBxUHtY54PGzeEO79yJF/g+Z+V
4QCtPKf6bQxAiv31LqgvGqw7PojTRZRPKsCefN3PzXA7wKWSF7WYqTtVcGrBDANYqItCoZLnWQcb
u7KuvPjBOZSCO7HuPIRxK/2Rbs9g3N1nssDkqdFsVzW9xFDnu4YhlykrzCprqGunBUuX32TDS9xy
/QD47R0PYTMKTtsn7/F83Qiz32NBPfpvWNlhSliyQ+5qSl2OWAIidaJ5oRLCu0bQEdJrFmYckgze
OqM4w7HQ+D4iEy0VTnMTBofZk5ukPdkzxHRxCV2CnipO1r6dT4kWdxiZKT7GXZI6PMLck//hCZw/
KwQmGdBqfGbT2ZG+jyvXjjzouLpyexSZIJPGpU055FWzm598fUN/EnAUYJZIEJMdiD3pEGQrcxxa
3vsV53Q8kBF/bJ0kcLTMcMWVkWqNfndXvN2dmhABDqhwbEJNUp/SeH1kt52VD2PGxyQT1OXbek37
IOJfhCpC9muS4yBouk4p3b8YY1go/Og7PkqEIXI3YHW3+PTXxUOHQlh/nWzfL3WhB6/vmY1ID19o
gZK3g7ByU3Xx5ZbN5S0RFJv5zcqk+/hKcvswTTuhxRdhIvflYUh74Ll2ytK/64ZsIzMs7KtmNRNF
hL1ff9HsUQiM0dqHHZ9ssgWRCd+TtRWNL+9TZGC/XQHl8L9haLjPo1QzVD+Cw8+nMpaovrfVDIp5
CThjptGwjVaKcdfO/VhzotKG1HbuHxHMSjA8wnBTQcxSP7Cipb7MJRVJTAXhnEh/GB43kUS2uNE9
qgdoytzQvkrBqjQI2rwGhw2L7zXleSWof5hBYXq4TudDrYpSLqj2eWSLtBv+2kh35UbfN7R+dplZ
VwVqN812cJYAUQ0NntZ93jXaGlbse3CcB1AKcBM+V8mzaL4Ir6E7LPfGFeiLHO6eZl7K0nXo81vV
VOYNco0OsrgllKqq0mXDy4pXqHOXORGyT84xEbSHX2zp6ppSuDCd7fpRFjrQzcBqho+VVVpoHUgU
9OU47lpZKwC35sn3QykrOcRvxvPwf3jVR+4mbkI/D2TBjTO0lpRQ5kpXKmeFuRFalvI0CsbbC6kv
xjjXs5gmO5sTcs6YvADM+Bf0sPmBnkiFprFN4Wh6A4tPmm0QvSI8cZC3/BRlpw98VcJTYZJI4CJV
cBFiPp7SJps8rH4CTOFbE2GG0sdYRZ9ywSMPZXT3oiCwVw9vlJUQlqyLTyfMXcGQnfsoFITnptzk
KwBQMN1tDikz7Sg/EeLWmtUOHelYzHv7pZROHYo6hD/GlJR58NL4Lkrf8b8ZudWjkoCPe5NcBbzz
8eqUZkE9WeyzT+PebPaZDHNZvhaqcxVpsYp6MiOQCCO+wCFy57vy7WhEd8tjeos4dz4uUMptUdE4
NjrElBrtXLvdXJM6L6/G3Rg7GzAr0dgGRske8EBwaYHLbLUFli7J7Km1fGIrAeKh+sjnZmS0Hlvb
qAgfpZuRmkDn1jHAT/0BKRYGqv8izk22jvWmOnx9NFKGjfwCIvGAQyivQR4PR7SLNjzCLbRQC9hL
EypBmH9qgmsp3x+bDbaNuTWl6ABeJQ8WmK8P10mwP84XMzAPiAvheR+cGs+jQe278JaffS0IywcV
VtzmsueHNDQl90Qp+EjPKWaGqOyxGLKgWbicTjRcC9rHuFWoCgO7YsKJZqX4WMBpURLfq04oFNBU
Fz6nKgGccVfOccK/6UFpk24unu7ExqNKAkRket6ze97wSRENMuAgTSiRh6ggv23V3ynkSy6x8T+t
RkciImkIem+fzgcUAnW5lI8YKUbXKEbl32Dn13bFlzxBWJzV01l4KBxjp5I+CeQcBWN3L/dwIRZU
AVpDr4wkSOuccrT8OONdHSXL9fS+AoHUhKV/ozYRuWqG+vhKMGN9z6ndNeEdSI7eR6CMvSx0OJf7
ERiLFM0AFZvZ9Rlp/pKivplDwtThPOsIYv0NK5Ce+/Z26/UumvwWGbzMe+0MNpgMrqgzpTyaK2Bz
G+qUYERkckudeY4m9YwO/BPq4rSCid77Wkko72p40h2oHhXMkERJStF+kE0A4cLfEU8xNX6an2u1
3dnCK7qEaY/lExCxWwpjn+W47nzd97ppe9VrRyKMVW7Ifj0knBR9T4f1I6CjeZGAYXQb3jrENZjq
nZ15DUtflnihZcegQh8972wjv1g8NJudj6o3vfAQil6V7vsoQqgLTFnLsJ/lKt3t0v9ZAq09ckGP
yndHYWMyTd6fUnl/QPqsweVy5kbkLNMVk0nCd3gHtnUTtp/plDT2787bcNQcgJWJ1A8+DM0fnhob
7c/X9yuDjteYk2KLdnIMkoHIMFZoSyOPStIVq4WSFngPf9Fn0zMyfg1Do57D70zai4eaasSlFrGV
hXBoUr/RB/7qzGgATuxaHSC6pjXH66Vvo0xT9+OBgi/tKXOqHdOvIvdq0hgLPtc4O9+SN9jXCUg8
DcQpqpRAde+SU4PNxHWEU2DOow4wN0AjFT7ihH5E7wOzaIQ/4/g50ArBMecrKASliLIPIpgMO6Ea
cOpHRN2ZHunh5SjEUfjypL3Pn/f3cHZKKk0CFLhlxBUugn2omfymN+bYMKk71QzAWRCTJzp42BWy
rBbgeQiUNcVUmCiTxyCdIW+TbixmiGEbUs0qkhDzfV8BreIwGXCJKGwbzcUUPBPaKZzyWX72eJeE
2DUFJo0eR3o2w7TIpJI8+llbSiDSrvGJWbYBpx/udokRiudMkIt/cF6EfhN9Nybsq1r340IpxBPE
5IDWO5kJB4jWexbYRDSw1ISggtmuDJRH5iarXbwZZX66e1RSRLJwu6nGLwbCwQgA2Wm8W5a6xCh9
ok2jFPNXdUdDvx9ZAyjBmJL8DclBk+Nwl1iIzSf1CZNawLd5msaEtCEb4qIjNjIHQtmNEznIM78W
hRRvnwK9V7mKyiPIss4T7i6uRPBY1Z6jHTEnTqwGcQQR6yl4JRdkh9pRK97vpiY/NeqjFFcgmKbh
KiqcEtXPje3jcocPXMvVECZ5mtTEpL5sJx9Lx+j7aKq2PjlNSkDQOLaB8+y72FPdGmSGJ1WAQP/R
6ea6t8CJ7jpIJAFtT/gvhX1E9PhlodhjioxUTacM+VO55YSJb1GKQa0I3Q4C2FWYw31JJ9vzSmes
R9fFtZMiXDJfHZd3KBYZPuU7Zc8BNP/0U4OR7A1lpgkARXp3b4c7FupgKQRd3qvuqlsmnyEdhmC4
L/eXlfsiHzT4yjBXj8McV1vneVfQhKe1mhMPUcg+OJrfIw/v5zKZMXOAGP8MCNuUJ88Cf0LPt5p5
kKiVgw5DVXar2+WZ3I5zm/SJPJDjPAkWi1fJpNelLEDXiSdI6fWqPy45oEjPkI4wEqAZANx05ydn
rcubvLapPa8S0zddwot6kR2J3imjoyifUsyZp988UqmCmaBlWRRX0bcs7Z/wiZFf8Cz1/JmKYcXa
jF3xBKP71PnGIzaHQV5pzAqCW2jpe9FX3l/XXI5ipTHNB4gHsPLNeYHsiZblLUcAScdB0Y04IRQn
fp717CJ411Ij8iLJZkDjgJIki8158Fu0FlIc1+V8lqOLuzcyhV/KYWi09eJS2T2O114DcwuAqWS8
5EMuHMBg8ihyQ5tC6i12i2E3qqXCagVZgXvCE8r9lDDRS1yMXAO3SHiSfWAeyG6pkc6vrfmUv7Zf
TryQ6LYGf+O+zmv05ZUH219aS6+C5gF29mmyP+SxYnsEhwutAxEy5REtbkqFqe68Qo7D3fdMx2n8
s6YB162OIH/LnvIy3c/8En7R5ASyxKQOC4y95NLda3WB4LKb7vbw/prNiCz4Ed4XziGsZyZ9Ycq9
N5gwq8BxVF+A9ToqrIA6yQbRI+KGrFY1XyI1hr5oK3GpEbAweZtEVoMdIRGv//VQl99w78XcKzE7
Wb6plbZuFcsp7dCTccQHFJ6TrBJNFXF2rc4UpVNCHwcVNIleUZy/ZrNEwFNWsRDJ39k6D0dMtEUm
FAETLEhZ3fyMx8YQ6UWFsWiLd3tyzQ0jZlklO5n3+yPPRwiYWUYY/ErriRBdMwGETGZQyuQp5GLg
kKMR1NH7jGyMz82zXevAjEDntpS16gEaRr9j8GbLC2Mkzm6yzDEsP08RTznQll/aibXWHXm8X7iC
zCCgq6NYxMA9PhL+uM5d7qrv3IcTyXOMGPEjO7liQI4vowco4+QkAk6C5Md2Nk16U1r3CI/FQGMP
ectbprGS9ucbwgcVRrHn46+MZKomcghnBm+78aEbXcqnkVPszl8xUNvxw2Nbuz55ZQL721n/9GrQ
sm92xfzh4JKLaBas97dQsL7bRTyUuf77eg8PP3OHitZ8VdElP6+4W4LOKckj+lTBrR8lZOOtPn/O
aCKZ2TmOSw8r91MLUmHxMaZwgZ1v62RQ2wcKeYj877qLMzzlwO7wETsZB1/tMKjEqCai8qAuwTxJ
8JoKx3wuEQXtyvt4A76i+5x9dCHOT29n5pDxueOWeE3ZOBrGHntnK5pVZg/5VXjALESHNZViiOeo
z1yXGUXDkFIPqqgdLM/jpiYWuBME7j/siVN6CWHdmK7Ea8cPteaZsXf6VnWpXhqun+L8CtXSw88v
7yxp+tl8Ab2Gw9sDj4PyQ6ZFDykxf6HlF/SpW0IwNR/3AhK9RjinuO81ySdF6FVInnq63f7nh2z/
QCp/2xztyI6pVDBRLlBfWIZc3x9NRshndSFheDzeTh5pG8vK36tF2r51/bH7lPp2ONcJLzL/8Dxk
1zlonvt3hFe4N0i3pEFXImOR81fPGaBm8TfNxW4Ll9AAVfgD2R+7xDGibXvum26Df96CXdrp9lq9
t7tdLI1ilvbVMWfLedbp5MeAeZNd4wvId0n7zSEhW8LdP+fCjH1AkbNghKKU3tidgQupjhsneZSB
Rwwcp/OV6wpdYP3oF26wlIFaRLHP0EVBRG+vS87bQ5ZIn81e6LM11BoJmLgMsLGDSEC1ktES5K9m
9+cKHPl51PSw87Yr62ZxdmmnePz/JNcabWRK+n34Wr4MUYyOJ0/1aSFKA67DMgMrOx6cZNA529Zw
YJ1g9iNRGQVux7AZ9y5hRCpPxwlOnbXk5W6jbmi8zjTBRlsVvI8RX5u5r3mAerfpwvboQnoU9JqT
ZEM9yEj7pcvfmMy/jiW4zaIjFXAU2im7GHq4j/0WrcrF7FxqolfV5tXHUlO0/bs0sA7vgN6sK9RH
pWAj/FArwxFhkJvUTx0OZ6P79goB+7ynevzMQ/x0T92gXc0RGW+enjp8qCmVeHCyrI23tjU5Mv0u
b/bfChUyglJzEA+X37CTdr7RoxSURtkIPRI+QAEO+Nf4tENRFs2JreTMrRfd+WwyOcxLIVt5WJle
iRAbQJrtVfcQzow340KNapcIzBSFbpXVZk4Bf43f41q3BETAB0KNPD/Mwy9cGi11JUwLypiiLt4D
Aw+wkHAi/7p7gmE914xy+wJz9jFekLAAHN6KnoYA0sRNAfe3wXB/bQ3AYBggpG59SqlSxTmMZjx7
ot1jjoszhPo7Qlr7OkXpfh92iJpSWhl4o6K923QFP3yw/LoTOPau5lDtI4cnNL91CD+xIeBD11Q/
Oog5KG1wSsQ7UmvcfYe1T/Gnh2TOG0s4yuu8iS17FY4TatXUCmWrzEXMQY0nVG9T1TCLiMozP1Jf
4GgbqQDE98SItVRzccQsYNHir0n+KAyOp8H/tb2ExBy3MdxxsY0INt/xXY2VkScQoGK3q9vBaBfl
CWytrH5HJckw+WetTZl6aH0AfAWy823wWQxvi56dYBHVq4GsiVJmQKaKzpveYAbByS0pL1BEwpwb
KqYXrC/NE74ksM+eaiCUDDf0s6ffgchGtj5gsAz8vH1VXMUIdObdyT+EZ1OiV/lhTjyeDu7707bL
Eq57nHfIEHdOkSmnxSavUah3F8CzVjsDNIFKDPuZ9W6zWBd0IYXPBUZORkuTtLiThAtnRxJU9KYy
5XCEL2iqeSzqFYmSfsOjLLicAxPLixcoUmDhhpHM8jcOU1G3HJwhB3IOmSpOhUU5raggQDD9YK5g
vq4QKA+G4W1IbdspiqoeOX6+/9hH8gb2lQC/TOB4ZtA32d8Q499AGqAOQadZNAI8JurzkTESaKdZ
GgYshbQDm9g9HqvySbsI0IuW/8+F/67qWHL6cot/D3rVhUuPPvcWtD5UW7KlNoemN4oHerSl4OTD
3IKCgKCUe4mKuqBv3xCJw+EjVR3A3bfdxVgT03V8x6/vHohiCo65Y8whgXNHJqfKWBfeBXt7MVhf
I+zXVsEhnIE3Lar1Zks2h+hfbHfMwbF2XQBhm1yJeAqmRjiWuAByJai+5W8FYiiOEfQ8Wl6NI+OS
12Wp9Hj7aQDihA+R5x0Ngpm9wjWyA1xstSU3QrnNdM1/Jv8RS02CMXiC+WmZcLDqU4l7UxDebCjh
BGQK68opwOu+hX83DAt/0zGUM2UJRHgf79Z91wwpOPdvl3/bDg2l0HxBQrwSJOLG4DP2xi7NkwBh
GAacrluj/Tria/qxzbHG4T7SsIX1eU3qTn8KC+izn51IA69onw9KqVAx7+c1V7petFI7sP8SEK4Z
lQQfPd5PpiESxVcHyKp4UvnBVD+liXAXnMOIn/MqH5whymhL0MCtsh9RB7k3UxG0JEqyv+HVQYuv
YMYL5FM+k1JLUbhJ5j5QPxH1W1Rd7IiAqfCATYQHMxGe5RiFHw1ClK0eL092cfwmJI/eAHw+rep5
5qE92Q23mNQtMSxg6D4LKCU0wi9nV+5khM9xAS73p5etPlnaPnRY2BI467kuF+q8xs3FrbeSPeoB
LjdlhnBL5+5bzCOsTuyg1eL6U+YANbKfBbCD8Ii0zmd7fQO7vOlzZUUti9lTvoga8UGARVojH/qv
s8Tl6WHwuoLkWYretcawp7YhhlRaXPwxbYPCTU8o1qS/v5fs1Ud64Tf3BkldP5klMa3at0BNTncz
gkV0Q8dwsaZHAPDrZkN6kfprPQWdiAXVv9j5zgGIvValpm/TRNHcekjLOdG1NhLTzpqN2dFttvVB
yvO6UmFeINLh+xZzfsvF5ItHpgCfecJjTTsVLKQ6Go1ZlCdsBWX20hsxae7glgsG9B2I5zQfLBvg
oj6wt53l8eL4FDZO4tASb6iyTP1m2c1nhrR8AeEOvx0rELqNGLBx9W1AmGHN9wsDRjxH9fvBv4/z
gELroCUhrM7ejAHBvGE7pc8f/4wrz9sGx5QXMb0tvO+bcyIHgsZGZSqMvoorPiJjpmWP5zfBj1jZ
Z+1cGrlV/2yD26/F6a1/LkzDEtgD6pOaNcaNgI24DngOIShk0B95RD8mtOo1ZvjLnofSYXQBkyCo
JF1TZokWP8PnIRe7nMMR8RDH51XC7MccVXHZyfCpeKIJbHVmPbFK0rPJlFSolQAorzpzyHOW3D4t
YOsEBykDfLdHUjRFZLJKaUJ//id+OfnDgs7famNvRwkAwutwjYgvCaWUGqaAsiiU1LyvmAAdUYF7
gC1jezIQgTapp3XOAe9x2zxKdSI7JO4Mcv2GtcfL0M8+8yClwXG1WCKuCT7l+sTAsX0HgAa6ZlLj
8Cm/ZKNJZilA1+bC/ot03d+xqutKoM/sO5AcLc17qNKDeUjKSL0NKkQwm9iSO7YUyddst/T1/BRo
H5Hw4dkgoyFXnF4FtmT2Rx4aD+VtCVSlx/xIqCS+kYrk6C0kO6Lox50OKcIvWGvtXQq7thmQ/YrU
00MaBwfwQg3BeGBFieQYmDWEcQAsdgO0WcenwRW6F8kn9Sjebeu+iW4EKUEMy86v/R5AE4kXOTYT
XtkQuYjyDprjptKm5Rn8PdC5cBDrM0qXRQsI5MouKAJXs0qwjqjMmEyLkn7CtZ6e7JOCyvN2P+wA
gBLcHo37zmr3wM8mt31eZ9IFMbFv9L9whezmF1wcn+U5T8wvD9Hh2XXMsWffQCsxikzc9he2y9aV
UndC8sHK7fkc5HXPuM2H5QSUN+r+XLw8ujzkOvwQRvXwJhK03qoJxPSQe4S33nOHg06m5SYJvyVN
Z1IeAjjfaxTWPmY2VSNB6FT0FHYFZ3g1kF7O+2tLHrsVKaPE/br4HiAgGt4tYz+avO3xs1rgY9BW
b0o67Z+xM97Zy3b6hn3fStkeuk4QNjRH47sXRXdexLTqfkfrJRMgb3dKZFuVee3lTYZcaa7U6O8C
XdEsyrtknQ5gSFfrzqJiOy796JQdguUcrhNwphRjtDyPhVzpmQUcQ+vocAmZ57gHKw8SagEl//PE
3wrV6QpqfEUgHRd9JsVFQJUdNNxee830IK3mubri9H7UscTlZzLVXYWVzc88u6ca8TmgnPjAZb4H
y9gDZiNwaFqtgeuZEWGm+0jXXmqTkLQVT4DweEfoBk/LS1DjxpM5TR8fvt2CxzzWtWXUgJN9+XvJ
gyNURBtGcRTVt5nFQ8g2BiELfv1ISoGMzxeTWMxVH7zV3iLtqtOkolxbK94zac0kHWMrpYsCqKkQ
kXBs2miMRoj8JYvZ/23dMBxsZxOUSp7zSQshOuUcaQLshHahEL0YP7FE3mw2JcEmpe/XLdQLf8A3
c4IKHF0xncwojuH7I+g82vlhbLWp9fqXqyeoTScyWxdOWk+ElH+lT2t/Sh3dAHoWCo1eOeB8IYhB
5Yn/J2OvJQGrbk5l0zCQb+ht05rW/0RHaUEHHp8jprm4u+57XDJvzm2f03gD0UE17TpGT5Cjus6E
n4oAZZ9ztaa7seWdLAgeN4lHcQvCroiJEUeTWx5qL7ZwGDXWGymN3P6HXcPaLV2EgbtnBU7kBwVt
5jiAaVWN8Yxr76BJud2NoOxldCGSzeFq9ol0NyzhzHzK4Eny6aseXFkPB8kYjZ480qG9/rS32c67
kn9B5uAHBF5B+ivNWWhKGAMi+BI+S7TNaMQ3+UnDoxb5wmN8eKEDAFppCA4qMc/tbqHfYr0aFUzG
KrWlwyZuok8PwmstgEMFYQFmV7KVWQcmSRw1pWsol0zKt6Sf0Z5IkPHTr3XIp3n+Ji/sIMRAdx8L
N5ySQdJsAr+DOsKRRcWuBZD12iytI9FXdyvObsgMC8t+NSTpQ78fR1gm4zcnml+5ejJNQW9Kh8vP
IYR0NGdCC5qGuRfDPM4BakvFELMgUFmvilvW/Yr8X8Y0G4JB2OgvjIwpnuZDLCF3W/bZLO/r7a4x
8m7Zr2mcx+K+Ir9XygNUy7wIV9+omH82+qFt5ySvWvy8duaX5peFhaLhDhMJjKXkrF3otp3xv/+6
wbFv0YNr0FBlQuRIMatPGMix1+Uj7lEaRkhr0ex4EdyRrExmOj1ftXSBRc0OMiKIflgwLEMTP4f0
+f2guBnkWCNMg8aywg9qXRjbvERliwSeFoMAzr1IZdUeha0qtXhdn7AAXJjjZCdW9zQn9gpGefYV
0qZKlNKF6R8gDWU9/krhhxBJRgz9Tuiyoi9FRd+JWvglTTsagxqMkQJxf8BYTGlU+/S7Jz6jaIZU
fbB1ywX/3HGUPydnpAVDooIPFZG7iRa4M4oHrIOzPd3Sjm8Azbpu9noKk4m3Z9QaFYrVgA+aTaLj
+MAo0GDYUQVdV83rizxFw40vWdj2KGf9jrkc5djOUwXJq8G4AxoQTDKDQGcUX/6l5X1PgXcLEjQq
JRTj1NG4S5qOZwH0T2lsdKmB5bi8i0fR99UdHNxu1fW55AWBOV3FC9JljRJzuPVYFXXEBBeSITkp
gGhtGLIHqPnnefGbL4Rwuy/CzJZBpYz0rTkrV++aemOedRrxT3wwNtgUtsyFVh2k00FOig837PV7
qj+9FbsqCSQdDymOxBCEC4i+mejabWC9XN3r1hImX3O7Y6jhAgjsbjp+KoN6oyYL0igF21Eb/Dni
LvGw2LM6dR6hNNs9nX+UHsiv9P/7h6jjRWZ9Lj9CAYaLvc8mcxYW9GEq/Wx+v+eTbK73mcOMu/D8
jH02mrNUk3Oa7qS94YJUZ9h72uwqtdzvoSmyplY8VyXikFNL2vK9WmaV+o3W27TH2pfkf0C46gR0
0SF1QQtwc//nK2be56jk0QxwEhklFmGVtPkbOZZ1nbtyxqYB76jxiIZ8m/zB8Cf5Hu98gHUIT10f
Ff7MwHg6U/WS/CoI0O6hUr4M7OGW21Qb6VWLSzJ+dHNrVNO9wigbynlAF66UMvKLZBb8VS4rVVZm
osyZUK1XYIxSbWHbDxZ998jxkx1mTfIk0SisPKY5Dqsmrnxba8sKvn1bCnd4mGPtlzn7dBz622Ws
VbaYWnPKQ6mzPyIkNrlb2fJAqB36qbH1jKENPGmbpSOmQTNFxUhwyu5ErtdX+DW2CNtNlCVswAo5
OXZ+8MVUIPUqRVFNG8dNXdNOlAyP4S2oJFVDARmx10VOCL/eQgoxm4cEhIMoCBCb7r98Pj4VKRKc
txBhTWUoLvv0h166yJjvn7c6QQI0/RP9bfZXl9g9Joozj/mc39ctyuJAgu9fjd8efCGJO1bqIDAG
G8mEhjuDFEG3go2S/McZLImrKYD05fnYVFeEedyOKM8Gh8v66oyW9V7Tjdah33Q9xOQdX5LbY0Jd
Zdtnl2E3P7Ov9OChr1lvREe6u5HCeFQ+z8MnBuYj7p+1mNoTb8MR7Isbd6xnBXqHtUynq3v6XjMr
OYTCwRcdHssE/sMLki+v/Jpt0DY9hLKjMHDNOj8+VyvXQztoHXbQF2rg1VWMZXDHE0rKDH6V8p0L
AyJNq3yvLVbXAMDT2BBo888tj+HnmC+TInMcRW90AO8Sj2nWgSSMxFq1gHKQvcy5aaQEwodCjFLY
twbeZmrsLezwyClRNz4h19cn05xrtAHOgV/H/doWDG0mxYpMjIAbf29aTWvTjVNcTet3YLThWLLD
kdPD7J11U5FWpPXn6MkZdqxnIN3hvcUZA2Lo1pmulSSPDlc25sH1Sd0Uk832ryRY0OI1uMb0nnBq
n12xeE/cf9sDQ38OgJnmFyvw1/GBPPw9cwttMvSzyySXjYCcc3omYmmff60rsA7yRjSZx7YGoDBX
mpUo9IeAQ97Dh8lKkjwYt1Ta7aqnCCTYM2mbbSvkPOv+F5UPiNEwItqFa4Gd7uCuqm652A4Er7fV
ZJUa608BpKu9BEV+QwRTpzbiTMjqb9qiVj4f3CTSoRcnTFfTsC0Vq6O/tB3k9eCSm22Jd0pWip4R
ltTwjV/J5QnxmfSvr9qXq7sHbxxP8LtHU4DSl/UA1cVsteyaSFD2FpjTgUR0rpEGgGCgt9oiM0yT
Eus5u5Qfs4ofiAB8iuziQdxpp4tKF7SND7gMTPOeFQDfjWC4JGBEB4bwKWktoyjvwAJFU5TKhZTc
BuJ0SdjXdYroE2GJfAxI013b06l/VIpdRhajJtjMCPPqfCXyzUhrOXpxAI9xBs6SkcXEsJ1Xn7lM
MO8/UnabrAhWE2AtHquc1OaKjPMOT9ql59K8tXgqlPKShFPRWk/qdesSNpJE7zaIoaOwQg3N1I41
9Yqo+0rz4ta0YXJ+TeBwP3p+x7XlJc+fPApE3+nxPsIjlojEjpRHPtx0Tz8j6dPs48cCQjsBgCFC
2O3Kdm1y4eRI2CI38r96Dolk5Rq7RLiuvnbaGpbf8pYG8Y0gdTctcy4J6GpVARY+mKIM08Ep03FT
ume58VibIfswsFMaNo74ert92Blks8mUKo0PqW6I0JX53hdMyse7adkeIiS5x3Ba1WzOc6Pva1Hy
8mjCydmJElhNstNjEGnAi/aui2RZCwKSiN5WXaC+ZuZfWCyiWa/z1p5xUsN9poki6fh35Co3hStL
pt3rMdY2YzB8sUnr5if3uUVGKirFZrFhHKPOLPtef5ecbLNVv1hW0RMjLTv2cCFJ2VZosgZyvkmY
4+C5dxa5+7n1ySjuWAyZE8AnLhn7KoKZveUoSAQz2DhH15IfaXPXbMgTg2CBN8nB1HGet5OqQ36Q
I99/YW62WFKnToU37m+TbBodVetAXttuEh5vu3IYpkKCSwnOiNtoA9lOna4ZO53ak9P8UZ4UPsxe
EpXZet4yotcEeallUtbWlBqAeaWT1Y581hRJryWC2rZ3JjcdMN1gGwb8+J7ARUX/f4jdbFgffvm1
rO8H2664RaqzD9t1jTEqg+uDyD0UqWDKLednlYg4Z7j/2MDa32l5XuKauGBCZvee1laH3mhxuF8y
sFdf6qB0LyQ18Q2iBoa5qd8WE0PjGPH1pnsjZIyCbQ9/KLpsoTPsmEsF7DpNDXEVq2ofmlMf1+iV
31DI+tMcnl0tSK/yZpR8SD6VvYjEzjOPqJzlFqFav4ASTM09Gw3aqug84FqtAlvl3gI4lbNKZuKY
PRhOJwdbX7gVHpHTdLasclnxdK3Bl38B9yS0z7xXFxQQtfUBuo4BSlpg9AjGd8C22RFIyLb8g/Es
+L34o0Jmci0B9a8VYXWjaYgR54nDa0esmPlVZYjDzCeIMtoZnels77fwLw4n5pm0wK9ZFW5wPgUH
DnvSj+B8EAh1m5M1Z1484GmeIcWO+JfFnHS+jCjiYCyPQ6EcVJCwAiYdd2TteBO1Ij1jt0cWJoqx
Ftm0MO+T0QZZl2S4Yz6htdZq8eUq2DQHGZwiLAdrMqGuXbUNW0YTPSE3YyO9rTBgvnIhL8E4zUOt
tjElohGv1DIDf9SSZWiOXskXVfnFpVh12Mn5jfFtLj+Dpqq8Z0Gbtm/HuDYsXrZIqOMieLraQapv
1N1F5765oIc1FvoV4oq/hQrRrVKmKzDaJDksoAe+UtqFVTqRpJS1DJyKIT+kTUIoHKK527MNq0Q5
6RMCZ5vmpXW1mDLHfv9ue+gVHCH6aa/Hlc2k+MeIQmIazu5bnoq97VrJel6AHZy7cvCQi76kXuoB
lLMRhIbFDFbnV88I6Bft8bpvqzbNuNO3YtUMyUbxoi1vZ128QnqekU/Fak8grB7vLn/+qt0skIzy
Ns8DATP7Y0eqh7x2EsF6r8ix3nk1XAYzi4skIIzAQWOq9ceZ95lh7KMKx0WLsQWmHIEAeU6ZMNUd
Z4sYQkSW1J3mA2Kj0z1uIimdvzOMymByRGRSEnAxpm9nHhGfzQcwcxFEAYqHJHMPZB56QVbZmF7J
znAx6Xa8M+sOd9LZsTNzJrlzbAWAQgZddXypXPRg8NHuu3zKtgfMdBbipGhZCghNhf4EGr/973fp
Yeh7xR2OWdDRNcYlGlwK3oaqpgwmA/spyV/x4uoua6l2PVZ2QVr5hJnSe/m3Y0rHTobIJDXWTwDw
Jf6F4uoEQyjl/v/yTk2Llk9jVuKR9dgkd8lSWsLWglR+s5mM5ePCv45xRMFU7NOrRjjAiDN4u0LV
YqGQ65ZmGrP6zVppD461YH/T28LmW/l7T+isuKYaUMqvRwvDahJ9AuPXFxU7AG15e+kD01js/SZ2
6LZoqJsAeHFq3kbIMA1Gsbs/Bh97N4DWg9o7BPQ2vLQQNVGwem77t+jbunZkvMlO//lFAr2xmfeN
H9gKrJxMZ2winWVQfKUG0AqHtbeOz5GVA3xOG5bBAP/1uKxREUFzOhdVgUXIIQWE2W4Pw7mySBv1
31VtZJq77XnG7Zz49ivakXY0FiJCTy4fGGeVmkiU15FnJkOgy/SHNYdOyIsdoAO5KJSycsVVrhgk
t3LRWwYGT0COgz/RjvQf2viy3vqwLmh29XxXpDazzMrDhKMQtd9aaM0VcNFe1P8v5cIxjAZjPCVw
L+DRlLgmsB5v2cTfE1ZATNu9FSTXaC214SjcCWw/E1AoxwE5onvt+7D+22cG8mc0++4DZinH3Fdq
mWRDM4pJFM1oZCYd9uaxe+PFxSCHbwA4jKhIDv/NQuogfUttVyFRyT2nhMciBo08ROe9pR54wbSL
6QAgTK8u7QkLLamZYUXvJGVnzHcSbY1OoojmAbc+dHsNXJZPJqebDFuzUHgYroeNF04GVIIYVhMC
JAJFMvH51ezsLDvBB2LUMGzAU53YkOqVsqs8qsiCMcuyU81jo7ArHIs13l/yqZ/r9QqOHwIQA7xz
7sY7tV5gEvskSblcNLQlLTrwQxJosTgUNKTNmLm1MjOTyHkKFvnzrtkw0Z9JLrU5mA4hdPDr4dMT
ol4IRQlsZBmlK5kQVLwOIZ69s+NzbfmsR/dclyC99/dnW+I1tR9NI74+YT0H7mKMm2ZegAMy7RrX
oTZZHn/JlGJPaGb20JFu/vcSatUWAG1sYWN3QrOM9fVsnME8VBN0gB3yreOJNtJVh7xclclkzH+F
TjKluWDDXB8JWioBpjXn59U7hj1UnD9oU17MgaT9AL/VkXpbnvbIRIghebcpfAJdsWpBwRpc6efD
qw/jfLs64gNgsh9qshfiGoeNFBfVwjlTZdaRW96++9ODHndrWtQ7EYvKIyRxX/L5xzhGLszMdRQK
VGAj96b0DIm9NrKJClWXsdlxURk7zBcBws8Zx0TSGK2QKubnLTAjDnmOaF/PhM0xpfph+BB7Vil3
FELYPZ2NGd3fPON7VRwXWwdF0XYTxyOacSW3S6bG7WtfcZAFLF42yI2k/1ax5yiaKiuOxcExFZEb
D/zH3ofgzt4e+E1CwOk4Ay7BlEGnx56mOb77hwPRUfUnXm5ufVaKC3cB0bDteKXhhfyqnGZTiwus
ltsty8wUnPCRFEcPxPnxk3n6BgviMfCRkJsSTfkJAPS0qN+vIs+t2d5y2QtbqwbeQoZkg6WHF4Y0
RSXbocGqs8AV4gP4kv+rrG/nQABn3dC51s1JIsSxb4sqEFZ3gm0qin1kgdWeF3UcLnIm+qknSczG
ST8mviwX1C/6NfRqfURXmworx9B+qn2s/qzrFXYo3CwWmpGvvcXUv0mK4BDLIpeYNsW1RAWTgIXv
GWN5mYMTkE879eb37Vh4tqsc1X99hnU95O3PQrdmZzmzsE39oRtLc8wyqJfTBOQHCH2tgXFY7hU/
76RCwCbdoFwnA116gRLEXCu+KvwhQqJMKuo5ckZ/rXRS1Sw1nVU/cdFJPzvc/naajsJCfIG4KNlW
Q9xcLdtGnUSl+ntHwAqzbtn8wGVHnIP6mz3G5j9Xqf0sWFXUpcefTYl35JEvO1GatzS/GpRjaoKt
diPEIcjTKNtmy/ys7H+SDpsYx63KEhKchOTZQqUJHSRAQAvuMUkLNR5N7+iZbPafusb82z0EamMS
nWI24o8YyXWjDe0jvIYWMOp6+pp6K7L3s4CYoKnFoHS0iIAZG5hQ/bA89A8UiEQNjM0aoMo2UlnH
mHIia7NQiVdVLBYMvcAeaE60I0Cyq6rLIpRlk3pQZ47EFdlaGO2t0AvlHGUY99HKXPhJ1XZpQpcG
xPLhpLsvC+HByEwaD9HJyexYKJrOcZFtQEvY0Oo0wZDIDurbT/Rn65nfcPkV5x0nofRYCWHyMCW2
V/S6mKro4ZRhs1W2wezabSC6ZGYNkK/TIvV1Y8bvqet8jNKTdSFDN0lEJzoit/5ExKM4Sf0uRDaL
kLBpnfS+7LfZDhzQsec6ZJojdsaN27nBYvCJ/bU5Vnou0mH8WjKm7SqhoXfTj9wPaMNjkKOa3iad
STpOH41ItNIyc2AJpqbphiHllwjnzKc0FMGhRzZFC2XVUpnL8pp7qaUYaPcsmAv4viGr3YNRNhNK
L6vCh/8h2Q3dzHmbE2iM6bE2AseDYwVw3E/7jKcZm4A4iGKfpIvLzf7mY8crzJE0iZZSXdNYlp8P
EC3x9YUYIdl/yJHoJSVPpkF+jVK/CKwSXJiGl1yU/qDgZaUKVugl7qMMpYAFehByjV86HempENkE
fDXSqC2/Gt/A8s1Js+JkzdUhr0C+hATj9y4lg2ZAbQSUxPxCjPj4WcZgqSYJiVA9hOZXVg8tquQq
xJpVw/wTTeiaXpJM/rxbBtZtpCTBQnHrSs2Eg0AEpnLMb0kLbTTsU252czlmQuy9cY4v3gK6Vu2F
/Z9SWMmQ8h9uQojfBkHfJI/VEmk7u+FxJsZk2XdqV5ypDTvQjuEPyPLZv62YzSNrpWzJy0WDviTZ
dFpyTvSkCAZOehNsYX2ZAOoe8BQdQLm07kaiXAGTQgaQB3VVFMrndUEoDCm5hE6Q67smVHMtXmHj
VCscfrlCqCb9jFd/tzeGzMV1rPAZg1QQkueBWKdNUI54pOgEg1Xda9wCc7PzJ0fzFq9AYtwGM9Y/
THVyy/wBAtdXduBdmwcAt/KXqfnj4TXFkBOj4D6Cmq+VGQzE4ACEw2rvOFbMbLh+WE3X8znRs7Kc
6apYtTvDW3NqNOUT/xJpGnpAt11bbRD7W7IHSaBN/47dVyGz/kDD4Q0Iy/jD7gOvI6ZOeyAyrDX2
g6Gfo9OpB+dZS6g+qqLfYA0SU04QsAP6T/48t/2y8fwKGxzltGJ0mWamtGCTDZgq4MDlvMRxjM4a
s4MpnSjbLRZfsXKcRIPICwOWpcxCjEHmCD/w6OKqkaPEsEXU1Jh0L4WWzRPl5PZBwOlL6i3dX2uA
l6Y2H/m6qGKLw51giUPj8vY3GpxISBmYk1KNEP2kCLGaWHkXbZ/i4O2ElFJp28PNxolgE3mcfXDe
qSsMYKWGO9CfyNsAyBOwie6l8KR32buDRRL0HR3Q+h6rsraIA+pDDwa+HxkDIVS9DXyp/NLDJJ9X
Rp60L/laPAaUhVAwJmkHxSM6CLx1+Pv+ndYUtJ3easP3cWKXIYP783QkohbDSBOwOrR6DnUfmYPi
qZIA1pYPXOL5ZgTt6r9ENw6RiQ/wKWATUKSytAH6H2nBi67jaXi+Q3TGW7JEvGKbm5wcmor9xV8S
Xl4brr9i5D90qRzJhgKwx5R3hbFKt3LwDFC5Dm6vvjDxEvUoPycxswbc4S0JsSusyKxwe3/aIiZT
TbOeVp3zOYxSYM826yKJCM2nKHDB0e6xVmmJzJWMhc0hWYF0iDOHtS/TMjJ/M8pIY6Pb0Cqq2cp5
AC5HyyZTW47IaRdpmGUaUREJST+HWWW92Kw8rLehChKfkXjPDuCwL3VBx7o1GgsW1vsnrrgQaDjc
DuXuyt0hTPPp5p19aETnZVf56WOKOzjmPT5Hk/nRHP5kFqxUGyv1NBqBVH5Hi6MUmSyU4ojHUkBz
piHLxyc4ELL2GkYSG0Q/o0aAvQ4cAMdZ0NqtCOLYJW3ZDyRdsn5RbkWDsHcv1p5v4l+1pZkp+DQB
awTtowKAe1eE/Nebv+ru3yP0xBY4jCz4HGmnwaJk65YQgEhLapelQOK6IYUVslTUmKzGqwxWDWL8
Hp7eOEZcFv6iSGosV8thKLHIl5hHwL+S0bwGiBQ+jpHDhZUhsEu12jBR+jLRSXyBtV3OXZ3FK7hM
ihZYLcLSmVlFidLBSCD9fcvL8gAHvHQH4if3J2LJAAGKNgjkNebtquOUMwBylSk50GClc8nkwLyP
QgP9TWPEsLF0JPknssvXjbYCT6vyLjWXrU0gxAjjoXOTBp+4HNAP5ZiAcQ4Xe7ikynexyKmD9uwH
1Z2aFDrUgXPQZFVF6U/Kd+RKOWoj1IEKJzIyFwatRSBHa+Ech0guG6U0kLUU7efV/cE0TNTYgrKy
UR0E8l2ncFMZw83lzCtrhoZLzTR8E/PhHvNP9+8dAGx3BwZaA1MFVx9b5fb4QJAnOwbMLbEXv1tq
nf3Vkaf7lWoBFi3YuUGN8R4A8NAq0F2zcnLW1wOFP9ulSlKW/49cZnD8Bmh6CWecIZYwv4Vv4/I7
DXGF1aaarmk629Pvii0UYXm/aldqkgpr+xH/PtVTbfYTaEetuXiesFK+ns219zkRx4tS5cO39T1R
56iSbJS3Rn7Gn1Q3qj6IKuYwaDWM1A9aFtaQwyO566WxQpO95xRVvss0QrMwiZIPrC6P6lap700b
cHC1+MgmBMwgUQ2sBBu0G8QG1ts2+NKi38sHo4S4RwKFuci86HiP64uN6xB38wloA2XBpKpylsAv
gDySOJ/V8wUtqcoYuTPA5A19LpSVWp3huAOXCXNsIVzWk6f4j4trlADqV/MKY0l6AGGawp73Hc4e
nYAvfpnDM9LgB4lfnty6Sdm0bn01+aILoVYqUyNokRD9qfvoEqoxbm0brN8capFyVuETOIfraiRd
LkiHPROaZYgQXZm/5+2HJ/CEy8xN9o6KyzWORumAq/a4d6dTfRK5RIKoTmSEonv2L60YdRv7G1h1
O53QQLjNnlgJ/Uov1yL6MaqXcsXooP27bPczpOYKyRP3YpUzCBtE37mRbSsd/RZOF+moSgF4dNMA
zAWLjjgYHEB7J7Z0AqltPnOj0iWKN4Oy0oiatrP+rgeyMm+gF+dgqUoPioQ28kW849oBFNHQTNAf
S5IcnmYVLveK5bT/Y7GYrAulB+evBFL4HSuKFruLkCqJgGxLUa4GaMcHPldSIv2jLFDF8CKFphbv
JpOzDu7UiIdu6kUwVBeuqp7hnURNxt+h8T8DeRlmdBsvoL8Abw/Dd1hTh/BzuggsC+QfS9LshV8z
DeydomkxDVhD04R7tSXxu/njdH9aOkBRi/1672q4ovCcJLYUdmNxKTLLKl4Ny/orfmUyjBaGQw/s
rTdQU0f18eC8CHXTzGEvuRVrmo4xM+y2X/UrkBeS777ssWqC2FAEUYfaljiKGZFMA77XiGiYvgFR
acj05C1NDnKtpwSVe3NhAeSNpfmKDvJe4BL79zLHe3L/RiWWKg/g444d56kMumgF79T2y6eylwH0
VGKDs3lRyHeVuNzJjmFg1rULVPUDg0mVlNg7KPh03RCkh1cYsB3OnbBWtfB8BidSaEohxGSWQ0oQ
KxgywbrOrR1KaBrhyrbqiAe2zD6rWMfk/Ds79lgeGO4aL6GuOl63kCg44nF+PGh0S32PrsAHhqB9
JeCi9sMIDnG333JhIcxjXcY4hLqLkm0RyFMZH2QPA8rWrqenjOpVbOYiB/ufqq2fSx+nl8fYsDmW
Ewbc4TK78hKpZxYuUZS0ho3xp2eD+CqFG5cM/tAOgHJadiQnvbJh1OStfNnjwSUtnZfi1kdXYxxK
1TQ41JtPmL15qRp/s8fjHpSgnLkBt6OyZeYZpWYaZRuIsGr2dIWfPcu29xNvvtTWTMNaafnSs3Xk
QxfQ9JvvCHc4r7PWNcVfL5/0uajZLjH11EhWdOeseInjkelm7xD0R4X5G5OQrzHYJy8/Y+6WMDIg
R3hbfZyfoASS8DwPTpsQC+SwLuc8MIQF9DTECNejPjGBvxc2cdxyyYTznP3vPuePyss/a8YwmXse
ZQmDXtN0dMv7TpC21AWo2e5WOx3zcutw2GgwNDA4uhTqUg1zQ5QwlnYyqQDOLpTjHOnvPqgOcEER
HZF/4nI+PPQAIxh41DQwjttTXtLH5npo87tZGxTCKuAKc82K5jWj5bBdgYfyx8zL6rCBYwgs98tA
Te9+72Lbm4YfUM2s6iTDHfJDVngRhQXNx4qp1jiXkiSF4N5Gw+n4bpYvF+wl1i5joxEN8yfH5DII
tZdAWRZXgEg8ZodMxVW8wadmBiW4gt4vrHRJKEK5ThFN+CTf+tnYe2kghhqXFWAzaeJNIJcE+XWP
ohI/4MOm5Y+aew2nKFVGNwxxYX7+ntH8ipTwEivvpNiAIH8ygHl6nzugNg/zadyorlhaue6yBQIn
AnDX6aVxasiqQF/aj70AadEVYseuNFhw0P8yKMw8ZlBcUMd+YpEKZ9PFa/6dwVvjUXdQ01uQWnNH
f2QFMgiuYqY9qdPJXT7spD0DT3nzs3GlVIuavx++k00kluthYt2ytrIzpOtP5IZx7cI3W3YU1aWe
KTybNKdRO7M4DLWlKCG12F6u2WxhwlcStimY1blySCIvWL/RhiwQxfzBjDeXKoeybp0EjnV/XHI8
AtYSriBGIlw7oFCq8Yf4qQw4qGXS7+l3yJrK809XJEkPow7tawN5ms3t3PyEAu6OhljuxCtjrieq
d2lSlFxe3xHEqO0z5YOBJ+x9K4F5BSbeqZ8M92EVXfJqgD9+IymY17XOLTqkytmu296QftPX4d53
T5GSOqWzjhTudCD++CzZIk2+dkE/QaHbb4T9IIww/GFA8IgBIJ1cwgJPLtMASybnDI23hNFVNZPm
g9zATOLGpl4B14a8o9zRUslrtBbUYUcZ/dE6Ha/Vjlg2nPs+lrd+dMfocgzc8vdLCnfMDmVR7VYh
Qkf9QkeaLVwQFmdXn7+l5qn0Wc1E9sRYKeV5XtIy1/hBROFUCsm7ySgO7lCM+Fg6PTNQBDCVuzmw
r9Qny0fXCS0OZYwjFKlGWy7gctJFiu5YbBaYYxEodsklT7u24lvinTw2/jvD3u3bY12ba/yNsPaB
3HOKLHKNHVIo3zTOUliSrl4AQ/BW9+qfLHnwNw1ix0dasSSbt0EMWRtD2Uh2bF2lKWWJsvibUE/q
60ZnqOrxwOhIz61GzlN0bXNoEQjPVWf/Cb+znzO188HJnQQs/yZPHqJlTI8/+lRcIZcxEyxbGrPI
2A1dCMSRZWiXfIOpLOVqIHYCY6AQzrPIdmlqXICd4pijTHgwvQU1ukCkkg1ZY5DsXc9uarvIsn8s
CwrZjTXeaxX33MVx9ASAsovZc2RcyMZtfMRnIzh5NtBoW+zEsfGQpea6MIfqU37iYg1nTbXoQ0uX
3ZIjpOtinwWnVnYaLwwNdNFrm6FS3szajXM4OHjSSJfVqFmd3XZgAPQEnSVbxcDNXR9YLZGPYWfK
DpzfBXmNU5lM1ELsDZZ282R+ZOJjPPuPyIcXaxqJ0Fwnfo1GPbokmUObU6t+4JKC4paJnSoRQ1+8
2UasQbbMwLX5+3BIZrGBnw3RTT56rmsSLlpL2RqKM5ngjcAP97v+3WC3l99fzA3Q3NARbe3jHOJr
zIlGfvBiLSb+X6Q8i57TAdD1Cg2ondOXPGQhfvnwFZhQr6KX1uLCCd2TmmJFtAXXctzTYqkPLh3Y
e2Adc+1WH5tIcz73MUMVif3Z6Zz4j6Q1wM+WARKq+9tlxRjqRPR5YKYBqj5jdd3sUcrGFu3zWJC8
m87uLv7s225QZj1rZtB1C3VLta9gfX10JEkyt4V32ZLUE3mFzcA1mwRG+jx/FX+bLU/5VyvP5eUX
YaTCiH7/NmlZthO9am+Mfp/0Xu3Ge1VquvzWTPgPAVXMXoOsukoJ9TdAEQZLYjaae3ftP6tNG7no
FvZaYSwnfFzAWhe0mBYL4yqLDnCrAe58k+sOGpoSUevKE2hN8n9n9fv4jTsPKklA2HW2UuYb8QWa
xaNTg6Cr6g52p2hQm+gp5DpHkTlBGvuTVbRDOJIs8jRzE7bLpXx/EFtZCLmB/ec/fcVcflKC7/I3
uqnJMXb8JURul67+UgDoC78vPwu/iKS1xb/11iyOsr6NBkXdlsd1KDiSEqg/GjMdcTuVYUp3cwN1
ZUI7ShmzngME+d0UuCaq6GlueGqa4VStZJpKWuuu+yGMK7I5W0IrNs2yHPicn9pguh1RxKW90VGe
LS2xn530a+2uiS2X5SBgI5x9X49HhOE54C8G/nAu30n1MBrAB8wWCh6WzxOQ6wEPYSzSKrxuEgcn
Cbolqqi0lR3f3ASOfEMrR6ViRMrbwK0nf5T1XEPwZau5DvsvlP9tMTA9IXJjpxKRTRatFFMSmbqN
dQ+pxBkrcDbnqEvfunwEo5NbrixTrzQPj8xyy3hsU5ptT8RHEBH5yjIeF7rQOLKz7dnf55rm34qU
K3+vQ69Sd/g64TFuWFAx0aw6fZ0EqmlLM/hAhJBIeJl3ygP1usIqo6MM80HZvGEXwPtb2bQ19STV
VqyKURIc0ltwkqNeQSEib6YAVwjsRNM0HD4vRTnuP2Lzs9t7ubpKMa32eG8t20NIOxeE9a1VUpy3
tZc7/vXsHaNoXHFU0abfl6nT1JodMkCj0ij9ylbEQARNg9CjxGNxlPZE4M01E/p+QVNAJNOWdt+/
XIQWFbOM5f+VITC7YajD8LcamCzlsp1R4I8ax0G1bBOElV+sO3YB+PwMw0+hya2+eLSa2BJD9swK
pGdkP+inp4OAfevvRknktSoOhoPkJYsMqnL1wxnRHajHTyYCr4S+EStajjiMvLR3lExDnkApDzgl
pP6wz7aVNhjuircY7/ThR8WYJNm/P5fjFb2nU5hT4d8ycabXXdqNqIDw61WGuMtgNBYNxHuQFpPL
OQFp57SX3AEwlo9swOMvYJnivV+7G8Z/KyV68sNCDUxK3fsCZS60evSycgpmxh/diYe35vd4gmpU
RRghpVKgueUDbeM/c2+GQJGbZV7D9Q4Z0PazBrwmVfD0I3iWWxPwDf4m5NZNotOISJofUaSTtwm5
l+qYT9XU2FSFTmXIltKsx81O04s5UTHftiU9blriLm+4VmXrh2xbUJZ7vRi+C0AmrXtXITLiG1da
HrXE2oRM0gYLgTL5xQAtpoUXz2GojdVVyiWv76qk2V262BNim6D7KmXjjvgfputsYeclbyN/uqwd
+Xz4TnfSDx2J6944QVUinLWFqH2sHQK6uwXt/B7dIeJTcXjLzWmnd6y1cP5wv4/N+xOUO11scoxH
yBswVDw9HmpunNIBtMaoqNefcrmKFhJA/lKDE7aiiqVa7ztZdGPssLHzEkO7PwsNk0Dnl8b/jJ0D
SjsQWC/oo4dAE5wUkRyn4PO3c9hsHkwKKHvKhfYf+T+ZbPnyFtrvM67WNTYL5ptuAiB3PXl03KdA
NKPOXQW5yLT8Z8b9rz++kEfQBbeZT93FGBLCekfA2g9F7muR4C/BeTthjmUfDUqUz9/ag028DWz0
cY51fSrh0PiaxBNRNk+p537GLlAh3p93ytehnh8aqfNGF1pKrJveoJcvYQz51bYXiYM7OY/xZCFP
4AKsNg2WDChFmPk6zYzuwL5Bf9lGu4w+O/IoycfhRbpVpg4hexpN/NTFuhCmpGkoZsAw1xa05bp0
MPsNii8x7KK+iSX4ik/pI+ODmMHo5ur9MH87VFYGQ0iPOqoq2CDk1S/STkU9CmYKnDQYjVcNOfqj
G0+L/NZKKlLTtI2zAX6bleQfrDxUQR751e4eb8MDqH0vJ2VmSb4zpSP5v8m677NbGN/bjpUfZUA+
EOi7YeiirHxdkFOWNTX1syIUcEdRdOVDqnCKbFmiW983cj+pRi+hx8nqPHaRqAtGGSsFjdYUXavG
39nxjU4DCGKugw23wxg2Bf3E99xDwPmlpxtwHFDQ8TmZAckWpUcprMmZo6kO2Fp8ZdChwkhyx8u4
32AS5jy9XAt3wvuppW/uk1GVF1Fc1GVYoYZA2ay9uyJTwrgeCEsbwff9R4N2nlfc8YiQouY/U3EW
rQrb5d6osGcJzjG009mitwWAI+t7rKlt4foB73YP6oZKyBxWLtAqr6PzJOr5pxYmfYI+1uqBV3RV
9LQKUED62DMIpWCLkd4hxQpmFJ0K97bZrI5kyj/uINfXRms1EG1grLXXIEE/dk4bPsyh9slrGZs3
QZYru9asLgWO03C0o4CzZjmaRQg8QVWsOyHnRqiHx/QnT7rCEpb+uSrXWT1Lsj1cRZBm9Eb98qXF
yBCZybV2XWbiF8DAHYa/bpehOeiCP+a2a/MOyA8dzvsL4AKmwBY9f5klQVN+ljwx1uKnXw9pPFhw
7aM5FdVJLVaGjcTVJjz1PrZ/D+gh/iykThqDKYLe/CCAwdD+JwozI1D30gFAERlcqaCEGfePVdGe
xmmkv7hBLWEthMv4LMos9kpnV6W9nt7Q4zlgOQRSwi7WOeiMzAUD2Qho8fqi9paEU0avXB5rLxxN
hNIrCqqx0NS2IkD/9c4mH3uK1hZPZy7P1h+Xu4QKAKMgbpgHseIZMgJPnthZeYB+8EjyROxSoW+L
lVlNT3+6hrmyl0L3DmN3MelVX7axc4DWJdH67yPiwDrzD+bXBI1Qzs6l4+UXzpB80yGC+7MNoo7j
ec041wkTeL5tKPcp6ZAHSTz444vCIjYfnsiTx7SQ4ljTkxxziDZVwWDWyO53oqcm8fVeXZGSoyhh
QqUK7kABPydZt6udA2FNlQl6i/Lw9ANyXZ0Ov11QYrAj47hygfl9X5HY/QVARtFDH8fpbsV22OtL
1Z2mtM1wxaDP5zd66OLViKXmMSGZH7JQ76IORhWVj7x07e1MY781tJDJpyDB5QkiTK4ymHQu3+N6
BBqoVU7sQl6yp9+WgGlTbLi51J/vYcnSuOWww4FkpwtK0ylU+qxfVgcQT7y56K2HaaOuOntFebAJ
fJkSu3xO9Ee249StKN26KSKnRCNSmBkCv0bJiBdqfPZ+xxTaJwf+k/JgksAhtX4ejt4uU8Zt8LWC
dAzowJG232LmG6+uwFIvAtvAsjxci3qs3iXoD2HT6fRIHFj6KfwsbJQuD4BgSvo92TyOhvOMwDJM
AvjflL312rEJSdfZjzSwhVhefepEcqZcgDxDiCQGJzaz7RKhepZN9KY3K6ZE9I6WmNSzoldEMVDO
OkKZ/JPbYwXRU8BUQNSiYIHjZSDyyXrJhR87LAr2sa87dxCPQH8n9Ps+7zsSbvj4p1Mot9+9Azqk
vy9ag6c96KRJto37ZXDiN4I2lydLKQqF187ek1Upy52Wo5tEOClDTzaPPu8/BHjQgQf9Qz4pdyXU
H0WrEP1sxOyKwxmrlSaFLgP/myUZJaoN4Uvk0lJh7Da7J0qsQadCMwqd/aZYmQFZt80Smqa5cwlF
ICf0gz2c3MdfnCKPrZ54y1tuHvDy2I5+GKpBpV1PY9HyxnBtrWIH7D4k7N/1GHDubcP2v97WEPb3
2U3BfDrbXDyoKsOR3PsuMwDnNHmfTQLKCIudWBbnxlaGCRC5MeWpR1leHVGxFHWf2eBv/ESqY0lv
xBBwcPKv0/20biargnOuodaWRRez0qtPde8/3MdF87yCOzCf1Z/BFxLBArohnziKikJCZIeIMljF
skyZC2I1G8lz/yba9lpxvTDaf1GuqVuh83/PdJcyexvDJoDCP9HBQmEPhqElpCM7EPONWfhi8yaD
2rO2SGs2ZILKd5gBygltUUSaf9oWAnA0oDyo4vEwyG110E/Ds6m4bmFqKizD0+GcVlJsel3tmm4A
K3dCI59uuYlUdN158BB6WbwmkpBEfDgK71SBdZ54UG+OtwDizxVnNqZ9ZGZNcovRrpRrk66t2b5K
MuTq33NS6cIcqIifWS8Cqtzc0eZ/uMt6UsNhNTQ3StJm54I9qHYHGihju8YWGDZGK63lP2z2ZSg8
jxbfpibgZXw9izV6NgLxVSU8jr+ZPcCAi8Z2eY/6BSe3EDCZmwe/eH5Ocnstu96q4SIoHJm+qFOa
7UfmieM96pMpwGpgGFZWOmPH5jdeTIrF9hexHEVPa+DxzmY2Nao7VNkIgLgNC3MH6n0OS2T27QOy
ES5u+Y6lTPi4LdcKzkQA2pblIGMk8qj4xkbwa9UZsgBuocKK5cqlnJG4K6y2IizsXGqmC/u43rBG
8PMEhC6C7lFXy6CZgyp5zOmcp7KNlczpdasnwftEZQTIMqRROYqtwcXL8km7CxbAGkn30fd/xkCb
kq+oNNoSQi6SvlJwh+4cfucfRKPdDpnp0IBdzy9zt8HNsvHGyLm249QuTeGHbEzzwjeEcriFvLAe
t3krRbaNBnf/9RDOo3OwblQ4TABzjHnA03rdA2wp2oMQRoPuI51vt/Mn9rBGuHR2a36wIPzuyNJP
WGDWXkWu3oors6hQ47ksV5k5HTQWAgoGqf9nJvoYZG7BQGB8P18j06CwumWuHZhMbDPM+geFqqaR
TYmja6wZad/UfaMZtGWX7BzqTx+r/OGQWCbd6lreZJNVjdWtPjtFIVBF7hgEuIDzOqRFgVF7RBk5
xgk6l2HmEMKWttlYYWsfeuMPq9YgtTBWzmL8inqtSQrkMazLj2g1hOzCUDSi/sQqWgiM+/fzS3CS
1MmAwFxWZAM3A8sN1u4Sm+rTgLGT8cfPitetiAj7htEwxZ0+L54mCJ7uMBmjRKQYKV1RUxtOlbYR
rLx6yUkjLA2N/IvSGtL6zwQqzvrYYxgNrjMicv0fMmARiWiuRnQ0xR0szVMV/nwyDvkC5WziaGjv
gpjNRnjPPkkZX7OLOe55VC+vqJGFLorOXPaExSOL2FtKgmG/fUnmI+6hrs9V/3uzo2SvaTtdPBGs
aKQgbKXJB+KOvCHJ5znkHWNNIDs28YPtBvOboJaSZg3/xxBUgj1oCEPJJYq0C+226NASRc0L6XxC
uVXMhLtQKD9NCowwr1rCOXEkc6rv4z949IHPCuelw8Z0U13QZfSEsOmNnNWhPLezAoqswyQGmKUY
8F88e0gESxbB8Vv+/o+GXv+R6zbskM6kFbWmzDaXfA+WNoMcp9XDY6Zk5/WY2jD3JLpMH55vwbSJ
L27ca2a60nKXyQXYKULFkg16bmH3rb40I8vYOtgtTq274JwSEs97sHHVS8VyANOmriqhupPEnN3Y
YGmH88SR4cVsHXd+1Ferls1MN2nkM7ejs64d0q14ajkfZXA9w2NHKJGrAEt7IOTiivHFH1URoJco
69TU4m+TFyK2CzDHP81NUARQuVTU79WOLAPjYOY297yjV71codzQ4OMPY5OW0hI9Tc9VYiIq86nW
bxBiLZ5RkmnnfZu7CILoI3Ru5UGd3QMMqvBk8JM/JqsduEp96Vl9AodZ9B2K+ylukqN+reHfh3xq
8XtZL3ehDUWklx+BGd+LudKc7aTzfORxg00d/3f2fbTF2o9gTss+hC1iHogXEvDfb36IVKhTb/Jr
YRKklcsRsmuOoAtaiBrIqQVgXwQZI6Z+PvY79JHR8FaCh+GVCG1P4lTFtolXjz4uPt/wnfhe3aLE
V/RlFf0sG5yPYiJurkDRTtijWQcewPpZoMKrGiUeOun4BE+jYgQsdP0zMzphH0/EgjB6UJ1uixG0
4wKqdITQSGDUhUaaoEpmWGoAlvnaobkB49KdYcexZOf0UOuVzLFh4OcxmaR8WBO7Ef8aD85a25zs
UBf3HGcdIAmX0iiaTF141+oEB2+5q4q1XkBCkXMstG9hczCpwAh7w70KHMS9aPt/HBcqVTsxR5xr
CITneQ1hfzB4PF198+rovq5NadqGaSFLVLQWI1VKO4xaDqLT/TPDjPlCgrSQpJ9f1CRNos6omIc0
2UCtHYES23KWcj3u53dh5GTMbtxguymT8FjjIE2Et528M2A+RF5hWzP+YQleNpOM+fuH+VAcwzsK
fF0cBJivHGa83CEf+ZpB4I7M2/H2Q7zjXyKJjW01ny3spL2675WXnOJY1GumUOgFBTWXrY+1yIly
UQHLfCi6cSwG8mWM0YLmowks5dZf8wutxdbpH2iaCYKSF7FwcV353+esGWam/umKWXCGL3Yt2yzW
sYASXyE260bgOValaBQZ5vw1Yk0sqEHK/q2LU2icniekFabJdl+hUZ3ABvEU22axwK/W3e7kdBE5
vtujCp4jLdMDxXMeTRm6+7scNGnxok2JABNlhaOKQitnT8mutJ1KBbiYsvDhfn2QiDXBsEJ0EK9F
iUNv9TLw+Ykm6M0SnogvAmsukqO6ZiCdiFeUMeIiRLuL/T/AbuVi+8RsXdOaeMZpR8bZNVN9c3+q
Yt6mmwI8xdCXRVNc3EtY2Ig6LKWxMFAsxIBBuKchSgODrTtNn4Eh+Bdy8QsS3JcDsoQHtUf42OJS
nZcwaHstGdQhNoInOhY9/3QZY5f8t+ZiTAaojzI+LgHqLkmql57vcfwkBurYE6NNvjgtOWVQZ63x
vhVB5ZchV9sp4cEHAur9Vsi8WleBsrOrYu3mTmbRpfMyCJ4pR+HgqhSFJKOiH2jwKxaBsY/lQ8H2
3DI7Kk+Jux3pJSPxjM63j+P6RfhhUG+HcR3+rcYFH6hyV0NfSKk8hDV/xdwR5HPK9WvjRltG7eXc
licuImMrGZfV25Og9vOQwxqsiPuat6IlIb13CM3IcO9r4ZGPqOixSsO/kX+9vSc0UZMVVsr0unAu
7TS/+AdEVKADTc2nOdu/ELD8GsoPFn5kSDNlt4TKjbw2DBvGW/43COkc9fyChEFy4RZPvmeaWz2u
Zjc0Mno7YCH0I/f/CRDi8AeNxhfts6FAqu31EKJ/jdwHW2XEXv+OTuBpMxLOfEeBGaDPWBE+G3gu
N+fYvUf4AXtn+1jB/3RhePeFNXEHzsg746ZQrNGcVlpOKpHu5JmwLrLR7IMr8vfnVVw7GVGoe/H1
wa4V7WwgNZuOLeeUOiv1KkkuGio7p5dwZnxfZt1ZVA4ylkIAJY4h7oVwdA1AcLnFDZQsGaVD3ShS
NXcULJ8/21R6SXqNKkKSXN34LT4XnXHi2G5+STZSVhsDQlHvYP+OjUntCoYMSNyCwEU/1HgSMNGV
4iBtxLu+1HayMjBHD775faZcYBLyHilENHNA3dKRW+O9mUSzIewzcMfnY02iJqYV9pq3X/nBtPE6
5NVZrQ1JaEb+r5nFb/Aoo6xXQ0y/8ggtR8NjoSmvBCZNi3TcXGbq9GuQkt2Bqn4kpZ4jM/A+8r0q
5WfSZnbPnNEQhip4GkvCfDUKPxwSfIOvsNSlTk+aIIo4L0PA8D4ofXn2vYBfISYYGz8Dvw7H9PBj
LmGF4HrXf8ncwhrHksmlcNXEQdiElXaEeV6kyR91jabgqUOtbyepbm0qwuTb1PgtSVg2On0NnnKY
e5i8+Cu0YTiVTtpuBydDnpk4oiK3QKsGVSRIhSGtI6EcZiVHKHa9L8Cpuu1DO3uZZ32TrOy1KwRj
ceL50Z81XH7Rt+V9lU2K5paLUlQxYtRzNz/S0w13ijgGmraZdOXARDH0JbsDe2gZ68SEcv0xYGjE
8KD7NoTAJvy6qf6BU6Jk0pcw70Lb8kG/VI+5gdMeOuKGXi7DHjQxntwWIgsQ4hv/MPAzbnTUf5Z8
ZYALea5q1FJqMkIX8eLzM2JJn3KJdl66ANE4vbAoQDPgLFxufKh6Fw1qQq1kjH4r2gs0cYA3EAKl
7/PpI9czJF56Tv1iufmYVaedNNiiJT/UyaYLJXIUWxSCcQ502Sn1u8LKi6hbvIn0I+pe/DqAilGM
FtrYSQacp8KWFIUdJhBdNEmtaG34DhLZ8rnVq+YMX1IEFObJTOA3VHmghZ1MqH3Y+F2SU2mY5/Po
QAQP/FYxbH6uNwj6Yj9dcdORJTPOFlMaXPmZo2jnagvsH+qZEgXe/Z/WWwWmvy+KtsPZHFqM8MO/
SVj4Attqod8ZNFG8NXoXipM4b/PNLlJWWMml935BIOI34RerUu9OfSfUVg3/o92hyMxaK4gsRar9
EEAyS2nFTvYSVVl96+mhwrM6ykTCBy60xuGCrHwbBDPNCZnzidTYLCujAUVUxHpWRuPUMaB179Tn
u1kMyn+NzOjb9lz1VMqmOqi0EmHVd2kpt/FwriaURQXQLYMs9Ps8e2z4boP0eWcs5fROZKpBiybw
FfOsS7ENZmRd4idcERuuwz/I8der09uzslXm9nYmKWonBNQlDRxKvoIYdZ+GH1vYODlCiYXvMtev
+YmghVf+aThudE7q5JuhSbt6KO873/sgI6e2kKjalzvuqGwAhrl+mTrd2DJdEze6YLe+9ZnXulSZ
kcAVMxvHBkVhYEhaeaoqY0UvRkaWJisnUQBYEl0JUOi99CKsYZATCIX1G+R2ius/3WGjoxK3TH+i
5DINC9+pJEVWVj4i6Nq+0vtHqpA4XeiKM9fatzwf43c4K2hMHwZfddiLxy8/b4FAnAMVHKz+6EPz
h5tOVJpd/gpTUjYHX7QMxxEY668gKGrevzFznU4MxEOmO1hIr7VJ7mmXm49c+yqLjpncRCSlZSaF
zNVul/DT7EJDwUKcZdR+aFgXSluW+v78EVAmQJ4OIgqO9/AdPbnVW76atAMO2WGaw9nPahczMrke
CtMeyapOLcs4/oM/8Ye9fLa5U5ubUyZf6IVqOACkMVHGzydhjkfvKZRgFutCusdbAZHQxqLyX+7P
Q2oKAGsiq4doyMGYRGw00GCpFo2u/HMx26aeq2XetGvWWJtsjhqT0fA9dXgncJxtlOXYU/LgGusn
m40HOLS/0x99nxhZRDV8V2F4+VoRx8V0xZZ0edXvpU5BIPUKFDoQCkEjrjbZFy+s6O/fSIVWooIx
yXhQwOqezv4wuqlSVVucBye+cGPvJcmuevB8xXmW7arPrLPf9USK/2+xewoqsHPaDaK2M483F2se
pXDoJ149XNe+9/43MJ2X1PRODtr1Y2nG9+pOk4OaP8PqYKWBX4BjvTRnxfVhA1CO4pix/Nsv9fC4
7eiHyn0YTQMyxufd3C8esWXwuRpYSlR9Vxw3Gk8tjzvYgFVoGEPyKkUyvypDH6Fz+QiJF3j/zmcV
qpaiq/TxObrJpxrDJA9r9SGYjBfXPj85ZRPS2rd41/pgBxQAgLJfySLVdKWKQnleNkkfwlaX1ter
ICix/Lz+kcl1mjQDV/cpb+yz9gLdlAPmyMqM6aRwolQbI/dAKjskvwg39QOzAHhUpXjEEscbH4G3
/PRZkBtRxUD7kfCmuz/fOkUTEyfYetdibvu3TGp09IrSNmwepIy4eXlvbuQyR9o/LN3nardbtKzA
CF8mYtgdV7jSPapO+xVu5etButJnw4SSQ9X6plglQt3G6qvLWi5ILlDh+r8G87Mc8dJlf3OpkfUw
CnTQPhm3TYjXgGVPqPUDnNsiNfGbiMoXbJZYzYa9OQG8IuH5w8eqEGIb4C3syvCej9ItwILg97if
YNyiU0MZTt8gzR8gHlZMihBIya5zLOCRXHUijF0Ynu3alSBL3TQfsppRMRcZvYnk0w5CGreVGA0x
lzioEXMeChq++D/9Wj4fn6Bp9agbXp5GE73DNW7w90l+HQlFBLCvTf7Elg5eKPHdSgxBCHU/8hi8
iiw1ZxbMccsTYmZHlQ0cSkD5s+aYgULXmDtUqQGtC4aIxQ4xm/bXl3UpCwhX7hvLU5SOMb2d4SBB
aaKGtPE9NwK0saBXwY92VepJtxIxybiIRMX3GVT+uq56TECANZe7gwepgcNfOvedq7EXC+cGYgra
EESd47dLpyOvmOo1McxUxDEmfmRlLqCIS9orjyzKJlTOXdOgsho3+uSopyl/RzLd4OmegtomJnCs
CauShUBPHSr1m9SBwhZejULxWCPDlbqx6XsMt6ik53dXdvQWHdh7VCTIzO1VYgJaWRnxCksdQj2L
Xfkz8sCWAtb3V14sXa8zpOALfCz7gI3ETMI5AZnmzk20Ym88wQIWQ32bdIk17mKuFRykzHezVwZP
hvjPOP+Gaq7K5RKL8+bDxeWV/t1qu+X4zSrWxqT2XdhQG5V9yZFr+9XBuiklU2OuWDkzDRGbnO4b
jLZDqaWc8eEhRHx47zAcPgwr54bTDQmQqA0xn3pC92AOO7kPMe5rPIU/daMzEVJQXOOrC444icPS
UUpimFqwnTLT3OtUxCsVTh23k+Nc6A2BqTK5I8khZYStvIEstwxNOfjwo8O6aXBh2ZO35wfbGvlV
BeuqZOeInrkQuV6A3I98PVumELkQmXeNdgd9iS/zH2EJx5PpgdxQHGi+FCAA+fEe87VcHyzEcCWJ
YaPgpmUZfT8ejx0gMoE6fGb5CxNVu4ipHheTBAiMKSDxvmcV0r3vKv4of4+X77zlLI55w9EB35B1
rW4sypBV4WdOmQ/5M6AcwrGCxwaZOcoZ4a+vt4GriYZX83b9/X7fRCk9LFJ6AX/AhqzQskfCHBh0
emz8Qt1viLUcAei2NnetXWUDoKi++aXN/1ITYhAGUXoxz2qym5V/QYeMetwOztMNqf07rDbnKinD
BOdeEFcMJAUdpoLVQwBBGpgsD7yx79LbXfnNUc9AaNbyj+ZoN2Um2X1UMgZT5xjrNabO4y4AdrUt
FOI+BI0e7oMOfgYVA7yo5urh2XLn7tAL+l1y+c4i2t6tgh3tl967eJiS0h4YFeZ2TulbU7/sicmo
sq/eW5PlD5SvIu77LyhjGJ579VMO8M9Yw1aQFIUHoUa05NJdrcVRRHBq9EmwNoQltI8PAsqzLwzk
nIXQoCMXqIbN3HnIWulJZCsuGAmkIb+WIeyzpkYF6a1L1nJlaiL8bXBCE/MBvLp5fWG6dJli7Jz0
6ENsinwGBJNn1AA2bhZ5obMXaP67kaRwpuM4Fs1GEABnHQacUUCwig1Kb2HyF/qTz1lpUtx/2QGL
7K4gBb6+yV/mVDxXfZwHR+27r0ruES5e3qEaqYgntBOM0GIIcn2AsO5cJ3FicgEsqCnz5oux8lRa
92o3OW4Hi1vdy0Y0/PSxkAJwrfigq/NyD2nA6xFhu+0cU253H7k0P71FXod9braQWJEj0lOqKaH2
kw/IWL+D+ZgSsEk//7Yx0QU/ZOsXwS37yjO0EZCXyPvLlyf8i0lf0M2v2cOOV/k6LBx1sxGMAsiW
ToNokFp+HhAs1PxcB2lmghFHMiQPtDKlVn6FIcUXTXwdzrjOK+STJt9CYweRXsQi40dD//K+Mz7w
lY+ntdaYPIH0vNLkwd2uguTOVYN4C5uuxaNJD2t18mHtImxej9AqgGBC/p5WLfqf69TtieWENc/G
+GXRagCLQMYhtm2sXFouBTkwMwVyC/s5CLheG9flyCvcWrLNHb2YwcJjrg2sipLCd1InCYg19a+n
CTVB002b/AlFmmyAgX5toXhdJNtxIv/UuabPucAoxExP2Ei5H8U3Y6IhX//kdx2vApOOJXWX4nrp
vUudAsroFYhjBJRdVpTsP+pNaKmoy3lTy1GWsqQWBkAbK3jIxApnl83ICqbSZQxlRew7YR7IfB5L
ds+o6EOP2wu5pf9mwUw1unD5bDzw/F2mM6TmJcfsoEHziqdFDbIv3nJEW72DPNiUxdhHY1VRwPyE
4oe+eOAO6pPquPkpaLVVJi26qEgg5b8mtFgkS7YnjU0Rc1EYov1l7XURHz0SWxJDaqQ4Gu0098up
lSbtqSy+V7BNK3u8VAAqZ47HzHAnMlYHReUMyBy+V2oOn8XohpT/NVO/gIgILM4AbeTzB9bSOJYH
oebAMTEZJKPYzkU97EKIWwX5YI4TsnGN6ejPum9/sGjlgNWmdqFHDzP3iNbPBrfTlDqCI1nR/gr0
RIIcDR28KSKjf/pFn/ZKWVntdLdyNdTApIk02DeIPTanEiPJ2EAN12L8UOrQ5Epfo7a1V/6ciFrP
P7JM1XNt+gtE4kAJsbAEu5LXwLBMKMBl2RNXhs1v3KP3tst0etLaoWkjWVVaU56mLVt4KXbmpGG/
jsJfr/9QqwIRsWt0iaeqvFPQoo8Wn7P3za1Vn6yH7yYugPcfK0/GpQg34CbN+jC9UKSYWDkg+mzc
U4eriHmj6RhFefqR5QW8gFDdAWc5Lye3xM3D50hg+jS3Fbf2uTy72oGhCQD0mZsip03vgeY7Rw28
XTSQV8+P8XiY1Yvxhjo3rPB0ZBDmBpoabtLVkaCdJ/oshOjLSL3Tg2WFVyPtZo9joeUoqYZUPA0R
vUyTC+uH9yxouGkz+CTmSugc5xZrwBkB3rh7LhcO6heGqq7luQs8rsDm6keWUFRNCn3JbEmSDclh
Hifp6I+Oyo/HcYCOuqAUm+6xE5zWaQaNVDY+dXl9wXdn1lz19Xb14oXPVsX3FYx16HSA9YAtbfuo
3n2u+HJE7P2j0nA2GQbzzjmeLbpgbDk8TrjoqbrEls72OBc0CElyCpjKY72dHGEVwnJyIZg9Wm7d
DGVjVVzhluRPUGx/yqZGxKqBXwQuOEWAT41jkSxJxQUi/HU1yzesXOcPRbufSKc0rRJEM1/4e58J
dHpe8C1uLqBuOM+nXp8zci6l3W+6QaRQWm7IW+hPQFC6HKSATDOSmHPDUoFstTeTQDdteNepKCZq
+WsVXSVgEy1Jy42vI0WBOT2YfC4ZXh30xPmnfx3tApci2h1oYxIazq8YSx6meC32mfWCn6K0JAuG
11ZjZQwiibB9RrCNE/pDxmKFQfNVADfcgCOm8ttnT2FbTQVproMX7y2T9/cL1WF4Kq2Fot1J2A8b
DOys+YAljc9MBvkSi1wtwRECalD1Tted+Kjgm5BtiKIk8jFlDiWbGQjSX46tF+3FG7yfaR227C72
WREHF3PHXEOLnESpZ9jJyc5JozCeU+/Bwb0AvzLeB8GHk1C8kqWkGWN/d2EvSSjaIVD9sQX5ENgk
Icmo4Cvlg2ZT7Y6dRCcrTkPJkxknoEAW60R3uScCZRh0DltiMYvgK6ArFd06AiUwQEOcwCesND67
vEjt5sy35NqI65sDpWkjCZAuy8rDRoI+XUyCTLM9kO+ohi9ASEYReH6hwo6aLOy8aw5okqGCZm0E
pPeFtKrqSzE/9uhp6IAJaJx8bJHocCCkQQSvnIxNg4vWLUGxjCP2q5bh42+yV6Ii3B8WA3HE7KwO
U9MNEhO+Zs972f3bJOu/557pH+YlfT/sb5G1Ype9wvaFJA9LKBVM7595fKGGgiUQjQTGSCqcLmFY
1XRsqSFS4TUQbxZQ3J4DRyfJFc7u6JTtTxgpsj0GTpPI967muck0tBqHGgJxxf6jn3j+P8wUkzkE
LSVapPBZ4GfaY+u0WXtJQtXAnCiXqNuhcT4aXKHx04vccdQxXqkRSehVeM1koHQ0HqNbPuJEKyBc
973k1tr5hf/2Q5ykKj3CPVfadp9rHEdsr3uhbhYvuPKN4GemUnrjqEmxnYjb1HGf6Qn+oANkUI5G
r/bgcu1Wv8fAX8A3XNSmaiiANYl1wY5qWHRVZVyuhuewaHd9/L+OXxMzHjpCWWL1gdHLaq7KsAif
TKlqPTEPrshXVB9wUoMM2L4MSmhxdDtKrlFQsD3m70/LOxbjNdPUbU2HctjYqe9sqq6fOAt7JDJH
XM7nj430owzJtli5L09LoHUpWdvGzkaU0JdWrNm2u2E7UiJggyNo1w1c3EVbIzyo49cWTZp4UMm9
BQ63npob6fHxvm/wkCzZHM7HWp0LUylSZatvm41sKcLt3EJ7qIiRRDniakpQWlEK7MbTCpCNXTn3
eyha4KixRg0ZFyhUv6ImMKv4Z1lgwSA2E0bCfe5Tl94lpZpZqqTuOyCj35cKDF1x85O0+IArXmjV
F6urQJ7hubjfaaS9FO51a8ma18mfH45GqE9jyt2voGujnzXzJkTDnyeXB/Jzru+zirM0GYz31Eo7
DKhWTy//1fOQORFfuWnJ0UTWdbzjQ3ENk/JtRug4wECTiWVXsh6eddsTiZAhxVuN6ml7MmKKeRTa
3gg2p/oBvNAE3l0ZjDNxChiDHPr/ioAbSVLg+5DZp7Iilp1DHT//lWg60pLu5+wC8wf/X8QODgtS
PW/OZj5wItmDqI7I/bOQSkTrL7llO+xfZiVa+fCs9H6Qq30r49JTB5vL2ySgTRhuQdRrJI9b2Hji
42GBOclv7l5FEQX+z+H0mfWvfGhEud2C20s6p4KG3/JrrMDE4NOiHxe7QdzyTCPqaq0Mi7ZFVQPD
F1ZnueyUNrFwFq+aJ/8GGfEGerK0Nf8pRN7bMa0JdqcWGvLwN9iBcE+r79ALzOpxpbR1IpsPs8UX
7udQ71YjFoFuDzpp1ZZ44TNIq/mhTecqcienu8i+YB6bfYY9IIr8NrPBwRqGwl8x3qzi+KEBg+xO
VwqtPtYwLJ1TEVVxl7ZIoQOERkKJCCFtD4wvpu7kEwnFMfB1jMsy4CqcKhlODIH1Qy+Nm7WgZL8R
tB16+Q1X11Uov1qzWRH1u3DisnXQUi8bIbKIipHGgKBSX2BRuJmbS0XsGMwEbbzdihbej2EYnQNu
nfMgU6BXAuvsDeGWb+sIdB/zRhM8fvXgMWHNj1Wwi55UunJiAVj0VTxV8k7gQLLTh8ntjSXp3fgf
TskuxLrqiUtQn7d+8EQQNwyAKC3Ynag7lndJPy+tE3LbcwOOzMAVIp68FORLeq3s0yjdfrz9vH7O
fANTYnsmN7F4LZleg16mNhSTw3yHNm2snd0uPh3vmS2ragPtO52b0+1M0o7gnkqmqLGKu14x4rBC
LYOA2NrJywkF9fMuj+HxsUGP+ypYH7NSDPvynmUGWQNptUsbawil2Jv+Vpc79MTdQi68ZE4HslGB
v+2ROJ3JQ+tM47hZh0fMUaAucoqHwjybNIOnpZqm8FpQfriIlvyhh3GEixoTKHm19Up08FHEku7Q
hrmMyHMhNDJrZcq5PbSVXbAqWcL7yst2DR9OiW4EJz3090/rHSHAC4tpMOBMiXFwTB+RjvPSyn64
YxAj0RZ4YYcjO7AbnpCMm3wSK5iPWIVDxh8X0Mj+MqSk1Y44+sxhp9xkEzeQeLANVFdCMu5qMCoR
yltbodfwmxq1Sc+EyCuBsNrvVJWPnExF0JWXdMVKajpANZQjwGhruNYkM+X4HcPoYNdEDYR0fdDA
IIVGcO0HUuQ9XHGoPXtbJEE4Mg5ZRrLeDDHZssHlmzE/0AEDjNk1iUcI4RZ8oR1BVjIF5AcqyXEB
+FVRUdl2pV1sCBQv29GQNdPx9IzrmWv+vBQ/32yB4wmStmvzx2FZEiheFhtSbBeEz2bnxs5+ZK2S
Lfr0YovpZDGAIxTwXqfFkZe2NUJH9CjeXp7is1Go9oeToX+92rGKthoDCsq+YwWQqrEGowV+HNdU
/uPeE6wu94jJPoSVR9P0BjWwENg+mvhpKFw/samPguiex6YV7DFEZvRWk/nbd5bFnRs2ie3H+nTz
EIuA0VF8tfhrC97Gi4SRVRu6qlDBXmIF+zZf0YvBahzZRpEUUMrpBNiSO8YCZRk7U+Q9rdKsEEGI
DjTeKHsx6QgE2yd46kLCroKBMTmx0XeUxwcVuQUJjwOpRsmgYJNTAqPJVDBl3t6k6uu+0nb1I+AN
vWSc3KJwPHgG6NbcjFpTyjp0UL6SPDkYhltC3InDlALd+Zck3ji0hYExgTMuGaQjV9Hikw77udZB
IU89LUnAd4kyJ19/90bp2L9N1sLfum1uKuxtxuKKG7DLnzn0t8lRk6JsuNNax0pdGzaky+Wpx9ad
gxJ5OoCGS82edLgYLJYfS4Q0mLw7mLFq/YBk9Lb+sy0iAfQT3RaMbNIJ4/bfoa9A+u5qRDCJuc/5
7Mac2LjQqIlNYx2OyEDeZyGNkI0Wcd2OXMsMuvEY0eG3OZWDO2G0dDBBsK73ONlcPYOX1H7wiu82
/PjN/X45JXCLRYro0Lm5oQCM7g2Xbgt85CdDGqKJm5AC9kCWqeYtK1eJWFqYz2N2QXNM0Rh4QHO3
Y2RHFRU8kvPZkRzmJ2XRjtwzCuWGvkqdEU3m97FiJz2omHPDj3wMRJn05AxmwUFurtGHkUj5HPU2
CKauOSnIxErBOA5TRxJ/bW2CDcdmDLOXbPqTeO81Lw0KCrmc5yGpYThL017+KzU0osJgBOVPPLie
wKMCczFb/JNDXa9f6boZLnFsDwif5NeZvelaNaizgkvG+Qtw+gccDXagn+2qPTrQfEzPgnl10lW2
4sSg5/e6XegQYyujr8mPsqP3+LiuV4ReHOhzT84v1hRVfkDMpJCk2e3fz9nKkIl3jBjF7iUwS5zH
/xVm5Os7SetKD308IunxVtuw2geajV4n6qTIj7+U8oVBE23gCBGS+tfA5JbL6VeFdpwz6dt1YjsP
M0IQHCCFLqits0ff9xVtmJfjjPIDuU/9Xqwi5m3WGEehdC1IPeHWX/QoOjP5jB/Ald/zcGSwdV0q
M+D8+fZY7QFTi+m+XPyIEGcaGjcDbPcSpN481gsNP+on3x4oP0/I7Fu82Jq67UPIr33NStY103UY
6TJ4iRmUECC+XYyLlJfHktDGk1VJSoTKhMr6dBEvHGv+exvBRHanNAMyVS9cH7ZwN1dmfZTG1kpH
S1kF47ctT2tZi1BAnxLLX0D73UI75bxLHBJgdcHxhkClqWq9IN1J0FsqWyePTTgOMWrokKewhjbC
jAki++pFmfDyjXY04TlIAx6glgzskN4Vk2QmcttSgHEFlNRwnx91n0hWMwY/uYrxIPBtR/cadtva
Pmhd/Gcp8HSpEIg1LbZkTdtfyzCxxqwUKzS3r7tuyvotzCP8m//OFIdke2oF/3hPgUitAHPT0com
yamFd4Ix28AZmUTFcMohEjQT/PGRtwRekA2KAq2r4BrxA79tuo4+4t5TB904tBV3YgmHpqCceq20
/Lz5U61XnJ2O/2IVbVy1R8ODSiR5NypFPrN9vqQBJek0OL0KL0309xX0MhH7NUUo0oa/sRbdHiO9
XVl63tXJmyytwOzsf3dq3JhgAPz0YXd7Lp0MWo7nSf7dg9FLEu6t8y4BJZ8KVBYI8801vtKoR+Zg
olLRLRxDYPW43l2zEa7AeyKYcwL2nL1XwqpAJKHB4mqQ/m3ntdrYZ9Hyhv95AAV1L9g1PBZGtmM2
HFBXlEhLa9Ei3Jm9SlFjh8m0VtwxIvcLkd9u8UXwSW7f9ZpM0qVCcD649ORYtJ1xAkKcsos8gvIF
hL0qi/cKx1Hy0RCZbYl5oitS8YztDbNmP/joPZkFLSOzQxNyPxSFcBWqicIjvigkzDpS2DFfIvxl
7H4d6djf72gA3JAs2YkI1q6owg13IJsT1bYzUQ/c3UbTykCem+aihrsVYcZzt8D+9wsV39krNGLE
RmOfzfsv8tx01S6+liP8nFXnfUGAyCdePBdvwTBxxTcHi2av6xgxrrZaPZMrFXp2HI1MZAN3p6p1
uYhUUQVb4V+7zI0jcS6wTCWY/MLGI8mNYO2ljVFm+gEw69Ji244w1BbuG7S0h0UI9YRb0AzGuMf1
Thg0fBBLESglMFwlhXOc9lzLNEIwmAovOWUQTvx7AoZGDLlKD5wZQrTFQRBNqpBc9BPOmjrtqKyw
Y/C+ia75dWi3HPuQ4fnta+T+g7iDsqgXUSNA7n2J1G7YKH/t0aJ6sPRk0v/VE7+3G1xydm0YRZvx
pTXbCxLAB2OyvZdIbzm6YoRFnxOoGjqV7FvuWjS8+Y4DygSWdm15JVC2tTFgk88+3LT/LzQKbdvd
t0jhGn8RinA3vxi4vJktzSSfMo2qdMutyMRw7Y3FmpQ0dHzO7IV7TZSyptojY5wGk/PFhFPA3c/o
WwIt40kNrmC+eYLqRdqkWSnI1nZjnzGB7XTTrbFX79VbXdKhlIZ1pGDqG6hXBsWWTJZGIECRU/m+
iufXfPl8qzJolxxpfGbwtmyWQuJQZKgp+exfiOWelouTGyuPA2FdMfqRxONks8mYYJ/yqjOC5BfX
UndNNassIv9KwH/aBYVq2Od6oAgysH39tX5/MQGsPBtc7dya2uq3f1UOAO87Pjd/CbOalTYWi2Sy
d/Md56b0/nTkBBreKkelMbl0zpntGRMN5iJWADXDt5mCTK3afl/EGYRkDFrBrYFcpoWsYJaPDfxc
DvoYNghGQMH4zqqd0sam2xsUbA2VJhQLH6XGGGpGuWNpGfuHFAQ221ieFD/nnnC8iacq/5lR46pA
rxpoBH1YSmbXQj5bIF5bgkxRrwdXbHaOSSuC0jTNdHQrXWSvAbySkG8rOvcrBpaZ+WCoG5kBK0/+
NHvob5ysG4SAPIKTsWp4kDuKoWOwxQsgPPneDaQpAdLtHLFwFzhtgYErLdYNc+0yu8rimDXDgkMC
CNxNd5D3atp9nfV5CxbcJXgZbXqHWobiSbHIS/WtPlOdmsAHFHbYHUu7rgJmvi3ZNYwlMtYf+rjc
FPvp0mw4KjuO+8TCKeFg0cB6ZJQiCmo3MtV/SvihcBt4zjjpOdsG/hCkpix/6sRt8rMC/ZzNNsy2
+8PY4uKSCE/FY4YquNBbjZCxzJwOHH79fQAJQ3T0mVu6sEb16PHhKdPKz2s2Ntv3GBGTQmLOWe1a
sEEKXHpWjz283yfla/5HwigSGx8CXOtDz5EQEJqcmYf3EfmaDCDdl0S9YVVfMT/WdwbAvDxrr4WF
qmzvt47EieOGQ/C+k0FDUD8C/mra9a1Y7/Ch+sG6pjGEQTf4OpyqYuL6tNTVB7tVLVj0uRzLxNbb
waQdiOvQ8uXdZBfwE8ZbutlErzvceWWNT8ivpKharzP4TrEKkjSxdq7VRaL++/KYxGQBlupj/eDY
VoUQ0Oq/JTRd4+CDRoARnCruwnlBmPT1e1tzzaS/jrJPJ5vForb5K/B+doUYhMV8py5xAwKCaUB1
Ti84nQMkAlKssrCLGzlq3Qbli8PxG84L+aXyOqF/R5y/LMd6aqj2oQn51b7U8csYoEgEPNsmwIFJ
B0M3sD787dcZoNQZZIpwxitfr+e4kB89K3p/Om8p1mM2wdao6nvnziq/VMuS+wMR3CweqI2FQyeN
MAQVEYQYZTHjDkqVJ7OLjDPdE8nbp5vDVYt8B5xlvaNwY1RNdDG1LrvREt5pfU0SQdaxdyU4Unay
zf3Z38xDw6b1YvtMrg8+BOKBsltADPIaVyoYYxo8QhBowE6Lx0rnSwmPeApwB2c7CuVPok989Ovz
BHEXyJkpwv9fvyko+i++8jcxD+B3ZlIYDGD/qunhFERjZelpSOsXZVbKktOVTmxEIzcuTlT3q1Gf
t0rQmEGZUjDE1ub7s5+urXowMbjHP/Kg/ERMp86GoR1MVyfQWGmp6qwOecuDrb1vGM3LmT2qZZpg
ioCnfcau+CsTsKQNFZe2/+1nSNeuFhYd4+CkFZdN7QLvGcISXUsTDoopB0HXohMZi9cRu0H6c5yF
Q9Hdoi8SXS6nKhUFSWO/N1SsSEqNCNhSruNA1Thys8xja4Kdcy7Zw3VoHFkPHDEP61twwVj2/gBc
8sfP1L/LebMxlWzs+13EFFap0UYYmsocZMdZKSkVkqpf5GXvuQywIyOkvpowExkx4hdPSRzDwqdC
C5qfQOkGU5D7Z71SJeJWZ97nehrS5eKn3npsCbimTG96UAcsZq6MlO/CAg9lnalp91PzKErkkroJ
0j7iFre2rEN2eYAWx7V5HC0SBeYqbmd10EG4wzeHeikgeG6R+n5/t5NIAICQuGky24XSVkiNo7Pb
7wpS8Qf56C3uIZuFoeIBTx03goPcUvVruokQ87fknrINyVRCSkNFlWqbvVziOuQmIhXhe5ZB3HK4
Qn1WZkZSY7RNSWGd5pal0L8rs8EGLQa/ycMi9gj6vfR71BGscmefnRMSnBjqdWomqBgqg4Y+NjXb
WT9wSaXTkUfwdGNkygH0rwTnbeA0onJqGnRUW6NlqYqhDFwWTnHKoNhbDMuZLt5EY5heRWNhcTaJ
PtYZ+evLm873NwJ7qi29VdNEaBSkTaGxwoM9WM/VO5uf2GRoJhkTnJMNxW+v3WUNV1Ts8zYbdq6V
z6RmT1Wg8JL9bUeLl8pB8cC2Mc9YehsZmTTtkAKsPZvADig9qr8xjS2nh+E3UW9fuAKJDA7Lfupx
6sIjlIka4AUtF1AoDrSgqpFY1S463u7kdGZaC3epF+p34Aj9T32nDtp+YqajTLfgo6MeajkYwQz8
JpU9B0I3wYyrc0rlxNaGDwlJCBg3uejCSgq/es4Cx1tW3LQh64EbYtTu6na+vPzALB+SoLAJxDS+
+8xNgIuASH8bailGk5a5UsDsddW0Ypmr0pN0zzdqnVZtJkG98Dag07Aoh6PKyRQTJ3YnEk4rD3iV
UvAvwDcgfbC1rLXLReXS5WIbJAIKHI5UuD+euD/d8gua+RaeFTO0jOeOqjeUiz/E6y0qjlHiVUTX
NCZISUt3Bhs2M28TXeDLz08gTOyR+iT8l6OTbfK6TVDYZPzv2F6I9POHo2L9bU+TtVqyE3MX7xzh
jpzoSXnLpzLd8eaUNeuMmFIPwYENcsO1dWdeGDlCH0dRjZKBhhg2pvpcxa2OfK2A9+Lfpldy9vPU
nU14iiv/rNqhWxBOOUrsWn8P+jSCeg2PjP9exqERMhJLByOR6OU23Y3hvXkKhA1EwqE6qlM9KRK1
3s2P4kql8KpVG4upuZhxd7gyO7HYhXoSdB0sAKFYFDWpXNFNYi0l/XLHHzVNj6w1W/JdTO/DyJfF
o3FMDx1T85C0zMIEHceO0oq1kCoGg16djTkf1isEAK93Qb/WthU0AHFZpLijGxZ8jC22izgpGbdR
+NdzLztDqa02UEcx9YfKNmDJDOqNA0YnOoW9KsoevHKtNy/jdsCXIEWCpOOWATlU3ZRkVG4YtLqf
5/I4sZf1SQL24kxE1mvvRKFzNnOEoytd+d74lIDGLDv79UpoujSuFjvj0Kcw161vQuUqQ1pYgPFc
k0BKNQlvWz9v+BndfwvVHFzPnFqijJU88ZDz4qJE9jn0h7Xc1Qj+d4x/o2XwXS4HlS6mlPT7Fo9d
7+f//BczDJAQotNRMR99We/B1fHZglHp0kwm02z6BNa9CfM5i7jevYqLBRfme5aUZzBvzzzDzYp6
LFDDXJ4slAfr59dqvumY8ECNYF5t2O1y9R9CQbrHeiihQS339XL8TcI7Ng/40XDfrIjTTm03nCVg
RFxGCW9NGFWsctDx8CH/zcuYCST7+LT5o4D1aPUj13jKodtD7DA8j0T5Udl7/jH31qVJMApavdDI
rHGVDNkPteiegfgE7ChO+SBkhYIrw7eVIdKouAixtT2MADS9WbF/TC8VQCl03XQSllgjm9YQeJ70
+ERb0CWercavOyTURMMB7fI4yk/1MxX2wRowGxO7B4CzJjS5hG7XGQGgv/VfeA2Vcw7Eia2K6NjS
9FL1hePREWxJlngiXhyQic6+v1XEEyjklIdqLiDhd2m/y1BTjG3+9XNrkfvUboCmNA6csVZcaEpw
JsTdIQ3zNBnsWAy1dKZGdtnGwWE6UyA7RIjNWs+wlyAeAWd/OQAU5N91lL7TDOp9XYcP78tDkdvp
3i/pUFs2oFm3SpdMGaUzSM+ZFxUVjnB2QqHOYFtp+EBqMYyWm4ZCnjx82xl9Xm2fcyjJvge7KusB
zefsFhKPOJKIToyu983n9pfpnjHIBADpKkf46gscAWMxTiHCDVYuHTDeRL40lCZe6ICYH08JZsV/
3daUCZ4/wtm9JY5Qu5luQIwWqc150jbbbquVNjza8Yl67VFD6HxK4AFYBKpuADTO1MBvqaXoIxHb
HIEMf0w5vgoigp6Q8MWyRIC1241N6hAFHFBd8QtZFXvASccOtiBeHRGsX+5+suwfC8raGazSZaUd
C1Wyh0faANp4pWjbybOjqvbX3EAjouZ3qz4RCLBUkNwOtzOaG695kJviqeXVm4BWEqBE8+RXZh1h
zplu8a6GwTUdGR5TrXPIsB9/xHYoOAWmauXi+FYFsxe2QArbS6/G/JPlaupWQ84xj8LFmPjc7LLT
CHTxB+N6l2hWmVL6A+i82AxeczXB/p9PAj6dKnEJyvDM354bYf+O9CNkdTg8aO2gpoe/qeJ8q/bg
DwbwHog9mJMp/nXGBYyq1vK0lqphUASaZHQ7ldFB7vULFwTPKiKiIbYB/C/oRo6cUBpglId9LDoN
WLlEIIh7M8XUGAmFlw8nKmLqzYNMnP6L71rhBMqlStlBO9g8EP8tWWM9tF+e3mqy57SgBqxVLbxB
RZ7+Cr8yob1qIzQqrufv+DBhFFrDL5FwvCWjDMd2HP1PzputvFdktorMd4cdbtfY+GnYg/D+ypgk
PojT5CDwvL+7GyOnOxGDUVpSh5jAjNoOxz/XqUh/0OVVWiWiO1iPlchhNQb4JuUWZrimTQWR26vZ
z+2QwGwf46DdUbj93N7mNeUgy4zw5/dJgxGBHVxDNkcKHtoP6lJnbJ9kiSHyUs1M1YC9NjwEsD+A
99GgO6yI40QflyCkljZu0PFwaHWhjCRQf4Y2Puj4eVMYt9omZbe/algqFPcAtG7OpokItDmIMpQA
yBghaZeefUGLjXMkLq/vdV9urvZXc6MmEAmu/v5QM0EjpSL2EucgkT0NjRSmklBhw0RScnuEcOm4
qhlQ1LOn9sHuVKV/dfDaKTOBZ6cXjm8NqjgnIBeKKKm7In5Au/BpzrgEGkqoZo0w2B3l7iqS/+da
9ekZZhiKuYxyndlwzDjrV2ijQATxJGJ78o0bGN4AndQDOyIu1WTt8xk7SgqwQKg19eOAMzs2CBLs
J0Rhph7ZoenqptSUWrUCfjlNgs37oSxsLKQXqCuC2211PLMti5Dkz3QQQolL76RzDMihM+P5UvEY
ufAJZqQvmB4xX85CaV7Pjt+fEUlrObAAC79BBl07iksUUU67Jj9PhROBzJNEOHjuhklWtTGw7Orf
FFbBuWOlmkcHR0dnqR8hrek18FLUr5kfLePQWTShK2G7pkKMqmuKB6axjZgfL9Wv+SklzQ+oa4KA
lJujXm295UhgrgnkRQ8lzNAZhCHlg3lCu3TiKeelKwctxyeY7Vu2w3Y+wPRAvtWOi7TLqXllAJd7
9QI+SoRlRu9q4pp42553McRc2iFC1WlS4Y7LyMhdnsABKawO8gwMyj3kA+uU3+Y7JigiVDmagbX6
tyBGphR4wUtGwj6gf/yNsk0Pg0Pxb3+lE3vI1LWAxiCSuEMl+uirEqurtADijRBixfSjvfvqCkVp
he/k8R+Znzcvgy2++yvZO0pQ54XRZcrCuwRKX3IsZPUT4/DKYTRYiKUWH8weiuUHyd0o+yWk/M7Z
KkEc2kQyMMFNrR+KeBf3YaJkuSzAI8f4aKh8DkwbEE6/woKepLB3UJNMpBNpG/99HFPq8ru0STOh
BjDTfH9AXrh8dJ1YadjIp4kkenesDqPr8Os6LZ3QECoKlKuwbosE6/NOEvvF+2KNsoGnVzkaOx2v
rp7f2vID9XXT1rKFezcfWAGMX+9dRtj4GR22RSz3/5+MKo1cpIhABOM9XB3nTymlaYsaHzF5h1iL
MOVhAR2dp8XLxqCs20tSzAfi2e2eGUcOw7ZeqEjPF5L+zMlsiGlIi3zQUHYLHjnyNEeP5c13jqrs
OOzGKk8euNlyIk5wXIpTYZxNEXiHYELegLUrrg2EaQel7odkuzGv73+KS7CFGaIpLeK+C14qi+5e
GrzAmQTldL94zDygVO84QlcLpiVs1BKJcH41PvZjTmLF0BdkDAyh4RSkEiTKGgdOEdXgHBaeCh6T
JRWDbw5UVeiOEzSzRyvu6AUfL9ZSnwDN0/FWE6S0Fk/1FHwC1XjuFUEQcyN/MtbDYqtCoDW+n/h0
iq7otdxehRDbkj0xJKoolFz5LocisZa0DYCeuwXPDEDEl66PfUH1Ic8Cmadple8o2O2StvRU4Wbq
C1ZMfQRw83SxZuLG+pxGJrAVjGNq+jm1JZVcJO63msxTbFaoomVexXoAimsKI2Rhpr+f5SnUzNPO
OmYOhigQz/gYIEg8rkb1j8XVChgoZ4jD4Dn+J/64aQcYlYUTaFw8Rp/Qa0fmI/oenp9DHiY/7FaL
lYiLN5Cr5aaYYPKa2h7kAGE2cKa7ga0MEHJzdYU1axjuaE1AUFRTqH9S66Hu1MyVABZu574MgqZQ
zG6HOSoNG/VZ1+8xWuNkb/kNd/5/BXWwXy1tVCZKAVKWITTTw1vk2+zooKBqHMgba0mGEprkQx2u
kjVancseWjVuCfUxQsNly6FytI6Q2GMRe6num99aX02kayT3Fo13LBrkQzhXn9UHoB0D5H67AJkS
e7IbAPwjS9ZEQowSbnHTG5jnj9dgL8vt91y1R7UaGh9vzQH/4vcNI5ZP9yw53Poxurr9RiKc0dGw
243vFDqdIuh7cEVBmOFZGi/EsHsOAOto1zE2bYHWCY39bmi9TjpXXjwPDIwU6EcmrpOo68RskQp4
m4sKvJVwDITyQ7m78ubT/2Q99RPrNvyJh6Gq4gfZ6e8yjFBMK3pgXMc5R5tj/nnB9PaS4fJQfR/N
i/G303dooHaRJXx1ZI9ryUfOhzFS5YKOHUzpPdkwCBwRRcb1XlJkMD8loekuEv7MKydSX5hE3q0y
S8ZfHzBaEUI9eXto1/MwSmL+QootWwSSi/1gARWvU+zbr7sbiS4K/lhw5IE/Z2jSv98LaP05/sNP
tIjO6AJEQyIZXQZUActGA0TDZWwVA4lAyENl6JcZT3KzKplwqwFawF5lLifguhj99UEeGIeZUd3s
fXW/jkU4YJn8oy8ycO9DSQXDfCFbpzKUSq9xTpi1GHkfnOUAKrVYeiIK0qJKVbL8XVFc87IMZQM5
WjtHjXWKTKOsh8pLiJnCIcTZZyBDOdICl5CtUad2TXfh3KbDVwnAo9tcxB9hy168OBMeiGvUHAjJ
4cJ4FM46qDr6UeQ0E/uw4lbs+tvE35buc06CNj/jqLBfHmWT8CWjw9jkB6Q7Usb5s4cfF1q9Rs0K
jrBUBHWFQBCAAx1poAUYStdqTnCMZevreBkGdVVQwnc71JDbf7IMMvqI7wF03UrINag798b3/VBN
6h9X7SYtHDuD4ULvl12QxguGhzuK5e78QxVD8Ka8FQWD7HaAbsRqRYa0NNMBGoK19/x+rbl5P4bN
+Bvf+Amuovjv+IGdalZIMA5TIbKRHXB+Xugg+w4a9gOfDf75lc8jaCHrHj1HVOCeSLOJMvfQwD5P
J/i4y7jexvHM6e+T/xCJ3DjdkbUAeFcMB7hn+z9Mt8zgLt547T2ex5pQMmvChwMHrmhG6pZpDd3c
XxdxQVPd15BCq2+DL6/EPOj3bdkOGkzFymuMfRHt7P7nsXWIhSmCzwa1kPd8AZ0z3P0JBJK4I5eF
c54FGibWHt5jix+gzX5t0SfFGHXASw8HHqm3ODwU7sJz5zvaGbaXHNFb95LwQmmY5Hv4uOEwVFlO
peug71IKCARE8MrkLp2bQXHYtepEqUS6zrv6GsTPABytWb0HHCzd+/fmMt4uTCNZJ8aKmbt6fBsz
jppE+p85QUw7AmvH3lR3ue5yluuJuB/O0ehIZLB7qThlsZRIVPUTlJnxXQkAm8inZvRsR0lizV6e
eEbv47SehtI+03xQAEVlrXdAO8WN6b6BSw4Kp5qHEWvnQNC6Df4YvX4Z7Fsu4mU4+/y58PLSfa00
kxxk6kFRueDrFWhg7itSO7qqgA5JQg4lt0cRwv5VP7EersZgd74StZD3YYlMzmWozktaSFO14+A+
N1Ky0ULHZBfi9bJIMeGGeRFEnR0a80WNls2N/1uq6VaOkOeIYT5z6m3hRXqdXR6Ok12yEt5B2EA9
FbDrSvLvYOgG5zaQV9G0mWsQ3yP5wVJOie397H7/M0ve5gW4xxcxkSoByA6KCB1ApjU/g0TPC2jF
g6OvkVNvmWC5IC78KOwaRPOkHnv00MBmp5uly84WuUATeBMjzd3EjQyczWTKwPNzr1JI3QqwBTf8
/xi2UZT48MqGphyXwDtCgYQLXPEcrrA/bcTDvzS6yvt3Qr6adlNUbGtGr0k+zwtAdnb4Q1JBCOhN
A9bfduV2VTXg3s3UhlwE0gIgKwwZJClYzcq2hY4O2osyyr44jNDSq4H3gX1VbYxEBvaJOda+JObw
yijV91SAZGgny0XPBh2Vd3M/zgnT8n4JyZsoa1yDRRRC7+dacPc3SHPX91S5IBZX1Q+STWYPdPRG
5in5ylzhyO46pRKbY6FJP4kLO7HTpUgBdM5m0zZTnYAONvgqp3i6LYnewRCelfFtSUlSgPNfCssm
6uiBZUwcTXscMz61pHgZlheF4eNkJBZ95ZwsPL3+uq5qJJUsOJ/w61GsjzO0IqYQUCozdpxl+B+9
tbKaNeXyhsJrIUjWh1gqXpWY8ppsY2qVZTk4doY6s5LrcVH/CLv5uk2O22q0Pby3vDshB66e4HU6
o2gzOXxToRNj7EgSLmX//HCHMnQ5A3yTLN0QxcpdueT+p1PVHJw2FJzkj8FEE3lvBOn7rnQ4SB0r
DTantNM+tnc7BxB/pB7MTLSv5d+SefSJFTAjELPL/gYMIfuzadLgMqLGcxZ+dU/G3VR/njnKasXQ
Uiqeb6eU5DeC7H9zexX7zqIS0uAcuWr4r7maM1bvIURMJXkiohLA0dfggDOesD2anzzAUl2CPllb
mLbM4SdB9GkmaaU2J8dLL2LGSFY+4DYOEhSkb7j82tmUz5c6UxBx/426SsAd3A+FtZvIXUfUVIM3
QKE6RNpPFkJPLuPCjd/cJ8TKd56jTowpB42zu/Bi+8pA+tYfMggjO9rMoU0IGvCiwCppmfwFgRH9
uqwxBRDOKcrJyy01QbrluB22IFap7SNtuRO8hLa5LVAHeZs1/GsAH4axFiDl5yHeCof6+2dPQVBR
Q3noPsbifNBOOjXVPhuQbsZHPFkK3HahffUbU4f+Zvlgb6mdiWtxU65CmXJ+pudK9sPoJPX98RdC
Y0rzcLbuS4/u7kffBozv820G+j8LHkbHDYLXqztPdO0vH514pHbQh1YGInCt43hfvYLeTJL1vYYO
4xta1JQqu4KPnUylQagjO7GA940rNiO7XCRVm93sVxS1+T0M27SRfdA8x/qfQbFDg9jpXDB6Tjub
kPo7h8Sc8B9sAloQ824u2SFVJuLHx2aYrsHwFHayE21y52+yYEt4cWQ12Vi4P9nEIKWVvCkvibEJ
gdUnZKiXERSw7sV9LqWSmWnxv7EYWdMhtSoVHfSNirkGlocPXZ1MV/LvNF27ua+vUrVFvt2SdN+R
BcXGCX4UBtlmT1dGkeucvFYwECWjhpUlvFjjwnlfP2hezs6ykBegEbhp49EFvdvGXQoii5TpKPl8
SHa8P2ymjJbR51a8erP8vPgS73qDYFRAzfF5hz7LgmmwMJmslJanXy8VKvHWQCQkJevpECggr1uT
PXTntek0cnJJ6BkHTVP4k4J2YnBRsP3vXJQRI4kHLGcg6SS9JwgPyjbryJYTqbuHChZ1g/ehhgYZ
C+gfiRrIEmkvtGcc/8L3NStiJ1a6A6HwFUKQIoXa30swF5XFvhdjWoEY+KiBMdRgiOXh8twYbLoq
WQ8c8ghx7obk9twTG1I/Uav3+RwmpGYDQ+pQafz1ud83tV/w3mxS3vxOB8qwhQ6miTLTWw5JV0Ru
Mxew97OLcxkCfKKf2uvZgeCTdyJmTx9rJf8G083uB9Mf/1VE3q4iXs4JLr/GANYAVhpD8W10aW4v
x4FDnjNUwTv5Az88C4nb/cLAWV8nt5vQ6O9HlfaPkXAvsKZsKguMy2OjlHjldWlHbwhrEmW5VVGS
uPoRnIIQtZVlKcJ4kWUrFooUWS+Lhd0u+mP2cNQr1GihZhPkFpn/IOYo75rR5Sj5C2r0Q2wixyq/
1SCKi5LGiB8v4kUvHaMLa8gz19myrZjWarjdTqq5KklVl+Mle/rAq/DnNukEtTHFE1KzZxj5TSG6
slHjeakaiKtjgVS227TifbpFZPOAgLj/PYt3AU+aK+xUtWuHSrY2fEqv9UhJp19xTO+hCBLT4eNI
DTQemmF08FDgK+xVhgdxj6zS6nP7wECKHbn+14R6p5iko0S+V7Gt6IXQ2xZKt6yxyq3z89LuhfNd
3N7UFfRo41890q6y4CNlkkaGq+FqvQvHL0GWg9WxlrJI7NBTObjijOSmGvREU1ts8L3293QEeshO
iEpcc6vv9Eu15IlHzvF8hRYupAF9KNThFnZdo/1p2b0bi5guEv00soHT3iuafSeNiuBHV6H5ICZ3
Z0xw2sEVcaF/cwPbw0HmCU6BRAkwMuKuW9ilzmMMNin/Ut+vmDwpQqPFLepZl5nTk4liWPlQq7Ae
KhQHbGqZ8lLfi8PEc8UvDIcTvyM1s7ypW00SJYSJkpRPs8MextJsegGvRGogEgX8d7VQ52Vt7Ku/
vsVM04D3y4nlEHWK4oji9k0+WLZlm6nOodpW3FxEWGZPnwXwq/mIjDTIL1BQgnVwY/aMHIU2wQX6
3X5FPxDxM/x4hCblg1WH/ho2VpCL0AQabph3805SLtV4f60//vScIYikd6TW8CrossSGUIJLvMPx
vq8qWyS6iu0/zqnzRVb+YD65V4xwPeFiRQlHTNt+jGfrZ5uilc1dVIDC5HtvwJCr5jmznpPo04D1
5JUZ3qiGlgw/BnvznzBCzj2FUM7tZTThlrgdLnuHKRIApxgSa+A5FCwr4i5p1kAHzYKVBBIw7RtK
Bj2+y0XwMdETeESnUTxxlpop0MEvzcRRvy6YQgVf+3kNd0koWHSa8cHA12kt9qZbgVp3PxrwlMCv
1w9MeVC2SQs+PDOC9POIEOHBZwT/0ZZ71uoiK6EYBHEJg4qfR7EvMIbSiJyiU2sLvKJAGB3kk8Pp
b3ke3jhNoXKtdKjC4syJ8Aoh8DmprGXRel8sYA8K/Q54GyKPwzzRO4Fm2gcbOksvzFIXIHalnJVl
n+Jl5dBispdexUoDSoob/+I+S/XqLkdj2S9DN7C9sP99jNYh4OSqNx7hMTSRKexT+aLfCPZ7/uGx
JhmKD6Z75wY3WQZx5MrC0coUqyyOLNhLjfQUlPtwACzGfN1fJz5FI3GwJk61RwNb1vTqADgFCnO/
Oqo7kSh3qF+a/l3g/iCEt4+89KEFSVDQxWNJLSQLfxsjbX26JMvie4yE/Vech1Jr7ZtOHz2ixbIf
fg3GUgFiEwvejQMNzd3SFrNnpSzp7UDBCrb9GbQPupLbUUaO7dElbCqX3jUz+cEsxMq3T/YnQW2I
sNvs2vhi67LUkOInUnHkCDStKZdSVsgezzv4Ldnc6b4oVyozj77txfv70AqJVLkpoY8tIeuvsR4X
JHT+6EzMxnOg8wONUrz2CVmnvpOxyVN42KRTm1zL31fY2glP0I3q7HDT8kPczNeWynp1/5ZFVPy8
URmZ0A/PHVgaggwd6fdvcyvj40b2HH+DrWA76Jjb8th9Y3MZ7zelgAxvk96vC8NolQageVNGLLlM
v4tSoWk9Qvde6EQGBcXQy3W69UjGRYN9XWHBdQtrvHl93ZJWbilbNQei4O7mtZmLYmm9GUtedOYf
T2hkgi6vNUlVhFQluL8qUJGUQERK5VOqXS3kZRkG9ZZyEtu4TAx+vpf6yJohkx0+xQlWwv3f+fhP
0VYw0F6z8grkXcKEiE9CmdYWpxz4i9hClNV5S09x/e7GxtirXI0UQND6mSTV+H7mbtOWO/l2L95P
duaYWFCKQgKR+zvdB4+Y1a9i3/VESl1M5Ky6aSjA+8dgH9/dQhr5YO9gl+tigQAVdr47zyK6x6y+
KiTiHL6jaWHwO6/MVScS7VnXjLOF7xXAc4z0rYsN61mJi+ZbGycCN/KvhcyfCFzBTfm1zM9YGOqo
2k3/f8P+JxW4X1YASTU8pjQ8jQpqXdbOmzoKOau4q8JKBy1b75XoEeCcU8F7GHnX0TklzP/s3wse
a8bYOywIAOklBTGoLX4vOr8MuTQkNCGNyuHyJAA74mmWxQEPKfHczoaFYsM7WtYgjSkEh4sO1szR
CDVEhKP5SkhpsVEEvpCo9rX0DtXZMyKGiId7R9VTZ9TfEa2ibabpbz3QWzw9ZWcrJIlHVvbeFSMB
esmQcbtDZbPb0P0o2fPLcCYVASkpUdma+dnQ7I92QK1eUky57gR9jVhXZA2rBO97rpurOwm8Heq+
AkbSUF58rmTZ6hMy5nPB6Dlt1KpCcrrcQC8KEJ7Q+4mTpXTu0pKsiSMW5VKpContJVrQAN1Tst+h
oFX8aNs58YKZp/Se8KuQx7PsUkhYf6IPky/mjvS+aE/isBGIdLcdWE2uErJ9kEZAXoEq4YISqaZY
Qqi3ccfavYxgctL0GmlzefB3U5S8YaJ7fcB3YDxwpjag3I/Iw98cyfO5J6+wrkZjRI70MBtr0IT0
QSu3HQgFymDuFCZ/q7vN/MBPunoaKfw/Iqfj9Z25dJ1ECR2x46qDlgtAA2Uk8SOuL+CILlGKjs7v
x/BDxI1einuS1yOxqkI7rAtSIhOwByYWk7Qlf3msuDg/BUusGahQl42jSmpSZ6833/8z24Fb6nIa
P2JFRGeOqY6YZnRaJ7PPAYYo9rti5SRI3xy1qOevITL+Ym0kI/pb7i6cyklnfnMOv3w04a0LhQOS
bUMTTh/Kv+yZe3ElM0VnZbDV7t4xEuxtz6vo5havczyEPQMBzeETsmUb5Nnn4aaF2cXd69IGFALy
3lE9N+B18L3XXblOxI8fy3Pm3AbBAi86TsdTMRspjwv7mTmDklajzixh50m47LcJ7SjdwiLUhyNk
je2GH0ioCvCF6UtL5ACCrhiwU1arT4B4W5oGdZsLmHF5QEk9KvNekx9NOEa7L5WDcuXS5nes1x2Y
mr5E7zUu8YwbbWmjRbVdVMRmGix9Lm+PekPgwOZvDD2o+tnj3v9GRkFn3slvPc2R+qeraWOI1qTS
ZhxK7OqwbvLxdBJ8lTloRpTkQeHm7XSUVEpl4xkcJZtSgMSgeBHqVyf5Elb62MT7KJTxCHGJFp1i
7duLum5/2BRcCLsq5YMNphkoI5rvxNge0dDGedmHGhbNbkEqotrUJEBSbIdBPKjTuKGWlG4ngxIw
qr+mwvc91Fzh78CycJ4QevHN4SPHVh5H+3FarrszNNSZ6TzKaV8F3u924ynwKAghxsgoGpOJpkib
/2z1Frxi3jPvTHGTohA5ZJkDQjGrbjQVUhtysGMbp0C0eFavcG7nSxo3i3ZwvY3f3JPCONHQH2FV
d9E6bJS7pqLFYrv7yAXgCl+qtM9YOtRRBsdgd40C4TXtzjiEptgVgouPIb4N6qmE7h61Ama5oBAz
u2yMhdZigQ8711joReQxkp7y9Z1dlGX800uG45Hd09UuBOcWcHucefNKhCHFxhpXGFrO7i3jrwZc
CmN0V+VumtBPBN5dcQm6QHpPicCdxbry45qEkE83/RK2dGskrz5xbSKpYZ3mdrk17DMyKsU/I5Zg
5tdi/tEaQbWRT5XdbSzdU180N7YAIfS4uDheE5yeVyASi1Dapg89Y+JkvkPQoxtsHo/D/4if/EKI
yxV+C4dZx8dUzdwxae4r1ly7vYMJ7qV1/yl7EHXcVSCUoQY/XTYAs+Rtw6WK3tgKYxmhVN989dI/
rINQu1zSwNVtXZOmd43grwrvAw+HgEEsruYYfmoCo7B0o5/wbd0w/Hv3nqFdO3ju8o8+svQ/D9j1
Pnok6K4IGWqbg1atVWIaJcEeHowhFqkAaKf6NrEROmf20Q+q/C/mBUVy1f3Bp3/vVGhke0I05Gtc
CeqwSIw++RU+PCX7/vvRWbY8Bi/16tRWmYoYUqICwnQ4IlMDke3B0tibLt8IDhISbWkv3EtG9EEu
StCOW3cFZxdoyaKIuzNRAbFlFliKn9yR5+1NFs5AVOccN2ojIKoxMkHxKc89/xCHYuXZRYTVmj/H
ZHfXXTC2H1ZtJOyW9HfWkvTCPcJ7UYsx+ZsJwbImHjx5Dr6YYOlHZIO5JgHe5tQ2l1lJYckSq5ek
oFbC9FpLeLP4k9uuqridQpleaqkKslFeBCE8bYJuKWiHmiFnzOjpWRChY9M1Yx2ULs8lEIunCn+G
xs+b6KUxHdFvLz1Dr5XEFG1WfvJnG5Rqs28++MHrP0OQ0AHInOq8jmphsjenqRe0xgNhbb5Nkc1o
jgT6cYlGM5wiYqg6uCf99enB1kS1HJmH5uJ5QnVZxJVYimUxIx+U3rqNdA1N8joHfbdemlLfkcqh
3Crgc5tOjbPKHye+JTP9LgWZWURgnQxatTq4pKrxQizC7uSLdStFsZ5U2fTo59DLKrvpfnA4tOkd
2ztM6D3Y9LV6u2fj01rfrmi4YsaqeYCPCqGoOFJwscme3wc605jbaFu99JKwyUNp3QEtdZBW7ucY
KJmm+lAJeiQelbWB1gUBZ4YvU2gWwXPgy/i6USTuhGjB5wLmtYCkvod1PtODy4K5E6bJNg7QfxDE
HkiqnKLWV6UJglmUbCSfIM+o92Yi5+XIbMuX4HhB4uv4YKhDXMmQPBAn8OMwfmueYhs8BeMSiMvD
ydRWYOui91LXaSacXp84oOfzj8TuBlli058bBNv1aV2m1xWVqEVg+Hr7yFX3eWAEVjyhwNWL7AWA
+/DFft4PQXoGvpo4IMV7QJ7dzBuWfr0IzmcdarwyAATR81SdaeBqvh44PkqTdLv+geCfAXkfXMAi
nIxOBvB0J4TMBrlm82k112gRTzenuAbI8dYoUR4w6Hy87R9EpHxGmW5nLP5iz348Cw99RipbhzsN
4PDrSV/eID+/LJ9cc4+1h/l5QUwWwiZUlOdDOIknWKUHhhurYVir6pB9kllIg5G3bJnlhzh0Nqmf
dLk9D2ztl6kLYgzDk0OhFzCVKJRp5dZzjfcFRLopr9V+N/iVW7XHxx/mL29kkJ1ZYRFh686T9t5N
AkkqydYZaBcGH35aC9iacbHz2KCFYzN5c/dOIRR4nRSjfwsrwIqT8HPaIfeCnIYDE4paMLRxULo6
s/GSaHh+Jq0Wy1J4IMV+wxIaeeLVTg1kyyuhvOOWKIuR5ASvzntXuLgpneNeqQOVoDDDvZB7exIG
EdFTyW0AXI6Q/Fy5NSrgM7KwetcSptf8fHZ3SHkkyfvq6m/J0C+YVA0vqhGUmpdpQJFxnoOZ1ZEt
hkPhTI6+9/cNDLw0v5SnVLeoDAgQNMrwubCNUKFuFJGVD2/UHSzZ+L4tDEJRukKkhnoGcfqfzfFI
mmcuD+z47d1rARSf2Ge+IUyk6k6ErdMvXn1DGFyWwqlzdhTCN//53N3UdFDFKLM8pV4muV0MQCOa
KzVXupjshDu013Hg5JT5EhnHmymhHOjwbsSFqiFap53mdk6QwOnAyjrnxRjOodLiz6p+BCLvnABH
Qj/IyJe76kSIf6xpdcLAVBeSmWyBeC6vbpOlizILlgyKSscgKZosamNE9/KOs5YrGvtvF7mUee2Q
U9ibrzHfEbkx45uzhXiFAilArBMoBJiRgQF/41SrLTTgkznt7QO0dRGEC/S8r4TsCbN53LAZGHWq
+wT77JXpWBwi0WemXJIOtpG4MzwPM83pcOgVzncJ1x+fY3CiqXrr0CkmW1HhF7IFMg/3b0VLDT1u
/5YoYGLd0hJZ3yd86vujjQrF6FidYLsja6MSvCTvqWfHhfa6QleWkxllgd+TMnzfls/rUJGzRTUd
Ulz/5we2cGGaUwtVHte7VGutRvwdwOO6QxtwnteKWSFXoni6wC+y/m2hHk8hWyAyZx0Vx3qASVE9
ROa1scGfZQ2aejZEZphoX3LPb2O62XMb5auWs+tkjMiCfDog5oMmgvxaqtIIww4wRpLaLzwaFRDy
7m/sQy+jWd8pKt/YznY/sAN1iNRa+V+sYs4E3xk1ifyYmKAAQ9fERTpdcz9cV7sqd9ZugsjoIYbP
nKhuuqat3YuPxjhq+oNmfFs/tdTiU/ze4JpjccrrSDFl2VVbZ84upsW5ZGQ93p9+KXu2kesqKt3L
0k/RsqXZfTt9cbUq+jy81jcQ8wOXUwsKSQ3LfWowc3/tePQZa4hdmPT/66/TIGub4qRq/sSRNSzm
bU1exO+MEP/gsa86UIb4Vug+lPQ+vh1HPRS+pGlRLTqnJeBPlBA5yqFukCesaoz+ShtaAeMUbUDy
1TbaEP7+XKKy8rV1i6h+OZbmbGbsT6/VZa/q0CfLDsuYVZzAsKppBtc5QIfIKlT9AYIGNdIsrSnF
Qm8mhh9qbaGvxAAu/oOPkIUEFRgSOQ4th+gpx+c+pFFKQI9RP6ey+Ee/ELVpW/kGFMfpt9EDAcZH
7EhdX0c7NzbLO0++ngR4aKk470Q90F04JnTw6xXvfV6Gsfud08Ns1IlrDZGF3E1hn73jOXGEm0KJ
hPZVEAxNiAZCfUSAIrOp+qYxsXOHpujfX5SFa8HzNbZV57rup+aGnU8Cw+oxT2NPRmFJmM4pOH2P
FcBVilJ9QieFLHszy8xufDyOOKfvzqnT5InD/hH3F5gZSKIEDy4JuEFXG/G8S2lX55uzHOCTl+N9
LlyLItc1uAP+9FoxcGbNibg2k5beG6lhnnQFrQzlqSGhCMpx+LyiwvEhtrmxriwK0/EbacodWwAg
mj12kb4USwP9Yz4cYbOwrHeCkaeyvYXsUhB+d5r5/Z7UbWSbqhxFpbNTMmPUx0Wkip9Tq0OOQtk+
R6AFoyTT60nviey/vqkCHy7z9Q7Ibg47j7/8v3OXRJtKl0lu4UmTKfjVKR60hnd1FM2wrodWtkSQ
jO7QzNO3t7A6xT3K+CeuL01kiv4eOUweev6UnjLip+zwGejm1M3vIUGYwYkp6vMyxEf0c8FvS5Dm
nKP4sCsw9JMdsLoDpNeD2HdLi/qvbsr6vILvOce/8BFitpwIYFDzQuMndpYvYBaWOW/bqcBHep/8
hM7ODGLUIGV2Frm1Zwp5ZgHMHgOY7IyXHv8iXidPdz79Cr31KJSl3cEWD4ZyKryK5ZTu/8qFbNZe
d5pxaPylOKKmLeHmcsJxo5DfMC35HE/awgcorj4+ZwITtgB8RYubGOWWeREKhOuXdQsiAEIy0sUP
MvzbkUYm4botiE0A3nphMl/0sqQwy5HMu/k2mGbYUttmD1kogkxdSIxiRYrAt4Tcq1YC6SN0lE0V
CgminR+RaQhyFOZsHQOK882+irwTDcNs6Y/lq6hJbWDd3TEzQO97kTbyeIVoYz9Pi+JJd5nDuM37
g1nNmSY8y3Tc1TJ/evq9Q/ymWKK8af1yhEnLRYgrR5GzDqOKhSPcti5D1ZRaMffREBRgbjUYHL1O
nQv5Yi/Jtv5BrSQe6m7nfZrYAdw1lmBS7FVhWaURvhW0qIL8oU4oy7a4bBtPSe2L6FP1PMlRxj9E
+BgYyzzmSi0VOj464VmB3URjfhZ4MtU0zxKdejujNzBRu+rpXcfrwRB0+nlr8rr0UzzglpgBPajB
EOVN7nGCdDnGmfFpWMFRQe7rkqcqGioCV1FLi5v+chdYaPSDRpMAavjJ1DIIC4m3iriPn9WxlkfB
Cc+WV+goLffQwmIetqZrX3FtCFRt+FN1ORK1Kgf6Dby4Zjc4gUd9vGndQJu/VwG+5LgPR3CnDHL+
xxGZHA7d+3hfh8t1YQW8UA/umR+ZvVCaxHzMnzOiOsGKXA8KpqKxXNuUChiEOVhZIsdGRSW9WdOA
lQJdGDt3bvm29UbMURq6E5KM0FnBjXqEGrjfpC//QGoFIIoYcKsGFzPE2HkT6w1fpZ8lu+AQZNdc
v3Y5FdIQYIRV81Hz/TJPacqgJCCVXtcorun18YQnh/fgmC95HVJMOt6FSp7tePfwf7KArn7eClY4
+gRxDJBUJaQZ+hD3WqT8dxZAdL+m0SFmHrExWTKR/BO9vDIcoHOdYYSCNpgLYCz/0I8d/Xy3ENto
V2FqvesvaDVJ0xkdzubIZbTWfYoZvrJ5u3WHkBh+vvHup+G8fePstp1T3nbiavHslb4Z4xauiU1J
Djqpr1jnDlG01+jI2zz0W5b9uuAnAhw7Whw3GX3FsAMiBhaCi2f4V5KOP0JCk1RbfW2LF3MJG6uZ
sOwEHDLnkL6G/8rW50WHw3bK+3MO86svHTploLx8JNlBH96AqbRDqKK7Kevcsb4G88F8oVFTbrpN
0GO2hD2P1TVt8N3GhDaPoQVLDTu//MjueLztBEAjgAA3PhOW5OMKpqyxqEIWUl3bbSGpSPqkFbKh
jgqhrGbkaJ466xeqYxK9FnDESupshYEmCuig27RtbYyzCzb48Buig+b0nVWw22ThXGg5xvMdVgj8
JyLnKu6xEW0f6AyavcwYEOGBhTZ3khotHi3m6ifMapKHS4s5Ja1cHIrdD1bZxlpmUypOv68UFBH3
YUXJhQ0L4NV8EmMBdBn0w7nE4QMedj3VeavTONdrmnGc0ZYG9LCaepQ3IpFTw4cAShyJlazZYaj/
S4++ecWgh3pZ6z834CiT1wmtOQ22RTzA6M9ll0RVisLPdWDk20Wd7ni7pZjiwSKdhpkek9ZmBlXG
vuNhgk27Bq/cchdMKOK4sIDpWoF233Hc5MGwy3nqHuSEydj0zwyY2Rhy4jZuBLw6CeoqsYWwY3jX
zZfBNKV8Ga747OB7198yKqu/VUFOxtNXEIyeLf1/0YqMiFuvKP0jJzJ+P2k10b9SWRuh6c0a8zrD
NGYpOGmdywfjqnWtja3GXFjpdFKxj5u++5sIkcgn2Us70yr0Uj+XJOJ+JPPQJbeO+/ZCKBNyWdCw
YJP61T0ioTyPa2sH3JsYX0gR1UbQsvpCosUNfNOUDi/iTfa75mz+vhO4Mk9L7jU1tqgUEXWJFh8v
KsBXPk9N6N1MAxND1LbVlUPlKqksSBt5oJuZSyh0KbRxap0ofzsoS62EKfADgfVfs3+l7iTgYKa3
AJ0b8DTY2DodugKekhj4Xf/va8SXUnMMQbPaUWg643x+Rv0ioYyFhs/Ihw2DHPJbguzUtyzd3Aie
gHpwVLiKC2nw27B8jI1ZCOtdaQJsSaIKICGdbDnvoQIbj9nIXx3c5jhAJ9SHtJS1ziyNCS2SOM8B
AsbLT9iTLl66heqhwrkc+cK3l+SlqsrrHahov3iWwkRg1T2H0xW4ZjjC3veerumO2ygdbPq27g7A
hKdKZ7bSSBvKf+0aH594j16fnF5K9i++damqiZOcn6QLoAeXQrpl+KVRxVZd4kUAI9cSoUE5swII
p1H58NMUdM1SkWbtTAcYrR4FFWcDv1kX0qy/CLvfiu2XyX9e5B8J+KY+0XCie02MXaYe+WFstIA1
6d+yJEPO++EejdI/dxl9fyKjsWP2NmjYzmKCwTO2hyMYBrgw95h7VzaQHu3NkF2D+2gLjX21Cwpe
znlNV97jWAL2xCUo6G63lroyCWwj2bT2UOLF5HbHXmYbkYo2ac7odtjJobcR79L3L2sT3Xwk+549
RTPVScHC2kWVFg7xUjEcbxpETfColUNgETqwPUGqLqPdd60Iam/wcLnbq42tefF7653G8FkQKHNY
2DdS0wBH60AN/cANUDjInIWi8yoZ0y8InChpeA3xOwxm73PumruiWTkzPHrNVZ1U/W9S7ez4n0u4
eX+vZdcjE3GlIb+o4yEqWbwPvHREq1HeL131K4O1W96K0igW/K/uszF73XOGFuoqXN1EwHN4l9GB
3rkjigJrwOr5FTDfpVFeQUFgPBzItj16YDZwHutWbFivNv76Mzy1JIEsUmjIHMdjTJwY0iDdwYyg
lc9T3/ZTCq1z37VpI5ZCqA6vDD65bCSDyDr7RwReFeWUFdg8uOYyUaLb0G9CaHSvlH2BOVOZo4hy
WRoL2PCwpuI1THYn5H7b3UNqN+MCFmvTjkCzzTKUUl88JOyLw20DmRUGQ23Oy2Q4xIw34iZK6xSl
dV92SAS52/l7qmaBpiB/vRU3q2N+0237WVtiML1PGdoVRjbN5VVxwPB8vGS/7ZhSFfaPLxQtMeGZ
sA/abfMUhU7qfdpemiwfUc1iFUAviRuaJ5S79/2r/1qHzT7wrOcipznxgJ5vSqpdTSiBgWZV9Czq
KXy32Ypew6Ruxi/Evit+GhdU6V5mpdiu5oBYRnn9YjPo1uTK9oohkvC+NlASTLLLTpO/34rgy7pE
9eVGa3dlofPsVumELrx/mOvmNJ3cLAW+Qe3wyWQAPmXqayoDh08Ud8hO2uYRYhieXXblypWNmF78
B1cZeSKfaZMHmtWKqCR5/Vs64WpW6kBkeTM28S/z4oWVOFVSBzC+H1bYivpmponIGWXjsj1Hhhnf
vcPTP38F3fv1+cxUkRMgkomYXSZhruwgwjx18zfoFlBkRbNDX7EYXhP+RdWMePziMzmorv5aN5A/
nSlo+xKz398uTh2uM2/+1IRa3tuMytXHLItGWve6orrGHqa/m/L1WjAWRUoBYH+Od3YXQbXeFusS
mYR++vM+mP0xb0OPnsfWxKpQkr+KCSTmuDzHKt0JG1uxgNx7ReKcfifKbGKbBV7L3i7DnYSZjgbc
IOq9bmdxLoPtAUSolend42gVUqybKXGFN/UqGf0H17ehmaz/JYuRplScrZ/EoNmxyJk0gsIAczB1
89ciawSDqACCObn+B1bm1BkxSdHAxCJ9We/erHLNiLV7ymp4v73zHr2uxlmy2bpjlW4G8cGTe8oB
UMT+YZLifW1QyfHBMkFQEosGUuMtrey05C8WLf4OCB5nX+jH9uehQAv77ZyGGyFH2t6b3kMMraUl
1E4B2lNl2sXnql9Zh/+rbqtIc/GUyCNvDzmy9i9Fck/8TqjzHCLf5JUJN1cexCPw4cMMr7mlHJXT
0hmYPRXNFiaeZ6w271xZCGEaKUmb4zjX1aNRV6ZKPDIL4zaBb4zD7BEN5b5k/fPiNYRkPZ236wC6
0S33uD7GdX101dkwCKJUQaurCDt/FunaescBeMGEW3CJy3rNQlqCJzudpAl532o6CL3cO0RqC8Nt
qLiYH7+Ic6/lJol/rjW+IqqpNoCMquBAaRLbk76HqmrTdlVYwg2QscglFg6a6qk5qwjAY2arZYxe
M1aikaDvBR7LsRIT97h0o2bL/nkGuw9BRUhAeMzzz0mSWKb4bBtFYGV/4hRVoEgUwqc7c04QzeGd
nQ8vkQUITeSfsjl0r/FbumuiDWo+pI/4uyr4T2OQq2cJ/hZzPe7plct7mIWJFdHWeKbMNM+2qSBq
7rGGnXoEeD+5GqC/ZLK3c4LUBYSWf1YO64z6FxDA8LPLKBIBJ6BzE2ifHMImdr2TNtRPaBHbRDKB
VQcbYWWPnVaT+SR1ntbZD3rX2lkmhulhTy4vRnVMV3dG/7KMBlITxPt4B7hj9sHak2IDfuyZEB4c
izS04Y8pHFVIZhswdhOXXoDDloe8BuIsDPl+QmIzE+ciXPs0TttLeY6ER1itmeP20ZIlvYT9Q1va
4OLPEuk/uEOUUEkK+ffJ/DqHI3/+qis8znhB5BbxLd5dgXlZcp5q3yS5dubMIY1COEbboZV8OT09
SBJV3JkG7xLQVPjQgQ9uwCRPHMbsPuYJNeC8vV8KKRyjvFazNEoLSKes3DKGqcA1ngNpLC10h+Or
v8oBm5boAoodCYtIVjXKPqU5gnBxQZN5DRn95bn0hEHVCo9w2wO02tCfmaSFtx3lc5LwA3TfsIpq
rwAJH3rAKPVw6rxANa6/+VcZ5I9OOZrZcCm7u1cJWrS7uUhPxqOcN+vIXmZ9ti9x1y/TDHVAwUEM
qdfcaMoDd/oUUWZxeYNIiga+yF19tP6Khduk3UT5LSGbRZ2YCp9bwFDhAz/VWh6Re2wPRfIsNxfv
xCALxmu9Y6Ke1PfBzQYFdkmqoFCH6SAorKshXqjepBJzqLZ+mfBkSa73EUOIG89x0KWdDg9+S8JL
+y19fODm9gTuuQZRg16XsA/px4oNt5qTb9H1u+hwopfUiG/UzXGaMMrowgulaOtxaj/w88kS9/o8
v8mjfVVu3SUWU9FKwvJ1njn88s0isiNsf9z+9FgMIeu+Pd+xTkWwGTdlCT5ZlrZeDh3N+qMWZf3t
tACyvpS4jlPcB5Elkcx+bskNAgFLvmj15uvee58hkTJ6s8tgcoMNgf7nDREiR2rFCkel7uS4yIta
XiPdLBJjsK7KCdxKXueZ08HXp3cy/d9DcAPZFzTVD+/QCbtRG3t/nFFJ/9OunMNtHaapJm1u5ri7
Aoq7ZQlJgKOiK7zRMF+hOYjHrqnZc9kZcpwQCZQppKJVuXhoeJfYkutKhMZWACMkk061TUgfo4Me
6ICthhCx7bxlntS71N2JbPyqzQj0SICEOP/PPt+q9CJDwe6pmREH+LCpi2SiG48JsSuEqhTkFUlW
c8bPUbjtmjXgTNwXDb1BuhM5NTfSkSkoNlPiIVS2stQcAmPGbYpQXiJnmI1/0PKGoqhKyVqn6fYt
WsljC93ChjqmjiXKrlTgIREipkY0Ar5YGzdAqtn7gv4g82/MFMSsp0Jvm8hXTCVKQdNl2hc1O04o
a6HU1DFZuGSoKkfnYf46XAaVJs0/9WWktvtW8andmyET6+kt/4j5qeDvAGf+xSEo0PydhAoQjrIa
84ogmE02W34rdgMfGgIgwCNlpTVBumCnQWHU7TphldhiC1s43mIao0PvpOKkrvMnqBAa9JnZbzRm
CGhkqv2cbgYV1ZlCbbQezXt49p1TbeZVrVFnOIVHYYUXSWiI9/G3bX9yt7OeJAB/7+wGFmbxTDzF
rgepd41JnaOFOk/4GC2NwjtV2wj8Kw4nZTvmckg4e8wyL5iOdHThJvNkGYNhN+elrblocAUsi57p
nDWtdItTlJaRgbywo8qMOqbQSRvjeGGVcA168wWnRAvSEKZmEwcIlPvrJgIamtwv0saiFC4nKfgX
sopnTWsN1VweTAsm9mOHX3IcPpuS5ijM9iBcGaWq0BknH7spto9MqWIk39M0LbIDfBxmr/CLgJfJ
JOU1DHbMBi9dYeku1EXyQBqt/T/VPs3kaJ9JLuDd0nTWK/BGTftv6KnLn6FE8aQM7VBL0JLjxsCp
jbUDvwJMhgFROLRx1/RtJR2VTqOfcZnwScIVDC9O22qdb0z+0/JyLTTMxmUFMZQkbLylj0a9fMk8
6P8oaUurnDWnvQ2+lS9IW/DFj469gX5fcCKgnWlhVpJCrwPCwvupUn7OsN1+eYJ3PsNrmMRFyVdz
iO6itWhZ7grgf+xPwx6UOCIwJQUzWOCy5nLeSW+W17SDLOmsYo6nQto33POZl1i8R6EWQdg8syvZ
Qc8vfEKcccZxuT6oJMEHnL0Fue2s9yBhGiiioIYmlgAsIk7Qr/PPCQH3VrnqW5EKfrdAMVpH7M9E
WTofuxfGSxbU0UPKR90o9/iL2bmhcdsfB4cWtbYNT3loyR0Xb23Xl8Arx/nAsCIgOx7mZh0acXRF
ry3px+q3He8pDAyGgzlryUs1jjaIoZtk/Nw3Y4bsH1LZnIlsPl9ptoJuSlsHxTUPCpuCM4xcj0rw
N70jXZoGqNWYfAKZmfKzPRMBmkN/oSULZSSazL9/wcu8uX9si2sMntWMx8tUq8YF5vio8HNopnQw
MijAENrTahAoAKkdYkvE3rLMsc0D5+Z/ZCeQtT7Y1fGLnILYZVStqq7mpiIFOoAaczC5pOjNjd9U
bnLQhvCvnrvGV6ZhISseEND0wWP4oVFA//KwjGb0bLKzq/zo92MgHEgTSw1gi08cCnloEDaBrZ5q
JIWZ+3+MrY6rPqiI1JBI+qcsIgXUhckFMmh87eUncfGyUJH0I8XXiCb1SJX5IJPiWdw6oNX8XYDt
/P+HTNX0xD/miQlvfi70D0gccuPISwKTenvDm0n+qwh8qQ5pyp88mp2V5bZq4jiZkxaDXFitQnxB
RGOoOf1RhW5/NypYIQIGJN6Sz7wFwLh8y242/ASbNFTJ6C7rk1Bcl0Q5GOQE9MY9thG+oJKrbgQy
1yBhSYRI3rxSDaaUPl7KaeQ0Vn/irtVM3OHLJK+S4cXX7jpLJsPwSA5XdkAQ6fwIzhxwCyAG7JF3
vhoJ43r1uvUVcBuofmL+3ISrHmp5Ct04dtijoBGOyjt/y8Q9kbqNFZjhFNKqDaB0Cxk520JkvLR5
dKacp/nALxIRt5KkQ75AlV6VFTJb0pSU9bxMTubijjCOsptcmHtKTFvVv23aPHD6r+UpSSXcPFAH
6EQYmnaisU6XJiaUZCfclp58Z6yCQ/BR+hFCnqCbT74KX3S27XPBlgVu1eUuRo09QIlVv8x8hOZk
mF5/p834zwIluegBT8s0pYCLOdpF0cdMd+mQfy5R7JHZPuLs/0calXTkV3rl7xDK+xIdwZPd53y3
BhHlMG+mcF38kwcCVdFrUswSUPHE8qwLXkEmxpY1QeLwYY4HWbuKXvqBQE4F+aSliNGxhd5SfSgT
9wOuXizSeZgsFWEpnaeIRCw8xN3U2znZ66RT3kd/YaTxzNGB8Ugfl/ORbkVvLZiu3y8IF6H5vJUc
qk3FFrX83eM8pN7MiApbvJw9fCKc7x3FRDhNy+P6ZWFo0XrxPZgPgeKbEAV+lVJfQXFe37liLqCS
5sbFbaEygIkbkIbrF9qWYFHCl6rel2mCCCLYJ6ZFLz7ACuQN81l/CkPJYp3Ve81ZJTsF/fYvUrI9
oc0ZlOwh6oWCYBCuZQFE+ptamoHl1Eh6STs2W8FzXTt0u4H9EMKEsOu26jhuouffTjuhZpQtCFOu
4J1aUQQbENO/NSc0sOC8EeoM4DzsicyiC9F6BlEkDtTIGvaFN5zWRfDLYTfDM6lWzsyJKgYbdM9I
kzNyqaLkzxvae+ic758JUqeQat9f7U3wzhKT7jfL8O5HasYWo4izSGgvcjyYaEZ0Y+uJREBvdZrL
T4q+6QnEMIFcSQ8yofPKlniR6oxeKD57CNl4/O3ttrRsXGS5ga3OsgpuHKKWSU14o4YW1bseDMp8
hHUWEXCgBJarbVSOhWUFZv3Zfv32LCpDdKI8HmYG2tu6b+zV2Nzz9lSRDPJ1Pa9eIzBnEUIwBt72
5nLdUns6o2hWz+Qi1hi83golAl6GVpbC/pLdLksNedpiWAgq6IudosVF+7h8uPRAZ3VsMxS3DwBA
wNPFJyr32Ple1nxMXviFte2313hi8fVIWs+hmZjqMcAvMsxo8MsJkY73qI6d+c+8iwrfaXeNRLuo
q4OB8jJe/Le1ciOQOdPsJjyCNJnz59nhixHOVF98cAV7G6PCB2K/S/Z2jl8ZNPkCxc+pWjZ6pIBG
1XUYrJJFQqpNLT6A0DUoGkesTONFanv07wauH/MolAFQVIGVzmDLC8KU+ex2rOAor0dnNPEF86+d
th3pbuCOYz8SuR2CdNWHNGD4IekNFmBvjmHe8IE8IMyYF/ZY01iyh9sCCoFqhbgw9ltW4fuLkgaN
knQPmXt4UzuYlj9dJxBM1VOkk9tbzbwkGc63wfyCdbvOwgVvKZwR8Qlee5lW8Gf4cFcNRpNWWuwF
tscV55Ux+OyGHGLinGsb35hjp3z7y3NsYIu43kZ9dP1eMeFJy7N76h67M4Ez2ch9ZQXADK+hsGEw
fh+GkcHyR+WMEfUo4+grPrYo3Tag7+eDRwrfxwcfccxqIqMm5g8x66TbOH2/Eq+r8vw9iXk+OLer
mWC9a2Q6W1OixjOETWq8Sovdzb1wvUrScKZ8DHI5vInOxl1hyYUodxoZ14/yoIb8CrGlAely7vfg
4jMdXKkmLxJdMEo2NDfWh0H2kgUQJ085wUdwt6ok6cYssg7luqXOF3vEk+br5AYt7ipRItykSSUI
K+nZihPPWryfziqfGfQV29Py3dFj9PbB8e3FpM3B1NJuzuYWxo2TB5el5JLRRuItnef701vCYd1J
AXeGdOiKMmczT96qGXnW7BQZsm07qYOKOEimurEx7OBWGh1IOGnakNFtabeMa+nECcl8Ui5gqRL9
NkE7tKhRg17APiPFrm2Mjdm4DwRYLqrUYA6OT6muDMXtnxTBRryGzid6mITtAKUz0n5K6/JAQDKC
ih4KygXSC3xF6uxvXC88xhfzi/db8xS7lPiUI3ox2KX+VR7cj4VnHlch1z5vM06NggE8CFNeQkFs
tNHFbMf+3fvzL+TFM078xkImxBsyJlk1RFW7LQo6WNC058oV4LX/1xJ38rHQ6BLa1Q08Etm3Tws6
JRDi2gvcKaMCFpMNW8FziTdin2jHOheSA0VkmH+MrDGr47pMsZTLPatXmEoaWB1T2wt5EexivYXn
xYzW91Ad37DY50VO+I5fVSpZ7Zxroh9D6WXjMT6AQu3YctXvMdf+XLAsz1GiNM+qEtsmxcGKYkyt
akMSyrdfWIONjICU/kM8hQLNesSmu7bF6N7w/gkcH4qxyqfQKu45JdiKueG8DBDokGQ3ZIyUvPTr
Su+TEYV3jbA0Yq1Cb7a/B42XKYoxSFIROPg6+qquOBOShMB7TBLYlEa1RKQRkRuVt296JX0poW7Z
/q+E1L+x3HMhUr+oo07Kmus7sE+hlL4rXxcHkWcFZBmP1DQfOo4Z+mUXmwaQhe/35J/iLqx0mVky
xnpWdQXpDPOJ8NYaUME2jFg8+3p1dzTZxQYzGd6b1Ti3nlRsqzBYzG6hstOfl8zdGHcKg3+B7SwF
9gf/AYQ9zMZD1/RnXedWVYpOvtk5EzB/yQZmQ5mUXZjB8l9O9F/amT/WwnHJ0jRfoTY2ZZzLUsQf
F79UKdaR29BVhUguvUTj5v33Rgl+wFy+sEAxldO7TrPXUfqL8/IffUUBZlzpqB/BaX4yvUuEf5Gb
iM9CgFeBtWx9HG+TzJSa8oAymKIv0PJQpn/Ygn3fo5t05cgw+IZuBQBXykSEAVbOAzZQKrF+lk44
p3Bze2wrquGIx4dgnmtkekeGuF1WaFZZn1DCj9ZpR8puysxQFqBd4tSQMn/deT/Ay0W8jGubbXr9
VP0Go6mGPl2gW4NkHTFtfOukZTIwN/CCteQjHK1gGNQXsAjpS+ARoTVVAxCfT3jp+YeIxGPAEw06
Cu4fp7BUdMSCp2vJ4qtf3HSemfzDOTDtMunXH+Gz9gTpOCau3zSdzu1d/wK9AJmArTpF2uUyO3Xy
nFeSi3iXv93RzZLScJchR6svbCN5wDoY9JTNJwrde1NV4jgfBCfQHOvM74ZIrDP5Rt3wcwbXxR2W
nHslDz6T+fqQXmkgFTPsujv2ijFqQHYTSSHUwWH4LF3mrGoYBHjml9uQxKeGu8hq92LI/XBRLcwJ
ufpHSoRk6pV14T0nWWqflRkAk8FTPzwveKXCh2cGy82Wo2mU8qFOmvTEump2RW3hF5VxFIoCPJck
aXo+w9Oa11VpjrdWqaBgjoctvNPoHzTt0R++zZmSCx5NhYPgVIYkayKpsH0a2iwKcBZRB+XiQ0pN
1fPGxzLRbUPea7TBbIRQm1lLpAktxemHfgMZcZ8hIZ6cK8gxBiMhA7X6IMCKXQ7xKlWR6+zLrCuf
jkfSYLIb8p90QtH4T+Dp9UZRs+IwOxAWYoyS+EzxBipvFCTmjWtWkSce9SFS3+ob4swx8CIn9dwP
PkuIYuwJ1ioBvrB/WSCNf8ZfNSrsBYRxKQApwpFjci//5pGhkjbjTcLh0kxTPqpgsGfG88dOih8H
JkshsqXgXi3K4yXy7kuvpYX/M+70mtsqJdr+K1Yu4xzbFJnSPfNr/z3kgI7d1hlIri+zkwZrq1T1
gDw2N42PZRVgd9/kgvelyZgFqL6eMhxrb1oEQoRfHPv9vE9AZ+hr2yIGM2uMl6KsarU/JHdxejK0
oxmAs20PHuc4LtiYHvGkC4zYSbyy3ShjYlyMBhlkzW+a3D/Jc7P5Q/ETha5LD25kkpPm38EQF+//
jW9xCDDt/Gw37um/ihBwdrYOOVsZDymL3eBVVa8THklNw2ilvFEGdKZ28E6RYjyIbI6NjHt03iwO
32zE8VWgiyNV3QITDAmEBMewZQhLWqW4ihDgNJhhqYw8Ovu+BqR2FKt5OoJ3N4dy0KYxx4EtC9uO
msi3RMIyoR2zMQJiJP7axooRKlnbxqsbo1FTmDaMZW+0k5WBoyFaLncEksX8hwMgDF3KpDJ5HAgz
6MOQ1X7I0ryoJ8ze9PaHbOAUoNBs3NMX67T/RE5vqeArJ5K49c2QoMd57eUwWfSLU6DpLu/xW7s5
8i0CV2oLQtm+ZfBrULmAJ6Nyp5PFzQj9vCbLAyEkJtsJTsY7wnkmIy4nNB1TxVD+uL2lh1aMWnQ5
eLF+LjIz5VKMCnIDWgdD+RK7SK88/JVIlicPS3W07aqOnY5sMB4VooOvWYjISsbMim/knlyxX4df
CuqflUdf+QdEjtmal6veMzr38GvwMpK5X4FKKckSbZemIyB6BhMboCOa5WJfm64mBpe+hwdAExp+
bPoBMSHWapMpiDz6ZWwetKwdJ4bLyNdf9z+G7qjEMq1sQQwwemKRo935RHcFTjjpn/LWF+lnOEjS
5yWppnvdBCJwyKy7oH/MNkXf6+1mvGhGGrzAqFQ+QDEG1PZ3lZX2EvhiE/F/6Pcsh2UPPgRhdAI6
IAf2YRzun+itdFoNzJDOLINwaBbcRpmDb3qik3huRBOviBudbes+fqitJASmFEXK20vxEc6mHacT
yJeG/cUSJMuGBlNSUTvtY3qiyCRqCMMBRbfAzY6r7DWZkLMuqvIaSIMsGv3D/LvIa1HFMaoiIYpW
aliuM496NGVZunOUXMCN8Ckxlq6RtjR9Llh5KkgRY0zhLHMTgtmJBoZ5OCxRB8SAOD+NVLgW6bJg
/Vb7yzyR3mCsj5vJkfs8DWazC9CHvECVyEbTwYQ9JFKw40aZxIxHve6f+jdBuPau55lbCrfCzcif
KdL+AlenyESXWBFepdLzJ8zuoWwUk3zGzQX36Xc1La7sUWzn72lmWTYadhuPKFwkszaBFK5ACN4P
Hj9My7bsJ+dzY1e+Vo23hY73R+xH1lIoY6T5gR7h2z52NSynpv0weOy87BzlbebQ7siTqS6tsOiq
+RZk1HBnhmxhFFOi4S7I3OKuYJ3hYEmQGR44p46zoX3y9zTNkBPE2+PPFx1toGtmHqXeCEebhmqd
YxwWJ009rVPoffGat7muU2lpQNm65C1KSTlOs2ZF3VEg5ZAK+Buv2chcSGSvXAvJDCpM/iVr48Z2
bCSQC/1Ynr6sxnQVcki1IPUq3sNZ1Ba2rnze2g88lbLEQDjQ6nkM2tN9TP27oWp+/60jRQhe2uil
BjaKk6R7g6ASfPugfsz4TcNGpDKcyx2yHmweFicZae+hW1URfYywyobBWZmESSLqp4CRmLLI4Ebt
PqlVjGxiNepTCn3wPbaiEjedSq4R8qJza11QX33Lw95r64UG8V4LOa+Fdoznxr9yKq3xi6S+KNJA
EuvdIBmBipdL34ia3rRRMSKURI0F/XZKPfvQHGliZ8x8Zxwwb40VPem/+yIxZYPnThD02NEb0EvT
3H0PjdnW12Sj6u88IxpLjgDM3MG6eY0XlZAGh1p49WeTOjqcH0OtD8vKIVQsTzNKv0ULCQSnWrLP
v42z5YSdJutoyPdP8UvTTFEQW7I7ha0sz2RQ6zEufbAB+IsQsvKWCH4N45jFDqtf40zcPQJt+CQm
1w+2MBBi/aLxFEuvdDjGwzxuSuzIOg027oIIxlz4AaOcnsKiVwKmtiQ9dnf9tac8eQsoeCW+b50K
0xXsvz6xbhq9hx77+PkRyUw9GbHRcsJ6fQCth3IZ+TRUiFFGY6etH9hSD6b28hkdgKshOykAqy7t
bydw9pHfNFPxzoO8O0rn19H/ouDroc+jItmOeibhEHC5zFP+OfgIJPGlTem5IrF1H5WQXNgytk7i
WC5lhqvpX0IaYWaDTVsxh10v1dVCcQ36vy2KGF3ML2jehvGT8PKaNOZlHOYS697aK4aGIxtJcKR3
U3wp0WlrOw99mNrob4oD4qMGnWThLXiorTYVRlBmu2ocNoz4coBvZd4eW0E2169PIKazWwlo4GGH
WbN9zICou/7LCI/XE0j47244cuv0de+UOevvjmlrOFB6StermFRZiBghTXjRA2W2BbhajpJg4hdX
nYZgz/95YizBQFfKs4xtht1uaOjo6q2gPzp0YQv1xr7B3qyMrJCCUjnQzHH+tYMckUm/CRayuh4M
CtbBE06KUYzLhsRbfKrEXryfF1ECpy4HmuOWOPb3u2O9KoOItC59xgnoLRQsoww7YcMtExtfa8pT
a1APudEcVurUCGgPoawFaYZhldCZB/k3uEUkWzniK2OJw2a7q5zzN3ZBENHg8lyt5mNa5vGHknAe
vBlsaJoC3VjDgOx3YFnXwKQpuUShMLAQo/F50tPhHrggRY3650vQuT9O5zjFjlRN+0TGYjEmj5hr
OErE5n58WsUE/6hzxCmiI90WEy03A7HxlCkMbUBqgR3WrIhw5DrQID/eCIYox32itLc08+odGUEB
pfr+cSOT+/hD+mDym7wlnSx66vuUu4mHIV39Qw6YoG3W1SaHpILS+0PpyJk5n5xXfMihsISCjItk
rusX0FV9sPxn/Q8hywpShFc6MGVlv1F4pGULWao3LbyaSdGclLNTPgLodAxpUbKLvpPxqkNEQ6Ya
eid12DH9IqimYbDLqnBooLgTfEGzDXRVvApZZicDrNQ7r8aoDjI9lTEc4k9Bg5E9rNIuZ25xB15M
P2IolLpgZTOa/MYmKkHuZ0bspdExb3tPPrp1yB9hfYE/spfhnnAXz7Y4g+vjuX//57LI6MkrQVJj
4R5zSb/206g4+dBhJDT6LpuoOjIp3hggoBG14OzjaiziU2YPdOu9JYVwi87P1FEuu/3mPlo7NABe
76M4P24q8ohONk25ERF9sdyGyIcf/a4DuMV9XCuJlV7B8vXMSywkg7OGyIQxwSm6RPDxPxadjlTY
58oRPw8JDBWw5P80C3pfrphKA+45mNOZz59CAcTRK1rmGQ+scC8Di64LroCS1pdWnbsWcRxIqScm
JdebGMEmdw9fl9pzb7l/17AbjCDgvaNZWWreZyeueeGHMR4232Qav37r5otstMOvkdrva9MlKb3C
roK+vyx6gKMrgOUQhy2p2G03IqBtu8lbfpxi2AF91GD8Fa5jidWYjAU6Ltt6e5J+3yioyxDrt9sQ
O1D7IIMIkpvhBj07AdBIHH5UFyitZKo1ikF0WaoLmhMIg133io+/vHb8X12e5tjMy7ER+LjyVJXH
0x3Vp8NxqwH+IADJigupltPSry3p41H+Y2qlf2dkYwgXXE/7x7+eATkGDuOaJVUist3BatAjPi2c
joNfW5DoAVbCiMPOU8GNWgi0OuaSKBpzusb8+vtkwOaJf5VVkZTynhQBdJBhXhCGBAPyOLtbTylc
AFvdsFVVD8tURzPgXXUUgvDdKSv9s+YULsIVzR/L4Xp+pLilKCTudOX29CPLZzkKmG/PVAdi96ei
BEv0K8yLQOEkbqkcDCC5HQgNi1LPBJYjb8Pmd2dN5LtIlkan2UsmHCKf1cOv6ermS/6QCjHXLKCK
SIv1NDE5wbjbLz1zxHAcC0X1vCnivNkTRmHHvqrPD3PO5/8VOgf9SHowBAUZMWAYBynfonZVmxFk
/2iU321IMWoOeY39QKnYAW141m5gJZU8PTFI5W7UcHa8Gs61uSNWU8A5IFLTJLdtQIR9eTLWfDCG
+i+4vfN1d2Uch7V0TL9tIryBMGhtNubiE7thFsdMw0Rgu8KQF/2yramSf98TIdaGJKthmw7MqS4s
ZvaeaYQeSnrBhcdfd5T1/VIIJK9yKkZ15OiLHoRCC2d4astfaZTyjp4kYidtIc9SpJu48SzvTuFZ
Y+HNnsL03WPOBkFQ5i4wDi0N+CUgtsdTXyhLM1zeVduEhrnwbXWpN5rpSV8iODYfbbsOiRj70epK
/lzT+XYUIs2s8Dvn/4WZFdazrH5HRen8fUJLAw2MY9QDWTwalA8ovQDsaCBF84c5RoBr/fHS/Jel
6K39NlzZdlUOddnB4TPwVqrTTCM1rctgxvrVUfmR+BQ47fEI0xpS3IlYtTk8C2ARsKaQz7NBA1/i
9olV0v/xb6NIAihDol+XMBGdlTbEBAc++ItlqRlDRUHIW2rwc4w9S7rmrgnZJRDsvfxHedcIJ8kZ
F3m/WsfHBM0muGJxblPw/Y09WSqwow391pXc53dxhhlOFiS6uIyrotXMNQVNpGoyS5yAaUpW6VhR
rKSHlh7pyPHsnrQD5XaCx/J41cwXRZcUIEHE/PmL780Wn9Bc/NRsxEtvv2RyEil9McS/O337B/0A
FvrXaeWoJD5jjZnmZdDGzf3DxSByvR0qTisegTToVLJ3gPutIQsnx2vNqXi0paaKGqXA0tn4dkg+
qNlFu2XtqEs8oOpL9K9kg2UlI0li1AZs9bhhVc+2HdsOkfIaCOvCSW/DYop1Y+nxnFRg+/pDAD9G
D1cb9uff/Bec6o3Uk0kVriiTWlqEuKqzgBPebWhOLWx1eMWwh2E7bYTtguCKE5fTh5+3OzzFsHgM
s5C5HU+E3rCoSXeVKjnxqjiMhgTEygojA02GWj1duATnooQTy8ecMeFbHI+sCclLupTUTEn2h75h
nU8ek9CiGSEYawVXufqjKhyiMILOtOw8QV8D0NSBkwPMoYTsL1aqKzaUwuhAHLkLtX10OXhHBQLZ
zuwDl5ER0Q7AfCpAuPUuUb6sxuNwWlOKBP70gO0a2gOzQP4XKMVI8mqvuz+iPgUvdvA2XXx6bU4l
qs6hFlPCdHHqdCwQSFWpEOhObywV3gw4TRXvY3eGKYqmwL+I1kWX+EgQbiw+fU+zmiLXpXkagX9b
Ub0ctjCYk9njjI11VCnoflMPaarSpny3yrSQywVINcfnxB6UJ4U0eCdGk0Mpxjj1+RMmYDIiqObE
j2bSBO2FhivHX4KthEkbv/3WBMSXwXz1yRN4djwVTrZk+x/1LXAnHvYI+RxPCN1WV4q6zhFHUCUe
j98NPYBrB/h0/AQ83OXzSe4H8t/RL2CF2LTYC1dwAFIBovoYXo8Xh8kyZHTRiR6pqwKQC5v5T9sf
lltXoEVIf+LttX3vtFA61O7GbgDleCthpGwjalYjS6ESuwgbK6TY5TlMOSBb/smNUawtcUwCcBOJ
1T8SA1QYKm6yxaY8Wn3j3TggyXGjutfDsNeuU8vkRAJfKOSQRVhJxAx/5dPomPZYW1coeuFVMttE
lWgp9RHwXeqEbBRg/dbo2dpCBkntnrEM7YJBttHENtNyk79UIsfLPi2GtmbhEawXLpJE8riYW2ot
FU2GjVgo2i6qQ0L85H2IqUu48+iQ0sikq8B8JaUv4XTw0mfRiJfdmYu4KWUNXXIAk/6ZDga11UQq
vtA419jpjWDpkNa9zw+nC+cGT0sSYbMpohBZ4Jav6D0wi6ZfcU9rJcsrmITjNLW039WxGPdT16vq
FY7gx7l+D/pMCoDNC8y/N6bqVY1rXPfV0cvAJEz8QB7tvD0sRRfdcouSozI3wWdrjWdRX6UqtwFq
0gG1VvpDEHRJBDnhKnz99GGMxCKsWxAeeMJbN1YwBxZdEFpCKMmSFveS3e1dS6GeoN4zg3/WaxKl
iDIuclLT5NOh186hKQFBd4QSTWLJWYCgwsY4TWgYOvZyulwlFtGvax0UUrmGjTT3SW4fsEbMVkfs
DFu1/EwfVmcG76e9J2Ue2P4bWy62z53hQzbNvpSsWz71JDLFQ2aZpCYkFjQVPqLvnrCRP9ecBTWV
uWi63gWvrHcORufog9ItsQi9r6bCYXxQGkmijxQJZTk7K4hJmt1qrnBl2Aa2puGh29mAGMvVEWbU
rtdooEeTwKxlDdCEMt2NfOB2XhEgC9ec5o8iKWwyH53Yj62/W5tEqnJK0UPgmuzrGl1LhvHEVI5S
RxBqk1/xiGZ/sLr2F3B/nbSuCXw5LSiLk4mUt0qAsKqCWFFN1GROuag7NLZWP/6XWTjiMnhquWN5
xAoHFdUL+r31xdthbQU1W7yTnO2vX4f4GMyxrvqRPvJZ+TnqivCejtHqM0LvKveq+k+sbo09w5VE
PPDS48U5Q73kgYJiJUCzzSMvCLk127WO5nVGZpPFvezVU/GuPyVk4fNrQsG/avZZFtOBJKCBTPfY
AQi3BtmT9qBbevFgMMD/YWtINbHTdd8BQfjMS6rm1gHEe8+E3/g+VuNYi91gRUEoXjWJFtiwIBDp
biY7Z7/QiCxqwU+MLWkSKYySndvGNMFv//v6kr4LBd73OWXeTKMthzWMv4hLShcUWAzkpiaEH/zL
aIzsVg3c7iJ4fxUY0zH1Q8NyvmBCJII+5V0MC08OuGWqlvrtc+Y26HO2yCF+L8MRbaDxoVrp7JwC
yKjKYhCmE7Zz3fmX6DY9ztklyscgK5WnI8/bW3FumRua6IASnvVGgbcFwwHynrCamS4poCpVLq1I
HD7s7S5zwvg+y5tn3IilCJtlRNS1z4rVnRrmJ8iRAL9xzFqJzgusLZ8CD/k0Qeioaup/f2tRJqFx
VLz6ISocEaAkTVoeeb+aFIEgTNhrIL/pf6fHxTETEsd6SpUkJx/2G29S8HrFOquIC4lrejbpeRY3
P36hd2wvORTm/T2yqwxYwIWXeCfuAfj084mJnXE4Ynsv6gUEXt4QURChoZzQ6IjIo1fHOOQCy6Sy
rDVtZBVDEqTuLgur2pjolZp/h/VHuqTjZ/oTHCJUBX0RUTBrohoefJGrF/PKUf1Rx6QYOuFxE+1Y
HusbaA3PwQjwNQ0CCyxHAOgthtaLvQ8/07Xsc9xPltiGXDzoOIA6OSUDR6g+oszMJyI6Pj6hY6ag
GO0wZ2c/gri71wR/8IKo5b5452gUVJgBPkpsqu7pulmHKa/MIfmETN5N9rECwN/6rP+Rn+Edy351
QyNqN/Q1c06Ss3nM3wR82ugwumpBWHjMniDUVwVaEGNQ5rfP9YzYNUGnMTxdYp19N7IvVyKdWYOn
eXODVe9Goutx/GPMZrDWBCXxw9mtW/YINLdUS48BrWYaeZ7pRsz2PYI3H2R9pQ9OjsVtj7iwV+qh
yVy2yS59cLa1qvTig6XYkjA6yIYjJHDOx4hc7s6jsdqrotsTAP+3l71/IIl1uh9+oDzZmmNNYiEG
ijCYln/+m7xCDMxU+cBPapLgakhGFCCKvdgw6PKvyY2YKJ+UBcbmy+h7VJjMQeRxKtw6zBDWcVmz
eh6qaf9wpq6N/sgspzDpTF3zg7OyXwKsrX4tPshxlQZNyHaV4Ge6uG9JmnCleyWaPovyuo/c1B8b
/hEtWIGLFfEILkwbm24AlpwiwxQ8pHagILkkiZG2xOe13CBLIHHkd67wkI4yZryIfzLRQTktqeRm
e4Tb5uUSA/rHrUS6/N27JifBWe8VhV1yqNAfkNtnGmK3Kz3sHAInBcC/jQ0/zER8mb0UdLUZ7Zr+
Xy/gijZTh230REpNYzXM3zNM8OcE2jGvss2whJVsudwHvXhDc3eFj7DjTkpMFCM57pwaq9J005VI
6G+czN8IcHLk8z7VUD28LAEB6hySgO1fDwL/Qnu8LExQhrwmaDId+7YWGsRzseOhaJhkjkEJlBas
94zvt+/57ZJcXsDvbS7u8M1+yc38qXcc66vVACxJN0Lx7UW9PFQeIzpoz2wGJE4X85G2/2dc9lIi
eWuJgTP3Hicy1bUoNahvuLO/ji3TXfXz+rmhlnHmhgtRnVnQgESmWVU+M9zk2t4kzIFk0yg4ckcC
GHOWDhZsRwMoCNDWT34FSwvdQCnCOscq8b7u6Pc4Nay0MqndoZeaBvOAZbC768fegN7sCiOCyTg4
Uhkoh1W17E/XV3WSy2qHncB3rMgx2Xs4vy6oowcEHaHlIr5CQgcon1nB/vkcJ2LiZUjop15WXyJS
AMM2s8CVgmP+OpEEUGzJ9KL5eoCkomlXX26N9lLvNf5GQ8uI7cqrHb8ucrqRU2rW1eSyGw4sW3J/
DWPGXGkzIsLu/RcyjzcDCc/pBIofksogwSxc1+OgXmHnOzpZv8VcWsx30GV6txW/2DWUPwa0CnP5
GdHXFs/eW7ZGkUGpFFk8Q05GvZRxgJWDwhHXRUnZs290dD/plvjn3M99OLQkEck8/hcym8hsAc4I
FLeXURW/exHoYTH6XmJAsWZCsWqQ3lwY/c8HV056hi8qxQL35NKuVSG4Qz0p7yL5RdDch0ZzLQOS
/915otK+yTfWp6nQdDgk2FUuU4updyjjE8Jx3y+gRlgHHAbXqc3VvHtPljfVrsEJvvpsem1fjt1E
r4Mx3afRJS0TYYlXMYv8iihg/w55+kLEoOqqin0ngZKbbgKpFGcQKNUIF3N8qg0otd3Exs74Rbnl
6Rp5mkgtZVt58ALq6MsNHWLNpGK7nCR9t712NZMOedNd874vSeGVu1QAbDNAK72puSgQ1b+Gz1RM
jflY/OmDGE1E1vCLlWLZjrQRBKfHvsDYT2Oi0UMlm39uVx+5kTRpn/Zb3vPM3lczzSOnzgVNk3TC
CmYDy4+KobHYlh+uxVyc0odOCMlV6EE1JYgksFEd156AGu6AYDRvgZfNnpROKZ+NJQHcaVFF9dTe
vwFvKcgcumYZkf4h6erBJAol1IdywXchgqeZm9SXO/r4mCxMZe5fz/B4yMGcwN92gZoovRJFrxwA
M3wZooyByWaDa1wIIl8/pYYBCuUbjManD+zm6D+AIf5oau1tvrA2IuthZLMsRa7ZzNkeWPR8Bywn
NAloqvsVBthd8uz1/TnKuZpy+OaDPYiIVVpOynRvNlgqLCDw2u/iEk1t+HRUz3stxdTAZvYr+5gB
iN+N68JfVMgLYZXkVGNVFjhbmoCK1n1Ejc1ArSkU7EleoXowXzY2166aHaxzId+V+mSuLGC+j9av
xeVN9Mr7sB0qO7vSE9PdczMxFeY5/PafW5Iud7JlhPfcbMaFddzXNWFVvgms+A+DBLEzkkZFMugk
By098u8Efi6A5vX6Y0X2A3MoLw7ywNMQszM4nt6RzJcikKvepFBWZoRXZIqIWyi70S0pQK+kTbts
4o+ehn7o6PWB6E+JKnUN9Ve3di57Rbtac0uULp+hl1zZaa521qQAKikxN1k4ru1vvZzW3g4/DV0h
OeDnGOFKbwIzoLtgaFRIgr88ZS7eFY+YOmY6JtLiwF+OmPJFquYS4KsnkW/SJZp+0yBBjzUzZzpD
Yx4GxVhkN7TEK91cA2YtZ/GD+yZp2nmaef8goURaISsKqYqn9Fn6VL//cHncqeMOsI9X/cNkAtzo
OU1mnvBQ2xs3sY3HXjb27XH1X8dScrvSI35CjC5t3by+cOc+DDwhGq9jVLgkIExhlPMvA4HXo7Ru
bqbHzjZoGveXrZkVzrxIo/9zfBzeHWLS62PCAZSkju30GgX7LBQ+gKtfonYHDxQVFnUbMyUrabHF
eUIjr72H1TR6YDACUl86MUpfGdrR+vaQBrfY9m70qaaAjvbTJQAtaXAxzwnM9MHdmEQ9X4s8FRok
YYw5tOsPDXbN6YbFcoXzFLInI6nz2gqaZpFBuyPsDEOruUkb9BOMAOnLNc0PpqUnfxdRzALVIRVS
/syTnlvGINoDfLQjCbAhGIWCV94aKk+Azpd5ZsokMc+qM0r4Ko8Amq4qEVfuckMDCd8gg8iqI7Ie
U8CSlVHMCPAKX9lErbRzeBRoEb4xZCIAZREU0VT9MLnV84foOhfixLmTXWsq1n+8PC/1a8ZysD1W
YiWFUJZUAL1Wvhs+Ksz5NqBrc3DIjn45OTZziqYFirsqBTXC7aRzXqzBKicltkNID2kLRbyyigG0
Le5qD/c64s7VEBW15/EWzcCsHNmcQ7WZ2ZtUNoIAmUqxOuCud1lUKpNBL+URZh3vktLCC04cUSwc
TCatvdinrNmtnEmSiI05I56an0kUWrXSjr0vou+MAcxerBPWDXmzjqZTJ1sJlas6UDAY3vNDweSq
4i+z5zdzuMm8GQG+cr66zfAV8uUXAClM2tp78iOK9w/BQ5+sSvZlEIZ746XVLsZq1XHb0euaI9if
GLkyJ+LPa0NPdJWYeTFd1TTnRV2QZuCPvDSMTnlWtjdKh7blcQr9oQZngikfzhfTvvGTlAIceD+B
E6mROE7/ydwMlvkhHwhIXWRV7xtPxAn+DupKuasnHsXvmjSRTxvuGBSTSRMrc1ScM1L2m3Ji+u/P
Si33WAh981ppvJW2+2G9qILRMYfZiXUC2XKFGk205EBqT+OaNI3Tcpf0BG7WcM8S9AQK6H536Qxs
mAQeynqHl0O/R3yKQvoMjqrSflBz3+FxCWfNLTe7zQrVrhulhXBTX+29PnG89Kj0zMNE/iTNIga3
xYc9xgJ2xAXsHigmDNS4lvbwbEGScBbyhfSitAqZLxyN7bmGiMws+V+8KabjKU6xJZE22U8vU2t/
tePv/P2gXGxj8jj28PluL37CsE0LobLx0SZYDuK3oCFT25JS+Tthq4RwQ4WEbaD2UJ5lA5Yadpr7
2qDfZOqt8vZmf0MIDGxHFDKxEuRyz/DW3msWlGlSTNhCvt6qONwCvcWJ2kUslaKqORWqP1d5zAKD
UjP1lPkPUzLq9/oQqOjUgDAX5GyvNUBhZh+xnRWR1PkaLwrftMn6KS0mgEDfYCvPsmBf6EMMSSTg
0mHLXsMcE1cZcteu1WudtP6MI2zcECGh/CGiiR0VcRvU8xcYQ5pm+2Osr2BnZhFHCX/lkKObdin9
i+QXlftqeuMOmDiCdbUjngSRVhW7xNIj0nQ/CdaG3vIzocLe9GvhAEWF6KmE3LsDun9EzYGm1vhW
NozPl8slxBpslNAdSYcZWu53/ScLzWbL7NM7W06Qr/OJe1E+EqVgDXY45/9mTsvrSBR7GadvffuJ
+3bPH5m35lFnjGRmpFY+2Z121j28JD9ZutfjewkbbXVvDmDfXLUIxCDykN+bL6E2ifvLGgBGAXIS
n86oAPwHC+szTmbeHuf7a/CCt2FyAbm82wv/4RiTG/iBXIpo9/as7qQYLpyIi/Hjgw/wxK/9BSyP
3pGJ9qEAvBTNSzHKFWUkBX3gsKW3lWdlmQ0f23eiIAUkbUWgD7K9CKGd/dydq24QBiS5Xy0hmmCv
pOn5NAzHq3o/OX7RsI+NMMiKfyrPq94oxZQc2ij89JBflMMNSrCEkpF/1BEvWYG3qip1V61856FI
cr1CtPIuUapwRIFQfXN3JRYMAQzpkAtSKA5KNrRoi8Fb2gPs1UF3AGBYUnf4vqAfprx70VC6zKFA
hu9WfkBpr3SnoRCMUbKLAHyQunnU2c8U1/hURc3YKCZD2Y5ISnFlhAFp+NgujHq8kcDLM+vhfihY
+U32p/eBd9ehamYUx43J90AqU6qCkgPYMCQ3CmSQ88MhVOG95nn79+T8X6+6bhGmE1HYovnYaw4R
aAkgmipgoP8i+K/l7iJI1ZrAgnEGfvmts2e6y530z7UZD9s2v5E/h5SvgAZqnnylX2LaqMcTWm/f
jAqDl4TcFr/ha56T3xYBdy3ddmZ1Dp2UHEZRsWPE4ZbVNMcyOmg8/1itOv5qkCJpCcRIDdNPDI0p
J2y5GU+aL3uE2upUuUjIH0r5+tgbjHHXzKYaNuEZ+c+0NJmDFCmdL4Yuf96s/v8lir8mdytO11aY
vMhESBjpCit6M7ITKRmioxUY9AeqyHvuAfZ0H6nr/+ZxaaXcDT95LQSt70/mNueov8vRcZdOJCg4
OF7nDbcH0O+yWr+77QU7qpJJ3dAKzBx5VvrsZnF1HRMOMfhOpF+z1nSlzj/OTDiiOYxbN8Ph9teL
oqfKmA3j9ExNJgA/qcVqNrh6Ctf/s8ANDGmmGUQQVT58r8HvWMpsTds8jgarY+RS6DFXlOWRqRSf
azozvqWn47HqgZejCuvF1th3Ap5OfrsxOG4jEsc0DOB9NkvmDxOlkKPEiYVJ5wUhWqIU57UtxTc6
+thbhPiA+1BUu0Qm7XWQbn3W+4XeXgqbYlMmZ4CKU4cJ2K5wcRm7oPMOAYkXcByMNYv5tL5lciPA
S60eFpLiJ+wSc6xBiYBmoap1CB/CSXnBDZF1IQNdM5jGr17MDQzL6rZUo3nhzocUJsXtOODpKj5d
/ABmHLGLVsKhnBQ2gAZTNLl/3j8e5zUOcxMl+u398WeNrwzigTmp/SO0ASDZIMVC+g4oJ6L0MwG4
hhepyM74exyip5357iXpwsM9LkNk9t7fiH1hNCWZIAY7fkDCM+YfYeZytl+CY0+fNeZawPb5LaL/
xf0323W/ugtl1Ha9WP68QJ/10YMYSGXJgUPE/JTT3WPF8LeGVfvljOq2R+fss5VarKO59/23eqpl
nfA/Dmai0MRnl04Tc6jkD+vR4Sd3WxnxG5UWP1sc2k/aw8ed01DvGsepj+uvUkeULOuxrLkPiwkk
3/87jM4qlW9bVLmAqSF0ASMDCrXbTFFlSW72cwnY66D7zQOagMAsIsBPSis53dhECJbPxtgr+ukx
dgCV9ufTNYWrU9iKNgVECOV8+T7x0aehZU+FjVgfLLl9WAphrI0xHjDqC0W7EiJ96WnZTjJr751y
vd2lE29zpFohMBvxDTEDikgGWgW6kqdTnQOocvhHNzbnB9z3H8UbzpfXLrmjO1cujqBykgTSJ8bQ
xIx2CgpPSKITR/IwWJFa4tReLHQVY+FcUz0XWY/RRCIKEtsvYLknJ/XndH8672jPc8gTlIqldz+q
WKpGpmtWZOzqxhTKFMWF/aOis60XAUDJYnLhqC26hvPGLFo0tevUZAcmMb+FF3co2UmwZzezOcEP
ZoamSQKubOXvnLaWQlsJtQ3trJcIMGHjJm/2r3cD/nuiyuoueQYw7tqpp6Q74yq7TQ3jr9kPlCdm
7iyptGWiNzMCYxkWnj/8MfdY+y7XXo8E/MXcvsm7X5RGHxo/azxwvzW9Gi9N8zzxj1PfVKXwVLVZ
7Aofg1jwchg+96BPNA7S/5PkEkX9fweukk0ktSgt9z+RNWHjEDrVLIikbMdMv0yTKvqxjkFKmNsz
Nbou4pfm0LI2TL2hhMXHId4blQItRtHeaen7DUKa3XWAZOCTgXrF4axZUms6EHP9bndRidJZusJg
FxAjd5jY6xglsAdTRWXAEk6b8QWa7MaNiHEHwBMaZ6JYsi4EZbzg+ihNteqs5Bw2eKbzbvygOjSp
5uWVokUmnfBelf/icbvRfJeZPzS0DLg+KnTbHeU0ADiglyGQk5Sp4mxgfCIhDtf/9/FEic+yhKSU
NkQMqCxnRc0jAhVZwxTH2LziDbc77YmBJJl3WFVN31RzNusmvTs3XA0ubOtKGvItx8WamWeyyhzc
At8BacUrHNFl+ES4PQ6RvQC12fODheEF7rOPMar8cC5KFTVavOa5IpxqNaC0iF3GLLOboyzaoqcA
7bAncBi4TTrK8DQDcx1aNtNUfj1ozMeEk2wDhDItzAzb3lnYW/XNaQGkE+Z6s7GPBphbmjh3DVjX
kILmQIJlJC5IBSzqZzNM07HY7hnbYNU4GiVGkeV0jgJBW39YmqRmrfQmb3PIIiYxP2YxcmXu9w8L
3pJyI7MAJ+dZql+QvPd8B+DZWSmBx/foycjgeizCh+VmkDAP2zmXJGXURvo65k9NAXyO+qRovQBT
ePo2zLrexwoWW317WaYLJDOVOzB006ORXrfe9RIerWHRtPCQPG8RMqZAHIemVqGaACzP2I5QYfjy
wvY5HbuNC1MVdXjO6Ax1tGGmS5Mpd82Yqb3twFsYxAqYNPEWrW7gA4KXSOPypQGGpvvM4ZYDD3cF
3rADBtXSd1weGfMmATej0w9632ILKaYRBaCimGTdxtGpccLneUZrt9+I+OLo9FPj3JS5nnZsYYHv
aMeEOhVX9IVkzZiJJF0C8TBDJoexmGCd7OCF9pWqhLtw1l5Vyjx1/ZRsmnyWeWuqZLSgYMTwe4Vn
Ev6sSxS8xdSXoNGb3reKvtv9H4FocfgNtB+NJbwjZrQNMr8FpenVuEtS52tkoscP97j3E+26BLcS
vMEKumd2E5QDEqbONugMAhW+wrDxaJerCEpLUR+igamAlR56egpJoSQNyp7/uCtu43yYQsI6geQI
KDvvvrcG2t1LdopfKL9OI1Z2fpk2XFfBxH1wzsdxukMw+EkjdwC3onR7XHxUbSbkuN1pJQnltArh
UAmAB2EVNzHtziL0JT5tym4FkXf/j4a977RHbXS1KRcllD8qF9Q3hN9ilFS9gMMhkw2k81yzpGEo
xtVVHIqqcniUOKfg5LXVmVHr5i8G7B+xn39ykMguqKGOhCB8Fr/NOnvqvJt8GAAiLEfwnrhJlhyu
2vOMkpAc2wlbOGlEQsuSroIJPRIXyKodO3V9YRppw7Qd7STylbrCH1GEFo+KRTssvnrauDo+IjnN
q3ZoUhq0RF1RxvCrWikTQQbNWlbedvtptnTL8k66CcXpDuMIeFoccDc0qdzmeiyE1N5HmFDOQjaw
CwBS/URo9BGPDNzd8ahy7VYUdt2XThtRm+Z7z9PMxoA/qxv0z1rt2xec3WENwCeHD84zRXNCnvB5
KHYkPaDInbqxDK3gV87XL94AIyNmStQEj6+4Naj8JWB1IUOSigZRT28k3ALzWaO1Tsgkoowvr1j+
CmKELNhLVt9RSTRqh4CPuFPBotAKptIMU18oKwLHuNJsWWNEalLxqomL3GtsZj7W918Jo0dT2EAw
qoSOtq5R4R3X0wNWJotp97w1vIERGsH/V5ZmG9sZbe7gWdVTVks3aYAOD037sd/z3ujM3/hy6I9+
/wk87gtJz6nZPYsuR6QaJao6etbOMsfeuaZyI4DGa0iiBcE6CG9LpU2mw5HvhxK7+Z9jBN+roNf/
qJcxxi96T42DlJGKTIL/FRdl0osFmdESno46UzCuiztON/MuNp07qmO2g3dp7toEE6F8vFg4M8W5
qMClR7AZJOJs3iaMcKr4dBL59yUB1uxRnLzDXqD2LSc0bfqSURgdadaNB4vggN5HuJ4tfk7lBKFL
yUqoE7+8gUWshw4oU6PooREyL8l06dEjR7DLIWHtlUtx0h5wy3OjYczMb/3HDWxRrEtnTM+I/hWi
ywLa5h55hyY/JmsB3qFmt0v/KqMgMhwwyorsFfSraOC4k9hKTQ9K00eXYGU1tFfAvlGxogxozfVx
1VKl9WKevy6ZlKJUiLMc7XsSFAoAjkXdy1w+I9d+qTvgVMpyioBsTFhcaakwoO61rWNk52x3P/WD
g7rChSSCEjqhYo8xm7rOUWRBQWMK744q08ECJ09xAfiW/iivLSsIRKqPQsgf6d0fkcry/mZwBJIO
FSxXxPLFXZtc7MrKhiqz4XnnhzbXIe0Is3Hqnz8lwAFyIVC4mbg2d9JdXFWxF2g1kmcJw8atXZmp
pOWjvS8eQsI4EWGSMXJKLmWCyzF5PykXvoLsBWYB3h3ONeRCNm09CE+T25ssbKCs0uiceyp+v+Vw
UPuci20fZ8nUoMi/M5NM6CYITKkZXw1dMGgYUvs7yJdQLeaQi/Ghk8YcaI2bhA/SlJyN0sayatB0
865V07YaalusTbhmHSmbJkRu983QBWZ73+hVZGJ8L+EkExmOeO3kVsWJbhj9jIKq2JTMUyGae1gm
E/QK1qbwqT/6wKIIvtn8i3elgXNmYwN8cmskH6Th8/XxTfPPnRgYMOStHyyxA1p7EX6ONgStA9xO
7yMPe6fE06OXSUy15Q8i9O7mRXSDs1brhEV3n/yKtOCmevkp/+HDOlwqx+if//lY4ha9BZHbcYvs
GSmfOUpei6HVIGZdGN6pWAXS3gVtaY7FHcMpbVLsio7eDn04v/Q6BEv+yTcL9UxMfmZhPJiy3XpG
jgaE0Ujq6swAYdv5AuDu5NCd9rFX7WDywJlRKdan2sIXe59U/JM4A0LV1c0U6DlsZ/RirdWtjt9F
4q3L9ESnGS9nw5ZYsUtzBHuPU2xRlp8KkjzrbmX1G/tZZDkZ6RTdbW7k/X3v6ZOoEhnaplugXarn
lx8NTzcmAyNlrmTLwVf5HkltHPwW9mTqPBkW/usqu4hj+7KDCZ2M5+sUSNnlss4eyJ/+AiV28IxL
kcb2NqH1sz4d1lGezipDrQuWk2K7yUEiGMdiXpH4TNCdh86zFt3NnoOxOASXLsFlGW72lJB77amp
JJLGORVGOcxo4Z3lRtaLkdV2erLqFEwkZfiiytbdDAzB+7xDQ20GwDfLNrn2zjfVak7Hzb6mlGEa
iSTcq0rzNVPRT3NrTlcSPqIQqO3k1/Kn0qUzkL/w8QqnQ4OxzRy2Do/LCHo5yB/hOx1XIvMlqqiW
02+kVllAa6ddqOViKedoAKFv6mKxXeQjN0f+cN+zswKpSdvA3YRpQz4k/EJDQWE95rKeyFAg6QWz
BqIvTFd9NNy4HQFSBZ1r4x7/UNRJX8VdFs45qDZuhSw9YSTbuAW9MvkMNhmLLlWg7zKJ/jR0crKN
Zb2M7L1PQpr6ZRh2GLERpE1oakosUn3+T3MFk7lX5JyrXkyajiSpSgYY7FMsS9zbm8tXbgZQkZwK
GaKPsKMf5MCMHjqVDAe0xIiNE7HMP4BL+qeMB0LRatuTKj462ni97U9w5Tad9D/SCJKSNtJCJDyi
Ie74W0JfjgBb6Kmi5i+Ta42covHJVl23enOEElbaMzIE4bMa3k7clxg+jTW/EbkYtaDJv003EuFl
ZS/sy1VBb3YE/D82WywJ3hmgj0O4v+J4B0WWmETFG5UrY7lWZoXSIjAu7Ak7YgP1xd52ZPSn9Dxj
NN0MCe0hxfpl8UEFD1CzAC5JVXCxoRnYm1wJLyVjUeHSn9GHwvN+TEZ0Rs4iAWLn5iFZ+l0Fsi8m
/4OxLiX5O+A40hsx5d8RF7jzcW0cTtTToaWA747LV8mUy4Onz2EhOZpdkQmJ1FeCb5xuAZGYmKy7
SsSHhTKJvV5QS7uhfYjDXVWz8bnAcDu5evoYQbOsmeKXHe3UIKMOhpFTdfcuukSpW+OaTUQWtRhc
FqmbCAv0UdLOCBTNHAJZHOyqqL4E381kWTR0x0efER7ErPb6oG2GUY8FKB9bOGNvPUGwxF5pjj7w
bgb1sz8mEYHCuiUE06Mu5nPBxoPMITVfJ12JsLEa7rHSPbE6euZiKPH1EoxkG0sqaPRd5e/8MlrN
bCuAXCCNy60o+0KQ4FQvgaNJquVESzNCRuOdUQNrlrje2IqiTDO4acio0gQsmSInj8W+YYn/4StM
G7Y9QUxxSWfiUbyQKMyWRet269Q6ucmllhz5+6p3uvyid6PstUuMZtTSMgWKK+ID9uv18oY77f6d
vwsv/TTG700bRllBuVyu42aeE/1RF+xWDg0u7rVMr8DrNc6Z38D8dihVfG/DFSHtpO56uqf2pf+O
7EVZ4kJM3NRqOL8MiiQlMPbNfdcNM2wRWEUFqZtXK0GYv2RmJ3OhiroZFVr4mNvnsHdG1unhDjqQ
ZBuyjzneuHmI8oo/gqR17QkC9J6psT8Frpa+Cf2Mb9ToxPPv2yN5pdlAE/Xwj5O/DHhTTn2YXYuM
6Dp9thMAthR9OFZzaV5vnUoO6a/TXOCcyeJlZo/hBLwY4DVeGY5MjHt0yReMu/ZaemRSh5nqfggT
Mt9AIQ12AnqfizGBoTYa5eOSsv8u+3NwS0FKs8KWknmwMPDI+3/jZ4/0kVY+8Ta+8c6d/e7m8g3X
VPH5Q4Gy9C4OQtPUwJFzw0ygYmlDtv3bVKrzO0LqlugIVZh4CleH6yCSbMJmtZH3sib7vwOjxd/U
FY2DVDQkU56djtKmtsBt1qCHvZGoLm5AhEEmK5d3dLN4eRUlM+HMOEVQVdenia1Uln+/vF6yPVui
BKzeU5mpW3I0PFthas7kUgoRcqlgdziAY7JG+WjMyHmp+zkNJpwR/Hhv02JnMcoCmRtk/ZVp1u/O
OGmapxmok42ADca5NaWs5qneeOZni3d1U6mPzvdhzGYh4LpomKNvcVCQDAUlbKTx8PQoNq0bng5a
M7YbCIS62qR77tyXr805FPChj2olqzmNPG0hibm+IAfqfncEY4V7ZE992/6wOX8I9GpRyPJaYbFP
lALIeJC3yBLXqv0gt8PO0wQgwIsfx4I1Yy2a68aZgUiREu/22BXm5m40ZK+EbhUJJ6rICRXCX7E2
sAN5RWgOXeH+ON/yXnyBfxZtySkbj4jUSdqBT5gWHYFyBX7xrEEyKPwW/DS3zQXVXfSry0juLnDk
UJmDCGZnh2lm70TwrDBUu/Fe/yynZ5h17dJXXqy3Iq9VSrtvHaTUDiF5WR8YdYFNTIzf9Gte5j32
EgXxAQCEk02YzaM/hMFcZkLd+OwC/P9gKSKJ7/SWJ2SSoPWJ4d1+Ui6cqAAlt6XdWndGJIdsAmoi
pAzvbSk75Q62Gx1EZh7hfUw4q3Rq1LxFnjzyoh5kP3lpa6uf12ipD/oovNNeG0t6vdDlCtqBOVhO
8gSpkVEhWb8Vj65PfSxK5G5bucJPBO+6ANS3jgzDZ/vkNFgoRv2T9aP9UVDvUnHtB3sr6o1f1MpN
F1xkoT+K0PjugqJAuQsW4lTqhmIdGUtjnWQ5tCIV9SegxWcNLcS1YAzg47rKL69czJQOqCV9upHe
U2No4WB+SYx2XNgTzEqyh3AFMBmJod+EGJD4z/hOVfrEVO9DjGdclFQ7fYe514IZdmDe2nqGaOxw
f27wP8lNcwiSmcSVVp4kbu6pMSWi+vNDPsJG/aHUWIhwKBQ1iysYZf6+TTS8ScxFdgG+s2qNg9Ti
hDyIE9WQeWjVVek5YI78KeC+qpDrGjvdKldp5i7kDZkAgWXNy8NlIF/h5gieUEAhqGmUpEFbTbaB
7obcvcg/0SESDLWhD2YnlAfzqOjxNkq42sBX2mn+vesCrI4GUVBAy1x5NefFeoDZ4p6VyRwMAgr7
bXIYFYvov/9FgSvIzwsS4Lfxx6DXYPRpeDZ8cC9WbzSvXzMKIRMYopMCI1yc8l/w5ySCX4hOwCWf
xZpgcDW3Isg+nxx1Sc5W7LLHSRam5zxcrTJld5++taVzBbsOeb9bvfGV89cs/vnmGYyc0ozSdkPj
F1qE1OZOTAjqWDNezefcWBI9mlAOnS6rME4G+WCMP/LkLRBZVnz5yczSI6/COxfR2mKSHwP9pyZ/
sEm6Nnv0DAgiZhlOfxn2Hd/xNd/ALIlRRFu4VeQqeop1y+th6CugwiiIvay3SIVwz/wGhwl7MBCI
IWLPLN0R8UxyzgUdMoluXG0kuUI+TULBz9a8YrlHgydqp3Y4/C1KSdso81PxvRyDAm5PeQYFYYee
Y2uCAfnymY5rH+yedEaOJp66mvUZjlkG/enYirnNFmb/OwgBdzpXqXRH+f7RcobwY8paQmSy398a
vRpW7i9VtjVp52vjfKvtGzuxRFi+ZS6c7IXZdHUyto6zzw1oohQgX0DmRab8CNkyOxFqxf6Qq+0L
Ie/apVEzjV4cKZhWVGyzOsKW0paDOFXtURK2su3IiOr4bOg3hkQCOsVrO4xMsOIHwD256ewtGPUd
dXD5XHBE8XLw1Uio9RKeaziUVL09VqZ9B6Cg109fg8WADUAl0HwOMYeQRShT0dyFrfZNjqXrRhA3
LXXdnonb9sIrT2OE68dn551sQS3nGc1419fq2G/iO7B2++L9EEvRgdQrl5zqZB7Mxez9NbiKa8Dd
Aa030gM19xEzUtS8SiqgOCikQpX01lEOd7p3uqWShCAVlOT/KzCd4gE07GZFn9ITcoFGQ51V2+7n
o7Dwa1GjULxWQAUBCOiwfqfDVQLb1thczW310M2lw2VmVbVCGKw6pzzcjN4a0DQkF6245sEUkh01
sAnzbPTiX1JZvnVRgg49Mb5+nvU96FOMoLqs9p1dVlklCFBT3JvyRAePXHuBb6/53le85HZhpY9A
EyEB/PAP88fS6FRfoPGaHr+vH+3Mzkoz0Ognrm4p1ts1ZMhPYvPKPRQOn3OQdJldvouM9LZs3Wqt
AftPVkXpC3Zuc5xsvEMqtRMc6gtOmXlSnaqBFs4Gv3SA+duVHFiGvtfls5vQg5k50z49hjFIQ0Kp
oAPXEO//w6VEgJVSo7AHRLvS4HCEWMYCTGWwXJ5G9Ll1CinBgB+TuvtFSr4ahzFmtBEz1EyEoe9Z
5+YtDn0O08r6ObEq/LiuviSoNGZmMMjNSB35DgxbyJ68NmFsu1Ow9K3AB9+zywbGnpLN7ADp0Nck
BX0cHNaX/RMavEKkyLc5+fhCXp6OVG4u/D7GbuHKPjBi0VhUM07sHqF2EdXkkkDm7/Xy3m4po7mS
ZtNo2pa/5Zp4ps3SZvmOPxO96wG+vf96ROhvdvoyGMF/d2dM8NJPC8v4LijIYZ7kgTWcwVtvgPC3
Ozvq7Z64StuEYINdc+Yx7jPiDGvtMKy7cXK+HUq1rszYzpyDLJzWFJ9xBvRY+qD1Yd2okJM5s72H
2/NNZOnKz6UeI8fa3Er7za6mM9SLeaZTQ/SfevBy21tErGdVu8s3wrvkWK07BuKZ93VVdtcC6JMX
AN7+TMj3eUxKVIqYhniRvcRHeOX2KFcXLUUt589JSHqSEunKEBJw8FAyvXzsoDJjjzB1MlsPWWuI
/gB6H/rGS7aeSEYeSmS8UWF2F/HhwxsVfAlmYsI2akwgjVxt+C3uRfi7k8/AtgHgoyI291rVSAWm
/7RasiiXWxTkuFpBIvIdsCt+IRBhP3+K28uZz6GMRm4r2vW7CwTsiLKr7SjGrPx0pCHS4We5V0sM
yNLYhmQ+QFinRmkoqECqJnb4aaaTqgfnz5cU90EPQCM0mayUWeLWUc1hmC2eNJGAb3JuauF5uG6k
w443VQW/Vfnq54bZHhbOscJqiXKyu16tQmyKZd/3qr5G5aJcej2u1u0l2+liBFboNCHorJmftdKl
Qlp138AI4vZd6d5hXl4Pyw0QvLYu3uh1BIr9aSBjYzYGFxHdf+g4G17IIH9AGnElArwQ5KKF72Rl
ulvuOT43kvVjI2UTw4CsAWHAQfctgSjIlTf86Tz/kHo5/kOUr6wrOOXNfi4TjRV72XNd0V6szOx0
U+37GbBqFXY1Rh2wIwDbgR6frs0jQzNhXMC0wRFTKumZ0ThiVjsw1deQSpjQc4zD9MaQ8bVhijzb
zpHg/6mZFRMcrkbd3/Q7JV0+e9CQdG8xKyea044NI8Em9oBLTR87vQUrur7reD9TFjI0MDsyp9nk
u0UzWCvYJaE8kfY9c9Jz2CiL0Z9eoKJ0PZ/e1PXWYZhV/MBV3W8xbkocaZFz3BcY7+3Z8Ipb1oDy
S9qHy33onNZ9pS7CnXqMc9oVHLmwDs4/KyCmitQpVLdUWPDGqGMZaVEzCYnMzPCHv+gLEjyn/UdA
XyALvpcPQAnfkP/WJWPCDrS/p9m6w3tu4WR9QD0NXGOzmgF2rS48O4fQMkRIWW4xkrKJ1ng0E4ri
4QAZeSHWAumWmMx4zu0btIvWgjVh3eeLbwVBYCCKkz42inOMFnh2h/m1rwA/C9MYkdf97y9Vpvlk
Nn0o1R777lrneFQblRr5adXNu3BlCWZBDXiEUJnGJP/+/YHLaalkGGqQyd31QcSSoHqS9wi/IOoq
petbqARiPMyUVqszemV9qtoVW+VbVRjXMmdlG1ewgQCpV7KyBcK8ZHEmkimxNHSi+khLevmKBXY5
oFOnaIT9Zg2oLqP1CP+AxK77nKxL+EtBDvGwUX0W9bnvaYFVvLoHCOXNSxCH+ji0mPr1wVXf1hAr
PHIr5KgCAcioZKXW+qh8D80YQETpOwTBIXzH5TTpWuY47xkTYWGwv749jMGTf4S6fLJVN+IR/FTP
LJPioYu0s7sgd9aAXnzUzyTctKFV4ck2uMtywNSqxHBgug1VzwudqIxDukjhGseh0o3BuNzoN2en
e8KnYB7ztUlz0f0ssRe0vFrl+NS/IK8vqtvDdQ0ZF0WH5a7R548fytsgKkjxuqWN7Fdhb5G6mtlC
svJrt73McEkeY4kUg5SOonpV9qG5zT3aYtD82Y8GaoO8gv7S4/0QGPf4fbCff8zWLaGEJG8YEQ7x
HZk4PCbCOtRcmUGypSGzqBv88B1cUe0Pnj993Lum2muWhCCJTq3kl0kMlfglAP6Efav4Svi3578Z
TRNqr2mf9PNMjI6A5wIuHa9Cwj2VtaBWlRpeBCWre2YnJrpsJ+Ps/UzI+4cFoh4CQUSsSt5ysmeT
9C+KVhnlDR42XKpPeGy4197ooc3tKjSmYWQr+Hp53KhEc6cmoNW3loMUpDjTeQsnWxpi7y0l66Ts
ovD7QtYBzJj4qwlRIP6lu/92qQ5jjingm9n4MEZt4KRMPRD6wjLWtygTEQNNIxK77ol5STPqGS30
6QkdUl0q/5TMLknmIOl5d8bziXjZuW4FtK2mHfVJnC/XwxT2MwBsp5tsM2dGZItgZ7QauYLiRxAk
Ku/iO+vhRSBlS+A5nr2QwlEzpFrIXsc3GbdZXkl97x5IumZglF+XFbpbDC6ncrx97tlGwMFAIhFe
l824TPj2wzBd7aCfuQviZ+tvUhyE/gjEwArHTxApxwBvWavrR1LNielTSpTtCpyAUrg4H8KARZXM
7ey4n0GVbjLzmtCxUDVfGcmkhHjNnZ1T5AfkO4qaLzALFRbxCyL/FNCExLr/wYCNNzU6t7k2lYVc
9nTxt5VsLSPJZ2+ituAWpfZ9y9ypa4bbSDlYmZ5/tTWFuOF+5cAUcHFcIbo3NAda6C+FFXAl6Kru
GjfOAYpRqhPusoeIpym3wNyjhRVLKXUIxt/+urcWdtanRUc6JnGRj96laL7BuG+hf218Fr+sujiO
T9J1CmkIkaa2Thrj0kLFuIm/GO/+SbjKlRkKL20blCrcsee5FybXYt31IKyeWyR4c1k5WSHCW7tO
SPkxLnVa6Kg4YHrX69721YG5rzhVl/QTlNmjez8EO+9lScrDW7UddILaprUwkuS+wdVfH+7JrHDn
6fAFhj4RXrvbLOTXcbJVL4VHWfKFTLSXniA32BecAAt1nS3+awyaLedO14F4haM3mNAaz5qxe00f
4xaYtMLP14beXNMImC7vPsJKGNp/aLfEjYNfy/Ld5jvEABWX8GLeFyBEF2aOzei6uzBDi8kl79Fh
YyEU+8P39QuhLylWER6mfVItDMORJa0E0cfHZ+WjFj6gi4ib+nZYXFcgD+JnWa9/SxAlrCMBb6kb
VNlTv9CfZh4zbIgv5/JhY+qG7Ir2Op7e4e13z5MRcvdXt/UbH9AsBf/nrtRGCIHTPMXqsKfzSv3n
A/i70EK7DGXEm3w7IBTTavLHWXivWCLll4XqQjzw+KfgMfag943BNz/cZ/IARXdDsxhaeeeThuYT
MQ8rPIJlYaHrZGokHammN28r4usO1v2GafD3+wsz438jGuYSK19t00SmB3zGnyGF6nA5OEO1LDqX
v/jvY6DinyZNFWUydOk8UJOm3wDiq9TbUoOuAx6vq7uO4nhuwztk9KqGA1A8CeaWDkKQu11hOdl9
WEL8RkfTuZO5kA4cms0OdxMiDn0Pvl1oEMwC4bhyQIGL9gJMJjWF48/2n/6o+AWsWopdqEHpvKWW
O+ZlyyjwTmunMdcouNzORv9f6croq7so9qQ9rFOsg+DHtB/PP+3cbKhZeBr9Ncv96HV/LIk136eu
AY/N5+ZpZTFdc7x+TtYcFpH9Xu1q9tVzte5+L+ER09vsExDzq0B2eOl7cGcVvXVMJNH/+CkhUEHp
Fijh78kHLVjNY6KwS8CJ/J4MP1qvt0VYsNUajT9+hvPQjkm5OQAfkAE1WuJvfadY5UdgIJylJWAa
beYpkPgQda+4sMaTZVtuh+vGTeQjLvVeDBI7TyrQGDIQrcHhpVG1O1OMDCgtClXQIdAR2qqZ6l/Y
gGYlJWvX2o0TK/xkHMdw/FFoOq3PQJNUcKIr74fMzD2Y2bToaTsZl/COTWlMH7qOh67+whgJSQ/X
NiieTz/YTDglrLv1ng1bszrchoOwH2It2r/tTiSYcuMHh6pFP0763wnzTBvUmNOV+yHQ+kqN3Itb
bGFNRIuDFW6vspwiHXLgpCBkFSuRzz7Gzby6/mEQYOeGiEsK7d90sTiNQOIdxXmeEYo6Jy7shJSq
Fo1PutTEOuF9HrlQN8AXHa/eS/ovBAuZrWr8SEmK7+e5wNYogiXMwEiM87SEM54Ckr1ksCTVSJDx
7JciZKMGPiMi4MGjFCq9AspuQzGU+O7d+0dZSFAjvvWT0pd8L49a0gH1N0J97MznwI3sZtqVopyB
6VRLu+VzoD5vUm2w9arvqljp/cJHu1DlyzT/iDmJ0L15cQkc8vjtH2aPhKk6YsOGwXnT0C5n6MaR
8xL4TJ/v/gaFR0f8soJ8YUVpwU15c6IF0xM+3KjlooSuDOcbmJeiqYXOxVwjIQgR3vkWIiFN5pgA
ECznWMjJHVs75x9kJsR84fdA7LInv5BpEnCtXoeCaU/zVBnl7iwBXvvjhSyJ/zqHgdVyfth8u+eV
kCt8tEmmQSuyJKk2Hp3OHla3UU/raK09L6yh+ekweye8wWFNyottD4BT4EV2/cSE28m0K4wLJGvs
oxZVDvd1lzhv0SiVGldUgcf9FX/FikeB5ErurXGszR5WXxXq6hPetYZHHDmXACsBzDluq6NlhslL
x95nvk3VdsTZpNz92y3cpEkTXRD4SsBAzHIPuGTmh/96lmckBrFobmsj9VA+hchWkCvK8axx8M6X
YAw71Qh+ZnNk9V5aMT+OhQkQ1RpnrzuRneEnH2cOP0XZSn6Y+phjAVOK9HpkHCS6XZg3XhnlvtRu
zbn01CMGXJ/WXGMvWKkL3pDYPRsW05ogqkwH1Dmv29di7oIb/mO9uKH5GJ44y2WDga8206GsaJby
PiVz4UE6yGXVzvCZKggz7wpTUW09LjN7q3yOds4NcsNrJWQz4pc3Um2968ZIZfer4FS15ds2bcBq
5ZK1c3qXe5wHCASFPLJCdXTQXWY7p0K9TvAV8QUGIJpLYXrO4CWVImAp8Bwe2JsTfxRnfWNqDDLH
QM8Kgl0xh1VkCxz0/SBxKnhHgwQWlKFjCK4F63MF6PfJ1P3Zm50pY3AOs4Z88hDdHQaGC5SxicUy
Qlw8eT3AMxNoBfbJ6PCLrYJsfVOgAGohH7c4vw98qgQ7P9Xh4nr0kgrXhXpsu/2vIw4OiujUAiAu
ApDQgo7Ivrmei5/q3Br2C+Lr2OVmGgnMeorEs/eeNRq2w85qtuX3D69LcdtdW23XpiYppnffy7nB
GUchseL4PoE76zfDPh+sbUGPif3LZikFz+nFa3MINwMuCf1fBjoJ10s/zBMN5DGIgLroPUQWKqjE
dka0XOzK+S1f8J2jnjPEgY1gXDwS4EUTgxdtN80VMIa68tO78adwAEicGn9d8Lk9dxdxhbBbZDay
xX6/1eO6+h9xzYSJqF9uir0YiJQo1CLPjZw16BiM4IXYoYgQFUgJEmHNa8KvCchmcFWQGAL4Nj4T
OxNNKuE5K024+X1wJbXyy1bmIzC0yDMk+fNsWUo3GobyiCpiL3yXoAkGKG/0IpOG/W+VI2HHr2RO
QZH1fwYvASABg6XPWPZhp185x3HOyQE+y6x1o9gHJEwDcbibANygmZNfGWzlO0k0fdzKQqz3v9KM
9agBSjLvvLrTa9bbMhBKY+zERZwBVtdpgZrWwgoU9QOGN/u2I0LPdzFe+4Sgrs9SW9Ve+sCksBXz
6Tufe/ElXKcm20tn2k9+1XZKwxAi0sf9CBRB1Y2mC1tP4T7c+wEdullpBtNEZnl7kkyn1qAyF8AT
RvKhGb43f4PoEAGq4a8O4jrNIJx5vM7o2mt6HgCeORs69+JVT4UE1qZW85WMPk/rW2riQ2Hkh2Ne
lqe6k4OuNi6A9bgO7HZk3W3Tg3G1bi26RfmultK65c3fABQ3d/cmJZ7bbfse7YSY1QGKBBZ9g47e
XW9sAxGPLGCsIehhyM0iegnPdwhVVeOWeMZ6LUf+cEczsyL3RWV6qHS7DjTw/r8ZN7Dp7ESxKEgD
6NaSsAUaCmnVhdvEYWMmc1Vm4Q/fOlJWQvHu4yPdHmTp7Ec0ihK0a0LzHNUhfKUUpQ0OJEzZrV55
ZqYIflSSUG0jvTLCq4s8OSZgujxuzSklNhmRvmoYj15d22KzsRN7/l8fxE1uR3X9nIPyVo6fB8+n
dRLlj55RrcV6c4GzG7bOdWtX1n7QmeW+QJHtXzJbxe2He525iGULeXssWBIRoKm4qzxOjE/dnG3S
v+ggD0mTMMB+9NP2PZXlhGubpfg0b4keNj2i4S1KYPCaPW3R9e0P6+WjGkUnrGqfFoUhDRfrBWpe
+MsfgfmiYvcfjcnKSnD74qNP6bAnrXOBxKRgImf2betAE8XBf0CrA0+Pt3OX5soMkyKx0HvkXola
ngw1qiFITzblCrxx1mOAPQVMgCqV4LF68mTiOCRYOColb6BfexROe3fHZhuYa6vmsosYmYVL4Ha8
2L/lY6nZYaMJCv+VJzrIsgFekBc5rnWOIO3yage8u1hq58mDaTEY8zo5SvfvSoikRxp/KoqwNv+O
nVcMw90Cc9EjF1+xu7QOehnpej7Unu1srX9wbkUgVK43qdemPL1B06fB/zqYSdykQ65g71HpIH80
Cg8dNmXU1TOe5Rf+V9AfL/5vWrPxO0SKH5Hn/zCjmcHTNWkwcWCHixPSO2Aid6R6JE/LEgWA5TXB
xlhgccDQPHFWPlsONAawcBmxb2nlZx7TYQyPzFz1yh+BNGsYYVbkPVl2Dn30uNxW+L7dRqeXVbPn
NoRz0Ai8Q6vjCi3Fs9vGEDD58gJ1dCUMNPozACyY/1Vc/54rQ2nrhV2hRP6LRXKY/6S/LrS2jWEi
O3XjAQqSJBrdBf/m//WdXlJqzbXMPvm4lZbnuYLrOC0Owfm1/t95KQ33Gk6tHmVLG0Lt5hACQmu0
z9JzgQDpyVT9zPqp59snG2Yoba2oWtlmJfF824iM3XYmqpLLg4ER9e7iVGy8ZfM5oRSZgtH72Z/9
V0yhB2bm/z1IOndeYUhN0POYR2ud8GrwI+xd+/mvRZBowlzgvcWsgZv3Zru1c4Qmq1SUDQvjVuL/
T2uMW6WzzYGvGvjVauHtOYr7pLcZia4rtmY49Y55Wtefpt2Du6a3m8J1ECMwk9f9jCOYpPzH89cj
0ymH7q+2TeNZ5PTZLf01+GVhhxT5As4MjG8QdrqXeGwFz7PW23xOkExD+kPWTS8Y+TIY+HvYJ+Td
eAcEWsxt/BnoOujDivCs1+0edzIzsWifWOKtX2q1OdWM61u5DxUyb/SVY1xAONkggjuo+ETPzZ6k
ljXn4As74lwVx3SES1CZuqZGdNhNrWGhX82ZbCt7j0ZL28EJC9CHPE+ZuhgN0C3qA8xtMLZTBXSo
bWMTStUmujtM+nYYAciAAUwzkotGldZZKcE/kjGLr84z5DNQcqn8Oa4nU0eMsOAjIt0F75Ebem33
hRo7fLBGgKDT18WN7AMwfV2qOv/uhJiuTjuNB1HLu7O/eNM1+DTWIQcpEo85ujZIvqxicb8BZIS+
mIVHwNb4MuFdCGkFFrQrR3P6PUtKCfVIjjUS9aMv/tKOemwk4J9zVwHuAL5PsXKT+J8DXH8QI/TB
VlM12PHRb9ynGN2VNETwvJ2u6qXmDhpKbdPm57P3ErcOmHq5UPghu+ri9qbbYKH3TqpF/HKGs3Lw
MASxty4Cmr4/eJJnYRQASu0k4HFpry1HfF+L+RL4lkROLj3ViQHErD7FJykON+M/iE8d90yV0UTD
ffxE/etIJqsLAeLXKHkvVZ8QVg3AZpal25hBg0gjTnogu11gOkjpNI2SI+Fp+SHJsBbA5L1dYjIP
WkCxqD3qipOnO6oU5EMXNvsnqNc5hlHbjquxleCbTH7o3zr7dlj2OU2du4czQXEaFHNnAc0XSgrj
DSAveVbhfqbzai8gdCkVRYGvOnGpchrghOUQeSYH746PCxsgGbcOESNhNSX7MkxMKwrHxOGnTlUy
92h/1zUK4Ozg8y7ApQhnR+hmcgZdJPcyAEQHmPgdfZTW2E7YwIa+/fLAg5lgCJwgnOUOZUgXL0hL
YxYfb7/NrYa27P0L4j9MMpkguZZ1GUNiW1kCm0ENYcURMtL8UtKR7X65A0D9CPeqCJUzwit8WN6T
E2zj4aT/TaG50pmTj/0xpgUU5yFxgzbpmXsf8iumH9FOqkZH/XK79ANsKJI7+eT0FY13sz4iHAW8
9+cQTkHoh28L0Qi7PUQYNXdA7cc1kOU+pYyWrnRgC4EVDV8i8b7fJ5s8p3iDxxHZAImcAwAwMiAD
Nr/NWPVkcukKSvCms7SVumXIt53LPUJZPyVuRaIqTTJeILVvTirnTTj4eSmo/tLSezU/NXpSCeVY
/9aOiRLXkyGjt0/+ig5BRGjqGep1Ms2nimgEY6m8ws5ShYVxJutoW9/0vih9QKAml3OH+SvSsAZ3
qU5NYrGxq8hk455tCesB8B9M0dFgFpDfbWhyU+DgJ2IR3riQWTNZyzWgcd4q6v0Cr6tS9lrc5lmQ
X65PmMFYuYFtivTIZrA0LKMNtUiEt6Z/moh2izS8vqp0F2pTmLvgnSsrvGJX0K3DktDnkzTAa5cS
81Xvf7YuJaaPTuG5Dqo/QJb24aP3DIkZjF651ddfBhe+v3/0GSD5FZNw3mLgMf9epmwEB7kSLIJ/
DGcrM259cDIMDAQ2/hPB7d+GAifzR5YvYR56mdpKxF6jHYO5Rt+U2H/Taw1BO8bH1NfefJh++Rvo
XVseStCX/GCQ2MIwHrccq5azuGO3rnAfocaZrfgl9VKr8ph+zkiJ83vD9J9tsi41icyx6l7ycV6n
GpiTpAkATx93N+boYdrQ/4Iz8Iu7GB9ajpl+kQKQuhnJMleoR9aQs5WU2B0H6qpLJSst4CoX5BWG
fGlX3htVhVh8Eel9R5KodBVWVSkWJg59GTUIKUzSb0S1rm9hHyqfNsHZ183KbP3kMBCpttAsEgBU
WhCo+mh0IF6A0PBhm7sJigsI7i7EYhTxDcD4sdeqvBytD6ME8w7gXxrquZdBv+9tV8NJ3ccCdEqF
dPlO6QXjQ1+wwuQ1oWeVaZS9dHetYtDjmZywaV+uBqZLi2wgWW5gV9dpwULDpmFWegt/ef04gt1u
XgC5on48UdH4azGgcIhEgNmnOSBhHE3rgPqlEdL1RD+xR/EZD2Bn/DjbcnBN87nc1B2IE0rbrVaz
2WyKWQg1fdldQzU5Eqz8iPq0Ht1fKieMiMSTGjsJN+TJ763NhzX9kUnZN/T03casr4WXdB7+6Wpx
Ep3Ekz+vUj+Q/25C1jt1wqQ4SoiGZ+1hiolae4efaIav/74dZYvBUBC+LVAhThSdibJ327b9aIap
76OFZLaU5Rd6+HNA20hGyM4IyTObELzfJ8PbV4zI/auV1IhY0kTvU/5gviN48FiHD/MZHBIPD8LM
ONO1oJo9zknqq34vhAWTiQ2Bx+yEKJpGFaaeJ6ygVrOTJ82KwqYAkWRV7egGdT6kZhRa0zC1T3Gz
DQTNJk6Iaub2huqEZb3S0rtPxM+F+Yp5dC+4B708M5sdT0in+JgCbGzBcLCuDa5Ojw4rTVUpRxBp
80Nh9qMZRheLwjsSI5tenP8VOccEqWubS7fHjS2lG8rYafJpXy51jmLdwkIg03b7KrJCf5IeNJHN
XBkhE9azRTq+kCtDXVIfhkWpvk7G+HDgSRHVHhKVI+0XkqB4gsiJpq72zxq/lKZjLrVajlcBSFwn
vUj06VHvc2CX2bn6Dp7EmK7HmIjzZvi0P7P+jvMPFw7Ki+CnqlnqxT8KfXRJR+ckUlq2hRyzXutb
nh5aZ04ULljbZx9kSuUnGjOlpmlNDjfVHm8RkVwPqST40+TlcHnIInGAR9GgBFOk/8bU9kCKJmF1
Q5kFanmGpCIXYqs1HGnATYK8Q5HtEn1CZr9zacbfohv0gAZYri7UsgWmmLc95nYGf8Zask2yvSYt
YANA6j9Do+05h6sBaTRNlmgh+4Lcf0ur9/wYl2ZpY7l7X0WFum78YB8rUw4w9Yv38KnPSJWt5lsp
zfyPwqbEYkWtY7kFVnvaWPsgi0jpq2BpidjIek/dvNiItPL14qVKoG4jnLVaeFz9o36Tdo/Vn1jg
smWZNvi6ihnWrCFwZioBGdc22ssky8/FRFWlOVmVByQAoRBJsQuAHQyQGXn2nZNC8Jp43dzWL2N/
6Vu6/Kx8mtTpFWEDiAr6BkUQT6Z18gR0pjYh7a7MogJbXznmg40EefGq96wmM34E72gsl506UdHi
NqtI3nWmX9aB8pKvK63BG3KbTxdtffKjPLRvEkfwvCbW5L6CHd33rIcjzrmMFt+E8N2vom62ds4e
9XPandr2IfeH0K5rSGMnMfLiIUdmSOAFRZX7hcDYPG7ZH/yfzecrUk51Gw2c2LO/CZTQPWzBDT31
OGhDUU+BAfWQsrbiDBikrEoH26xW+rW7bXNTq/Ir+LBG7AJyStDtE9J0LAIfJCFLSY5JAerthZyG
9g9osZE2qZrv81iezW9D4a2si+KN/4PV1/oGXOI6Z3EbccTjATzcAjb0/BCmLMdYlZ7opBpuoKV2
Xk1rTSxy1JA514kuCz7GVNqy0qMG/Xth9uw7cwDkeUEPUWVJS8z6TXIZKT2dL2I9POLVwxZnzmWF
m/ozt9lxBBJSQRkUuqAT5n/h1MKNsd0u4PJzIEKRbz2L5KRKvU8fPKNluRqHo2/8JDvsbToTce58
ojHNKvo0oBPODZ6qJvnZX5fmi61sr7VY1l9fq/QVR7JPpz+viE0w/dZT8AEs0uBe+o+A2J6icH9o
2UB4UOr7LizvbDTX9QHhpE9lsaa/NAmN/ynXGdwN0nzwfSbfsIGqBrE8ybSuGO+Ykf1xKq06k4rS
MsgEEC2lzx+a0L/FbkjcCHKBrsmKGvsF5fanpB1k2TM37npVdUBktBOaHEZ/U/WMZZEoE4X5luZi
FeyG3sHUpota+4kC3Lf1+nuzbwhWio5LE6VCVcA5r7Ac2lhNLJRguoCmLp8UAHyeHFKp15J1uy0i
0/o4ob/wraTBBt35DRJr1EpL840CN1GJ/jj55B3nSNlXVfVVRZAaB68DFkSCS66Xj54k6S4e9mcG
4Zx66sIZRaLRKupbeyeESgoecVfavFtVR0RErAbGrRUkdTniCb2+16G+hai1Z9J6C4CChSszsNm/
jVP+GXe3DDOPYSC8naI9pQGahY0KuK1ktkDdW3QLQSYJvJXkdC3ULjE2XuehCj9CtzybD2hJOSQI
Hi4uDowXhoeyD4grpqI55A3HqCChPsS8/sFyE+Jpw+x0K2PKkjk8q63IA6WzPXmzgU6iz7smj3Rp
A3AtV635scTS+QyjR+UMKrFx8jqXf7E4ZK+fHsDSRrXZIEKoKQo7sV16kwZAHFY1kEbP+bLJWaOl
VvrwNrB74k7KnwNPXqidUoXqGtG6NrWi9fjyxSfLiTlPiJlTuv/3VdcWlk8SPbv4zYXbBh4O1eCd
5Z5ALkdi1ld/ne1JLXpYZB4key2uSgHTjL+2X6J1Vr+L710Ezp4pk+pHJAFXaLUi2Uvgxfcr8vUI
BaH1809/za2rlFlXMPxaVjKYU0Op7yuOLOHfclrRM9YJJ3dh0fgZ0AQsx287E+wFTcBRhY2dtS5z
useVOmK6dFgvI669HU310Na7spBuOPEM/SraFPoOmX0m27ju7gzY62zGFBdjbmMzTNABqgwFgvzX
5asj6GFwyjgiwoUNMgavHXKUd+ViTBYPnOCXS5+y+e4qpq7YK+9IHT7lgZTezw6wMmxENZQcGaBu
KrGTIBEfZafXjtgV6NHM2U+o8J8Ga+jL4DTzKSH2cmWLVwCU5/XNuHbcpcOVWPLkQmAz/Da/Zenx
jp/MMDgF/fBy/aqJynrZvWjw0OWRXVqTipvImVviiJ7/nFg2A2WhrwVbUDwZkFxyuKNrwbRMlyDw
PgirLUKtAl+F7iuqj20vRlM4FuKnlKLOv8BcyTf/bmrIBLVE0HJ/z3dZ9SXtqkA2UYyjkczkFHWB
RhPc7k5/QQWR+CvZNZvgYK0r3oLD5V4/PfzyTN8b/m6UC5XiFvT7V0epccBxUVRjXyf6qy+Q0XoJ
DbkCTb06tclPUndxnHEuwakJxhzvRlUOav5foV2jYHu6Y9ypPUiP6aTBcJmSjUqvydwwcVLs2xEq
h0yrQ42fUt0wu2RMXweGgWBgWbOv88usRsT6vtQDi6ZQu/xHt2tPuVPyiH3hab0b2H8H+X1liwXg
cra23cgaD3HFyqkUWHzpf/OOQ0SVu8islv91IPpVFWPx98fX/UGpid7xEIXUe4y9usT+ZQiBpAGg
3iOBTZkMTgCHMzKAQ31dGGZcMM2Bi+rokPXcq0XgayFqio2xpWULulxQ9mWDIm1zFGUYVJDTYA3+
UWckdsANJic0/6YPmQJ0O45BrXDqidHmfejoPWgrKcv7fvWC4003GgSbvkD5Skr27iBQk+3DJKBK
K4Bwmp9gRpwe5XbIvAKBkKHdSlNdyO8FhD8d5O27IeQHXQxdIksmjsVvp/JMeljG1dGUVmA4tVkk
VEzxKfoAfKnsUnkfWjeVIwc86Pb5iW6rN37TeTrOifQII6RQ8grauV4oywtSRzdkp+/xXqYLuR3e
EDmeUvewEwc1dHQbD892SIGn4UjmWA35es+WUAFysnApvHkVqlHoMwJ8DUUenBSL2QfoZrED4ogm
cXA8ieckNL3Lx5Yr0Dl/vGFUTpfFqDny2m2RylQyShUO0eeuy+EZ7lDS2ths4xsJPN0Zscxetv1z
xH8MVUH9Bd0PH6JKqcaY9VpJ/ywh+w9POmHyJneDEJcS2HjWJRBzIiRMxBx9m65H8iFy9VoCwreL
HOQzHti+4wotM6fO+hCeJADSkINWG7rwg8FWzQh//6yfAuI7u37+w96rtNSGQuhUOlXa3sx7sTjW
e5L20kRd9R9jKFN5AspFWGVxJWu3CURkOfnPNw79RHPQ+IjlZuhRK5qe/mo0Zfr8V80nqwO5+JV2
0hMA70PYhawMLfnGETcVutw/ETH6NShtwsM4lvQGDKMNkw6W1gmSwW4iWc/WjZrCm8yic0MC0eOc
NxA2EUs2isb3fqz9Kvq7l4ocyknrnBskdKTBzZGUzIptCD/R+pFH1Nz4kk9HR5AIt0qqDv+kbsFN
SRqmt7QXME2BI0OeUqfO6IS/DUpFGo02VC0aqJ27hWasG99QFVayuZRdtvUL3KJBKLyzTtR+9x+j
C/HlFm1hLvxzbn/XmQd5IXdZp9GfAJjQZ7I1ZS5CQ09RqP6bTGvB2vAjlrGScx+JnRV07nE1m8WC
OS53kN3XjEYDOy5lFfBpeBD6h3qVCjOjB4fjNdm6DaK8IthebsNiDK02IOW/ApIYN/U5WcvCZG8x
9OcAYGY+4A2nKjduCh4zZ2Bf1ZlVfoabTbSrPqmOlBCBI6KGxYrrgHnlaZK7OhkE+bH5/LnGp6BP
klT8MwgFGgN7hqSvu9xfy24mSOgKXPhtD1ubAxwd3shzt3s4syI7fwoDbydheNwFi8oiT3qukIWp
hH0pH+D6qDWfhv8QOBq56GPMEZRJSTwcMGYEhtw+2xc7JIOBnj1vcq/m2YHfYNmgHAbtft/SZO4p
ouQKLP9gUpLVqRLjkejOLUIFfXvwYW2zB5EHS8khqyRn1nn8df5vIeDkEqMOr8tVwDHdQuMpD6wi
cfZXKzIrAsza2xxgyt+Xc1fDT1ogDyxS8MdM1zpj5dhya8ujQLBQT7+8QBn7JqUvfg9IBt9PHHct
R+ws4xj0D0QXB73TSjxcBugaE2tHBg4VrC0I20dj+FSH/t26rihC2pZ/beGugvBgwNdusBuyymUE
UXBx6LCX7FQyw44oi5+bFvRZZY1xMhS/o4dI85peUiLBV1RAPHVAoG0nUuC6YqTRTS8PFhTwBcZE
2IWuNCWei8tGUuVQ0oEDY/1SjCwVSVChv51bwfcIgsjbRuk9FE/KPt8zK6ha6bu7bHm+ei0Si1XX
UoBWQpkV/xqIUhMrlqGt99UL3AApdq7EyfZEbNLvXBXT2Mm1ePOkhPUAWLu9gdZVz668r9CtkhWl
xxdxi9GKFZexpziboFIolpRWilu5kCPvIAWY7cFbEJBwW5HNsX0ms0TdWXF4lhOca/hha4FOCSS2
3QaG21P1r2FpxbHaM8Y+t6+lNlKb2BZMPpyGtZqe2jtmAycBfkqkgF1W93YTmgReSgDIjM+zZypc
hN+4kRwq1isD8JCn4qBiy4xYywg4bZKnaZOWvKXw6yjN+buIpiIlPcTyhUne8vjkVJQe3/WS7tGJ
xg6aQxWOitI6wJT9IRqGnM+7WBhv+BITw6omzlvV2Ie0ywgprQKvot+NDvwG9qIsSI257Wyr4y8S
U7mTweq0K/AHkc56QKiIlUS0BI0qiFMxyMBfPOiF8QTF081CbxqJXvoA+2r2caL75VdSYPhmVbKU
F5+vN7JhJbAg74HCG1JT8r62O0TLeCf6ejTmyErM4c1s+f2xGGvNa8T102Ll3N7sfIU3KUzFCtf0
1P3+LiP/e5HoHdm2YK7LhPuvzs/QiN80l3xeAw9cyYZ82Gg36RwxniX6YJ61PWIloPozJBB9Nh6l
xEFzb5W/MTC47OCGaXnAKIISGVRKyW6cB8yqecy51fNAN9LGYuhnV0A36rWXMEdjPMw0o2CmsPZu
fYClrYLNyF9Skc/Fn7mjQo5rnhrOn4Bm39chVqUOZm3HMbEGjXEP+ULyITxSPmeZI3YfY7GY+zbz
xkIlFxr/QuTQ895rQu/uy8G9xFi2cdKHetnutFrHbAmGzCp4ilGCXjlvLVxELuF0XOTplKoxHOvL
V0F8RGbOZ0SyDdQOc00YVXOBmYpgoVx4awzFZd6paq0CAKbhTnFA0BAHWeAQzvnhmjICH1P+wgu6
J5O8bm6Lqmc4caYDdB4y29jQETF9SLgMqB19XKS9TAmHf5A9w025L1cqNGhNrtyW24ddQJc/d5+U
UGdpXJV5FxRtTtNcAVr4B3V2IqU3srRFICxPUDRXeB6zb7UWiXymPP8odfh2HtqHWaKNAzLAbhbx
f60yIwquEI0TbZKHXeZy+kP+rgvtY2leRRdW3qwhcEkffLoYG85Imn/JXNjbKNyvojQ7BA+643Hz
w66+5FF9y0KTdHffsXlPqgslIrAEoHo0ps1m4DTuvtr+01kIJkW2iLzWX83jKndhdKexTOA/6v8l
fSGTvHJLOpfiv3bvOqcZPRBBEK563Fo8YP+irCEh2gIRmLUKUmVe6wxoPtkfXVy5rcbWGqW3k0Gi
S0h68msWTyHTxTwP4K3+w+Ac5pm7vRPChBwznrtpugPkG+7onuCctNSAANtG2P2bf4ynlLvmiXIJ
/2+Rz9J98oh9i7uCTE3v4cIh/eYipovq5h5lBA+X+gD2Z4SsrHEqrDbATuLlzVaxZBHUMHZADO/v
sH5zwR0euyuptk1UwrkKRqR19OSiaOiHI2Zj8LQSjrGbTlmjZxpGqgsZaIZtvT6S0u1eq3pdnl5O
+uiUAMz3Fzb2j8Xmgol0XzjiXfqLS2yV7QoOjgwWEMXMXn/Vr1iGXBXgWLSUExPhUA6QRtLugrz9
utwmqmDbygNBz9ytOLbpPgUzYj8JpFXwe/W71v4IWjVDSUeSBZUwlnxr1XkMUuQsyxcv1TCZwCMu
ht3j0DGDdVsD3xnj2zTqWo35MlLUBtdPcfWddzWzbgrWUxIqkCT6FLz/0xIbPyWgbLpugppeIv2o
x10GAfnEbz7cZLIClW9ShbiGcdePy1paeRDFMMpEi/U4Dd+hhJqAnhCehRooKt8olxwih9D0vrU8
P9Oz6s9ExFIsc1EBKcs7QEXMqzVl8RX84HZgHEZFjlnK+k3SrAEUilglhaIWAO+uJDULnOAPEoZI
zatUt6melT/zRXaojXwAH9TPL6zA7zc13OhHkcGmoYcwtlQFJPbnjablCNGzOCi0vYm0jAFruo63
9y8id99cSc/YcRgeYcN9rnPVZ7QCwtzFkV4dPfIzc8z1AiV11xhIylFS5QTJm+yZ5l9vudrxO0D2
OuSV7t/Lo4mb51t2Mz+zLdcPAvDWI125ffVQvdPtiClYhugFCJ/plp2ZSkTTqlhh26/BYEZ4qbrq
6QuBP5NuCpNTItK0zqVfa3RP3tfTXUoh+7MXajcPuGtbg2A3PDN5cKeDw7NUynvWt2m3KTDVEV6f
2lx98XszJKsHGdygdDTfVkwLkE8tgB9U4J63eSoSoLsswvoi7C0K+cz1W4ReQcs7i7E52xMS/QlD
cVOyN40b6iu7w5lLs9XsK0KMuWb3/lBkGmRWyUM0SvuhBgf423xX9WAuh65YyEJ43kD6PM7q+xjP
ws5ea/fMBMG3pMHahBx+0nHmHzfny0KDMHVPuBGZLuTynyFYoM2qodofNR5k+b9u7qbATTCCq+03
h5HezSNi3tcySKEka7COg/oFnZ7ttPFLLcww1B0YoJqMawpBm1XYuzs1F3IT9PVlCn8dZ17DgE3X
2bX/uJ8SFGf52BQDwXZArJlaFP/rm/UpPZrALvnFnXkd5nGDJVwIobkzTKaRsiIay4rbtUEslXyP
4vkdnkkTWeI3PM7JTnOm2wqMdCFlScKvtOYOaIm+d4kLlYv1MKeiK342NTzrBW8WmkjSe2CmNL3d
mhN+FHrd/ltTILoyC3ul/xIQiLLEJ8E4eYgH3YX3gfNZNMpHVBM/Q8NaerKStNCSanNvyCroBnpa
8YL1dZmBXYuKjSa8fznEhDnpr4+91RHkuEHGH11RK8x3BWpkEGOcFZ0UAPXcr6VypNuhYA5m+48L
DeMuRXe3p26Kw4a9dB1QsWYJA6I7eRAyYKbM4wAv5he1zNFgwRTc69RdDeE0N5LqdOxJvk+a4wwh
NSAOkbOVIxL0d0fOfkpaeHvPYkdq4qNH/74wXQTVJ3QHowB/X51vMF5gzMog8VdR5SOXkjL8DsUl
pNT4p1UH1ZTIXDKTnobo8FP9W1q9JpHj/M8Qq11AwTgudUsB2xASLbrdHW3EsWfDGPz7j+wSG/bB
S90J1+7LikrmTcI2IRWHrGIDQR0vUrsnP9oIHn407mgjvz7O1pXpjygmJpAxf/8u3VTA2KigLnc3
tm8YWWy8eTwkmWr21FozAeUBhKrJ9NDrNxu8RHq4ZAA8UWp9woiX5b2igYOAV1k69dknTaho14Z3
/n7DC8LqxZRZGB//fYHRoYGh/EL2VCuWzBe5hfVJw8LDqhCYw7ByxMRPw0Bc0xTpguZk/Rzvnr7w
RooBkIh74nly7j6Nwh9sdCQ/lBpzrTz9YjYWJ+6Nrjt11fH3a+H+UPj8I2PfygZwh/R4C/VJS4Ci
FNu7QKSalwM8E+DYYBAUY1CRC34iJnqEor2LFkJ5nUZaBwJ1Msw7Xq+j9Xg8fAmt8gRxYi2yUm8i
UtPaldIbMrvK6hcoeQvGl5W0RN6gaIXbjOyHYQirOYmQLRBioplnAoIqR09oMzGrEabCTGovGqaS
X0HheQUdZuq3ttTAKIxEwHAfTkk0UpTVz+BWk4aDr1P5Dpzyzno1m6ohS/2wvtYafBl/AxWE1grC
0awPiiUFDWsbAX0ekT0yVLs8JEFrrPjcf1inthvuQcpP9KZZVpKv0QMbOkbJZg6AcHvGBei0XfOb
W/cnMbmnA3SYPxiw1j/tATqPQ9gaBZYUadmgFqY2eUNNEN3O5Tdbw18ZMou9z3ncOkmtNd6bvob+
r/lUqMEJmdjEMlZSOAwc2i6r0D9uSUmkowWAg6RxGkKZKkiCU4m0iPxWVd5BIkq9RszPnu8GMYpL
9R11BuDDnOKmOWhv8Hc5Cwkb0nUizM5EDFXb094uDuFlV71nU5rfbaNekxF0Tl2NAUWqzcfPHNM0
U3M2NPC8zMgaxFseBiArqY1u4oowMXeqtX4YJ6z6Yul7S1OTGU0DHkmauxWwZIbcPNeb5bqyyMLr
2S6jHzBRJbdBQaCyBk41WTVSLrh7y69Pe3/S8p9EIuH1YrgaQD/FmsXcb9ElnG+scz724F1TJZog
lXDUxonlfb8+WHNFxvulbLs0VPaEkP/GkA3M9RLwTjZOrU7dyIOmP26kH75xeO5EfLKWzBM87C7y
7MoV2bFIcDspZTk+KbpmAZbF5GED9m7exwQLhI7+X2Hnf+2YZSyLT3715Ud3TdK+hO55dlB+Qqqb
giDS/D+IYvXNScNVB4m7v1janCdsrb3iknkY/PQA7xVsd7tOd7XSal536ykg+3LB7+ULUu+NoyRG
JZVDB1yis10phnhkU2t67R6r9BzJZln2nGzDSfPFkppxVLacdIvuXTcLr1YTXz3kM3vyOzw/rjA9
wiBOuc63Mq9wNArJtRTRiV4aTmCSml8wGQcm6y1drsLSatMvQ7lyTZjWYehIfsodKUCkkZrW3qpQ
beGuu97vDNWpf1f6WmChUoPmJUIpxRbJqM17S+t6gAaOzuDyDDwKJMzAF0DtXv6jDH2W6ZbUrOCB
Xi2xNV2GuNjCG2E165r4pHa7MEJgjFUW6+Ha1NUA4dwbyjxDnOZqigN+0j+0bpvj3x0+su4ZlLWg
btk2mVyxVOJQ+3p+dzl40pXxg0nqVlBpde7uh/81P1cSdurSoxUPwrS8unswgfPlwnDQENYupOQu
G4osc0EkffkCBDQcx59mcJC3Z4rue04tFCm2sp+PXOyWlp845ixmwz3SOM4SEQqYCFh/rF42kz0Z
9fSil66vFiG/dmfegmMaRht6yWh3iQnX5ZT4p7sPXw7pmkB4ZiQmnnGvO6T0qkP1NljFaLT5d4X5
pcMr1TjuyjvreLXQl+gL2A3Y8dJnlSq70Mu2tiFD/BDRuh82Hx4MsQm2d7/mQIsn25bil6Z82wMB
aMAOg6aZtoRJ0UiVebsCYT5RVB40xRfioZiWxs8wi1kXG4z/mfo8+/UnMzFDmCcZIbiQ5Fhzg4WT
QlBQV4h6nHiqfq7mOmZjG9upMDE9TDDU4EAP5KR1VEDywEH7HqEqJjafEg6QMDZ59BHvJgq7afda
2O3XYJe4OaPfyxwmS6ltmUuzHp9fXQb3FHvdZrMCo+yeD82fWbsC0MS2A8H86WuZ/NPNOyWS0qH8
jCLOqac4izVkOL7GyOXTnFCVqeg3gMM5JQX5WE1L96ST6AB/dCYCIUCZT3qtPeHl8fP/7Fs10viS
QHkm/T3Z1umsphHLF4dBtoGdn8z62rBFDQ19MyajR5z8jTooN15JkNJvSafD37MslfqQV3wxwz6y
O+e2GadO/pSQVrLhCC/8rqBttPc++FvzVUKzl35YIssusBmoEt7dBkSJurPFFpen6/qawAvIfgLv
9OHEHSOTzt97h3mvevC6tXcRm/tpHkShV2XaLKyZ1a3dQnf56j5za5BRDjEKaou/REVT9ljwjXJr
P1pudectoormVWmHWEfgD31djAx0fzsWxBL8KoeseP0rKFltSf2lB1X/sWOP6+qd2Rl2V+AklIKd
KKNzSujW0LF0UMKL11SUID/dgtMT+AWzR7lK2P4aPzaW24HpFZQ/GQ4AU+fUEyj3V3MKxK0Lv3Pr
AW67C1M6K2EqCCIXjCK0FGQ8erWw+7Y4D5eYI+AemhsCoWuTs8vnscnwU9w3+CeF+IDiBj9YRmPR
Z7pWORNq1d2JvCOvcfh39ejMu4I81E6zt2vvc+ZZAtQL44/3cu46WTIy5C0wM6ExQLraU81/bUBZ
bENwb2Mb3V06Juqzz2WLq45d3sm5WdoeQE3Rrh/q0mpJV6sZ76dCyDLYJrwSHtYCOL7YEotywL3S
WVCA3JYXVrZgqrl+FUYL9BPG+8UMRUdDoWnkXG7PXNZ7WN1KMa2xlX2UwE+iKjg58kRpL4gnAh+P
mNLhtTdQfHLrf+4mi3JVZmVNjP6vBpoeuKGtGRdSdcXfJ92ht2+mvoz9wCpOQSofZ8wKg0toNDeA
RXeKQLCyPvYkH1Wm0HfHoMFf5qZJyAxUV0c4bs3ChxdcZTS3Q5AUbxZ2/UNwcQ/9abdsKEPlEin5
n/gR7J/Y5Yp7PlNoUvz129JlBqAV6j7ciQTrH2qu4Mk+3le8sHX3LjPHtnWSHiP+mFIECeFvomEx
+ykonbMjKH9vlcjzaseWZdqZb5SD9aEZYJj9SKLBvPYApXhWiuccsuE3PVL95/6aYrpS77et11Tz
PSiWz8XESUcWWO1kctLkUp+qbQ0QJe7JCdgYk8BvGSBZH+H1Uo+Qpvm5Sz6AGjwZCTvylInRlnSQ
a7a8PECjrilXLapEu01PW5XsRF5b/U3WTHc58dNR7JR7MpLY1MG7mXaruEEO/0TrtAKkphlZFcj/
5t6jmHFoa7FqusUdVPPcQLYaLQHP5sdAkyaMdUumNRcXtJ2S5hOLOyV38n0kEpR260EDcaeyOXNW
0KKHxGz9uCYnGBzVTRtA2yPyJ7GTjjLP6dxraBrsth1BQ+Ux2SncMY9SwMiMEvLM44cdU8Bt9utk
ISRME79VYrEPE21HaPXjYFvqlAWssxKRUdPfPZ3xHSL7rZXJML7zvhH1cdHkCV5Epy6KmMWdtRHY
rF8T1Yp2GGJUfgB75sEvagFC7OuwPYJa6Bf4q3Jcu0ZyJ/8j0xDNN8sgEQEUgnOxhkFjFxMhOuCT
eXjvmPFEI2saeluO1g0MdJY+Dz1zu7RjQaf9Z1iAJ7r07iCO34uhkU6XVbyJJpQkuItmKT0qweMW
j05Ytla7eRCXGxXL3tbvbYKSelw8H6g9hPqBmSjX/ZQEmEcYAGch8+4AQ+DZC0Q86itf2MqGVEqZ
5r1DDid8p7Bbyh5NfH7khZ3DMphl6JBoMNdDCltMuySzOpgvFRbgHFb0AZ61dUsdW4d9Ucy6IJkV
KWwCZuUDq3E1AxTDGTHFDNuchAbbTm0cxdI0+K+rNDa51J2jQjhX0RbVzxMFVTX/3TX9ipKgZI7O
/3oMbeKL5E+YThd3IAHqPPZD0n6gZXLJRnN2pmnIbfo5fS1lgY10VdBZmFHCTb6RjoLgktSiYmk/
GTeSKwJ/kbmQINl6fDWscbMtrhDok27fXkIeJ99MlrvLyWs8wqeyLi0SjCbvqrzsumrmtRX6hG1a
4dxoSOHZaEUfAXHqhLbO7uSI09FkH9yVYeaB0aTdPz5QR1BhBXYteHy2NB0gg6g04S814RqtH4or
OGMiJz6l4hl7O743Ip1IVNcoYmizoL3ewH2Xca5m1Lq8iwHt1Kfo2BHwLrsNSB2GMn0LNHQGMK0k
MyM382iYbIQSnW0vOFFqc89PiHmipNu05yFbsVDkLOd73spD2vAizGH0Pgp2ruX7wkC1+O8MzwYa
lccq6OzM0Bogktfa8huWfXofJeWiGAY9OS7b2p9xnEUiuAKk4zqKg+rGgkNM8kwBzoOqdErlekDg
iKDBkBIrkxcnEYtCT07vkNSnnYhw+OIokiZ11xA4PbJubQVA+n5vKlW+O/Xomd3UhvMij276NNlm
6jAYKaQ6mUUKEZTER9KxdaO996rVhAHcXx4896rCaCgZP6tcxu+eOzLrgwKaqN5qZUfYq+eoB8hi
U4C3vuGDLul+E1yRUbjto5lsWtgcA7PBz6mE68z47e+uMPbwc9vLFC4vjmpZBuHY3XawHcVEaFsk
gVyRL4gYljbquK51FSTHzFFP28AqtG+f48qx0SG2W8urrzObr6eMfNzPZlD7ltgdxZczeYjuFM+V
xBU83XyP3xws3/D9nbkGETt9SVdrt5+0n8QsS6QA8Xr/9A8welWlp2R+7qokmASxEh3N/jTiVz0o
vKfG25+n8gHatkVAqmzB6X+GoEEtc/7G/yWVug2LfEIeqHJiav8z+L15MXStAk1HiEdGKABG6/Qj
0i+p5YqxTPhUn2LedBoqStI3HaYKn0x7fdZ9U/iektZVLinqrdqTFy80DthZunnUtjL7q/StPiVI
y8FkINj4flU7QmtG8AQBQIzVUS0RnNVXXpvN6AKFGzWJnlzefwD7xotIygjTwOZuplaHwIDsa0ay
zgOQi0j3o0kQyX5uAUP95+HgNf9s48xuM+wC2zInYEMx5VZPzF36jeWLzf2CO6SzQsdPzpUukhFH
+AqixwTeafrrjZtr2TKtPcM2pztM1DhQah4ZDJlGYjT5dDMoNpn8b+c78m236mPpdYBoD3t1JYIB
qGnpDVApNXXw+SrWViW50yVE3jYCpV7xkAfBom29YuSrRe5UOI0e/zvZzzkcUH7odc3FDn2kl1Qu
gMA+sKmCoV/jsvB/bGTejHiHV7s300BII1L4mG5Qxv+M5c8XE1QAzdDrc2k89TZe4a4VuPAyI74O
rEHqg0IvmmC9Vz5gy4Gi7/BCwU9FJaSsuLu/VLz53BbOrJuDQw7IOB7ZLWCazIq4Rc+lK08GCDOL
RiV2UczdNrIuZ9ZGUIn8t+XaE2b3+3he8Fg7391JDzWXEG8feoCQqD9Bul9DH6rKV8isG6bBlrTR
Q7KBuEmHRrUIwd4eJohdZ4dRxse11dBQ017t0YUn2d5CqkFqggLbT4/gforAV/f5LYYZcDU8Kr4P
lopGzNdliJoWVxP+T2Ldb2IQBi7ttd8CwlXfP9UR3LS7eoyRJAwGQvGLkaTFsK1IevKO68i0zHGd
Nt4wM2/c13nK4z9rirX0dZ3fbuGdinARSIF0n9N7qoN+HZYSoacgAVI2SnLKpxmq77c4HEEQluUd
l4NhLLdA+VYpq2IY5FUQnbRIhhJzcE54asmd1Z6A4CAMsem2snLpcvwLVU75bTwlptA5/xiOvfQQ
iaFEA69IaR95bMQTnyA0vldUntpxAFNmHClR4lCtdyvR6lBzNgvyhod8bMjny6aTi4EKsigwIFxk
Y4XX/kUdPvZkTXYr3mI8mBEwN8ZkIb1eIf3OHDVaFTsPIWspVgIb1/7JbabuBautkd2dVs/z7MPl
oFFav4zMISZyJWtKhAuADiGUaq2i8UlMg30nnW1Wk28Zhr9iqRUhCeUG+pyagABcDsYtHKsoPf7M
Vp/F9L0ZPAIcKvXNnZQblko6wIRe68idTzAyQ5lQf851MhWcvuHF63Rv4jtIDixvT5u5GbtiGhuI
ciZD7i3Q2WSzfs5lSMcvDc2Z0FwbYpiaCi3pOwbJymZk2jiL1JtKnszZ728qrhp7jv4PC3qKxHG8
Y/YR/ImLcX4pR4JeuMK0kC+E0RebrVkMzF6me7G7YfCZmkkNR/o13ZJ3w2uFRcktPgwcMqa6kRPB
mtVe29JH0V4RXtr52yFCYOyqVX8AMgstZ/UYHdGASfuO02eUXNgmxoIb5SwqWbr2RjXoI7Yr/4o4
RBgK2BCsnWY9UiljvTOGtBGxeVX+S3DJfvwH1WeIwYDr3T0+vUv2yrpKkZ0XL+Jh003bO1rB++Bd
/FMbMZYmhVHKKX0n7gCxCzXWJ55cpxUVW9afmNNNxDR1w+881LqiHUB0NIm66cYbBBj1IJH2duQG
mfSv6P2t17iN0BFQKdhw0EMWTzKnupLfS3naERr3qmQFOG51F4tNWuoS+M9WdZPGQfn/Lzek9hWy
dC+ClWsn1s1kpyVUL4JxXaymqeUlp1x6lHnN5UBpY23nmxnKrvQTlL4Hg6AGgWMQGNS76E4H6wtn
cKLfxSOgs8xhKMypaAFjGt93af8jWt1pfCrP0bvwcjYtD8T5yhPdtZvlqPPOMx+P5IbWRc9vzC2u
PGkllcIIUgJn6VxoqTayps1Mr9aA00lKeyB+KBnCBBqYh6YwtRA/lyp+DAKT2HJH6iR3ZDJwtrlk
oGTkS7eKfJtmK7C3VvJteXaGXZZ6pMxY7yufhjXXuzs1+nYmeFwD5KlYWRH7qfiD9KGzydCXGuOi
74ixKdYWzGK/7ZPavmMH6tDGnX6eBzsmgd7ogR4mZT50ulaaT42/tWWJ+0FV6ZgfrhQXNm3j1wCY
J1xcuT9+GABBEWUGKSuHOY65yO8bE1n9TwTdjPxNnPDegxzF20VPjVVm8+Yq4hiRF7WdIvxUQ7dW
J4114PbZ+9bz1fQOtxn/DL6dhGXmIn8uvLe+CL+2XHnPCi60yJKwV2DBSacFK2TqfL3ancWXoVBX
tCpTA/kHZiJhXueBSyWfE6IkdFz9T8jdHyTWLMdEeK4lO597Y1Ztlo8qzcU2Ry4wy7/hgO0AjPIp
8x+m/hcsfjJ9uUJudIEFJR/HtCUsUFnzu4quQf02Z2lPC1g9/pV3Z4/L3/9lVowyOAykknFmg69p
NGihIQ/m6asYOyctqB9Ws3L0+JBp3/kY17swmBs+yAhgLMzizkT7DWD9wMa20PykslQBfB+Yp4He
iK4vplitLFNPyrECc7gz5ho/bextBQ+xkXJ/LyCsargibnR5IfmjMgHOueVx5ch0AV35np4ZDTCw
eUOktovGtL2Sb4YflNmv/c03CikWRJnUHJ/iCqyDvxciboiesckJl5tfpWWWOXqYY+bHKBOPic0E
YU0ZgfxdImBMkaCd2vZTtRMtrbGoHi6ttkLBzHYKry2uOyP4ARzIlf9Ds+FLY1VXb/+6Wh0SMjJB
x4f6p29cSviWJslxw2IL066u3Aoc3gZ+/b7mQ9MwTqn0edP65iiBHWxyWZNYtSL29YwDTEbAEZK0
fCufxoVlQbGI/mstk3fImkyryq4De0TvMfzXeiQd/9qtLs0Pm05fDeO1NySu+Ucbn6kXi4tzaqeJ
KHSySk5aWK7GQ0i9/LlZBu2UdvSAjtUcZ+TQ6snsGmJdaZaDJbNOjX+lifLouciMP0QTIUJ7EGCC
xP5OdoWW1VkGhArZwqzjfaDHEXqm+2CJ2uvKqiWq1BKLpJUdZxuYshAElZI8dxKSZRrNFPnkBYL7
P+urg26Vq/LMaXAXeXcuVCKN4qpJgOUZ52IktOpK4hR9I9Yx3eASgzFGHt6BaCAtkh7sHgh16SjQ
9Cn54fVNF8PzkcFmCDddN4ZrkQTpORSrEVEtbF3ykVMQX3kD9/pF1eWeF3dEn/aYIKKfZjzGKZ1E
rEKdjGETNneO00hNixI/o5r9NAKagUySaLI/0phtewyvRIhxEbZhJXdCafu8BEP+XhsVhBP/KMbM
yOQ/zvXcI42YNEUdd/VA11wQdLMxeJYnk+sb3Fh1Cfp6btDGfXJzkRo7iSfw5q4+l6e17r36FfTv
Mx7JrPm6k0ng1WbdOc+qAz8vDD8Z8y8PkfXwPtJ/L5JtdzFLy1OoSFTN3NY+bSRkJfMtWZ1Xeds/
reekYlpFAovxRksXJb1MFnDQ0hvEbjFQ0hg9XUVo65A2H4/ZDas0YJw+jIQ1EmwxiLF/0sItcYSg
Y+2ux54QsKrM5MksfvgYLXKBfJBiKgduGK5/TMI/dMjTumbt5tLQYT2nKbR1LPRPKKpqBkzqtL7F
M42lrXhMJVN/fYxLEXGhz4OrvOMkDAYM3DrOS0tFtVdDxA8FH64ZU1Xl8rKS+5Dn0lxjIRNdwstO
a8HdXVLfa0FM6aYdY9+twPk+gj+ZcX6eIj3cmM0Kv7cbtH5NJWZ+cboTgDVkUFqMi0ScGaK38Aio
TklxtLXxEIVRr30tfhpL+gKkq/JTh02KOC53AvVsoEB1rjJjCmVsJ7lBNObvuCoNTisrc4wBPRV3
3LF0Sikrrod4Y3KcOdA4f805fPDJS5i5HTX6peO2YjqG6HUrzslzsDBWXOoxJZVqnTi0DVyesv96
1dnXrpKrC5oJJkm3UFEpl5HJ+eNaG6Zx+zgU6Z8iFsu4RSwn2jB9ZJw15+iFFjnLpYPozdzfeOYQ
+4uechjuG7Du2WbE2a0yTrsa/QvhFMEF1SkgFg6e+hXuOiY/B9voEVCGVDFZp61SsZA+TOvtoxcI
Tu0IWON7hj4LqkPPtRHJy+t1g3aV5H5dkpYK4DB7wooZKn9TDeYpCW86swMwTkK2DlR1gTRkbvTy
lLNi40U/Sfj0S0UPZKuR0d4udnt0Xift+oNS8E2dIEC78lwpqQyEbhZNNxqZXC/7rDdEk3TZROXY
IsSHB+2aQM0jmd/BwNrp1muOTraokOIHJ5jjF3k5c49SSEXVUe5pyt7wG+WvJVaKnmePR3swgaC2
b1k2j6/dr42gWPw2THy1NIgm0w4qRI542vMVmasLu6OlFN1Gi3ZsumpN6XA4tKFzzppbPK4xB2JG
SPREUrQa/zn9d/xA7IQymfanStyPM8EG71cdBgqUED3aCggDrFUwn/OyWnyiCQwTbbvvRSxnU773
nNclea9aO9BLQ38vxvbMTHJHhdQbaucaSO5z2e05CI4a4tgzrFbaYnsitzXB0tQKFvBuMSdAcF0Q
5vqv4bvCCyFCO50hIwot3++pa82VTOnazZ2IEcmuwWMK9fxWnTqvFDlaf4sW9HtejZsZDsSbL8JU
tHzABkB3qVAwgXkb3Tlb3dqvf65Jwm1Q726j24YKig396sY18q46hebgLN0S5gpjiOygpfLYVePZ
w8O4LuVVcINt74ost6ZBbrek2ipNWIrr/hAYIa2AC8T1TDbYrAxU1C1HOYQ0HYhZFSKPg33TLqX0
56v80qH40DmQZ8PPIDRfMB/Qkklc9nNY1zmL0ae55n4Pdk5X1mix2wqhZPdsIOSAfgpW4yEd7U+6
yaKT16YpK0xM7aJoZop24TK4z2Uf21I6qXHt3USNMYgugBYBUyaG0v4RyinCETSrt2BRV152iUf+
EAXCyCw1MwsRDg5eN0F4b1/z05sd5ixqFebF1jFH560CIfngDstA14ZLXFwb66TIR9o0nmZuuKoS
YmnW/FPCRZrjhR6+nrpRzZvZfakbPNoJkoJasYEA36R28nPwno/L/umGTEJod8c/GzWNmqoKGOkP
GnxeddV7spV3jqr4tvi8IoyiLMzaVUOA/GdMJgLuDi55xcAhiYmEblKcLyooz4Iv3H9XRk/ZHELN
w0kBE88n7FkBFu35cVx2sn+t6QRgd8T3zjbuyaGQuXhGXw769ydt7vzBXIx4N8DA7vqm2YULeMOB
N/bb2ZoBwanhySIdmZSugrKI+m16JBL+gXeKvqhK5yUQNs/nFtHvCP4fJzu/O2wIJFZDuD3NSZIe
k167qhPLr2S921iUvj110AeEB4QxBWDATLUjKmV/7UuCqTVCw0zibm0/IYUkXso4XTY9qlPE++Au
UCmmzCcrV5AVsJyCSYCCTwNgWJCZHDL9ItVaGjcHp8Jr1FqGtcQ4dvcD2rFLQfA+S9T9sqkQubDo
bWEOEM6tneqC7r6bZjy3zNK2U7QeThhF1KG3ws8Qlrgk3C0CPEbYneRTaZwbi4FNlkdG41z1NeYB
G57sl39w2BtV2nBp8AVEIYE5QSnIX+JRJFe5WuaeerHn8hm/awuTWxw64Gj1Z1FwV0O6q2JEpjCW
R4D9NfRNHDI5l1TZ7xI6fz9LV/GO/VyjRP9yaQ8/2OHcOzRliAaVJhoQVocgwM9CVmukUd+wVR7C
NVOiEP3kM9I9V6TbyAfFksGjjVjB5lv3izRdD56JGMTYm/f3fGEeGCV1Bvp80XWf4eQil2v2wrPK
rj2yOEaThJC/hzaX04yInX3EP83U7IgyO8thuXvWxKYr5YqEG6T8tYGYGKfcac1RfV4aYv9zWkYI
z5VOIA3DfHx+f0ZVEcdDF5M5ecdTPNIUJGJtbkTIIIR353mNbyPuoW9C7di8VLbHI0A7ZkWNELX9
jEOiU/yacQoXUkLZxBIiQtStcnRPMPSprn7dxd+PwCSlsHk4nVSXyWD8+lU/1iMP+ltL6I9ZT+tA
Dd5RLDqTtJy8ze0kzdKTGfVqZ9xeiYhd9xQ+4t6py+wcp10egtcF65nnf9Vh0EE7lzKpVxPMj+nD
0eT4LYPqcQI6gHp3Yd4Fa2TUrdAvqaVWl/oPsD4rkCB53g4yy4jU7AsYrajH6ZB0b723Y/T8x6bK
tdGNJM4BjGLifrhgnJs2wgV/grXkEl83yJa8EGQE/Rjq2YGJKt076a8r5nvcWv0hKeDqDWAO/tbd
MhDLrd9R6XCKwleEPZd81kiprTDyP7RVUAlGDMGBZp8VevEbLkSHqbaGEi+r+D2ZC7s+m6gT5Gsn
0bD1j2HDT9siLX/qRJ5n28dpvlxG+axhKSjo/Q2L0sa3gx62SIwfOijD2RM/aHfR+tyDeVHLfQV2
xUoN2/xWsLIQ/OkESXOm1kfKElQrsr39aVSrhePHXyTTJUA9eNVAnrjpG+9t9qvqI2qxvGmfBxEr
HRQleuoCPc4IDKmbiTZU8j4XbJijPFw+xTc3E7KmEkI3gA2nk+buwXp9yuUaQcSOg3p0yjxXZVwv
u10j94Hd0ewVn07Ninlr7l28FvBWgSrAtXhENb/td6Hpa0QscmsfZq5YJA19L3+8ha8nhHWeuQfe
dooYqhXV+NmJzm9p/PedB4RN6V/qTJrF4M4ZO9OJyME0klIrYHGrqbHVbl5dXWLM/tIwAjGocu+L
bUwjh/jR3HpCkBXJLkLQCsQSsvKd1AEDU2EsOZCGdVc+A9zAW+EILGtpNqvKuBDr5rbw4GQel/Iy
iTs15Fwb1QgcJmHDRPj+KezWMYI4FfmLPwQEflGKN+b/7K6bg5mnGrFVL5sODhdnF0EmwSQPQ1v2
zDzq/78t45EW48JmDJFSn62nLplg3KZoM9vUwZ9IAc3vpD+9+bpFd3EqZo9hdqGomHXOa/W51mrM
d6UKjNbSxthI3pnHs/RRII4K831dtyTU2BBZVUpYSo774gxM0HUzmpVsCPzkkJPnA5POMbf4U5l7
+BZdLaGZ66AQ7IZuSrxA4ZH7to0KVHOKLFR+nECiNF1MPSzsLIYxKBvWjj+jiAbvXnyPRi+Pv9uh
qO1euD641tG8LPctkKrTnDp24slIqtFvaNXUXHStjwCj6ah6QIIaWwRyR28NHohlbzslj1mGKfAf
aREb2z8o8Oyv1FAP9x4X9tp2PCBSq8U7C6TvgCyvUjo/hjY9KTtB9hUl8jLyLbkzyzAxWF4iPyfo
criovuNx/fI3iFtAT7ZNMvZsEk3y+hpObv2N8Fc7U1DdXRVcvFrckcEyXlKCsYK/cgYYWMk8FRjP
l1Ko4wmLyTraEX8cU1qrnbFnF29qop7v2LMpC0bAf2oXCpAq8gpt1teRvQbY6oT74+FWEXDOvM2/
A8iVDcB9wWdR00lK3GQLhmy6APAQJuUCd5aUYNTAghEfeIu//HmHAmUF4RK5Q7tZAHGN6qs23D7W
iMJe4Frbqc5o1akzg6HSvxcjtWRBQzCE3uzYuyl7mBfnRRvdaQLI79iDf0txrNghgi03LdRcXJDN
XvqJFS9eF2G+6jiQ8KktT2gElq9E27NCNlZfpWgzNEh1Oqlt6dxQqiA7ludlK/bBUwvldrkz3WAt
Aob/Ui/2ldDoVc+qrw+x3+h1RRKWoRRY5PK9pcZ3KSqruyZnMgXaBCEZNyWPE5WOWZPCdw8DQGot
1SGMK/YPvotCu5/2G7l6zaz07t7puz/Uj/AHpT+1JclwX1hqo423F1sPEbI7gHGDc/H5F0abXmII
UQ6eaZhc/WGPIOeipnMIvh2FXTy7EI7KHUq64MA9zI4csiZJNH9AKj/S7H+EblNKt+at+KfPZfS8
U5K6/IphxSI4n+ilH4o3mC65tqKX+rfdsyhJa0T9EqNLNBStLA+KHnNutRxb46rR2fB64fNAYRo3
8DHziaK4ANCzVCyOK4+0Kpz7+zvbErupRXu8ytKrN52uXUbrb4YzmW+mSLpM9B8F5V1lDx9Lyv46
mEYi1Dqpx4BnUZu2fF4tFE27hD70aWdwDIzd8/v5yWb6IpLByUY0DBBjLGo/mDLbWu4GIOx6xnwI
x+n92UtyNyO7Y2ZQgOxxTrywrcMX1PXPsByo4DK+dUgiO7gt52aBWZXXJBa0LaQOYNb4+58ihb5n
vUD/DFMDw6VzrXMGejYMwUGTfdgxbVORjZVrt+EwuOyLmdhwhc5qNPxXG8zYF2Z2UKk/KKvW+Zw3
aP5nhP/xr290Hh/B5HKdkwUaUD2YWQ/GHOWxi3nZqEAkAjwkgRrqhJsy4x9ikkll92Psu9lOHWe0
TJn9hq9pLMRXyiwlFkAla6G2+tIeFOdJ+G8lNlwTytd2DOsSrQDNPS4Jl0oqtjNyZZy6IAOqEF8z
g2GyBtQJnuGIoOjuce2Hr91mPnFEVOdf3BL1RE87YVIvfpamMmues0mVkehNYdSC5Gq3WiqTlCSi
MpCw0MXbUjdKV/39t8axJ7hOjC/MF2WAZuHTQ4c9xgTEc9MsCWn4pmlxIGn5vHpPMraFd3pBc5Q9
MpqpQJ5l6wQvDgScOFQS3peCI2czRQnLWkpg0h3QMTWZjd2H/pjhSdSheDYmduGIYfhU3lNC5mkO
F+VRR8o2SBT7mEoSKHdApZlvgUdPLzbQB88dboH/vTZu2SAUgp9BRMnZVmVwyexBqfbI5YCEUvIt
0hnz0jFdLRTg0RDlNEYPyfWtYjviQhpmQOsTz7nVZijEDf7E9cGXUClV3bKT77Nal2F2RfK/5LNp
e3WxDSHUQRP4Hpp5+MtbiYPrx+9zCxTaA2/SC5q9cm5x5QTZ+oGDbXDMii/RcyviLhy9S1ap2ABj
Sy8DwYYtTjvjespfOvoTLOXGOtLwkDFZFn9vdSUeMeIIuOeAKOocXVc+LzXfrOZ82jgQFjMdonGf
+1o+/onepBSDkW1ZqztO/VdlZaK0f6kx0Q0mpTf2pekdaTVnd0YthstW4T87cFKp1WzJjHs9767g
kdw//1VnWZ+kJaO4FA8o3i8+E3mgWJrjUZeFTP2QnAg1avZaJ6uocx4RPug6VXfESW+7gmB5DS7S
3qM+jzEvHjTm5d6WE4R9osEkT7WmkGvey1kJOYw6N05EP+5L0fVto8veZaH2ZUz+rLigYLCzu/n/
PFON6HkKTc/WZfNyqVeyewh3jCdFJ2GSVYamnig6CLhjnyZsLU5dYMk5c3XoUO8K20yDPQ41ZHKg
+g2U7orO5Nf/cTgkW28/dEiMRMWpLUzCtfYdOxQA3jyoP4oIe0q/xIOBfCdbEMaK6Gq2LZBx5D7w
aWPLUfGCqbUaBuNkzb4N/aj4EUV4d+7F1eJi4dY2YjEVaPA7V4Xz9n18x9sm4xSYmBoLXc6t3oad
4SMlYpcgFSvr1Q+cPGMbKW6igdXbLkU3r8Rfc/kQZMIjEkGxzwp+7Ft6YXgv1jdu6JNxM36wprva
lkX4Zmnnmg20sO376H0C9Mc09lgWfCWBN63xDmdxtxQWrbGlLRiKeO2mLEGKd6jtIzKo+cUUpc+I
FFQ5cn/Rp4cuxWS1J7LBzaoos6acED0P2N2hmYgIPvEQldi2ezPDVqAno+E1YTrC4NYci6lSETo5
oB7Nab3lni2ws0dw6JerRAWTYmDTSZmKp+yf9RM7PGpnBH70I6xScyVB9pdnKJ5hVKj+LqJgqEQh
sQj7Sg6HfA3uqXa6RLF9ZsQYT7HXt/cp5AzEnnvNnvU6ZlpP+1VNVNzZM4aB/kuQ+Wyl39OJsExE
xNA7tpOvj7GPrM55WCnpZGEjdsHjfEmIKBFBpP30eKz1ep91mR54ulDk4Xi2OTekGK82iz30ULly
e6e7EKsKZjNAZpTwkRqaOv01T6sNVy2BItz91M+IBW8VN+aoOXu9sMhS0OLqVm+Uajcrc4KroxKZ
4qwp7UIplbAwJJGGJwXIji8p8GS9wbkqmrdpDS+AzBkKoJcpxLidJZO8t6iny9JMTz/Kl6c4Nzio
z/CMjL63VfXWtXblbZzQWAaPE8TeifML8WlWD7ocfCUNSlR2KGZiZ2VQl7LKFX7CR5QcQpCU4KRU
30h+H7/3sPPFvFj1RrLyJ+CYjZR+gjcrzpP2gD9j5Rfcig6ET7pFnCnPsvCL3LSUuRF5NnXyYtmM
urSIcEXvv/oxNfI0uXjGejJSn6hQGkTl7tqYNZ024vuQh/NBelVM98Knwdf4ZUbnLQdJ3HZvy22x
ifOAx7U6UaRZIjOkknX0HhxR4cRTZzRSTnlVteBDvJjVyFnOnGfo8s152ssqm93UGWIy1KxoH41l
kahxe9ifZriahQsrVwdpL76l3RG6X9lRe7ZlU+0JfTyQ44ee3nvsITU0FWSNDjZkbJt7iyR2ns1c
zuVoflXG17Xz23TX3t2Pu3Plf8lcqfUyos8PjHAtKZcU5Nvv5i82lehhqHFrhod9Iq28svqN3/3o
NutMSgYQRoRg9RiQcqgbozWYo7Ss8fN5AyGS6qDBsJfOAaJcUjDx9yJ/dT3dlZ3Q4bHg4qK6GLfJ
tp5XfOpCFZdt8GlVnULg5nBinb87/YabtNGrzQZ7kH5moME5kZF9JjJJc5cZ+5pLcW82dFnlH/NV
JZKrleDQ+yVW3F9mv5ASmGILJd41vndvXcjZK5M9b88DSpT7b77XIoQPxP8Os0hD/ZHdTnRbLPOo
sP5wcIWDGFTHhrqZ/klBWkDcX3aX5GoysZmdcqZ/j8P0yBz0TNJMR9fdAs4vgAsXKbDR/R6MykGg
AC9QDtt947xvBICaYHuT+kBn7H4kKbHHKatEfK460yxCoObZK0o3kMVmo7/ZICKoLIbvbnGAc/ZB
GY+z6xa2bqxcv7b5Lqj5ncdsed6cJjqxiOoX/kAUn5Nzv34Yo+I0pLHMKiaicLqXOIj3FGldL51a
hckviYPhuIaC2ksn6p8aGcGTPPUEqyMAlCYExthSONwcNx/bH8TsCqkK0oNSU9TFO32c4TMWgcr1
N/5IA8JQS+B42qdHv6TX03QaV1g1aFyuFN0DwFWDie3SdBeXV6S7RNlOH+cdShEDotj7Z0cdrkUq
PRhwZhJY+WZW/xqDi24oTegbkvCT+4DsvXb7iSXVV07ksijncTuQKFNpvwPNRER64Vz0KFGesg6w
6nXdO9CfaxUfkvcvQwK0VMnoIzsn5mp/WOwBjbCjjD8zkbGMrqh+ngMQWv3V2/vMTtP3LRfL0kXE
8k+AxdyoCCMd4YcNyyVc1HymQ4l0HDgCP2kSGZ04pjBlDd29bLRih2lPpaicSrvZ5pYRQF/dxCO2
AnvOKGtbJtXK/lmXPV/EH3Z59JmnxNx1xnzatwYiRNky5VyfeTPAm7dbo6JI6NlqU+xX47IXfxz5
WC1r1jkwzdu0NS3XanJnsLw62vb/dYhrjX8s1dnPZCz8ejtz0sJUdw7i7dHkPB8aj1yqDC+tru3x
tvwi/V+UNBOY1c4T2qhP5v08pjEvZ7vsy0EjTbIOlt21cvT7wMrUrm1D84w3NgkX2ZjD2sAgnOOj
sYZiBhcG2V4/9bzOMEi/NXeAOOlROq1hfI47D0UMgpLfh7cIbuL+aJa7BaxWuzLxgUkOgMk7XFbz
NO2NqGRTAj22p48jn76x7lJNzzJgO2PvawYtovuz/gU14QG/ehzEb9Nqpk5nktaVOS9f0zE3DJqr
1Oh7sRuLb/L9UbR0DEKUtfBX2+wG3UUraIcanFlUYybOt5crx3WY+jTYiNEaLMskCVrftuB7MLOW
7xeX+1IsZZUaiFsjYUvLK1m5ai7+8ASBvyD/RbnE0M4yNX7Q5a2yRr5iIgPhN04zsXhX25QIHlzA
toLh7GgOTfYlA245jcS8Rc/UgGcaMaPNPBLfhG3zPvDbiBe3jtKypn8R2nq8IVjnACpVpAvuwwef
PXse+cjpQVhrnpaDP0JBCcva2pBCR7PWxdBBSzlNllXOaccS8bj4b5jMZdjO8m97hbuL0mrrLJYL
iVb9KbCV/dONKrDuMIYhi4t51Nq0gtdizt5bz+Olg6jYekOvMIg9LJbcZbEL9b2I+h+AS07sivxi
8EFpncSpYtbEbHc6w4s8IJS08yUQkrGXRleSKRetwYaMbszTBMezdKX3YZbsAUjnO5989dQg4+AV
mz8AnMdGfWwjYvFpJooNvrtpjecpqfgLAEPuXNf11RjGZ0I2Kf8XcU13oncaze/S9cn/rsTuksRF
5Hbl8lhs5W0FiReehy9ZV2H2DaFcEoCekyqs19VHZygm55kOxSiCsd6EaT8UJ2FbmmDilsbLTG8b
x/tgWhcmqLA9JYiRkMNCr14OWtCJdsbCZhcnTLCHALW2R7uf0TOF/2gL8c1sladCssVFi1WTRkRj
Dgo0LldviRNRAZHnNIwEQU6dtI4Oo19zHyPPSzmgOvMz42eQGzgliAZ2iOWrZE/TY9GFwtyyjkO8
EDLztHaQ7gYV/BmP7lt9yzd2AUTi8ZVtJO0vYrSwZpGfL+cgQwyXmuzDkJWT6IA+tOk/lFRJRVfF
diYUgGeTzezSgcQRnRQV4qhX7MenKo4sufNH7Wj0LQSRtns217xYZ7WX3Jhnl4jWVgSGxlPNVmuG
V/LET1vMRRHkDzl/I5KLBhnuI6JxZquBIIpmuXirZw3vTpZTrUiyEWPZi8cFCEqjIssqw/WXq9oe
6PXOtWaplja2LfYIKeCaFBGogCJ5el3XIz1lpCklYHXR1gVDxDQXsiwdfa/Qux8pca81Brmuepd6
VzvBss5nghmfO9uMHkxD3nb0iBqj69b3tbOAK3JbJx6Obz11X6e9EwVOjS2v7/OtqCSwz5wYom++
BHCoOpPCf3bnaEoW9UURGpsGcNDpHdLU2hSKB75ZqSIue3ucw3R5nApyv8OXBuNa1U7EYF+wpgp9
8GFOqIkArCKSa9HaNF75n5CTkC30zts/MzjnmeVEpYoGeI0qU/pUfqWHG1KExdJAHoeZGHYgVO2d
NO6jBFMsh+j08blrkBNcdfaT58E4gAlMhPPX1Cm64qlelueWsEdZ2FfzNvnvVNf1fKcp7Pxf+3Yw
JxKfDEOjMGntbrYVPAfzRxKl2ChKZbG6Geesd51n9RjCp7KFCi98MwxA/VxZOE9caiwLwUubLApb
rr+cNqpi0F56jqXroZafI1V9sSzsT5sPLQ8snQRBDAAsBkKVAcZ0uceEqluT6C82a8yayTymwYYf
64pgGvsp1mfRdrzB+GMR8o5TcVgZwhIwDWSAx1D30d1ijkZ4jTs38EYWVsA0KSoxDxLNYUDzD9W5
VM5t8kElIRTWBbMm5kfjVJn3wvpOnlCb4pH3Vz2DwxosAkUJUE76u5+Ky3gXTSE1r9do6KqY5HWT
oc+s66lgZ46hFaDqkElLCQQQtXI7t6ritAXrpphFB5hKDf3rZIn1Is6ErbrTgKhK3XThaLcHHPB7
xsWc3kXPdEoYU8SGT36CkYI6m6YD8K5/l/vMDT0gAu6Y1TL3Y2CXOMSFVU8pWLfm5sfX2i2fv6b/
XY2F0Smr7nW4+DJx/foKMIWC1fqux/FkXRdsAAlb9vlHMRdSb+WyKLGEQMt2JcuCK1xn9YbSVSCw
0/37t9itA3xePGTo/XjwpThNwE7QxKzVE5TwUlJ8przVBTJlmkpKXf9rKuezNgbxgu+hqmh3OFS/
Nech4Y96xBOKkimyY28kFWu+m8/d3xaCRMNFnYL+inop3huUnL4tpWXtfbJAsq6X66SpcfV4UqlP
ab9vCZ5Ug8wLWIz/A8n3nRdP3cXxRYQrGdLCF6Lu6D/4ddkIRsz4vIhV/XbX/2qDsG7DjIxFNhkn
zDulHTem9Sx/l/r1rHq3KEH1PIPxL1JUCKeCDlOHmjVWa++tjjTnupobiI98gspM5N07h0VWWa1n
JiH5l/T6ZbnnR2VcvruFn9PZvBZ26NF+wQo7flnfux2sjDmKnesdXnKJ0WNUH7e/t/Ry+wJ5auxt
zA6tArkqLouNVioIv5BwE2dt/gwDcBkTC/yDrbpt0P7d4GAuXjTeZEHymg3sOzyo4fYhSRDubmdn
FzuRll8w7XL3HQYpxOVCFEX2QFS0lu9dAuBiWL3el1ohT6QWaGjLcI2Ilf1eDTj9V7efWePDqW9o
OQ5KTGAaVAdLmsXv2I4F+lWSJ33fkvMNSWAXguH1vLCZjSntN1EmXI3c94CPlTbsdBCDug6T6EuI
xQfji2V06tAxVxlx6Es4lh3hT57EQHKS0Y/IMaGCBZm8HQdo12rADnVGkbbHQv3TUhQQdgVtsjNy
hzgTXiZ3yEJjcR913exePzonw6+nnaYOX8wa/qJ9mPkZB7TnRzmsrT8rqvjZMEOK/jyKKBevZ9lL
Zsb0qCNFRbIrwdkHNAKQn19ILbm2pFtKULUt1Xrj7twRt2+A3XTbGt19X1OD3dz+aEZbj5ymUgfk
ZNs+ShGxnaF3aGIpyuafi+0K/r1HYMv1KBJcAV1QnMNf9Hg5D8cQMFHZbq2Wqoh/XxveFi9qGoOZ
jq3MvdoJwPTzQnqHSt16syXldQi0QTxU4cyoKCVNqyWVMhAAMxkwHRMMtkn79tDdFwaGa8t7VOmK
qUtu4c3wTMBhMiah6wLMi/Ng237ZZMY9DoNOpez+NvcHcRJW/Y+b1xCKf0RQMnoyhHbAEXpH9dzA
lltv8A2I8qrb9yTzTCDNlgrMDLtjRbD0Ua3MFL/+CrVfanAdLnFEdxVSulziPsiDdMywJXgLjFo+
ilRcM/mlxwrNjSVMIdMkMD+o+sMFTdEg0uzifVbhSoaBnuqp9rW1IGKcd/PLr7xz028FKTDIaq34
Qw0ICOFgrIa8tcK9fx6w6agspGzgOGEor3F1EJMr+mFKw8G/M6bov7nJeCNPFrjrlDmvat/YHl0h
hQlQGzG3CGoG9J5V9Akm/de3++NnZEZBduUr6uIdh3KUQJOyA3DNDKJkVIZiXmZ8VwFTnJBuZHFy
y+0E98b1sBrGD/uhcyAfa0Aere6yFcseoirw7T6alq6Ya1MC6rJ9bD4p0qqKxETRiVGL6ynHo3Kh
NpKIa0zZvILD6IyBDREOljzqnOXRtDp2W4L/NOCf3CcWERCFlyNAiwv1LyCWl0NnaMVTMddjeFqh
1t9cy1u+ERa9b8/54qTmKxO6SCNZd89AY0mEhB2WzIg2RsGPbry1hvPq+EXvU9552yUw1HBTQahY
sfU5pAWk1a0QQZF9aBpak8awiug5A/FPftvRGxaeF+KcYWRsvzlLdWiVN8NwLiXB/kR+47tPt1r6
fDRriAvH7hiINKoZS3Xa3WY0KG0lfUgF8+Rc0F9zx9H/LMHfSOCQJVzQ9Vl0R/o1+S98GcT5gXVC
ZhPGQCFBgtnRbDrTwhD7IezRA3WPO0MGm9A/68ZNak4FCNeZ6HQg/3xZoDsKaactzKQ7IhoT0qJQ
2n8Zmdtg6a/iGmuLOhpQIExn0Ko1qKRGcoJliznO+/mpEg1b2GCCAOkDAVd97/4b5TvDI1KcrWKZ
MikmoXltjRTPsDBmr8MJ5t6+UPahFnGy1RfDbJo4SQLpEvQCVPw2Acvj4UphjOcWdUeQtAGrFwrX
4AwJZ/t1c0jZA/GglLiJgHzAatigIy+q4xW+AlH2xn4fDs83MAYHLPwBVxzjiufj9VeVRZZhZaEy
Iia+A/hPdmpuoTdj0157My5GbYGwbsj5qpRfrEm+/Zfvm5qeHncQKspH8ATC+rMuyUvYWlZ4wdcY
ohnVG9Z+hoBuYnFRPCitqphvjTaFD9eXK0uLdt/GmGJg30I/dbTtp5LrhNwWQ2qRl1oAw6IElCo2
T5mnwTSESceBYQhjzBL7wxg9Ji8AQDrtkOEW52TqLZdq75s/NzYYel1mHKZexCdgr+ST8+IUhTzA
3rmg5dIA1WrXW2mnEm8YwLRb/gcvKQgpO6Cgw7v6qt5FVifQEXkvi3ImlKup0NYw5XkZC4+UBGYm
+yAQ0xj8Wlu3bS72lX/AakJSp74VJwa68DTZqju55fwe6wYbhf/zp5sWsQrRaxoLstjC5dL6DDRC
b1ZGr+/Dnl9MjuZ/Gf48OhR+w50wiX2SrPlpu6nz9gD9pAE9lmVhHXN5eeTkTl24Q+JS+TxrJ3UX
Dz2M62MFgX00MAkeV6uxe/tXOSsa0oPKdfxJrqdpLCT1Fv7xoL35XeUB1wYMciHiOhgcUNPgn/Eu
ilfjeYvkWXZqIOxshzyPwCEiSCFT4iLT/XuNvoA1qsjvVDxwTPLpKwJszHfXNE+2otWuywNqVKH3
1XWTUZBaEY+DwPkUgie81Ky438plsLbqgpox93dGKpgVygX2OpVT3J9S2OJkeSQiUOHKfE7tfZji
L9VVAhbOl7aSOtmas29eTR/Z91iWsURkrA0KfmRah/OteNWKXL3Xe1ttQj55+QztRiWsq4LO2Gvt
v2hnziSggNmvm2pUkmENwNfGFAoRnTMFHnMcqIf9ExOmVz/r9mX9YKaZIGc3/cJCBn3yrA7a5aV8
hzuDd83DikcvFHT4Rb4s89Z+wrb0r+NxvO+ZrujmcelfmpsbekGb9aJbiumHnf/XsUWg6P1SYVpf
Uc5NStTPsGSVUjFDR3Gon2RSuAUO5rKw4Ko5MQTIq5vvCGGDXlaX5ahzrA9FsO2hCoclsPTBgdvi
Hb2HKFmtHbGTBX88I2hhW9lS/9QuaJUXDVhsY3jc7RnhCuYjz61CJx4rhDshO54O2TSrkoPuF7JG
3zimXBoVtfZKmkHTHwiQxMqYWL15QtmgyV1OSQRKwwNKu5GTvJcvNDhObISbj8Gk/lKMndYqt/zZ
P1PfS2kacz147iGbiYHE/QwKkoyDA5ekOAwqnCYkoslSi+HJJ8tpmjcFl7UPxWyGoS5npIwrk+0s
NvVuUGi+NHwBuia0l/nBfBzelykb5di7OGEDYs3GIuZ7XHueWMC349dcXcwRy8swVGvRYWXtxgml
SOLe8vrHadveCoJfLWdZPRlb08SsMQYZrkVQjju/Y+8VVVurpCezskbzOAJxZfWF2yhQg4QPCqp3
pkLXutJHhpiyRLVw2Cd1FO5S6fD98WmRTMqyHGaBkM2e76lRN0u7/JX9Iyt2uw28ZmbDwp2dj88T
yYxkSrLozy8c50RDqNvtM54PKXE2Tiwo871P7ol+koZChVvcgnvI2OajCGZmZNfVhT0znSxAbCYV
GfuoNt+4MbXdy1+cJdyVpn0LNmDIsD/VYR1ho8EGaTW2R+n8aLBWbsvlFgosnFwr2XuFNTdSHJ2J
eWO9TxwGaCUstwbek7x9J6vMMxVOxUaUgjO5OVYmxXcNmVSjs3EuamIC0GF6mqdcSmBCpns4J0L4
kmZ46ZVDFoVUzfRG083rHiMOlbSAtxAQ4GaYgJkIamI6Glljzc9gaa/mSWPoKx0EbUKNMvTfO7+3
o5tlbSiMWVcQ485bD/5n0dWdDaQksJ6ySFzg6PAje1yzLl8BMB2bIH986haFaE/VXy3q9lWAW7BM
pK8JoghqbanYKGIjhpaAbpco9/AdSqWuGxPVAbyIwCctmHbacy4exzklJNZAfY0//Wrc44Zw+lhd
qo1g8VXlO1411Jb1Teau1Fk0u34Xvdx3hcvkTM1pqefv968ozDE9jlTNzaRvt35r9HLoxusAgF5g
Xicfn8mRw8Jr2U+NGbx3B4bgo0uTXAbWrukldOeFHRWBAKvBPGgkpUHG6XcXFa7iXrCPLnB1WdK3
goQCJXAsfLjFZs1W0Skuxvo/anyst6fLOBQXoDe9s5vLekfJJxwnOfn8IEU3SkAW4v4ged6JJUzW
nOwB2j23BkD/G75sasJ4Sxk2/vxSXl232lg58k0L6i39q2pljzq/Gw/7u940koM+vPoyWvIGkf9c
Yac/RQoHF/wquqm5MEXLHUPFmCS9Xvq88ZLWceyPJanwtGlHfVc0rYyq4lapbHUdZDuCp8r1NH4+
zEximSIPIP59lW1HHdL2Njig4Es+L6LPERnHe9qQ/fTOk9oXsnctQhTvrjCkg9nBRlKANamVA7sg
pczOiowvMqeDT/ZhnqM1WHfymL+YuVxPGQIRccqYdqCQeuC3ufXoqbqmNRwYf/ChI/yD+0Wj0mp1
+V4pf6NC+0eCGm/QfkAIcxzTDaZn2AQuTnDNau4TlUQdv2CzL7wv64ZrW2ImFfRX6hIrOcSvUPDQ
da+txhOhVI/zxREvPGAGSaXH5GIOKcabmcK9m63Yl5CxBfaBj6Cqx1Kc3oiVVqqVQ1Zu4bPbI79s
52duyuuadP0C49+4ieI1RMYUmSzYwW8d9DiFledP6vO7eeIvt7Ook2oL7NtwPrx4I3HH8C8RT9dx
A+vp7Nd6i1NLv9xahuG1WEPoCjg9O2l/3UcgBm3eYAQNZ3xtez/w0qRvXkv47WK2d1hJvCbjB4f3
2J7U27OvfkPdEWTHAo0ohmMKB0nhQFuOuwrCbvgTHTcl63n2MJSj35ktsXxeodznJ3M7vEjA0rBk
uHQd0MjPdUkoMQ9U4VDfyNANBJyzU/kARXuwGueXZGd1RBXs94PZjs8MVCcK9+NPkYo+AVZRQUln
VfNslcV51fDVzQkdLM6gjp6faXjE9VQArrwqIF/RS1QXbr5/+9jUxVylZX+Klwc6YdOjGFAdgjXM
uDK8FZzSyMkaWVX1zmgcIfS+2YAMEAymGItjklJUo9jBy4WKiLdipR/5qNtc1v5WpfBSQPr5Z1Q8
kpHb1AGZyWSdr5qrrL4XpH5CqglXGOYMLH7NBIhgv/P7uXyIYT5mwoMLS3w1BQBJbreCa33KOJYX
uR72dCwftmJXtYk6qQJDpeJC5QwvmyjmV26z/+SmocMq3N3bCsA9FqhW9Eyt+fZj2OGVPe0d8Pqo
b97VIEYlOeaAd1rkEbyM/V0t/tCuA8zpMlzY3FGTn3ISrBzxKvTCAvcQUCjWUh116wL8k0ligg4J
fbSYTIiH5X0RlJiNCrom2fOt7NLD8Ps+bZvQPBv6lnPFvzuGlDu2iA9AQwgr7C5OoALpgChYE0tx
6Zp7oEdX3BeNNGXrInLWCzCbRW4yaXq9CshELU/qaK56Vh94K03OwoyFDRjCpTNCr5K4buTxWLLV
/1T95H1bitd8VKr2Lisjulcf+3n+Gge3n0qNdZCTddHd2hhXNv/54TdD0gBLnLpxIy1lucKImYhP
PFG0jNO7+tFgKqtwK8H6J9QPYbsCEqMNpa6Z85g0ucuGhG5/q49v4wXObQiiy6VygOiWWj4zLrzq
XjTOSq5D748IZP8agxkQreKOVCU2fV4Z2AcApr5l+sfo4gfw+2YdOSjnBTDH58qISznsGzEEvTCX
kFRH1NvewLKCffVNLwz1UZxqfkOzia2o1ZoY1FinAOQPcg3rcSq0bqTWSglnAr3gC9uktpuGvY+X
2UcyDFgWWj41F3bQ7amg/LHc6a0FqhgbW/fY1vVDN8mZRStl+xQ1+gXUmu5cLbQcHO3sbh0UKhJO
VUUsfGa7tYgG7skB/ijy8kljGm4uQTnlx9Itr6RQxYK2ri8/ICaiqI4jPT0117RYgAdszaR775I6
7PZugAt7tN3QXm16zX0psheSgN2BKFlRvGzWuZMg6w1QTKKy+BdB5d9T6o4jWYu83/ASSumluNAI
QHISX8CZ+IDcR7Crt9oMWahFixYre/twxhJ3mFlL48jGxmL8HdtzzkCJMZGtPzTwuO0ONFBwoKub
rOOaBx9QQvc1xqr1UTj+gttUj18KX66LluEQlhEN2mGgS2gmw7AI50RCWPpuo/zn//UEYZa+c0It
sXUV9ejyQQuLt41EIDPJw2vbuhDeDApEWVfY9dZ85bx5oIeCPDiQXgdw3rwxk3UR4u29rLslpGnU
M72/c4siYstPtlSdQUWVcVVA8Aj+2b3KhOiYS389btj4hWhW5tOrRKo+6bnxPkAFtxP875LLhuAk
vUJjErWp6uZ81vQ4chH9Bq9ayPjBjNijI6pN8+oQ4r8kRpnrV5g28XsqUmL7V9mHy9S04WggkY/W
7bSnBtMeMhn9k6U64dHsuSgPqDmK9fQSKXEN37xUBmnwd2JImO5I0y2bCCZ0+hdYMhviR+Iao5fc
qzTQVPL4Gmp9XL18V3cPX1cjf+fxAgtWjEQ+eBGD1kPJpPt10awifT0YvJgSqukUhyrk7kq7HsP/
xPlatVMrexXLXEkZ976BpoC64csazraKN8BcyjRBGkTKSBZLuFc1iL1CH61jE6is4jjT3c3xvC0A
Nx0I+cKIZ4nn5YsiTE8fpJBoCrXMl60mlna+D54GMM/ylZMifUfZh8EXWokVk0p1mH0pUday4ho9
sDMniItLf4gC7XDX1kjNytVq/pAN/mnJ9eVPShqY3A0TMfXxICBs5WPMpTthJIhd6qeyYmZZ+lQo
xbD+wiJcJJjnmXaCYbC03Roqv8ILt1PDSRD0CDsAXfCvKifVMGLwhr+sf4ACRvHmlqn2lAAzFO2Z
LicumG1XLn5dDWTSS29D1h5VokSIvZqym3Nw/g/HWn9hFdBEVllpyFy79S7RLb4dISXUuNwk1sol
C/ym801pm9M9uJpR2EFapRDQ4NydFe+uMiYsFUvAHq1HVuw15DL105aVxjln9GCKt7o9iHC092Qa
UORCmy32oKQWbVRs9aSrQA6hd1S9cSsoM0IHLr48zpCkV+hSXkQDNAx1ibSKBzHBZTHwM9IdTftL
7HZhVHjOSedz/LDBQcvXz3P0kJE1fu73FjVvsJu2yhSvwY4AfBEfMX4zpvdMh41/RQKE644CcV33
6lxFpLV7dj3xKDwkTWGEu2+BGXKL3M5dda/qCFA4jQKljV55pEF40dYE4eyC4Fd0/TJFKtHHApWy
kgcGMkAyz9o932DTZz1kDMRaxcA+LsT7XL0jur+c0Vp+53sTbhEPHebJ5mIMKfOIzkvgDHKF8Sbp
r2rARMFsaF5he34Dhd6+wonthmM4HdaMLFi5YI5oWD6AznoEf9JI97P2CqFPt0MeWn19TaQBStna
Wy30fa47Z01kyAkPN49l/z7FdpPvqceYE2hdBOW6UhJWlkVRGS4EtdT0Jo+pY3N2jHxXEKrl5kNI
KdUdsJjviyivOrBrmcnGIJOQ2ouOpMQU2jCMWMvkDDkj2cVtEZcYNTsutf/vve7FTlyij+kwO3eu
XQ897YbN2csCDw19YykN6B3pqnSWAGFe32qJ/Rs/A9JIU3nvgDNaegM6t06/DocmFYqzVXiviqnp
PW6V7va+IevQvSLWuAB7aJum1hwSiMK+y/uuZBgakMee3hfR6BU/3VcnPedGPtGFeswP2V7cEUjV
eb4lzC2x5r97DjImKczRMqUQmp7DGyC3nido84yyyKNwRAcArgyMn7c782ksMfeYqtl690VBYuzK
piZvXvF03HZ2qbHT2XRgg1SlBCvjf9bZAWDnd6F7uTIpjTOQjb1fVt4cVbheYbi9OnQbAqTtfHDi
R3mz8tBUZ50dLnhiR7paJ0D1rg4OOsLW4j83H2hlO2tWhDlPRNOCyzPHaDMcqHh1nljerRsSLJnm
OAs6m74aWT4A+EN8sIZ0aWdC/0caVhgah70a6+UvtGS0j8/2aqjKa71/Hhxedu4rM4B71wr5tUIu
06qvxUggzBAGRTGpaJiLpFrqrtnZG9SJF9I8j7a1wgF2BbghtexvL7U5xGd+aBczaA7+r5oexHad
f8euL6C3YcUB/Fz22LYSoFEltG/t67cWdjKdTYdzlPOXNfHBvgOE8i3BudmYMuDsbM1o6t/GiE2G
BCn9HYBlLx4JxVXhnGgt0YyNmlQ8HjmL9xm4LCuj/Z5gAvlYkqQRZks5vTIhy5LEIgaer+u3ReZC
xI/k+em/WqSFK2ailYzgyUX0yC4461m4pjJ5WdecrSoHwM+tCtZn8sUL4zfFDifuv86GMj/nGhGp
Nq3noHyQgrv0G/lneZr6y+HsovTHQR9Uxa4/JGN/jATEb+FazkJ+KlPDpTOE3lJJu0MgaifYotMf
Nr76Uh+8UqjOUmuD9s7H3Q1KZpKiDil1YAGnGs42RLC9iATh2x23rbFn9WdOhmtV8UF9Y4ZZ+z4j
qRtvyDS0qS13x/NT0JEgYn/r1I6o1AFSg18oY0v6zdpZskALCV8WGglssrj+kWo4dcHXS1sTA99h
LOcfxj2IpRMTatCLYHYubG852wx05ghjK55OdP2L709rnHd95Zrfdc0CrcsUyuDq25Yxn5mmFujI
rYMVEOx0NAk4cIF3BGqfSR71tj8ZHpY4ahmjMDzvquWAmoUZPP916e6WFEvDTiW6IScZtq4jBtGx
GQUyFsLPmLrzDZ6uHC5f6AYCzthi7phVhEjGV+lXtdpgU8MyRFMcP7JuIPwvLxuh8LkcTlxDIxCe
WQqK13OPpZa490XjkDksJpoHNqzFM41Z+w/CyfS6oIludEqFjG2UXJiBOaEDjJyE1WukgaWjaf0f
2F3lgfhL6uyDEYK9hTH9Ay85x/3xp8Oc27mquvu3jMUjSae9kPl5TdyQuiPCrd1dWPX7rmk+G7l7
oPjBZaUX3uTeO+DOOQB/+KrdEB2qJCOiB1DRSIOBRdpkxP+NG5NrIUjXEIa038gGbBxXke4fXi8f
4YO8XD++bn5lZZe/HURy6F510NemgteoP5qlVQVytBraJMKpa5CP0BV9Zr4lLtHCUBJZrRSvCQmF
A2UPAYHD2ykkPAqA0lbXPLoQ9DC+iqWVa0K9TKBNu7ume95oaOMs6Abtz3vKr25rcf+YC06z7M92
H4Qvhah97nvzbz8PayCJsyjY7fvmX7XMZoKiCc0eVDR0fnIbhF4vQmvo3HIcrIZFa8FX6GFK8072
OcwT1ia3f9+Qa8Be3NwjnztT9GawbVZHWTLzTSczPcjtOd05Nr49QWJFUs0eCXFWJvnYE0U+0xIm
PInbiB6FDTz1XBqbBb7MYm2hySvxpcvf3a5yCNGQDFXy6x7V1j6oa07zpBXO2KSulfs6vOitMq6K
HT4Rc8Rvu2oBdIlkApQmVz1kx4KoHQzK6hrwye8qCRLaIf/SbWGobwclqsBzjEVHIfS17GpSO0mF
gD2npYwIwodqxBNl5fyFkv7J0oaaTs6MRd3VXq5tlmwrgK7cVhQ/ryBrhyrWrEzKejses0gOaOk7
DeAyFeeKdP6OJtCM1N0d0HAhfj72kLvS5akKVcdQno1C9BKdLy6x0DaQLlSPJV84w6vnSuP9Iegg
L5wqDQtfaj7Q1LBBooXRSQTti8tIQ1tfn4PcX29nesu4jslFIxubIehKV9O5tkpkWrtJNNtEHCt4
XqSp0GTg0C/P8egyjLZ+K1KCxhIs64kEVIN0RGCgy++X8sHoJCKyOF5CzrbF6qOXRHF1+h9Z6PAm
X8KJzOg8bGl0rShvD27RgkK9niql29MMVA1q4H9vFjXUXq3MSdqMMwV2Hu5I4jiyWjIXmSpVaTvm
n5eVeHnUzWtri5NLhRQa1YIlh1RCIzz64zrktXlFKnBr4E3/4Z/HHPFNIB6gBJqreVpbtIWjAJWz
hGGd2+IbEZ4uypIl0vtwd69eLFaPZbeuy4kj24oeq8EnRBfM1uuZoMTHs5rpXGQ77mQSexjPFebj
dlQjTCQ2A7z/q/bcn+v6JTN5DQZWNqoMRBLGqXEf7wZvTTFYhpocm7aSZ4z412pW6CXoaf9feKIt
FVgYGGdeV6ubwxhC2mMiaAV0H73nxTz5HrveJvNPUhUEJYXvEOH+LZAb5QpAdfTwfw6JcmeMTBdD
6H5M4WiZNfI7jIwE6d8UvxxN2PtlKrQfhd1fbsV1pFDajQW4CsL8KYB7kDqw70ac0Om03LdBLXGu
kQagt8jIvGMTwx82qlpKoZekwKhq5bP1OUiViv6KM+2AfzP9SYuv+DLLvh3AFZJPPwJIL/lWJ39k
TNUDapR3dEAso6a+oF9K0ItzdwOM/kJiEXzVFILyU4NJUzmaueknlDPwtVJltpe5DA/SQ0P50rBN
/wtDeUA7m9aQ3W3KqLRPcsu4n5tRAb9RyIrxtEMDfaqid8SJmqDUF+GCScb4W8OJpRBR6mdwIFl4
3CxjVdcNqTcIikJ+kOMbJIFVXXvyD3qlU0ozrdCphgr1InEq2/1VAeEmmaQs+VBDTPlFtJE5eirh
ej6pGsX3AZggM/72adJr1dB2kQ2AN1yTyqHRvl61ibwMCxxyZSxl6BVtO9nljE6ssMaff8BMhr4a
B1jsxRbuTSKx0x6H9ZViLfZ8V8DTIEX9knvxvWAjmOHjY/aQf/arSmM+03jS/PSq4IbLjmq8C9SE
/2QAR6WuDwa0MzhGamER7AsazhDPUVC8xrm5hbr5fmd4CLVyFAYHj0cKpctIg+z1k0sxPnJmYtb/
tzzyURbvlSANm1eNBdAvyq4dTpufDlW6iisfdjGn5qITerIvLQHzNOeUgSrbUXrXJed/oskyjA7h
IJbQ8/AK6KV14aoJWL2p2dGO5Qzjo12sw2/CRD03TtpUzBpBPsO3D9YwFap+XL4yM4k936eQn6pR
RLWZbhsIxM8Wi4aHGplZjkL74UDqGnoL/Knf62n+whZriYWA5tI58LyAmUzzfrQyfkc0v66jNNug
UrO4VbmSkPxKNGDtzcoICG4cL6pG6pSCaYMLwKZIu1AEwqB8TzEeWCVNcxUtb+94q3TI/dYFlU+H
gf09hHXMojM9ZU1e//f0FxQUBebpWg4xb7wi0Pmo3gx7/cdHMzLtqsDj4xBkb0VFn9OmLqLZTOR7
57HHS9IPbagx1s5qOpVQpK2YeWQobsR84id9d/uK40u5Tr7+Fy4rtjEN1uJ3ZnG0DpZ9iih6AYg9
NIm0GCq0RFmV6QPmV3eLkSDcQwHhOv0SWhn1CKLfXShDuX6aNL5azXu9NJi3y6GOv6KwkhsH5JbN
lEd3JUFyEpXgRWEqv5/V8FmxbCVfB0Qt/DgP0IQYqDxuwntN9lXLrjypVfz18aKDNR710QqEiVkd
bsaZ2whr3EsQhY90dIw4EnduyUAuer+UpO2LaHWl/Xeuvkmk4VUNRE6MJY2bwANvjTHEGia9c5/c
2kOWoT7mojAKuczkgYoFUkrgzRyxh+Tnj/6cgEpkbiG7+lFNlEc9fmkp/UVMstBkOTS7jbazHlCY
Wdq3lYAIplXBeNFra3G8Yfwnlc5CDq8USsNFKrEMAIFPDtn0V5zYYMtCNFQiiBeDC6HNxGOyBazC
0e9sVSrcA0RU8KfRbTws3EenC0PLUbFaq1vDfNOF9/OERPM0WOGXr372N75MS12QewqnlGmgblHd
BWjOA3AT7iSxb8VvloqJnVR3RQ06RWDGzym3afjoksqXWXxiuFnCXuYEhEmFBYiiwyFi3P2LMD1S
2JE4SrGReM7H35+t2VMFZopaOAVhLTYk7ppR9vrBghh/bVqpxWPAO2ws3RIdev+3ItryzcENzIJo
Fo54N3K5r0vbWL1AgIoySU3J+3r3h4mGs0tBxuCRYc46sC/d72ZtFi6bklqzJZPoB2Tp4FD2Mvvl
LTBmWdUbMaJIzJw9Vxhyi3SoL9V0XeZP40eLzNgkenN4VbjV1ZLrYSZc/IRXCdtfB5UHlPAoTmpR
C2+dvnc8VXCFEuHqo0pUX2iVL9suvcfcqT7cqdyVQT6j2YMmiGssB7WEnokNrdTEMEuhHzC+iAPu
3/vRuKT07ugk2tci076pA0LitfuoslywIu47AIexgwD+1oVRs+Ox29IimrT6rlPDDvdz/tx16X/E
IL0+wELyZJTZrTxaNyQTGBd6XShfP4a8s4GLzSV2ftVMafzdQKym2sChbAMBp3RgVStdYrL2lWH7
3NTZV71NSvZ/ijaTYY7kH/uKXtiug/UWVyxrZBAwjD+qhB6hEoqRvXJv28/5vo8GeXLQb4LwO8uz
zNVRXvOuN3epm0ZzD84ks7UiBC+F+GJSy3QLa3FSXZqOKVIWzWGJtIoi8tDcuv70SRmoxdcxG3RJ
UeuqaKfmosgWoYz96cF/9umUojuG8jgPTckIlBaZNHXRCdMdk1KopsKWB+vBXSAB2pBlAVhsp3t5
X6woWSmxMvjwO7yCXIh1EkjHLc23XetGiEyLo+2c5awqcxEutd9MQZE/BOdEBb7cucJpT0ubwpWp
/T1mNLo3zzfrQ6NTjjjNucsSMcpiRWmtQugJwQhk0gWxRGzs+PtXm2se67f4qzTSQqN0Wqn5Bvm9
FD9Tx5EGE4A7o2eDccrQaFggdmZVNANmeE5i+EpjJfe2gBTqkByxybT38KyUv/M6ovRmQc/ZLN1g
j2Bv68O4h5YxXrHQ6KbnXLq4TETkWzI7WCbcckTNpzmUEofHlJLv3V6o9tFrZ4MkP3OaF4+AEQjh
lH1uvf4IeeIslCrLtbOOwOLPoQn9fcV8Gz3jBgDKTYTqbVMItL6B/0uxGUKtYqhispTuSXSwdp/c
awc9+u5oWlAjcQjjs/fiBfgQLKndGoFlMH31NZ8G8SACTPH4d4bKJyXHnNJ3eTiJ04aaNTiCzExY
JSImAptim8vUac+labh0ZNUOUl0cqkcZACMup92DATzSzEmSFRmLyH+X/aSULWyvwn2A0HOLTLfz
4n2m4K8AB5FfcLoLNU/h6ODB8rJhLqjtkjgVVkj8Hg3tBIQdDP1rhQByDJ5ZmU5khz4qJqs+hfa5
VDUoTmPFwUMQZyvwYIAtE4UCATcaQc0i9ymjjgpY/h31GBFHaRq5kt44cR0pm+/cx0EoMI49ZsYy
nTrVkttAmVcAl/c2GqZAtEpeeFVKak6fIgflwpHcJICOElMR71B7F6vxKkiGJG9hvKAcF5nrOpNp
3cNsyOTyws/s9CLn482kK6ulf4Y2QvkCxRVxD9dqXWk6eaPMIkYX6i/AV7AUyWE1oa+CV6zdPo/9
J1HeM3vQz2h/EEpnpKHRBAxOTej9rtRXrGtJz8jyB2L4bDXCjasYR5ZWnJYBIDEzkOnpd9bzbYpD
azWyG4uLuwnVrl4E/6QPHH/xS3ME8FOr+o0n0jTjrib63fB2TfQQq6Q0MqjIppemAMqbD2E6nc0P
fCnLPb+ZJ2ndpwtYGxH/PS8hqjvnl8102B2lEVWYEjY/wtzX1BdIxg5C2ON1FlTIBV+3CegbqHyC
royo3M+UzTW8ARyVX4H85PcTgUY+W/lGhMJHVUtuppD+Mzi+a8gHUB1BkFNIxZ3Ke7AsAKdoG4Ii
tBbYr1amZN3TUJPyM9iUQDDqJyt7W1zGPmhKsEQduolXF+2KwnLic7pLCtVE0t6fDxuB5kahrO15
yc9cjBCT9ObhdxdGfJbpcLCM0kKlnL13SPaOOSs5+2kfTYljuGjJ+n7myHmYeZZV1zdxp7IF/Xcg
AxD5corThZzwrKE0iSeWIwOpAbRyCZY5jUEnZ3A6vWezOHmybppzGwyeVeVHc1Nu9hytvwXKBXRd
bNgf71YFFpJpKmIQMmeGocNJ7oujt3GeSvgzNRe3I9F6G+sTG75A13wZaohb3ka3mWUcVbX4LQXm
l7cS9eRVWk2YdzwOMkOvFxsLOqiCPs48+yJxVzLaSeHn1vmBV9MV0VvBH92SmVywPRHRriRaALqy
AQbGUZbx1LE03UiDzKL/vYV6Mn8yuieR2JH8Xszf2lo8f6NOujGzZLxE+Nsxflbzwma5eteQdqjc
YWmI6korig1zsjkn+Za5K+vbTUHxITtrZw4qN9DygvWooePFBkwOZ/hZUEtZrEhIeAijxCUKcXLa
5C/+oSMA7+lxbL36gspHhaLzb719zXwvbEoIXgf3S7ZLDiEylIB0B63MTaPJ0LgdSB88LGoZm/aI
I4IUPdVXiF5dNgfX5cyHEo32Pxnq7KxEr7cQ4XZe062MdDErPa65d62svX9CsBbsjyk54rAAvgbf
gSNeLGrGnN2Qp/SWp25zxd9uxtB0rA/vzLYwrRgGXH07CQ0nHtcxt5GBFMubVcMbyvfPovYrpIdz
raT3PlX09US8Hkn7Pk3yvzm/u1MnGRGeBwNshjSuOFyxfxsh1Zwu/ue9IrFZYbh1Y4yC9O1H/l3I
PUyjmigRGJlUT2sNSFAdH15xitw8MrckiEdDZsqeHJ5qLpiq6ajLXFHctDrxhWldK7NuH5hyKlsB
+waH4rvIXrhcqG7eLvmoYaibwYstNdHQXg5myXCCjbfz3HG32k0dfi3Y3KrNiq7XpfMURSx4kMHA
8GK4jdr8ukzJpYjOBkqT75JEAyQlAQ4EyMrjWKJypRbB4rmXT3V04F5newZRfGK0pHuV3XOMwKyR
btjQpe3VeiIucneIbhFo5IU2mZcQFHIRofesrpbYxR79sPNrQpLR+bhJ1dA2lTnY++mp8xc2e5SP
Be1OIq4KxIH5co0jnum7/15OS8qU2eyAlyydNGlLUjwplwYbb8lzC6Y9h41VRBmbxBRBfy/3QCgi
JgihP/4Ci8lHOQKeEJnMiRXxV0YLWa/+N47CMHG1nmmIUmKOmUYfYIXW7akDcDeRZgxFyq+Jz/c2
nfgNLkyUOlESHlOh4JnyJRK9+6+HEhG5DRvv8XXaeR1kK7oarPFgRnLcI/ZisCcw2HNtK4Zgki/+
pU61nGewUiQDy9w82q85BimUWAN2Zu9Df80tSobVlkVzb+o81sVxkznBXSv/2BHu4DblB93QAYN1
vvHetncDPeCEry9R6wDVf2isAj2p2+uyhwjQJDiIpnroung2mfQXbbHMGgs6EdfveiGyJkQYOCzI
HWXyI3iMQQz8L/8L6wo9xWDCrRIbnErOIJKCMrPCZcodZn0nIgNh+fFWKU2d1/Uc7jqJbHCaX+fe
qTkdmdboM8gUlyNtDsG22SyPq1E3EMnaprA66q/SEks/RP3bqSzm4lfnJqNIvh3mK+3aoPtoGT9P
WozxMI+QU9u6wzgCCdjDlGfkZvF/qITt59InKrjgOxgLT5qhoxdKqBnJ7zdsiFqJHUqCHJbUV6MP
WheDnJ8dMG15G6oYoyXuOboTU2JMmj7BuMJUMnv2IFgFat6yMGUotQVWIR/K0pcB7Y5MsX/W9YUk
X9Zim0hMkFyo3y74TsSMQTygk1VV+xSm9Cc2rF4qXKdfKtZu4ERUNpVMZHPjfjJva4VTpvO2wHMS
kpdOWNclZHBEA/iNGRVzbigLmh2LtV5zSrPXjanOtPBciJ9h6awcOEb3EOrbsboqihnzePDgdh02
p++u1zY2egOxakKAT6WXP8UCj6UfLg6Ct2Xwyuy4EIaBWbiDDgJXwKRnF/PQayGlDv9wzib7tiy4
bebuH/o6aZVopZSqyAA8VgQ7k5Ky9l2ZHt32Imk06HTmXiQO364uaink/3kz4EIUJ1jBCKALeLUL
Sazsv2jlQUsuO1yJew7xSPO33sh52cH+CLWegt8w8wdo1WbAI7grMyL+eELSQkz0Fu3P71Ij6reA
woXf9jRssi5+swr8Po2NIv5qK4YSM+tNJXwmbmnGkMbyHNrntvahzO8djvczHTGaUdbCSDCo5oj4
lSraUNLzGXVPGiOveLPwjNr7phNNGFixjtQxugh99tFoGyIF2duvFRvBFp04TCKzMEKuhctkUDsv
sj1dfBQnIChADrIpIIHRT7k/CvPLK5l8rF78thLMeHAWnFix+ZvNg4YDBOyFTrrj5QU1uk0C6Oi2
8YE5Baf8TKwbkyBmph+dkH9snEUZC9bp/R2/A1j7iJVeE+W1k9bDG73TUduRZ7aRZT2JpCCec9C1
OJfgiiKHxlmDNLsTFbaGCLJq8za9oqc39J5VWEYNEHyuw3UiAWsUGXMiAYdDsftcxp4Mro6GnxxW
K0LWYVIF3tzPApq3oQXmZM4v1qsFB+FpBZQAt5KlVOID+8paXPP6bvlS6RV29S9CFo9egRYoXLOM
0SDK79ywAZb6U0AQYARdEeOkFY+8j4ZhVpvgTCJ6SMdjAP/ZfeNOC2iBXPhQa68pu4vgym0JPhIz
FwR5AoeIWlDkHTGsXlTPXF1nma8iWSNeWC7cvO0MgXX5Q/xTPqhDjl9vcgssvViztlbxHQfyFyKi
tg/DKmR6BL4QUVuo2pjzAutSatK+kE6jcTKARWpNqIj+Mrhg/FIEGKSaKmcAnc6i7D++iQG4yxuJ
dh+iDzrn/oH3sH9CVUhevP4ZKRgzw7CKacTF94ebcaze8RCduOHpBCdWoVHcu1Nuuv2Om/kcv/3K
q2Fn1+bn1BG7NMuvClyMXPBU0dkZQe2TC3JCfI6vX+wi1ssdGMO8WPDvcxDCzWuhNLLxv5/nBW84
j8y9/ZJHkKlUxPEwgbCBoSvMTrWXDjGLE0csJY79AR6fOmR8Ndh1RvTh5BfjeaY0hs5y3HgUNI+/
Ek5qEE2/DYSFwhJgnZcuQn8yBTCZkvlwZv8jcOHaw52D1959d6nVEd59h+9fXi5Ucct//c6zalAw
4CvPEEFY1cBpuIAbRwII4Gp+l3jiCyb6Di4Wmc6uA34HpbTDZtdr9Dz/0CO4ji0GCa3R+uJ4pej+
ZyTU61vlAl23TzROBa860v8beW6yMbx1n69x3m57dqkuYdHNsWWFKrFZ+JcjGkMDbIo9MF3RHcnN
xF4mBtNhtAVwT99fxUDGT389AqdVO3Ru8Gyie/sNpDJUQPYUm2sqaDoJmA3uWrT2SQBBsiALZGpX
9oOMp2mCoxK7Y5DyPEE3/Krkdw3mRAvDxpuMVObdDIzmxYJevzR5BkdxUuIvnxxX4CxpsBl77TB9
uX7PaVPPYAVn8povve4lx6OG3Yc75oqZZCNnxY4kj3Hj4bdJWh74wZ3aYZwVLY+OmcB9ETOZkorv
Z/2he4t4EgHsg57nkUn+Ms7w+yBkOL57giaGQ/Y6atArNIllyvFEbc0HInriCT7+B7oOf63akotM
QyRfAwBYKles6QGdP4L3Vw4HaSnceFxcfASYNjhZ5lJY3yVykW0hgh2iSymLI3pExv+7oOBcC31T
OpLVMb2p7DTTdSYtYmF20iKaCpHcFmFZilwcr6tH2SMGsO7wTR0dasQo0BjnvwLfeD8X5Czb2n0k
a+7I5lmQaZCUH0B1QG9usELyxgRnj6HAe7ZHjAks1h3lDL/1t0larDr0nTFIWZ6Y8+6qaN+AR/6F
CH479LgFIWnlQfJRASi2Dsbbderi3c+aI1XLYUYjiU4bZ4rMcS4NTWUO0T7Ox70hzj7BnF9lgGQJ
5dJSsx5S3FLG1qs2hFfmJ8RR43B1qQcWp8q341caqGsK0RgaSN7sKsNDcF0jKUimKVWniQd2Zpcr
CDSJyL2Xq7MwSX/MneKHvStyxtbrcnLg72XAmYwtq+lz95Qh7pvShMN/0oqmEgWqSJCUB0rTzX0/
XPQ3FBNEjqug7kcbojdIzBVFKHGPu7t2gjWne9iOqJOpZ/hLXLo2js3y0i35PH5ik+Kzi9oBIn1E
wqO3mVCJExQZDcm7mEJudZ1VRxw5/w6edkqBxkJr2ZaykqamgOrEbS0Ef8b5sm3tsp2fV9lWUEEX
zYWccnzmvUeAIeSVA0kTg7NwDWk1X5NKSf6NDTaHEgNXImcW28V7kFUGfSfGv/C/W1SvKHrqWqaH
ifHuBZTJW0+i+XXLCcDV3CqYObuUH5vik+ucVDA460dHHx1F7rPc1KfFetHmRVNRbO0TJ9t3dmYR
RUtCQvt9VT+ZqSg6hYoKYqfS1RkDGcIMBtiry2L88zVSOugm5BKQZ1H9QxOO+jlG76nPzM1pCXF8
+ychLdi9H2BnQ9p49KjCXgP25Q5KPH+A71armjoHt6KQv1/zcIhpkr9JsPffgxiJVXcd/9f9yRhy
b/+Jr4jpmQ8N6W/2UbwvZtZ8qhYUOWzLXP4eRjEkz6hjv55R2YCcNFJn0KjESFKvFN3AYZyeH7zC
+5nXmD3pT5ImacsYn6k3w00Ug4wV87PtUyqj1CeN4ZLqqqe4Oxwdr92kJ8GHSecpJCeEoPaHkcJL
/0TwcOiKMaEqvFavLfFxLPbThL6lAdrEhXlPO6ZTIIQC6/4ay1DQIeiNthGJqkUco1TNEIcWRdxd
VMDXI6N4+l8P12Ccu0FAZJy/zTrv/98dNX8J7fskgy2CuPf9x+vuyhaOvLFsIqjNtUNH9OChBAA8
cEbVRKMGXDSDi21/iW8K0UbFDnJbAZSXXef2STNG3vMlYqIkb7suDCAiQjSONpn23AN9BYtCTPm+
gVdG5S1C+zJ6YdtnX4Zq6j/ValVFvDUj7EzjePCPS5QWyjcGDyajZcXhCu3qLfMbUxPTGM700COk
9YjvVHyTwZoib7c5TbLcU9lDMR6N/2P2GRIl8Kb4yCNj43zdUjzBMzyfj2YsMUiaaeUJ3YDYFPHq
6DG+loPq4U5CV4JZggHTY87tcPK9e1EYLnQdyH25lozThrEtLgeLaMJ/epWQBxTq2EoeLY63miEh
fpxYei9e47M5d00Tnqa9gnZebfhabXK8RQ8dQLS2cpVUa1HTS1x7zlFVAfQKI/H90ZXTCzKBo7gI
Npli5NAJon9zj7mhOJoFGRzO/AyzHdBxDMZ/FXGDBNxr7b1+7QuHbeiz3wGiAJxQbFBc9RgMtQsb
ZhvMIDnwBiHJR3EUF4jJ1oVsGIedtP2dLgwikZzzEcQxgEoO95Plj4qom1sAOwBRTdDCMPW0CVR2
0/2ZQCGp0lwJB1l75UMvEWW/5MLXrp4G8L4I9lliIleJCraQULveuy8/GMUQAGnEntVEBpU2EYwv
RUM+X3NsevGf4/N7/lILfdCBPkSV2CqssZhYRtkmV2rFG/oqDtFBHDNcofQ7MMXQbKC05rUKFrRd
5A3Mszilpgi9Z1CAkyp+UhAbFO2DwBupwdXiPTTtPh8rRSYeZ3zNuSYk3eyfEJRiG0J8fVxQA8/a
TOtoTX/UD/xAwgoD5sQItE53guY9i530DmHEMGXQ2uJI0VTcWSBkAlvtrDJqd5abjlmbh0CioLZ7
A6/CPI1Q+f5Tpz8o0wE2MCfFNhXDrkIaaMIrrOTFDArWLuthrYvv+9CJBk93Cu+yi2eeEDS7Spx0
T0Ey9GZJ2AN/wp9LVYOPePchCkF1NRVNsdgIN1SeJ5uTWZewyoYT0Wzavk5LC+qt731XQTkQ/nMB
2gCpi76JiU2ZOkKX4O3z83oDGM1hIAaJ73LTVxjm41jl8lXU+4fKilFdKUnM7OosuY5pvDo8GKrE
VDR5H/srimP9SPDCcKOegbEQspGmdupFzJf8nycD39je5+URRsh77Q+B/TIABwI5woemAe5G46ZJ
YBTpDm+z6Y/TMN7flZdsAGtY2y0046/jUNfFT9MbUrt0JST3n8gMVhv+0/o3OJwEhLbw1efxLURi
haw4Ul7KDHYb36cZD7sXa4bNOvTvwkmCOgtdaPdtq8B71+8Z/+PUB4wydSBuhqW/8blU+iwAbkGb
XmBOnU0W5h5ZlJ+XAXWZWY1I0XQbyu8o6Shy2sl1KNL1SnLdRlYanL/K+JEJBTQnTvXXn7FbKZc6
7aL8C2Cm8Qf1qhibYKVfVvzlm1QBmeR32UC5crt70MEx2p/tNdCuEGxFKHdMJXLGhC1n0ajKbLQ6
fB/k45q0NbPi1tplK266R9dYMJk5pzNt6W1cUpwfx0G5aXKdsRHuexpRTvxIjUbvvHUZNAOyBq/9
YmLfkn+DY+QyX7PuvRtQ5THhe6vS8ksXPwO2YrYIIB7LiIW35ECW7meSeXb8AkLKUR1TZsyDO++G
4pws8sSPGXC0EQvnp2hJHwh0bULLN3bvIQZGAFdTUOqUeT4dtSsKsiKdfxEfOnUUsmSJj+lETkQ2
vRd/ycBlYc7myxmoH+IP2ZPnHBEHajuiFLzBdWvaUtdAuswtHKYU3Tu9J9aq5cEOPq5WiwD2O2d3
JMAyoYfhAIkNiraV4HujvNU8koJJvasqjWTHwWL8MpZx5NahRNinn9ByL/C4wJcCzDkCEyKHJPtO
URZRZgmrSV4HLBtuNLWS1t7MkbrZ20brvgvkIrMQEjDpUuCGPctLiNUMH3gt9GYh5Vg2MalRpJ0V
sQMx3Z0d4HQPL7uMmF4GolFxVLDokHI/XMgH+Xa2ij3ICH572jMhTGNOg04VgYTG+GdICMGlT8U+
Nvd89PWtM9dxV5R3cBYi5mSgU9b3RALKPxn969wz4519KUDDxkl3Ty8eX+FxDwqyKVgv5vPlRzDs
wbQysfTMACJvJk1GpfZHINy3dbFbuGpSNecdVi9odjj3XXu+bycUdzNG2lD3LoM/6l7LlR/QOft+
vbcpJGcP1xpjRKIWCJVgG9vskQtJLLDXue14cSd2cv/a6+7w7+hHQNla1/VutimBbNxib6HC6S3P
kJ8GUTzDWe0SqmhqcRdeqODXdth1bPVyaDXNCYTB/BDUoxU4KJugqXz6pTNrd0f2HWAuy3AGK0qA
hnyfRIoChhBo79aprJRQ1cdT8h42nMl6R+E6Jr3Hw64ONCHO7wn1DwN39F21jl6Z3EqAG04a554G
b6Gfu0NM6ZtGWWM2F74R7J8KmzWQFI4r1y1ShhGEaqu+XuhygONTuLn0YVpHUn0FPsHDRsXZNRcA
FsC1WAV/kLcVBI9500OHbqCEKCSUS1LfUdBZVs+Uwe1ls/kFZr9cL/Qq+yIV0ACbDC4ZpuSVZCMy
qxSf9wgt98W1gFSaAQAdB9T67dczkl45OWXTsStsS60yaCpb75hHl8zyQYeU+61UxaDMOEUoJezL
vhl79zTXu33p39JY7079zz/N0o+DYSv66J2nnCOeWxNFzE+QVxAlMhVF70LViPM94hKXimFt6j/n
7Q0ULwgGO6H/cFVvc9TY/z8Ym3uj2LjKH1eZzWBG4CMkpQyvmZbAcJ9TjceaCGr+Mj/Ahvapme7C
GOiNDhCyuBTNBUW7UuPhAg1qbtfA+SYATx1lv3L1EsKmE7R253YLjlMXFI0foevwBd98fVFgl6OX
go/NauiuRj+xwqsods0JIpBDnAOqoMVZqCdbqoQvNpzkVGpeWMjBfjCT+AQAMEV439ZUllE9st+a
UcfUC0yzfYFYajiT0D5I7NkystVBBo/+6BL2jASZsLshr4QITOuSX5hKUOJa9AVgs/kDwK+Pl6uf
lnK6WTo5sbC6xSj2i5yzr5IRznVF9VZu3dIFBFXvRBJbJTqKgllVQkLlTray49dY9EIlfmNghztt
oWo9SBGANYMc2QvFhT3P6T4NzWjSqdY5NmvkyPH6692AE1Frj7814LSzmsoabzpYB9SjEfIzzDm/
uFTNU48ifoqG47DhmwTzI+bP4vW+EUfDIFtzt1HMdsM2pS0cFYZVK/Dr9kyqxlr56VgucCkYGTWH
Uj6oMFd6fm7SjXwaCinawn7Iq3iOlse1tJdREXKcPXe96kX7V6YjOtrO9N4daWbEqHwdxXmN/ajv
gqU3N4lsK5WS5vYWu+YjIFtnp1dR2pD1yn6UJ+LPvyEznbCPGfLcMK2pcSOhk375MFgZHnFyohbx
dnWumeNz9niNnPlYP54BxEAlperWtllSmbR2jVUT/mxBIRBzGj3E5ZKlJz7dguPeb+Y4m2BwQT75
CFhbJ/s+bhzyb7MgV9/tQMmNwt9nkuoS6NHVA14iTJpPI6dPFgyYJPr6BaquaHzN4lvaa9wIr3ty
uaUmXVFm9KyyVVYcHP5zG2/kezTgFA7bSkdL352arvDlX2hKHD+0fIintn0kqKvJz4Xf+Om3to9z
d+fFuhBSOuY6O+LOBHWTB18wHDBB2xLcKPIal8gQsFRq8JfuQwZvy8T3SlJqti7AKzFLctX5FAnl
t+iIGJUsLXpwYlimpanpb5C7i9TbMS6ZHluSDqzdwRohFWUfglxDDYfJssaM5KseTD0/B0RGDFDS
Hhdwr2DNGEwT2svS8WwI5UEBj1XPbXvqbwMhwiq7n0IiXTpLr12kKiPh/Mw/jDuvP0mXHsEvaY1G
mXGHK5+HC7XXvwzHD+6+eCo1X6AZT2SJKNh4l2XAa24bmiykk6/L3DHV3GOFM1duQmkzfag4GBDy
QS3XmiuL6EOkrBACcdvL/n7G1/GNmDPUjznA1sMwC4c9GkRupw7xop/el4vpefzpb/M6GuXabYat
BVNg8XunY1pw20kuf3N4/gpQ4ol/Sr8ZndPxreR6NttBZypDo8n+0+uk9xBkZviG07/gCyK4bz9G
tbSgB7jes5S9S6rfVIVFPp1AXTq7C9iOvSM9j2gLpSD8iFFd767BceeknkqbDthFpnix6w+UGzCg
22dOfOd+RkPei3X/Rsy1J5DrHHmk6cfpfSHfI4J3oClRZOfGmzB9PthqV3NXopEiJG6Bboun6dpQ
KgV+YxkAYC8SX1wfpUvj3h/UayKm644PDf4IUkjThJjfkhHhhz9cYlOTrlyFd4RQY8qOmG6mNYYW
T73JcoB8N5y1GGJlrn+3Cb9JdyMnoxeILL/A8z6D0SkpSujcctZxw7ln5KOxKg7v0cjCDcnN3szB
bz3Wx9MvZl7UoybHtK1XUNaB+AVqaFfCNp26aKEiJja/SQkcf5xPopDRoxHIoLN5oI43BhQoPufK
neyL2DHm1gPNz27hIWtMLMV7tNV2+U7qi9FFtTugunyr9o/horeuGS/Mw5ZE2DYlGjQb3URqrRKe
RxGvpyJiBlXBDQDhuwHIJymLfKtPDs4CIaYAWWfFsCRETL8ZtVeiaEDix24I/7IRPUyOPo6z1OYF
EGgI6ofD4VfAA1MuKwAnzwRm1dLhJlZK16DgL1jpzsNGgnMN6fucVyzLVV/rGOlvqHTiwsAQX+c+
3raV0XU2Ydh4RpHf4spzXODp0ETEstm9/iyYUv9jI6JADEYSYM5HP3vAwmnndSpvGm+UqvnLeKVU
2AuBgyXt87a+xRp0u0lWveh889Joo/MWQLov503M9jR9S+UbOyUOd5sI6PDcHE7tYBTXrJs0qbpu
T+itWwCH8l72Z4p9BEAQuxF/GZ4BlcXfan3wdtioofjqnxSZobtTAebh1FpuLRFA8weoRuXMLWUT
hLEtJ4CWxyF6Fc/MrB5/4DtLPwepzHPTTHQU+hP6RMoS4g61UfQy6hL7JRPr6OPNHYIRvvHBUBpP
RL0MqKw2lxN8aFbzmJvOuYkcBgZGTqu7l6hbgxc2bF6lEhDlGveC4cdGBB4J0MxbkFNAQ9gmZXrF
3fOeJUcEetcNSrvYdD590qD76ndTlNedt02bcKmR/3K0+Zo6Oan2mXZHd9TEyU1Ma0I3FwXlDweM
KCCtRwoL9PSVfoRUnBePZFjoQfSwmwLSNq49aMfxxbomtx8XdHDDbec4HWZlGBBeu+bjdbbNPzw5
G36oAY2bj6NaZCnaeGC/B/R6+QcHzktQmhCWSx565C6M/Muvk5ER3RomMWf5WuqqE6+ycx+s4lSl
lVGRHb7vqx9I3SnbLa2kMxwtdqjFqzBAMhBWovAY1WJRLZN4QQ+6wJLWhEtNq1iov0wP7PaZU3nb
mZ4b6O00NUJc7oetOiS0vh83NYBXEdP86zbsLcMflV6daGpxAf1h4MW1bgBTYfbTaAoac/1DAYLx
4wZrYq9kHrPmkOiVNYI61n44s7knnCFwOfe0PhFokZIhrDFUQCyD9gvqwMX11o7q/ZH7wqaTDr0/
hNY3Sh6GDTRO4BRBWaIFM2EoJG/mwMtK4CDiUzv+xUOKrDQJHpqbkRmsc1IAEDFmSUHVPNbGBfjk
tpmtBIIowFTTxrwJAOfZAw/q5hLXIkWWusYDonuRvRNHEzB8dHb4T4MvTwVwKyhBq15H674Gzq65
oKIcKYTAtq1Adhpf6FFJfW3Y7DJX4n6WH0maNC5UZWSntGhASKmy6qpPs9+cn4CYJ5IpL6qUAybC
lFFMYNfJkWkhJhHoWe2Hr+395qOhESm5YJTgwcwdchsMZVfmVnofY63vhTXNOTh7/TGcWda/4+4v
0O1OJRjnQdRZ/I97Fa3XajNMGkIx4WSEjexgJzN/imP8PNU4K97okeet4DVc7KVxG/wZbJmWtg5X
WwJ8ydYDsmfOtA/FVrkmwvrSwsuLr5hWYgztfvr/MDqbcPGLrYANkxP8neTGmq2At4Z054kUZdip
cucMMkt6n3PXr00e2rz+sEisuoyWQwLjQRCzZHL97CIO+KzvA4yxh7HKdDYoRlR5aLqOxWTAMdwj
KSX3LNH+p+RTVPyItuj9HOXav8RlSPSUc2bV6ntV7pHSPT2F/gabhDC87NMu5U1NWkvHHSqYXEQi
9MbGdA8iTQOfPnE+xgXM6RPsy9fW71cZXRFrgGVmEpL3WnW0s6J/MRoMU4nVXZ9Db11RA7yScZm0
0vSBZyGHyUb06vBUtsaAkCLBEZ8kH2+71nbwhmXFv0EubgaW91UXDnussF0hyVTqe6oO6qkxF8G2
hOAxtd72l9So9wTMpedfre90MxAGC4dyqCgbNqNExPVWCBMC0Xl+HrMJms4tAEw3REZ6/yeI2vUv
co18NR3MMH9AwJWT7ZAbmsMDkR2Uou+cCvBpbPLGNGm/sBHICAaCto+ucM2sC3CHa6tLas+J5DQj
TDDAaiPyswDDTu7FythiTHGfqO3ZzU8SCgcjsTo/gtZdXlx071C8Tsqg9GDRQ16f+EjV5QOFL6EJ
8DZCh4FBn73QPcPxsDv7xqk8kDKvaa9UKmf8LIpHqq6/oXYCLeYZIFr9oBAa0YoLAZEh1WtSaJGQ
32WYh66CCHJwlCW51Gq1IqNQc8BgWwEkXu6DMyR3CsbPnRywZW2qZYVbC2Ekb4v5xd7aD3CTcdJR
idYrtjmeBDGVJgEspG8hCf178zOD9cSW+D+ylI2cGmN9ToIEdtYwsltISkeiKMP+1SBwBkbXXbOj
dyVnfVDHxP2PNfm97n9BfromGktITVpHbQcAzpjo6rLtdLV553v5ftzyqr3bpUo0ZKsaprLkeAvM
sxxTgWhUTNda7GNgyo5EAE0sVK8bSvthHv7NEbQjI/Bla63YnGIZ/EsSnenkCzK/cMvt/QoRlO4V
eLKJS1Vwk5F8j3jjLUCOgNbhdbdYcpk1mDrW2XvAuvt3ZUDOjx/oX8lc2uCwa2KroSRQUwTkAcj1
iayGD627sW0m6zd2jpGLqpfCr0xd6qHXdI6NO5psjrFANpbS9YJd5vXSWQGWKzdAKcyzqmO/ekMA
RxiJmZCadelXa+/RHlmoERPVPq5fADfB2h+SjuX7ndZSsnpH6lmSTQF8uY6uxK3+SpP5IajXwtTb
yh7RCnznUyN/DRD3j4wB+AhouSOBlPbh4TWXJjH3z+3NNEMI/Y2t+8h1ibZQMReyCKBJXMfUnfj+
2Bd4FGoYDPsBqEeE+W8rwTz9VqOCXWjStoq9gvZZOw2YjW+gv9KCzDN8wGin7/uqAeAA12GAJnCN
gR1pgdfkRvsJSuOFQA65+oqDitUafcGRdybecbM1e44ZZ/NLYHJXOrQaYqQLHuNfX6Xr8IHmZq0F
mCcAKUNrBEpNI32QHpuRZIhzCMnTea1bQsKPyxPf0dMuoKZtVsDH2sOC3BhtSWX2O0+2vcH2+Q5S
ob0VWpykiV6NMF+dDRR9xWPjFS4CGLdiqFxfDoGk3iCDReAeW7/e5mocQhEHGyzZFnHtttadF/w5
aQWPHhEFa/FgHYmsA3mvKFSe2sQc85bum8vnA3HSM7YGSSmhdtDTSugPVJF2qHzzNdh9+xnn1ae1
sZMsrehV6AWBllcwvUC1OKIe7oWfBJKlFel1kwYZVAz2XlSRZsD7RpyXSg/kaaRYyCzTBYMyp2lW
njtHxDWly+PwHjSMHmmE2r67AgWGC65qUCVHsLs0yVVzJbH0001T30YlxBiUZN1Ik12RpuUUaFXZ
0nIoi9cVro36B5biFtkTPmSJnolt6UkiC0yxyyhlXYzAZ22v/yshtLybWihteCax2ylj0/k4oL47
UOOL3Ojex7U0sjm3quPaHNCD49B35z3paBRxgusfZwxgmhn3o88V8xp37PG+xQwNBY6IARfImsQ2
C/b93oiS4HesJvKe0FmNvU/T8GJzkhyfoS0d/CVTLvkPZ02AP1dimkdr9OotEX07qCyIaWTaoU9u
KLv83Vy8lbed/KPse/sG+cO2WBYyqSl9kXr+VLVBD38kO/raGKh8WHpuHHXr46AgXDonYZQDZ89p
lDqT3xpuAX31128VGLsD5s/3uyhIc1CGhANdIwpls5eCt7FHDLhgtVsR1nTgBIv76a4kpjP9hbYC
CRD5JxKhvmgL3Z2z5hVnukkGo0R4HAmRLJ+/swjke49YdaM/iNoNycNYGlyvBgrMmso7NZPjOpjt
jO6JpzSYq9+jRhgf1lYdbSZhkJs9y9xTkxN/zYHLDBZoR8PZDEeWgl2kQxx7cnCnJlfEs9aLzaQG
6HHB7d+LvXKOWR/B8qetKiSOcb7Zfv8msKxcTUbKzrR5//a/AmTp5hY+MIBZn4+ndMkDApwpgcG4
fKgSrzg0ktccLwwHjpAgLLpi7MhYvJ1ntkMBFwhj8NAxTc9USu517FiXUSru9JERoYcv6dEBWpKK
8schu3jiapoaawX24pwxHpfMybuxZRemUv7aIsGVVg0ZdZRxsQm13XhKUSt69XafMINDF7PfSawF
sKxDv8kxIHZLfVurTTl7q8s6RnhbGemB5Or/3nZsWSCA3jWtpCH2hM825LO0VOzmh/jkw2VLs2Rc
x1HnDLRbsok6jqoOcNi1NQWRN+1Ip76YL1JSd5uRiPvLR2NdosigLxlJGEDKu4XQQVrXp0Dnp+Ew
1JgHp90SWjQc4Nn7b3lMb/EEv57ZEzMpQKxIujYEk8WsyGaOqBCH1JHK8WeWqb3IWCB8Iadn2Hod
ZjGISkApwyk7xvhc95xFbTLZyiNIl0rzjwl3U4++TSvobH6LGLYLZYKJ7vMhPcgzX/uvwg1TaWFd
3BALM4Y8PUbfqC/t161o2DHMZO0C3MaboTMOAQfyXiAw+P5NHfxnzPXGXzFzg+mrR+NHJTBk7qb3
Eea1PT7J5z/Ia6ELP8tL3tHDM80SScFzKrZ0XVvo5m8KM9FPay6dOr2gkV7PGX6XAM18+IWNqCPf
16VJkbYn2Q2VQqPSzS57BxYzkAZiqafJ/ftrHaMrVJ+cHqApgiRUfIgUp/qruQyHiwHtBWvQboTa
s3e69qmiPI4fNqcU699ka47QWFYT00vCJOWScQQt0WlGRGzvNeR5cL+kTA6qPe6xcv7j/qtbjilL
R7BbJx2CDoIdee8Tk7aJTZWJU2x0X0NbfbGWfvLUFK615yIGUhmcjBo2id45XW4+nhwYMLV1wkEi
xFaustODbt3YHem6BIXXrWvd/SGdgmm7djlCQPE6OjphZuZ6lQ9ZpfNQ6gseh26Lf0Gl1pRuSbM4
Wf2nToHbTFBCvbxvwirbB9XpqYagQnG1j4i+hYP/AlK+tfVaTdb8XL/8QidjBlo77fMP7lDFv78i
vTtnubtPkLbcPZ9/3VeuUXwI26uqMHMwhB43kBXw9q6C+h8AfoCSW2bBosvDtjOnuYdUD1dZdy6o
RHAodBIE8ktCcR7cPK5G9j/Ad6vB9VW8xrgf/JGoRFb4wq/z2Wld+qS9GtPCpyynXu8CWQ4S5J4H
cPVbgwg+Yg/bPvUbPvuOvoj1U1gBXcbpXxFzvMnokB754fQ6qG9M/Juje2t3romuqiVybMulABmO
kAq9SI1uU3abYqCpbv4HR30MRLM4rxlAbAMLEjQSRrLHlIIt3N66t0gI1/i0tQ80l9StrhuD72jA
+sjx8822KFX4dPaSwCTHlHHRG+1pL+AH7NKgWr/88Yz6QF2Oz5L4UiXV9TLE067gmnghlAe58Om3
k9sYakYW0q29PkKDP1zlqTomcny1Ajywc/Ho5194qXevHfV1UCgKYGSuoj3Zy4mp9NIvvjtp9omI
ISiLzuN2yQdRgQ3w1a3ltVR5eMGCow3vvD+yqutaX4nZDkUxw//67rwS6AeuDwVE0573agzdpKqw
T8v52IqSAPPLt16NC8011ako0ZCGnwMRGXi/X1OAlbFNpbaLX0VWlai7wtt/zpluqEoEyhjGelG8
F7dpQtwd7qJLtWQFKiAnR/+fChtwh/kMHozsyh5G0jVIaUHabNSN9pzbcenAmZbhnPqa6J9+Oc06
qFsVHHcQhH712mkh7Xh9CNtx/8IE5nAl2iNqX4obllzcvL7gO8RuIv7G5TfFZPkdibomCXwIcIS2
2RZ9hejdUX6rGzGFTq4cy+Ko5ATQoapH3t+5EB4OF4Qsf5bcXoTGKfkrqllFZGmF9ohnaycz/1tC
VP5pkYvgmska3pIbOBJHNSpodJpAHifg+sJMb3lWSxCBOrGlJXYd5br3t81b9716qnPGHzvf2krh
X2lUMDjXRWP+wUCKlvN+O679ds0SDNcKM+nZkmMsJFCpHwOn7WG4XgwpTfDTOzs9uHxlzeaMpEFR
YL6VNo4JUoXeMiR0D4lj5qVOTo9PUYC0HKT9xZEqM2VOyiygNYjVOZMKRzNDmgToC3QsVmoeIFmu
X83ztZw19iceQxvAZsTgtk+ns6sUa2NT2hZr8PCb3QAffHB30zF0yIH6aTKl5xccRm2ngdZF0n91
NwLkTdF4OItUL8Z0hy7930QXy/+XY3wt9378uaR/MtaW+VG+aZ+eH+TMk17trsdIy+nrSiclhljb
orNv8ZFuvdVaG3vQwO7rg0kSkGnyRyvDFu1ufmMzH7K97R5JoPai4CclI+yMUR7ntrFNO0nOtA//
qLR+ja26V6rPxHsF0Dddsbvm68jJDYwiSL9NtSdiBlFMLKhqF2WS7s5ZRJLpnauwVrvTRJnxFwkw
S4dfW1GYvJO79VVGCkYF1kHhiiOglzBHUD9Xdgc98ZAq6yOURsfz8iVR7FKL3R2rW9hvYLtrCmwL
eWhLlHezEGyyNLNpo4FSSUdgNtYzvNXjlUW4K57TAEt0/e4qAmIPr1BeXwPcbGp+JOeR5N8N+4Q7
iloYtdRBO43YUruZ7LZb38wYoErwXAKhDMohzfUf9wN7tPrHB1Pg/+GnjcUidAlm4vBPz3ngxKw/
Q+moss9kyGFa7hVz56Z8n9d0uj5Gg6iWvzt/BiiCsD/yik5ed5d3SlyV+bcw5DhB2nhX+xLT2ruY
SqBu+6/mtLViMvJMDwPwDQmhCmWrB8wlhSBhLz9LkHNE1X7TyIbuOtoMaC6ZWp/kCMFK1UGrdP8m
OeAe/JLiAcACj5FxlpAdPaMnihomDV3gytkKektJN7Wa7lpFdYwtBtjKFiCksJC4BEASpWNvLjFe
nHMNpRlBr772QtT5tFFk6CbmPHHoGvotnZwjbCNjkL/NzQW1lLNU8ijPLnRvfnNF5wXZSKz+bPcv
BhbcLKSWqnDmLd3qdXU898M/4ckIhyGC5+RJAwEDw8RNyLSAZmivMcb6wvwB6zPFHuez6JEjrdRg
n81c22rtYYu7vMImVRcNhtOl0Rz3Unmd3iAzG4e58Kirf7RJ9coibnxfypgO3u+S7ei5a4BUB/J0
eZsiHKSFEdCf+oUk/15TwZVOlwx1rbuhQbC2rP2ZrwUr7KsIAb8EJvvxwvBASIylMWXYADo2MRRD
XaN12ANQaPvMUXuGYx2hvjW4/3NZwKUeryvALcMICu4LYgr95yu5dQ5Q6v5edeVP3L2uo71Kypsl
AHg7yT0Fq8Nf9GnihpgITwhd4/R1mq/lgUe76f3YBTE6i4FFaC/DAorHWDEqMpibl3QZWl6AB7Zd
0mF7j4MEtV1tLJWUb6iGUd+I4UbLOe/6E1Xc425pr1kBFI+hD82WhrGGFuKC/BExnVRq6ifZv8pk
Mpks8CZwg/2sQFolsOOAK2k1OBYPA2X6u5MDhdI+AdWpWuzFakoAzxfERP4wtpmcRxfB43PDWduK
oe5yZRprEhpSxPwlg5p966QsTjkZCW6NQZVNn7JXKZoSGU8C4x3RjpecuDVBF8lIbTtSU+BUK5tH
lo0pkFz4pVr0+kcfZtxkPGXo8GHMquKkjZwMfvgnDhC5VGe5vxCKnG4OofIKC5Xt3w6OWDigvTv8
sfNuiQB/vipD2eQasMjm09CTuOs+GiupSMwm0XOo2ss/vA6fArTTcu3GCrLeQ79xJO/Fq8So+ve8
9KvWpBkKfP5mqLZlWMn1r2XYTH2/Tb2v+mnFqAG8/gKknBHMURKMPSKRhH/WSQ2ueDd4SWRfyVtZ
zdLie/6wy+u1KVBQs/4AwbjbgaqhsZQl0tIfBoZUJg3S1tGWjyMVPVdDW1rSQMJTJBagmQsKgbv3
ah7jGUWsUN7lVn4g1qL48rf6CBv4LpOWZPrugwQlCez+fzag8x16HiBWPssNNfuPE7hakUghwSOL
+DDd6AYxKTECtEleB+Aug/WtAONJ4O5FNFd0F7qTDuKkxf+C8fvb67JFiSb0/hR86Vxk0q3l9rQW
wWgIcX8uai3ygxFmK1WytKOxTj+yhnhm8/ZzSAg4eNEa2+bc4Hvd0CrhCx5m0YQFCVfXg6/HCHtS
UddGQ8qH7ASinIydh9rMiHY+eqN3FpHn8BkeDqUVT6DHn8wmZkpBVnUkfySlR/y+UBFbD+Yb2Oqr
h1/vTkrncvlaOm0UvcrJRJCXc4BeWlJeDfwsCpJi3FEAqcIEeGqKwC6AiFOCA3gFrPC8mMfDI/61
V0oDppsZgrra1oDVq7H+3MoOLYTpK51aWoX5fUNmfN2kDGa4hMX4Gsa6bWzjpwtDRAtBmQZZ095D
ro4/hxktt659vc3YL8e2oaoEddEKGvl5GmJRzHHAqwD4qp9bZtbsqRVpMTrP14VjZUtbwLh2rXUz
mustmYN2BxBh08PIOg5CcVhp5hn89hDdrQ1y6i2PbPtxVBqOxI5uJ3zk99eyaek2/HKRty/9w0Oz
OB4+s2hwnP8GF4Foj5ds3p5H0IN0odarDfptnIqvP6sQYVdyvMC0ImJWUT02ttvwjhPjqEo+Lv3d
kA5BPlcr+35c3LLcWwCyMzLW01Mhe/A4tCv4BsNqzO6qtWNgWTdDDgPRbeT6vFBLqvnQKlQ77qKD
psfMK8rOdwed3Wx7VkqGPH+tM3Et2m2M6ZkEEYWR+/7JB6Hee0urqphAh7khIb4iqMlunWZ3WWGu
y47uFk4XpI/EKWNj2Us/RLLHIlKRlrUh73tk8iPL054nyO/u2lsEzA+RT8fmzJuYLxh/S8sh1WkK
hkrhtn1qbGv3qnJYxJTR4cjGd942JSFK3SaeGA1fDETuxHakCnmcK7Nrdcqmf8aXyenTTBFYOwzC
MekDdgpnCBxnjkha5AWtCMR5WhG9FZVL9hFzg6LaKa1LqgBDaBxgiAwFXMH2L7tV/4KLt1BUjgHE
ZOrjbDQoClSFGUO4d4crxQMkSRnl6C/Z/yb1RFfxKEJZJrfk95CAjlqQiyzR3RapbfLCVMH59weM
fcerEeclWUk1rogjH7SduRrFGobhGh4/GFApZOk6xkSSCqxBbH8ED8sqj50QQt1wkg+D5QZ0npaz
pKmUqZE95nkOoQ9bk61rtzdl9iybAdQUkV0yD4K3T9SOxj8qxKKsWFZIPg+V2Yf67GFPxDQN3EA/
S9Lq03xBu5XoS4kjU+tif42G8xJJcfExir4kKy4h09Frlbf7fsHqQGpG9JIkKSyzJJ3sHqXsk4G0
+OHUXiP6cR+j6HXddym/Vtka0NSHPB0ZNqlAS3Edi0nFAJoXruuapUKaoTUWmPLTnHmuTFrruqxX
LpGLGYvnd1lsVsjYfqVGve2cgyaMvruK5hH1LlMayYX52QaJt7aSLzaDvTHU8dCb9IigLM7/Fkct
5lMQKRpKLXYzbsSpAuXwKq3mHNk2QvOSrMbjdy7QIBXwhZTAPwrvghzfS1VLzhsInAS1lrCz9ne+
AiHZyfFTiO36650MQHFOyPeXrhJug30OyWSx43nzH1f1LvcZ4MygCA5SBpTDVFm/zX0OHpJrCNLK
0MpL8Xq2r6aUdUbMM3Kd768L52TMItdopc9b5qiox1gqnVnhIlRP9IjyCza4yYVt5H35L02JAHJ6
sJDSMoKthCJXvnOIHyCSBqIM6vsxUKPANeTFO+HhY3cajxf3psisqLxX2pQDKuebU0c3yFSXFvtn
izI9TxkOo21NQP9A7XZ5jKzO6u/MWprKDayRQzXo+SMih9XYzyYsgS14zUYRMwiLlqXz0S3fYM3Z
ZJbqrkTdLCcRh38tVZ4TjWh8QipPWtw+s0kwX1nZnhTkG9y1ffvjMCvv+9U6/m2JU5AUq+uOLpS+
fZtu/ECs1Zbz3POvuq8Rb0wDZQaoOuyYn9U7Ffr1UuQali+vUrh+cgfOc5PYoOS1aAomdLSGFhZg
OcSA0AU9EH3TH/XHzyuWFc7b4w+piDWa8p+utsTa8va/Ox3/6HFhpB696O/fKLuAJAvVN+mSYbEt
tb5VkaGED32/jHCWiIaxMyiu6sIq31Zwsn86vsRPQrj8M8MzU4TRliPHayKHZIilVlTnWem4zwx5
ZfiW1U+0UHptMgB7Kw1tRwX04nWAxggsg5WGLTE0p6fgwopu0xaTgv5wfM3riJ/uL4oejfx4T+ws
CHTBROpJOD5eHcK7EdrV/eEsmrsAcPUzvVb2RFT/TkkSRYqvWjFMHMrtiDOBAsvs8qNDE9CoQPj0
+xUqlcWqgAvV2mB4d4+d3TuucuMcLbEudvV1eFt3lzVjl//2FVGWISHi7GizJBFVL7smCL4Xv7oj
W5xrGZlBMDEqYZgXh1hawcWIN/AHBczxtSZT9yqw/U1drcG5qmXAKkAd+oxfWFsd+PaZRKmDGJO5
hYZi32Mq4zY8FFv9EBjPZRBE/Mzh4cdCuWonfwLz2v8jaLZ8TT6+JfVK+fvV9FcB8N5EezN5ecrM
bXGMvbgcoCadHgpehKTaFIeaEPtoW7pFwAyEgfg4dTCmbYTI6WhIxecDsDyHZLLsunWj6lJv+oTf
TM/AWXhj0NJ31ZrL03COvb4IKZuGA9mYJV6qYc9bZT9hiA+h/9FPgSvxJz5SLMCbrd9DG0Hn8hOd
qE2WQ1tu3YoiExnrw1+qSw0ARixVbfBDXQnnb29h9AkMP3zyxQJY9TnEHUNDmW72Gwx35CiKFPYQ
h/n0Zk4L29H0n2sd2MGxoQ+aoGlufzYRXxJ+41pzF0uNwLxmBVgWWTOf6hakZznpFxUO8BUU51iJ
JQQgjNrsXlVn7ZiNaDYIaHEtEEjFTebDS5cG9ptbH5hj8XczJal9L2+ORkqOrUym0DPCN9WyyjEC
38VRywA9G62MYRG1Kl42hOocijKFBBCzY4TWjL5uaZr6BxVIHSVhkukMdjhDVQoqArJ1GMKHDwgH
rVeoLBRh2vcbDu9t5MzVN1QpxQ0HwTwsvPCCc4ZatOhvFrvdWhCEsgjfbcfyft6IkpXpLfhgPUmU
KJGtulwLxqBEooKrAZK4OPvGiJ9Whco0Ah5Ogwz7u3A3s+3uh2kk6eMMzNEir6O2l1QQfYo9wCOF
IKtJw+HoQqdSGIbkGdMbzdrUWcQDwgYNtsKi1qBkx66dipkhOoFiZ9kiFF0zJbwVDjju2XaQP3IU
4GRjETTR/WEma+q4CJTHYjj8K1Q0lQpyQ9ieCwH0H+NGzJLMC3L+XSvV+JRqZBTBv33pTjCzaTpb
nQdQVck32P6Zl6VCh+/Gr+9F62+KKD57vLDsTWaCnIDJLF7CvcoQXvRNe4raR5JiH/WFprMM20Gj
h4QqVjfp/cbyfYh5wuXX7rkO7QmMPVJDYJI+CoNUFY8tKLgMXq+XpIRxsIAqWyVeKuoKAOWOic4j
U6oIO4PgUowPl+VdhJd3noDcWsW2NP8lEpOuiUvMH4DV3smAwsjDqRxz9JeBBhKdCY6Jmlg/KVU2
z1/UG8wkxaEAh5Jk6FZV0cZVRqsLWtzAGfbEGB/4UbO3CAzRasowYEzTQuqHpiGtZd6gKmfP0Q53
0SVu0UiN2kJ1bXN6IRyH3IgEr1Spj+b2zltkU/2+lrh+ZqqtrOvMOwbglYv2irtClGcjat2PhYE1
OclvHPMvM5+phUA8e+muuggFEzLKm/XrLyOOJ0N3jw7JlMBzp2Nm3l4VcZvOPbuTaUH4Rz8lcBD+
ICoZ9qvsPvwipqExpMyxwHcooLHlOVBO8QivzrDID7HpGK807/3JeT8qIpg7p3ayC97WIFK+Nmgz
LuEgUYvakdjbxxd3jvbUZ38GwCOY3n1il/MlOzGZLxL1gOajXl13lmfxcMNeW1v1al6RS5iGzlnV
1j2KMAtFOJJGqQu1+6aB2t7IdBbRHWx9cZ0dKiwVCRSo9oXwI5vEBXqjVEnkgLhfKTC2RAl5KMzD
wLA5kijWAbRKuRUnLe8/vufS6//O5HVaPtPMMVbsau6br2pX0XGJaKThydpDPXGPnusxIw+G/+3j
stdv6kce/kRJTaxs0PWtFBGzAhPQMJyUrWQOeu00Gev5bmarRuxtxK4xTloDdV4QAUF8orCNlLFk
4TrRU+j/ZeOfVjpqlnvnzBaLoanC2F6sMQxWRl16Iz/kfGuGigmU+zMaM0P1PUJB86u6ahYz7TB2
CuM+YYfmikvtchlsxra54AVvEkRBci4SZR4He8NKg3LESvo4pJD9x0oywKFdjApXvc4lfrM5XpV5
eXTRJ583TeRI7m1I0Mir6Q9kwzCKXtph7fFIv209e+kpZemXCxXMSc8zj/XSx8/hxmeM7RrUYZO7
J+5E+qpwUpwQD20Me5EBpTuwtKj9O9MrvGRTE7TD0EJhp4Q/pKidr5+5H6YyUZlShsVJzKsgJN1W
zt1UXSKPI/zJr1wdo1PoLBsXyqvZM8OEQNUuKXoHxuHvdHFkbZ+lI8kvRFEldCnFS6Wh8aRazCkK
0tTkPf9crqOcbW/c0cg+v+SrvLZfhLtP/BIPwz34quyqr5NbtCN+n/5BhssBzBJx2Nyteo4BKvHP
3ogTchmDPctmgD4SI9a+1DnHWafVvgjivb8vhFpX7NIFbdWL6k8pNQqM9ER5Q6jEnUGJzD4FrW5C
7xDcVRYHxZJBbmOjyD5rmGdPAKFfqRmM+Zx4A+OLFL/UyT+cIpfZ/8CJpCCtsdLTko5+6YZDEbCD
hCp1s6xb0gn3qsWZPHc5DlKoCsVssoi8iCXvm6rKhk2+ocINBz47+gjHjwQyM3NWXkR03SBSJXoe
1KYYuAHmFvUrve8u2eHG/Uj4uXWP0CHujnOXbaIfureKOzdFYpdSYL65+nUVWxIqqb49JfcTdU6o
PFo845LywGaoTK9dyRJr+nE0KOQK6DkBbanW04TednFKOGro42wUWtZAwfdZQwgI9b0/QSzUqKHA
L3WW3gcqpFO5oHcuhsdbtkKVHKlRVflDIQVSyVAU6QvKnS0KnVSAyfQOnDKHMhGqz3I/Wxdbc0aX
L1EQw2q2FcshmxYcxKSOfa/K6xJ3SbJfIGxAkv0z9wpc/e5sgjwuLMAvENKxJ30Qda2PhQPaku0j
iGmttrzEQYDxWz2O3GtS56UqLJJBo9oIry/B2+YbMI5XeRuFPmdh/udSGWGktOHGtuT9HRlUwOJT
xFRz99LoMW6ZF9RGfBGwo23kMgjfKP1z6BLbxrxKmGfa1VfeyegyfcmLZglpppHohQzf7K0IzN0o
Oow01tQcXC4hxR2iik0qlRFAuJqoTJ+AVXQ97D4MIEJU439TNVKSclMA+qpDe/9tpe6zO+VYYVSc
6dmwRZJc9DWBOFS9s3EEQmVQkCB0Gx7HB4ffW/D/1oJE3S7+uYRYd0LpkOxU4ET8Mp+JHgrGM9kx
jDJ1tIQz+7xd+fa3RVwy/j2Nbt5DcdUpYbbQZ26VHVhLpgODMwdJLRMPMtat7eNzjj/DlC0jD/T6
viVvz5pcpsek9TEiGKRRzZyul4PDOA/wKrl13JtJr1ZMzkZhMLkhAUSg3uYYw0W0BZ9nmZaBkfdJ
Kvtr7onfbjyy32YYSLTM0gtRl6e4Ke0pT7XAt7ydY1sSsXFFeznuO6EgztCQ2RYD/3+3j/8yydPU
hmKlUy5NEd53rfH4aBzho6RGphESXe3qMh3u1fcbDPafz1Y5/Y7G6pVSjHOoA6VmhqSdHfB5CkWV
hNTA7wCgj+5dUn9rep6K4RUToDmm+1vZj9RbANn7Lb9h9NJToTBSTO3wWbnfx9skgDvGlurWYY12
jMh5rh5IueLDH2+mhkXWSvcXgtTD9i6cTTgyBW9rwLZVHOYh9+bM4oh/eRfzSXIcvxaxCOw9iurM
K/WZ+br9KWShE8+9p2kkLmR79tiaqCXbZzpovUjf1nDfvu/xlcly0ayi5ll7jNrfZIVViDl2Opl+
HekHiqW0y1EXwrNbyQuI1Iykw09+JY0ECJwMuWlcGNkJlWcA82kRXIvEjFQ0kvgrYrQhqlUemdWi
nrfj0kAzNXUWG0DvkM89hfWmsS36gsxaHraHzhh5VSsaAJsb79dgNCIvBWs5M+14X7LOtleAWwxs
Z4ag+GT1CFRATEF7hDr9uwObgfRWRgKlFdFBKDcVRNJQEqzmuwBwDaVlz1bFSYdTto7k/k4uCiOw
3EN38823jfy0hfo6vRKE7xZWZnFoYaWs9PKH6l91jDOwIqljlDAnpEH3r/Z+184P+FRdONNad2N6
9dwuIhXHvS5VSidz7Aql9fsPBCWuBc97n7DwwflU8CB9MYDpmNpc85pzVx0rUHJqpgLPhhDGMHuk
WsjaYu0KIRYxobKAc6qYddP2LXSnXgSIZ4kXOaJjr237tJsNvJiggMQKOB3HJ48Ov2VMoOAKyJXx
PYUQOEzerIUdz5RZXTGSvGhmc/c3BDSCqsBZ2HjUYGgRLNIkF3gkvx2TQFPWgGFDb3xerej/UStx
Fa13TFgSK5fNuBTiWALEgbJGGPR7xwIsoGI628vlmOpVFjwr3yu97BfnL3iw7ccLAPzg2958e4IX
xtQrlq1r4oHscz9Joc6zpS9rJRN+MbE8i/Z92382MyQ7lDWMfeXkFBUwQXFLHaXQ/oWSB+BySKhl
6DWWhLi007CmWn7vpPXNrK9v8FH5U2ozBYa3ir2vp1LCh8x8CxCg5V8T8/l8HdJpzkdp67VzWrET
C0aawM4zTqA85mGh3V/Pxzjp0zx1EUZQkVV4681zkhcDjBLFwgBUeYIsW/Ik25KeWm66fRl3YKah
YTvo04mUFnLOmCDhOWnzaV9uWBImliBsudwCyM5BH7hRw0l+m+92iLjjSSo8TDTSvIHU7FtH8mYe
9ofh48k+XPFyzSfJj5ZFntdQZmt/gINydI+d/Pw2m43kDSIzl4zHwQWjTdMgXyq/yaFNMY98gldP
itb0DkW0+Wt0CJPYVBF+92+L4OZr14wfKsmDQI63O5hg+YUs8PnhSl7ljlylEAdglqH4ii4pbg9p
GWjb4jYseIHjWjA62hMhM23XRA79u9d9vWKXw4huyarV9YnvWWEg3cFf3GHeIWZg6KxqHNWT4bKZ
jAr18zoqotLUU3T/6WgUIWcGIeYILS82MlnHBDlk6R11CP9gNDwDlsNIWHQwA87u1Ywq8PSasrKi
c9SBOW41vBCkxREwWWTbfL0mnCijpl3Um5Yoz+46hDVe5ZQhLs2U5E739nan8h4a8inHheNK0e+1
ilEX8BGmOjHXxQt14MwnOay4FuI2owEHeZWPoIYz/uQfNfCbbAt132vpP8w0fEBkdKcCSC59hdzu
p72xe/s3kth1OiAH5HoYaCcedSEAfrZxm8G9fGNRGQdhzVP53RO2801KtoKJnFtFACrYZuWlrwxL
Wc5p2K2l9lMqjOPh9ZvSXtlpxlPU2Ey7Tm2mlNVhcCfCSvE650W760pTWQ1r+iX6U+hXXi8IplwJ
xODmAV4jv5fzonQMvCJbW20kxOwi9qIiX8ck2veippPwLvdO9vsuLhD+CWVgSXrFx/iI+QEepFiz
ojm2v27oUAxIolt6wBLR6VHxwL1ua8x+tot5jQdyytYZtS+5d+Redj+8A/Gk9Rcgnwm+k+8IbFFF
53yU8+Spe4LAMv7tV7loQSHxdDNc2udnzgHuN/0RyuE43FwGhi9FhWz8R4qG7KEdAiuZKnpxo1H3
h502ZrinFmisc+YJoWfjqnVrnRotcxMG+UJmKHSmv4KuUbCcEz5hLlg9aUeG4Frpe3zaJd7pPzHU
X/oXcbJyq5ttCLqkoSDLa4waCfQ3kSVen7HmRRDKWHgtc44VcyJAOqAvuDBghWdfR9gVJ/Y9UX8N
FMbwSLK5ZpHrraRMbT69lG/Nb6eFmR2PWESqZzVj+z37JQX10oSbDttJsBZo/MwNOPLL4P9xIE5S
6qx2pgLCvjEh7khGxFgJfUBB3DZpTTs8qwXp4AXo3LimVnaO8iixb09W5qB9sipSlg40mlaxsBK8
FJbvpTNB5OXBIAn4irCqyxjcNCc5eeHWbZsw+RFq2G7zr+gTeoLeVVTSahq9TOv1fOrEHcMyX/1u
kcU5GxmZ8UON9E7EGURUSIVp3vm5frOQuyNYMhReGwiu0RbalIuj9PXDgzyYKB6K3ZgsRR5WZZpR
uLGfxxK9/8BYW1FkXiGbwKIQ1x0Asae7MTGt6kXSnDN1RDZ1lGpkM1nNemHkEIKEdrLVAyHKAGb2
jQZVhFo2bnM+eA9+NKlt34JV1i/0ZLccdqcWdmWNOucT8178/WYB87LIt6ikV9vdEnacQkMMZPs6
z9X4X86Qv5UJIP6oDA9RMSw00gZlxZEtyxed9MrXIMrV3hOGCNsU6Yj4bXyHCNrxkuVFfgbMmHIF
iSbPeGuYUNAZqvUjL9KfTHb9RaLbJLiMZN2XDJjHeeK0a8EogsYA07o9tCSnwb7Rv7OhejAlnF1C
XhYIlN6nTqfv2H9eagKwXFvVjPGsiqDuzqljKQql9URzJLgNmjYR8YYTLi34k79vlLKLT1tBrd9b
s5qU6DFOsuU1t6dCiPb6wa4clzsvIElrlEemyvpY7MUsf9yJ+hmrlx4BLvTz+k88cI3/f+Fr9Ta4
NXtKNWPhyg8jt1F6tnOmkfWDTJgP0rOf2GHtkQlk4+5LK005CtGlwr5439z6xkY39QxkxDx3NmkY
ZR00bwinnrij32IGnjXV5C3L7kgW4rgY7lQNUslqvGMnFfCCJIWlzunJShfhPliOFiYVgRjF6G/S
h3hNvdtnore1eyyuz03bmx8lIJvKqr4UsgWCDHxygUcDkVJMUN4X//N9FN7lIOwxCs6VCYn7Cz8S
9dYolkxg730Id/RqPdO5cB7lBJAtvyRD9xQTTKVMVCKEGdkiIOzvpkHxK500SsD3BxP6tzEAg3GW
PNJ5iv/N30K2Joi/77uqBgANjzcKIHg1k/m3OhHFvlfD9w+vln16TjlaxN6d70Ng5NsjHba+nsZg
TOAsZkAX6eXBi1PIV5c9bQHl28Z20WKMs2V8X0kiBC8yt8Oik2Nw+RvDGkQoVBPIItxBsWJM4VFu
hqe8o3oECP6ijMda4vL6tD30pa6dQ8PjofSrZls+ChRz2mCp9O1DPPvwc1kPdGasURuyIzDgAN7T
GphzGNTrV32kpLwoM7ijw5pgG9D3xvuNeAlMPqcYdbFtqsTjZNi8J+Bh8fWFMTUwrj/rypBTZddD
AXVHsMoqLWknqYVKHlMgOmm4CHDk1/jDApMnoOnEI2CNL6uZqUtOPh1bT3te9PffWbZIoyqnhrIm
Il2KK5j/CJWLWg+xncUFSl2ie+d2OhzKqgXF5HflV5MLREa7LKjVxS/XMdsQRN4+ACLNd7zZjEHy
jrsTLpdalwzHUwGYeBnys5sRacYUE1NVXDpHdQpv2V+9s6VOlj+fcRPURqHEmQtbAte1fhstuDsc
fv90E3nHpcPC3N17aURQU1XQOJDZUppe6hrq+FN/wm+b3Xb4RK6qatX/PjnELYA8cVvx1h3UfUNR
k/B8TrPuy6/6WPzxE/cWNGK+Dk2CHkTcXmLntum0mmUNKTL1k21blCS4LTyscWDkEEj/OUl3HLVF
2nD43vkdOmeef+0czme8SI2AL4p6OESEaBzt5pP2Rrmmqe4GJKq8qmhMBGrC3htXL/Ht+Etw1r0/
JoInajhBhyqf/d27G7WPqsVIJm9pdN0ZvMaskLQ1hob3erYDX5XLe3M1fzqSw6wGcI7nSqVEP4By
QiqE/CZjEpDM4F142OZmEmVF5TslNB20TNFbFVE5xlbtdZsiyPUcxM1PoYXygNYHQ9ti4mMTk4QV
AIvBJaHSnShJLoYQv0hX7yuSt8gS70dzHKiDnU8Jeyoc3xM3lKJnmYASY402s6heO6YlKvmP779e
r+lHzkopDB1CQELo/5llKbFEQrUSwkJZFs9kOiZrF7zSizfEwyuQn2cmiQEDvEZ0kyJiMrZTiwU1
KOYZZWGy2NmtqA2iJEg9INAuxj1uF0z1S4wST9r5EMuDEfpQcg9S650oT4HZpMv/hkMnbSCvyC3f
pxH+XgiSu6/LYRq23jmvYr7Qikvg1SGya95hTQusLqUWzCCHtKeM8lZ1TJOqlGbw1rZnAW/vMffg
hcSMW+B9GGex1a9sa4amm+Yujo/GCcFeDzzB2zXzH9uftzBAKuyAbHJAptRJEAJ6/y/4kpLMrHbB
KBXNws/Tkhun7DVRK6wU/iYXP/rmbjNXRkhOUxMLtHOuDeEPjFPP0AsM5GcPGMCHSO/Y4CCWbz23
fnUghuM28R72aUi8LScBSWuOeavW9DPWRKk1gcPY1PvC4G9G7RHfjVTKgb9Uj//W3IU44PL3tzVf
Kgcd1sI3CKGaDUfzgkFH6bCaEj3HAkWAtyCzR4j/nXmzWoNT5p7KE/DQkV+XEYuh/eLNm0ZLCJSn
RuSWhxiW3qYKDDjAIi6d9asB3cYwSqWz/p54iyyPZGlGqJEEhaO1U79vqmrmp9aJLQx1C+nx5Gs9
uQQaFulX1kUw1PMrbnZjOVjh0ijPeiah+vfGCcVKEkeofcQu+EvNQWU2+95tBLXItOuLkeUeL0hN
nNROiRbgPpmYH90S9tyx+yGkTJ7jMQFEB+7RDzTk+ZRr8FxwERWauePgUIGNh+kXBWAqJZx2mVir
MIKaEj/mr+zSLRuqSw4cnQBqDyVuwsBqBknhvZQbj69iGOI5o48kaBrty4gwJfk7+MSKFq904LH7
DBZgpeZRg9tSC1f7LgT1nOkoURjVJV8zxcfJGlrFlfz9ur+e36nsqqcprP44Hd19U760toElb6EO
7VoBzk24tFJ1Iatfthz1DALUIurwV5fIO1pB0LnUOdRV/A2nJNJ/M0MiI1u/PjkcXAj5oIxpdjMg
JkQ0Cci60rF/HqGOGEgNpgSEnzvp58WtRQnqetZckEU/QO4hrUh6zLopUT4x3Ny3j7LsKOR2+38H
ZUpe5JOH4mmTEzZRFdq2AmaDZQp61y7GQ6aGJjdENnrfeEuNVuAtGxls+VPa0GscUfCz9gTNlBRx
y12hVqmOBKspYqwlhAy8zVVbIiYnGlTiBzHB465hg7FS/vA88WBlcBxr/F22cNE3Epsdvpbr5FDa
Cix0SmUTneMkdjwE4wVGE/D/W0DLJ+xP6Qe0knxSUPf641xG+mUFbWQKO3KBoIJ7R2xQBVm/li7k
lWOj0oN8vCqugpHADJR/p5dFzfBeJA5yv4XUumITUGMZsVV88Hb6IOVPlB1i4rQsXIE7GBQ0QO64
uYjeul+lP8Ping2fswM5RsYQe4d8Di8qpsOq/T0yMZ0XpmaGxFmCJk2+lIVug3fwSXlKQr+cnGvz
Wbm7f8fL067Y+WjoL9y0cG1xqWBTNp4Z3jI9ooNpbWFqcBRVOEqUjbki1Cabc+Hcxn21NmvgDsE+
0qCNTvyu8iD+dOSOckofvAk9mTcNyLpfDOi/vNh8P1NcDdjsyZqenghGZyTlS4BLzVY3JehWdy6g
nR+k5GJlhEMr2r8Xo8qBmS1UmAKLqmAoPYoBL5tmmB1Pb1yhaOYORMRGTE4k52e/kDIHzmvrsEI+
q4fbZ9yOYNLrjnO4brVqVpscOPFUbjACIy13etA4U9Xe3nM33YVF2utKbGSseZE4M2ZFenXSKJod
cbBvJi60PCSaeSIX2lt/itq9ks4U163m0jNL1Fh+uJSNv+S3QUF6DBvb9QCBJoMJQdHsoqsjDTxP
UlRQZ0BQo+5ws7svuV8jvqpxpvclnfb+BMARv+FRfGnHwo/OPLpBVQjp34EhTjZZUNRZjaQUo5WO
sebUml/Caj+5yDPd97VYPz4xnGQAo4SD9pUCWgiKYzB/pEOD7ofbcdmFFZfcdVspeuUVA0x10QXg
3Akia/e7OgMLSC9OqGq4TTyVNiy9uyyoR3vc6X9sImRAZy+mrMYnbQHXhU5I5IP+duaJVMm6m6K4
L+bJiBQs/5ZwGSiE6BwA4tICx80yApxR4Ztjvav2tSU6VmMpl2YayvHaOxtKBJPafE/Aabm8N1i9
e5mindgoIvIJannmPGTKT7onWZ/3sdo4FQVPrmNyey92SoDjymtxhB9pIv3MJqVLE1ooBT2Hzi8P
u4e4Y6H1q3hJP6ImxI+t1PN42IWbaUtCYDxJSl7pom5288J32TUqEd/0IrZVYdWuyXRcRr/Um7mx
Y7Wv1BAj57cv4k3Vj5955n2eQMvQ4jsD4ysOgpHCNcD/3hi1064QjroGqrfCa3NKf96W6oAm3V4j
OFRMKsx3wuihboVmHp7cp5d2AIusMdwLGm3Zd9QA85j6MG6NFbLy7bdjm1suV6LXbrJfaGib4enC
QrYI/yTAwTOG5ZOtpjb7ako7sTXWnnNVYdmTOPNd62LKTS+kr4Fhb8chf72sDuFzpKzQQ+uzOVNW
QMlJrSE+z0bqpT84BfHnfcYEDiT3KIdLkjdn/N1ErKi/JHjTes616KbL/pLWGQLJtd6AB+xWY3mE
4Ja04SNDHcWp1YUmom66w13D0JwpbA3s/kmOM6+fqx2fgsq5UlFX0Nc0dHntXdY0xWDfb7z8Ha7+
hiOEM/w7hyVLvqO5tmy2K9Gu/1Jn+Yk6clZ9v8Rep2cHZieVG0+PGcVM5ezS+wrYMsa30djaVbrD
IaRIvCXyv6U2Fg74XXjcLMvJZslBe6qN1X+NlWeBlEP1tNtLGTDtV65iNjTsjmD9r4xxPutgeDRc
jvl9voqd6g+Lmnti8rbryCQ0lI6OXOXg4HQaVyKhr+HIQw0YmSTyof4mUe2Zk7DAiSQgm1EjYTFx
5VAI30pZX86jD2+YbA/4I43wlOSDmmg71O/EQqIun2lovIi8pUvtUFcpZe43pz4vN8bstPFN3cl3
YEN76AosA5CicBkwxRpIZOxx+3YqCb9nOm1/SjpAtE5+SPZuCgbXyFFfSEzU+w7191QVTe0Gw3wl
ggTzCSdiLiSpAhc2GfssCsRZ/DbuRYj51r2E5UpC+qrFh9iGyLamg74Oe5bIgSU0ZNqa1tRIQqVy
R6MtOQYf2Q/3bVrmmt+3WY3zdkSnfp/ChU3XqT15lmr2LYMV5OrGAsecKLDZnv3LQ2Hk1gBsWgSV
9lDCNhl3vrkxhvAcxdo18c3yEUsD/zaOIEUuxXEmUV9ZsS05JK/HawHrRqAX9t+Y1SeZqxi0pQJ0
xG/tNMxXY5MzddcgUIKIDniOfwupbwXGfo18W16uusd17KFcjNnNGO0fTUCrkENxylXvi4NsvefO
4+PH9WuqKVU9UFhTCrge3rjEahz+ftJ1tUWquennV6Uri5AtUnFKvbQJ/4vB+ba+kAi3xxsCMP+y
ccU9YaQd0Ck9Kiw30pmzaQBGC/RSuwuiCYRwcXQNJ/mzqGzLScSvWdG6sBxtncWMrSKF4poSft+Q
x4tNd8jyEPtPnTu5gofN8WGAH0PUK5bRksBocbuOZluBV16cJ2wnHWO7e4o5B1O77f3h5KlzTo4p
ETWZL7TkfCbr8m0a04SZkdJ4uVKf+9k1/bthSuAd9IXs/v0x4iVE7H5ablDSh5m8xkOf9T/a2YaO
zbCbSXsobOTF/+ejl6f4uLRG3FIzKxOnVHFmO/PVnHCMtidlyz6hPGjk4xMPrg6VIGYp9sLLlDA+
s2PJXoeUIPjXQ/efk1vjDKYn5sgLmsUQPX/zqXdp8X7m86/5dNFTym6JfztBKqOTNn0XI5hyX1Vk
ZPeciRic8Yy1I3IbmS85h+k6CVqsdHcqJhZ2anWe4TmC+N0MNe1HdJyAQWLhc98NiDp3jMiSxM76
ZRthmFlPsYGpd0/1DsshpLVgZv+zleBaYs7O8CNWyFASLprhh7Hc8F2aEUCIAvd6598rk5tJFQdY
Ei4mqIvq/IpfG1v8NLepYcAlIJrGhFFsF3TfsvIwo57wSfEjDkuWJpgnmUk/0oUCIplY14/PLMJm
H5H1ZDTlzEmyjL5Jug58tre0O7A98RdYqFAzGpiZRhtDpz1TfRFUqkxuOni5bxMgA2GWrW2NKqns
gUr1P8FlcwgFV7dFAxA6+lbcu+YQF04hRO/jBnwS+GS2846MdzocZjIwBiqGHgaoOrZGpTArufzT
WN5WfM1oFFH6gdF+b4m3QLI9X5bIA1sa0c6HhVQHIEvhOIA4V2yhyFdA0v/iIJg0v8RDo+vxIknd
YtML4YWTud05PWz1LQnbDzT6EpP0re9uNJ7tcpKTK1P35arvHKw4YDidFnZMrQS+1gblsHiyEK6M
FHyJDfRl4cgdBgN7d5h05Ryw9I6O3GxaMcKaNKmPRxExJ30lqDa2zrcZKp+i0sjiWH0/qcP6H09y
sHM3PAWmp/Fu5dfKPiPa9/Y7r7uHP3UvnCZ0LIYkLSrxLQzoNgVOkKW2nPOwyew7mX5UdnhFw/5t
cRUgGzEV/lZL7x+pNyUCoxl2IajtFtQQtd60IYU83yb80/za4qxxCwx0zKvbOZvKXWWTujt/H3QV
xZF5zI99/xWQrK3mNkeSVfv+t5w8AjZTxdwnCXcF3cMYo26zQ6Pns4yOiA7+Qk02vmViConJlCJT
YpweoVu6ftYplaAhcZIT2bAUrvgT9Ywq0fzg8bdni2Fs7A9Vt4+xPGIfzHHEnIOaizOOUjO6EKlP
M6LcuD5GPPrbEqtf+oOeBhBF4aohyecw8xOBjIU4CIp0y3QDRthahzksTLe1lUbxE6Rxm+ghY4He
BOH5dCLtCwPSHF0BoWHSk2EBPPHbeGm+KIoGMWQ3d1rVK65JydnKvheq5M//y0gfK3VeueLO9ewK
Ktk9H9CRLfUs+8BbSOdEArzrbb+x8Taz69Zy9py6XEYF0tKOba6g/x0xvmeysppk6DqCx0Eat4Dd
V/7iuWvXeGpU7Ek5GyapbtlpE7SwChJrdgnTPoF9W9vaDuWd9zzl3uxTGgX4k9SX+eJHhzaHq77I
Boaf/7y5kkhVfxcRzsEkdrLcsljYaCrxRWBz6m9LxJt/t31k6xerAuQ1YwBm3+cLbEZzAEcl2QVI
WQNKsOgZK/mNK8Ml21q4x4BBQswy7xIs/L22UGKRafLoKRG72md05uv5CPMledrPmBeGA4PTo1Sn
gQ1i5duD1cX/dDA8bEp3PkRENMrIwM7HAmJ+8PMH9/7KO37K2EZsoLOHmXK5z65XOYzO8jh3SuLE
fU2qeJ/lmmefWt5fxAnRF7xTpqd7L10peaACJHlZ3NpgvteruZtYHtubo3+tkh5aB86aZvHpiGea
JWu1J9ZGRSkxSdu9m/XEiQ7WBv4AsnqyX5prpMaeV+JRGFvx830I/v7l1QmDVtnBiBh6KJ59k1vy
VF052gN6VY2JjQmKmZG4hV7NpXaQCqX8CxvACjEilNetPPzaCqu7vVh4wDiKu92kuR8Hr0dGzPyC
7x5mtv5DyfDQwYTVxB/i9WtdU1+4STTVrFcbgsxcQKab6lLHHd3pJ4XS4jIf7z21Qt3dljsS4WPE
Xc7GcaqLwXcByTFiMBpov1MRSv1TwwwyoPbSiaYsEGHIkmPVHtAUXZtLdC7X+um0fXC2Cu5mJVar
eBBSiQzx4XfO4+9ij32FVEBFaX4DW1d/6SiStd3M5MmpWtrjbEHchLW/lJN3JV9bCYwwkXPEacM2
zBCLeuTfKJZbJwwbhhk10qPob9GYuT43lXly7AUKXU5VgS7+ptZ4jQYBF3qzPoSnD7kDIX4pa5JD
XfCic6fW7PqFCw09IMGLU5TEqGjrn6/rEDFpjSJJAjGQtz6OLwWU3LnuNgu0SGgfqXa+hL5Kfb3e
RwRB+KR9hlkfACcpEzGaPsv0NUGP8vwiRq4B3PIEYE8jxDsKW7JnCWDKP3gFpvU3UU5UouUC546G
ngBWUyEunUWm/2Ap03TRASHazy2vIgYTI+kSiWTtUYRdXPrhX4uXMMa2mw0VrrOKNU6v4qaYN2d+
aPTx0xu4uAFh0VT7+tG45KrbLeN1yRoFFIt0Frpw9L32U0Zt7Zd7bGoBDf3Pcvya7gX7CF/bhbLv
M+hI0W0ac1glgC+iO9JzeQAn3oW+palEgOZCRhGhYlWgTIDeNszElswbJcrwuCca6tnNd0TyHMEr
NzJktClzKdj8zCy1obIYMjLWO+LVg0etn78NhVB2AzFfMeJh+byn5ClD2YvW5sb4FxZ5rUypbDiA
SNVe8FAdzLjtTBcrvgLwEta/RQ20gdIF0CPvzEYsW73VQbi1AszXfvbt6dIgdAkaBTT1z17ZML6U
X9IQiEqP7bIAeTlaJI7zOcWP953ISVvvZqu9tliBoXGfGgOHRSw3Ms5Tc0MfrOaufXhwx40HYj/+
440HwJcSIqspzauLWY+j5igqWFuf7yTbSZIVuuw3hxqJgLg8qqW6ijuZWVZShbxUHMAPaS0Ig3cN
67JJ1XomykMEAqDrURdV2ZtaZdtNgIOXeTW4Di2IHmCah0mbqvbm/miI7VrdZPBK4z6S2zzklhXE
9ers+Z5J2BOPBcW0fWVHf+gUnrtM0tgNjx0lnlG+HXXdRzgRMmYHnGFRpntqC812vkYzXv1k4zQz
J7BD6WLpB9GvBf7lixpwIZ2YpJ/r0apWIDEP9zUR3alN6wd458uOnmRD7QkotGYTKkCJ/YblSkOm
A7aqxjTKRHGCVCraQYMMDywWX7xE9RRYI5kmU6BxNwkyi2L15UbkyzYXrLSPtGm6VriMqiJ02htM
Dy6HS0KeqSrsA8CZntnmOtPkliJTgCSIharlLeP9GId5AkBpjYwk1pNuIddJ9+tpm8UJfRIgEoHT
5fSG6NfbEnhHdYKTWCgFynuK0ELT49yOIjgju6FzTUibcztBHFtjI2l0Y3a6jtnEB9NTCEDVzkmW
21l/6cJ3uBrPtDougtTe2/urPoo9/jYmTAkDWGVgrckWu3GY/FafesLfUULkVMDzsrVeoV2tZH/W
odZqeaV0y53awLZhXeY7h+Jmm5jCob9Tz1Jl9WGbmLb1W59pUWAdngx1WgMBSZAHzqgpUms/B6xB
QifJMQkz+IMclL8s7+WhL6bBfmv/GXLcHeVGQW4Ea/ewbzsvq43yfNp7o/lO/6GCoDeNjVLVXqWf
9jhKJ1ufHgXtHOttgTniXIr459T6se9mNeu+g08vnC7Dwhg2Rv0QOZpfxq8G+YTBeYC3PDXq5Iod
BxVH1Pc+38sQ35fayV3yUvpN35wLgBHQJbwPf+rcep0UHJLNXVTXLPFRVHZMXOSp3mVMVa+T57hd
MfSk1rGBtKrZpZT2cFF9w+b5ZKnTdELXBt6NYAIfliOa3uEP80VYr74YqBZjvzxooAiW5CQ9kASu
7shyZv1wyFJjWrIR+HzJyODnkEE0AeKWI6gafGUxVzE0596KFOYPUGWCcuWtvY6ZWVcMp1DnHY7M
pXXmmoRzfeH9pj7XOCgZYZUPWHk9Sfv3OzDQA3zVuqP6hGsGRzZKxV+0OIQlVulJkklEIAUxkUP0
uok91VNvBaTouC15/GTPxIQ7EuMnSFkyGkTwxo6pPIGF+fEQNLyMABsrLftNFCrAG52XabAh1LDu
NHyXIWqwJaxIZgjswJ0CledkXlzYLc8Tac5xsBCbetYgOPr4rDD7yaXYLk9hbA08nq26sHb6Wt52
rMCj9a+RgI0mJ7vf27OKv68zF3RrxYHFueF/NpAgcB/V87polGBsu8TSD1pZSYpLOzg/a4gx5SrD
D6tf2b8L5vHt8PugQBUew5fA7W1IjJRQbZHiZMy6obDdiLSMMcEVGQxweDHf/9yUmGBeWFK7qjg/
i7pP0MJbJG8yc3EqZd1KxDV8NiYBm2t7Xb4mBk5XeJmdprWmlx7DNRWe82W4dfrCXL9DryWhqS65
Mq2ha3QHJ5jEcrces8/AIoFkssm9dFswTJ9LWU38bVZ6evHoSi7TpcWKKnW/afJadw8ncMUhgpIj
m7mWIsUar5anf6gD4lT53VPHJLbUoDhtiet2qt7hCCvwUZCwKAfUqrKHetNT6EddMp54IIRaRGis
noEfPH2wO3AdalOoF+gOaJSnKTvYDDpN5pdAcr1CpWqOvfWHOYc8/H7PD+bAh+6dpuYLE7/dXpsm
zCldTitkifI6uZ3tCd9XVZZ4xcaDZUgW3o8cQjJ/XEBxtvRpCLuc6phYSkoc4bFfU/vCVE0K5ZO3
CYbg8bMiGc4b1vS/cualUEiQkuV7GShtosvv+wbZhPXsxlS/K+wTKglMaLk8x9qXSeG+zG5xcs7R
L3WpZ+9kE8jSY+oEc61EqfKEfFq/O0DS47jiZAzaaudP4EXa4M50sDtExCIqY9F/++wcdPzpYh9l
MZQfFl1su7GyUoxhX6vXOB0dUkP4ePFE/VLymSru8BQsmhOKI++nnUzyBWWKugLL+hUXtLOFiTt4
vOWF+Lofstv6muH5PkHQ0Box8B0XughX5vCcC2K+DPhV92pmIs2Ef15Z0BXHbWtPbpX637giO14g
ixIxRlTrToOCLglGW4Zkd/Q+3w7xXHY2pUuu8iwxpW3cN6VB/PM0KmS1Lff/Z5ITyAh1Wu22jyJB
0zJivipe4agLJCGForYKhHHTtSswHNFJGLzDfk7p5wNGV8FBctVeolgXEMkASGWPiRDepX60DjhP
+qYz5vv8yRfzj7LQbGMjSXmon7ZFHT9mnDpk6z4JeH9cEMmDU0mu/sODH1rz+pTiuzMevC/vQn6q
nIBEN2p9zCFE70MYb3tNhqPrIkQuBk0JqYLROdAisrvr8bngFsOWISDjydkM8Eq8HiDlha/eezho
I3DdTlsGyUW52NRHBef5Cw/PH0SvzDsS/f+q9fOHPecWBfkwOMhfTh2mKHCtoWbIbo14MBo85POj
Wy0Blf7gxMhizE9s53PBe7wLMaSPeTzV7jvm276KHLBm3dSaZUjF0tfYw1PiKdpuraj2TbDMkIl2
k9eSJXWI3+YaJQXc2Co5xMProKe5ICR2ShZiMgn8hq1A5iUzm4hjnmckDNw1DxXbm+aqvn4YQAHj
p3TFUJGqTmwwzT3hRex3o+9DmqxQYVLurfVzCYIQ1fJ2YM3Xwa/lATYyA8b6FluKAlYk8OXurIYg
lXGhgBiRySoBjSFpdu4VA1LzpXfpaBF1Grz6YWlb3J8KR5rK7ouBPI/meYfNTnV68WoZ2mVincrI
oKccvpQ882BgPiuFU5yB22XBbaD7ShtSFXdL+mk/ZWyACf4F1sijNSOYvMYp6VB1sj/UAXdkCimp
c5c2qKRgyggG+zO0tywbt5ehZAoRqKMmohT28Hjz8JHOAdl8AOEtjZGKVvfGe3+/6g4F9KEQ1rrA
bgVvMEC2N6lrQ0wWptFH1mbDijde58uIgrg19W3ihsXlFHaMjpTCQzkxlIHkDeEOVuaegF0Sa6vL
hO0yCL/mKnRgmVwtigQ6dhuY1jkigRxCARCl23ouq6hHETVaUwikWAK2YrcTEbpeN6xUaHgWQqvo
jQdVmR/0sdmi9Sy1isqFlwkHm4HbhcibDk79CfSknQHOmfUmB1VANuEaCkTsBubn42vo2VYOOv1h
8POALxGDMzGklR+aKYRPic6B4oPPH0f/VqU6uWgCOVr5eDMxS2+NnsQd06OTCCOiEGTDVndfTwqy
0bWIZQRnrL2bKrCn0p4zAZ59cvFQZsafR+QmYI95P/8qSzzeHbZYcm/T0mRRl6GDOvA4mBzgLx3G
FpdSV32Zw4iAqhYE+Mov0M47H6XePIv3L+GJRRlKQ47Ylag0kx0Vk/Wvx0zgOMHh2o27SJ8MtBgm
fiBFBCyspf9NMOOoOz3EWd1mMyJkC03dqQDaicA+MMIj0Sk44i8TmJQ4k7OaHoOH/iLF3idi8EsO
NfZ8u0sz02MxzwWAI0ZTWex7qHc44XRUBcHFx9LESMLt0n4cBtxL4n0CVi8ED5/NWpvaSdA9guIh
M2avKVLDyzFjh3+GWL2Jf5qdN/6a07L/gwbKUizVBTPJwHaRj7M1LTImDuvCXd3ZCijkzyvmrs4B
yFGfKBaL6DnxTYqpWNCVLdpRXzdIizQZT4YUU/qWJm/ht5gE4ZAWAviHqUJasKII4ZOFYplb3WMb
EB7r0Aq04km5XvK7IT9Dmyz5XAFeIkwCwpsUwfhDC8RT3iToMw+efkRlk7ejezn4T6zxaSKQyPC0
ccr5Aj20kfrm6pn6oEZWQ/XJuPAoNC6RD1qYIGSTq5wONAnQoeQdRieCgCLhfseBpUUGwHQaZ37f
T3sI1Vdm93tF6o5Z5JGHUI0aS0RmtlXUXgqrGm4KeWBCY+Ek+fsvSH2BfBPiQqBHkoTmNFYsonS8
5kAFA7xWYPCiKrKHChqnjPDhwGpDjvRRVTLsQ299sbIFdivnd7FZXA2FUmZwpbobJ0VeVYG231Hf
fj/YT9LVWjNvP1/WHcLrVVeTPbasW3XugTi8F+OY8+TrOhab0k3Y214xhFvc+PtZ+MXjJyFV+Y6m
n/i7rqOPmsQc6yWSlwTzfxPeomluJl1mQ6cMnVyBR0dqo0Lz+6u/YPhiLV3PmYLtqzCijennoNxZ
ydglgWh732xhcD81pelP1nz07jmyoQWtmv1LP8LoR+9BGGtEGCMM+lQEdTu6h7CsY7UzNskKp8N5
l8WQxZerCexSLrPFReTUUShhlDnwDZrLXnDRcd32SEK2o392XvO7cOo+YOw9yRN5aeqIicC2yYgK
LMReugmFwGyMxfVRcIFzJY2bDG/Wz2qrT6IO4o+3vsoDkzLVGSsdJxMYWxcnP7sw7fnVD0DHMDKW
6e/It90bYQincxWCdFqhHPNxahw9oaE0wO2CBnrnXKnBXkmeQVTbmC3IkGO0kxNeJajDT7VZxOOn
5F/ll35wfYgUe9ISdHolJSEW2UoFtpDYJ3+zTIt6VxM4BOrtss+LRe8SXyb9EPWr5RXqZ7I6wgxj
Bz/RufYAqlS/7OUdMwTTpVXzip3HX4e3WrJZ62pKhKl8OaDUm9DpACuuC2gE+yBb57Axun/ZGxKF
tCWndtmGoIvnniJmCO8+Hf7zvLk41jCv1sNpDH9Sp3Y//6es/qhAAFPCeXSkRCFqeOCfX2jxqhRt
hm1oq2enAOH+VRP8iFMDp52l681L9vQ9L19wFxr/ThFZczhiNiz2OpRH2UcARHVXYzkSQcDv2aEs
8Q6VJqXjej9ZDz8hWj/a8w8w/RncaJYD57ScWkHgRRTQRneWhC3qE+kwgKJGskZmcSdclonW1yhJ
YjccZGTzM2bzPNh0YlMXIPF0KLNznnOa6U2i2lqhphQ716s7E9miwuQ5Q4p/6sxNYHQ0c7xxC1ca
xtZJ1t1Z4SndUppq1PZFfikRJpuvBaxmH2mCCvttgLZdzd05aS/R740t9+dnTcCs1F/CflHEa/s7
P6gK+h1vsjkDxDI7y3JMknPV1ZBPjnYux6D8se+xrn5M5JwX4mrax1Z8Wr1bGBnmoIxh5tVL7/yE
tU3NVl1jvdHRdoPA5YLVBFqId5hGtMhRTwVIpCulCZ6lonDUu5If5nnuVg4lWyW3OKCcFvFylAyY
cbBxDFom6389drMt0aqSc3ovaNZtlIRINYno3RC4nzjUg2NUDVoOwO/u1eXED5f5zWlW67QEVKpM
YucEKodnu2I76yn/BuK+OjGuLGkdaN27cCw6dAlUQjU1e0zdOYY3hoDTuC5bpMuA86Y14HcdKEdQ
tW1aRvcdG6gnaCh5JhTEjYuNWzvxpVlR/MXqIH/fF33O55lDHIIkw+/IUKDFC1WSIxMMsDHqyHpD
sRScGDmGRlBRrBFsrDPaPIh+3Xhso3s41Ac8mL9QM1zTkGz3h1ENSD5L6rM2Tf27Yjp7bb0LHkhy
527aJAQ+CUlKaC3TZlHGD47GuFihKNzfXukr2RHcGdRmwOYzHikap3IgW4VZLhve6luRLlz/dBfD
3zzyvFmWZSs6b0iaxadovzIRMTtsrZroP7cngXHTKLrdl5XhSQSWs/+6w+ICLF3Pcep6g5/zqbvH
G7oXkaPpsSeyVdE/FUYPCN09xiJuJrmrJT2yUhDlddwE2rP/tTo3wNi3GKr7TvhUG2mpsTb8JIF6
5DCrs497SRiZQKzZq1MNlCWWz44ZMEfZOSsSR1OJrJnpmFGTSRF5/oYlMSZIpxm5N02RIPV+ulps
mwb8IJ3wpC4QDumGk4jQvcNgH9v8os0vPpiuaEoE4mmb/hOxNW6cKVVy8xptpikNBz7vy7pRSGaM
nV8w/PBiEId0xT1y8iK1vdfCMZQ9/zV4bMix8FxfRnqilGtZcNFoyDiw7hLFJiKxxh4H1x8KYPhW
lVG4po4e9fiuoe5dWyjy55ozsk7SG13/y+Q5ut4nTP1xsYqtp6EmlzSJ9LMC6u60lXhLkOB6/8TI
du/5hcpWPa392OgNYDXuiu58AudTpzvpqaNOt0jsjNK5QfRoLxpHxdBMiWOFFMkR2TAhG0UiEt2K
uE97y01OhUsQ+mmUOV4pxyYGJnbfvweMJ7rRgz2hma+IcjRr4oL8vXyvgYcyqF3ucISNGWPGDWR+
6ndNOf/s48F8L/iJMuVc/ByEeAxawpzOavkGGDLL8TAKmtfAgpwdauhJYWHdlb9ZkhqG5cUNAFTt
4ONCmV/gYxsUqMFUSqS0AQjFwNzfgCXGuSSYsZoEh6MRGh7ws0dxQYm70kASLiAHkbaMBYgRqO/z
3vZuJ2Ye6Ho9PohgfUPEwgnzlLVzjN5yR79zXZelurNRREUs70RmN2CPPUx1Yohr9Vu8e1zi6jPC
j3Xx4mnz55a1CIS5MX7UPOo1AHzFjkobOg1+tysByjsApa0In0f3REvzWWEs/rhUiC5hVr5tbzTj
hjoo8eTAxEy4AbCugYobWDW8mo3B1fy/YXAytLqWI3L10bb+j9XtzG1GL+1c27oUKY/vfGTO3r5Y
ht4MnIaXfcKMNTy9vxaW7LjwwDHg9diwFeeHrkoR4glODet3o8kJQGGCw8g2pi8uY4pbYg1UBRig
P98f1KpQ1oBhIcKJ+pBKCev+k+ojJx3FvSa8+BcVXm1qVmEnVQb8Lt0Wrr2yyNXLEjSq06x2tSDF
QEL1Jak7k7XCx/jV4KfkgPTzFQvfIUQzN5Lp6rJU9CcZT8lIdojNN/1FFqcF19Ik+cCHzNNzPY84
Tv2/+hYj5nsfscDjkfhv77Al/rbvVhcaeu8cn2HD6hoj8goEVsslHy0eznnfeVfhFTl2S9nGLAn9
AhVSifnaIRiq/voCgKOdbOBQgdTkGgMw3clXE7qsW6T2qmuXfwke6rpaZ9AIDMnW6yHbV0B6R5Pw
kEGeKgGdUCcHAk16YHcg6TMpZqVefQme2ZP1OjFPOfirln5vgp2GYQEGC2H49mjPPf+zGvmVHmQh
OGUpUyfV5B5XRsc0OaGIlRq+jRnOTL0xxy+z08dYcwet1SJmkPgmmfnlU76DYunZAEN+yaDgA3Hr
0W602CkLKmx4q4LQJt00oGymyfR0T4yp20SEWcCZveBTy9Vo14ebQDnyQLdMj40yA+pRR+NTms4R
79EiIOHLb4u9GfZKr19h7OrCwvAc8mH6Dbq5yWQPQHakc4hAH/lgeurQLcysy/mfsmCCKzV9qiXG
Y3LcNrNlLjRZmRgM6lX8YOoG59U3u+8G2SMZ2U6D33Cuxfqka/zRNdsT19QZuIltIKkpqeKdrvZB
qMpl6X+G3oFpfqszrQfuhvq/r/sbs8TOM5cu87m5i3OPbK0kxmZ/WA89ZK8MIp0Su2jvtv3dik9w
T1059nguNV7naFZzzXCOOdNSxFWnN+OqZs6drr/Z0Mn8Rhfgj0tnItyv5OjQUCcpeY9Iny4CRz9a
MJYeJaFMdjeweIxhW66F8qImUoDOLUHZxWZUeg2lWWnCoPrG1eBJMDgxd9TnLktdalHfSxj1WFbZ
rqzGOOm09ih1q7VIiWr4IbZKUsp5TCO/e1lf9QuJ2304aR37Zg6jQ3HbtWo8C7VKHxn8WZGQ+7mU
7/2AealATBFQmmVTGIqv5BFUWzamDNsiZm/Rvvz1PwKfK7vL+s6J9tuunHL0gG66E46I1I2pIdGw
w1g53u84uJNiOXQra2YYrg+s93K+ZJykB3G+Jkfgsujx2J7zI43rCTwY2d4F+zK+NxngK76qfZ96
kp4aSPG7smqf8FeDhyWtGa959iTQmbuvpVEsSxrUOll/hhDBCcOFu+90Uh5JUSRoHN4vOle1jyo6
NpaWIcZrDKfDHb8GNZc3+altgeO8WmWnxBsn0jy+Ezza0vkjQ8yQHSwZ1b75NItJEVyhrBCsqUVy
CQNT8jB2rySAGo9p9XZB0JvCRNQQ2ZhGuRfoxHBqnDPyitOmN00n5f5zPaufpFVj80B1e9PPWqbH
Z5jgFDPp7cHbxo4FG/S/9p5Xk8+HV95w9nVMiyhoBKvLmcLQCVRD7fKyck7Kk//hFAeWms/7KDML
9fmxZBHZsbh7lbm0kq1u6NHaL6KJ1Z6riAGr8+5eRLg9X2YfMRxAlDKPQASOUGGApk7ghlo3G4pQ
uDGatdZKWAg43EcKZZoU1Adb08SWQIDfKfFQlRqHxAojBVxLIsxaSpdCbI11hn8gsDLWtxqKrnf8
4xl3UibE8XSYmoj52tRx3YeroMbS1NU3o/Uj13jXyA4Ct+lmBWbqCZB6W7Y4o3rvo609gyYnHvNl
xOFrO1nkWEb4K5GJLNhCNFhYCH5fcIcqxod/pEMs9lzfa/OLp0TpYhqK9hOnFHr+ecX4T7oGqkhP
8UQLo+eGHn1E2JcPGFC9ieVmKchWZEbT8YE2GdkbAiB3OTDN0KFRG6Tzh8oi1vsQJH4ixW17+CGl
UgrcjLRof4wGR/A9XiORByA/MzvjknC8iLT+wIVMAx9XcWFYmbsrjHCP6ct2fWbVQvaGImpnNXln
QCjjIT69rL+if+CXgnvRnSDyUnLxj1U8S+6zLtq2O+Dm3qrLIWQbtUWGzApKxz7MhkwIr8EoCUrB
em6VtLVH3q/jz+//0NY7YHVs2B1jvEgA9nxwjd7LrFW6bN8TIscRI9n9/zHcJdM01DrCCJ5cD2wB
Gtx3QFpoyKzX0qMgylqmCBZFkFAAF3OQkGoB7Ti+KW/rDNSDwMVizyhV33ribit/pgLieykxUBtI
c4/3dAMwh4mzQ7qd5nL6ZbTlkzHIJ9lfrf/NOmqkBnhvGITRl8hlUbu4z9MpZIRrVWrKCzheg6I9
SPXL2lJ2dyvOTZX/o1Eo/aammfR6mbGXQ3AnrxPCpeDicu2n134fKkl9G6Yt2U3PNZdi1NngUnX9
9vR4DCHXzpVIUAFmj8DJ6wenH5lT4J1eLFrK3vnESNc1v8jOU6cygdGJ77xILv3fgsqDWiEpf9Pj
q37Wq5DSsiPOmS32tBo4Bc97xW7RQ/q/qAaD76hK1CrcnJ26day+Xb86zDt7/Gt4si0Zy0ZVwlhT
4taJgbwENC2cF7GGVAentGZdZ0mbExmeK32+Y05Ljtgqheuf4/qTbOYzCW6NaPtdV2EEf3uJOvID
8+daaBgCyhsR3w+cDVfds3AMRhrCAXy8QvB8IrNfcFG0aqwHYSRdD8ihkQ3do/KxiHMj967s1W0W
tdQqilsi1tssv4nuxliirwbIG0Gk6Z2DnPqZFSJViSLbnEygNHuiml0A16howxtFWXSRtQG64tyS
A8yX2S/ZBsy9bBDn1XsfT9iHvNb7BwRnHpNPKYdIdgPnbEWVEVq31WtxAsph0rMQgbzgNAffysBw
lWGOCqr9csRi96TkT7TA431mq9cKxoQF0V2PQnB9s+TYCJY2baTsxAU+6mIUwuavv7kMCWGdgaSO
mpqIW/DngyckzZbdsFtTW16gv/FfP460ZJD9y80X2g23YYq0ofCHei84hYWUvyFwD6adIYXSFSgr
tb0ffGgp+Ww0nsgXl1kAJJyBGa8ZFc8S0JJK1jBOc67OqK60uJA2BVVt3dTO4pJP5OLCXc/GSR7B
X71Gs0Ttckii95c7HGyYRw1vrX9gGWTigXtP3VLhM39T2zHojVhoSR1Cn6Z6t6zLKdWDN2B4yGF2
aWbOEfHtV051sztdzTTXqYxfb4jbFVuzWWsfvIG5aRfzvaEcP1X5rPjBg9aopjnn0bbaPPgemNZ3
WZukCewm1qolkgSqXViXjih1t7kQofRtw6J7Z+cP1v9PYT67AVanKGbVLenDwK45Wnesny0VbWtP
PJdZmHWRg77O3cEEi/vV8K4hUXlz4k634cZvn5hUHAw8tGH3BmTLsgErPGWgbVSOx2sl/qt67W9v
O6FNdROQ5d94qY0wYl38ugQtkNurBHeeHlN8GN4qq38v2JKE4md6LitTmu7foqS7j4ZpKLKFfwKN
znVACAD8ldwadi94JvJGa7JXGzKa37XSIfYek4GmUDOgY3NokyMypcUYqxUH5aVUvQFEtvi97MO2
2qW09vf9fumjhA5RxW6HJCXH0T9Sp5GbMS0yp+s10W5yN+VUtg0EMEcudHD9o4aq4d+vMDeKIusS
mZ6iek7XSh0PAlc1A51CHGgu3xjKqVKwTdh6/dnw0YW4/+FI2EzoDc1b7T2TtYp80tdJWJ1KHPIQ
rgYDPqzKJ8iyVyee0z672qOpb5GLmgHqPVNT9Zv0ZHN5sJodbDIVcA4sWiE0TOQEyS/TsE53YVVn
lMLbpkmYoZw1l3RVghWswlEFIl1ZxaBkvlT0pMYv10ActUt9/VAvbAc0wYIC9wwbSPzZqYKdDD6T
43nha4bB8HGH1A4sQdSc6/SL9iIZMOkS9jlmytR654tkn0Kwx/UlUKt+SLZs36JnwbQwBD7Xi/Ka
sV5fi3nTsiJAhUQIg/X4qCavlYs1o8gvofDd9whFLxetPax39hQKhVcDnBIgN/AGD1OzXNBrmTRp
YaiWdoKOOmT+vTCtbyZzKk9EjW3OJyJ+EEtBgxhzxFpF0KIt/r7OCKjG1i8E9dIIigaOh51nPJyC
MfQfFNPpfvvwDNRV5f+JFauSSjAFk12yv/zMY3SggNU3EG1FxtpH6+jejvD5YH/MI60J54U4A0oj
Ow14kefEF7YSIPv5H8hZkGqFD0PTm0mSnr4P0cjR/8daFB4lB+pzLy0pKFkpoEbvFxfF+OxXU+GA
N8uU9ZuBa8S70IRVoBlzz7IL+P5UA8EEoBuAz9hb/pDjbgRHt36GPp/4hgBoULvQDa6S/mCjvVPa
8xTUKMnQZS1m9E1Of87X1iX0gdpuUVwEXqnbR2o2jywNvJrMpLpJWURdwNUjfEojafnoprxNqODA
ST4Ap20azPdiIExzoZh18Roqu4qUpSYeMRVIZ7KtyDhpTCOsMOJ2K96iFcO9ECHCsQ6zjvzCMf3a
0KpIuP62ZAxeu+Ahc4FJpgWjCJKkDNN+yLS62qlEkVc5uBgHKS2pFkBtJcJRpkfx/9+H9OKgZApi
kS7RmFJroEJ6Q9vigQ6LWkEizB5IusNuFJAgYOO7UpuQxHKSbgBxA9iham9yskl/nV4m2e9d6m/M
PxRWhJi5yUmeS7fJq70m0nak8Apir3j2S311eCCMGVvj+Yq2jcgEwmn0nRMculMcENctAkWXkYbz
jSDCfg6f5z/BI6/WhS03fXiYIcV5ShRIGsGDO7J33R64Wb0w6gJ9f8WUmBDVoUobo2S7iWBMcBn5
u1CZjKr5pureL6yyBUJIe3XkEiGQR5eWiHLQQWax9RXSuhsxTl/8kzefSe3pFvrDxV5BEpQGOk+v
xmMzLuNM2f6atAOy+pbYr4fMGJGh4RuaomAG2O6uOLxj7L4NxqjK4m7LLTF1FbId9irCaocNXk7E
fKU+SmRo1LgEZpxh65k2vjAfS7XB8oZsbGE6e7YQqYjufZDBtYqVG8RlcEiiNxdy9YLa5UKckfVE
ZAahwKQxQ1QsnwMH2nAsA75hewff/JJGpE4QPNy9ncTmHrfqvbIxFv5UGYHiTwuj6IMKrwpQ36Zu
tbn3TgxK4DG6u2ofpIwGbzLEpcntnxkW/z/oxTGJmzvdTEBougsLpci9eXIwsXMdGqv+h8I3tnap
Jh6qDd4vZU721XqgxiBisbi1vSyqsv2OTqKJBAfptXzj+7BEXI6jkiKrDoyFZRepdojBeffeX4Q0
L8pZ7X/VpZB6cm3Vl5LIOcShhh4XK67YzwmtdFw/SO25BMTLAczguUPUPW/QaVajiPSGl8EX2F3h
QLb4FX9YXcdUHssyReD7JpHVgfPkxyJ3SSX3rPBiX7a3cAeyBjvGWlSK37MeI1j8Sir6cETM8gLM
2qth5DlBgJW9rNFy2V95S4d5CoX6YWb/PjwOXhexYMj2ebpNdGpjVcSiz/YbWWF+/sHLCrRih7ux
St8bQsOXR3eGYEwvEzS3zJ3t7ktJaRL0VnV1JxERSQLJdfTD5Rl5cCNjqD+RQD876KysYThBbse7
TygwJ2qNQ7aaUKy4WwGAJVzGrDyXiqeJmFlveI8c/l2K9/dmfnbBK4ieLLVjEiAOR2/oonM+eqLG
CGXbyWN3LUVcYNhLs98E789WTvud4ZLh6sSMNJFox7fa0qCxCPQoa7ZRIEsmaLS7ykfgXZ4s/Ao+
zR5l+nnLYBYW8KXkdxfC6KrVzaifUsJaRqGwr3Ci1C1/xhuh/0qpgl0+yNjp2hqyyiVlU0/Sg5FM
BKKbinU6iNPx01XccdElexka2OyCvynHBdsIenx3MGSYhwoODm2Y05Bh+DofVWMv8mH9xrxqPr39
d52SrNE++lVUtsl5FrBh23Q+6Pvny+cBJiw1kbCQtgD+GeeegntlYYgckbagkJcwkklOHdIrs2my
ZJRyZWoJSClvnFtP7d07HFiH4UT4Q5vUIkqL5M8cLIgdsUCmamMP698DnNtllANm/h/lk6TAWUWG
M0GYH3BuP3AHidTf7JwkwpI+zb62bOEbFMnPQYKFg7sIxg/dfc8pNwYwzaVw81iruCpGe6Eetq7m
eKMmjdheZ7JFPRCgnnQtJwCgBf15qVTdM2GuE2lqnOC6OHwhNDh2gzYhwGKqgd5m4hdtpOXVNZR1
FcH5Q+lP9B5irRFanhHR0en/i3gHrzzoHclJPjDJhLScDnIKWNZeh/34gHdmJ4SuW9NIu0NPqUl0
SbgyIcFznl0Wwnobn1MJL4Ow0ujSnOqGfAiGptBu1EB4T2idgCi9kX6UgYLh1OPXPXqGbwM3BAFW
cS0W4zd3AlKxaqRRf/RgCqI/ZRsp2SsmI8t3smNTLjw1p/yhpRQRKvdYxtPqjtNqjWMUJYkvIRjH
I+8CaMTrvY0GgnxFyjy3QuLb8M6DLKC6U5kWqmt4jYl1SPnyOY27/PvaLST6aatvair6NP1Ei+ok
dx1LO1Me/CW2ep2WIM2Dug2QbeoMLIEcMT1+kIEmbBur2HppPtg8VzV5SB9kwV2zZJ2wdPLKeeLl
mddkDNG18y7c0fFViZBQT+IZ3lHDHYrHymAcGnV9bz6qi1Y7kLdPmmHGYxVOmMn5wRpP1a1AsYgM
aQSvrPuQqnqZRu3ZtmewlUQNFZZazaQWkDFOJYxW4efvpO1DEcVwCHgLdcnal398+7AEbB9icPJn
xzBB4aGQyXXP6Ka5824i1cSjvsxUT/ns/6Uk0n1iOnmDwc+sLzcS1IO0e2bWS2lHX14l7pFKhoKA
SzIwzb/Y97z33KPontcpjrRsXDRxKx30wCYwCCoElAnSzFz3cUWQq0uegms1XkcQlwo26cjtHAcW
Hk6/Y/m8tzCIqXgliSdoI8bW9XJPXN7k60ttUJdHNSHmwgfYlg+eiEM+kLYyJXB2y/o9/Si2MowV
tSX8oDYlVHJstid2Qka4MDtznlbTImarNY/evjIQwyMooZR2caLUvDptY6/wz9c5KqFZwdL0Yk/e
vEJ3FkKWiociPWuzCIK0fEUEWbRRuFqf/Q9EBXKA7FCmOM64MmJOeDCZdf1Lfc5dZUVvCDMYCzvm
QA5pGqb17Fqw7iacL2ipkbUKJclF54DO5D92e4vHRCLxr4wD+pCwGKKhZ4JPf3TSgV/rWlxtHR7z
hNcHLeuBSkn8c0dLqEPtHz3HBsiSMb+NWTWgzATAuYb0M50IW8rBggIN9LK7MF/MamixyaygPzyP
MLpwzHzGHgWC/wcvJSJvKG0W2AdCIdgoVGRXl63wwCs2U0d/PZsM44HZLK+kY4V889izhXB/imFf
u8oC+HE3fbglADJs6P22LpYSfG9Y/LJ3Th7cbvjJ80AKgEq9Wj0dFjw9PUq2g1anZfuPEuhcergq
e4WDUw5dEvG6k2pFLOgl9pX8uqElCyFMFxbpbnY1dy/sJN9fq5QKTKj7q+duDwNMYnek6CVp9a7d
eM7oiaQ73OZ2lG8zkHpB9QuyN5XP4oCDPdlabvDj1vHDjUz1lT3NTPceVy29SmZYyhBEraXsQN7G
Wz2xieCDY2sRzzKD8887JeUFYBo+Pfzo5iPVGXubPHv+1twDiUcfaYjQkT0egeGJPKzR3raxpYY1
e/nGPanodMri9YboXnwMdr9K9JI+hQE7sO5enTxBrYC/mUHvGclFydPPGA7LQ+lIIc8D3pB4yX8U
BTk/MPSeO+JHSyP77xug0DZ86/saEdNJLFdoFASgJZIbSoPLZrhu635liirwm7ETOXnwceZ7nzZO
QZD1WDJ05gAGiv4s2XOlKdHp8yMUhKJRL0KhNHrbgasWzgGmK39SCgNAIkHlp323kSuTHfXgnFRF
x/S8cRl9v9c32tk8ZeBsxGe+5K4Zl/oERI7LmZ6fRq3H+zdwsc90RCmiYqtxT2zeamnDmB5bb2Qz
ajnicL13BLortepFD3srlIG8yk5tV9vhkdHT0BWJbFavv1W7oWESlI68RsoKzQJ0RKRk/58Hd1V+
c5nwhluOIQh3dTYVXJzZi4GtgqloqzPIGkRX+MJmVUeAYRU+MAcKIHJCEq2rTzCXNf2FSNEVY7YJ
cdB9S4c+jaor5/8C85KAIR/AdiWpRPXBXB+QWjc4R5bQMqz+X+pmyRbqfrdSt5sLLvP0Ryyq3u5A
4oLS54i9cZebCK69UkJCly+cdOySIeH1y9Bv84crSGLA7YvjeZtAC5XVuuOrQLNSfCGxc9ZsMYR+
IXihrzm0e2fpPOj0bOy1I/KSTLT2hyjOWQ7RfB9B/mOxnyIdbHMvr/8Bg4izqgP7XvtD1q9kbt2t
BWpchI3cYdrb4FrkQ0g+QyBa7ykS97JfxfpVl+OKe4ECtqJLIuRPYEiHn10qHK/2PFWb/QMqCqAO
KX+TMuEwDNb+b4PzjDWUFGldPL4jUiloUiyDGJpSpi7aVq9h+PHJD1uftQt4rHNBgz8uwPfwy5tw
5aa3AQ2kuIEihMX/1KFEpwgV5N9AsL/jDOSEWQEnty60dXQ+Mhw/5W1XGmWbM+I4Rb7jmEclHAfa
YSTt4+BmorNlCDKyXNFKDTNwIcHWTciKhQMVx+3ky7uOdRH7CcyRUef4mP9TP7kx+icwXeCcNimt
qfeF5E+7dZX+aPTtNd8gopCZZWixWfFjDvoUphFO0/BabP3QglSlIulbGC1kJY+kZA6ZDrimI39V
dUDVfnNak4Sa++pIYFqEUaCvg9XEbp7yoKI5rS2J7l3VG9jDm0r6KbxVokrPhTjIDqjbZUBn3Omr
FtaAC/U51f7i6o0SGMbXOaTDeprSSYpdoW+cadu32xnGax7nt4dE3DJJQjGyUxTd1dQ/fhx47/xV
CRIcvKs3F0Zz/YuXBliDiE1hkQlHYZi3mUN+SMFxz3XPtplQWwR6yGhA6JaaVIyIDp2edm0Ji9aG
oYImLevL40rPPQuOtg8FQQ0dn0TiB6oGzq0MTEsKiGAzHm5FCqawUdHZc/f7jTWXBEigYR5Y01f4
+8cV1UAbtACDFMCBSOZQDcUYHvfwrwb9bW5s2GK4OaFZgVSQZsV9O9EfmXLNhVTmXOhf3DTLf1Zj
yxjpPxmlzYrt4rezPp6VGZOCPGMaYKPR+xQhKKmtIYKjPtdH1egN/OO8NkB67cL9j4yZVH1nYMGD
znRPQ6H7d8JuCQFlWzv39M+d3Dfs/26M8yJl+l0m4RT1JVwlXYrujzr5Jg/m0RzstwDl/QfW7CHt
iGrtHQNNwfi1LwI8iD4dNFejyCGHaxW/V/CvLdsu35A/TJED2G2Np8aLN1TqjnzpeDyTpNTsiT1t
hdfx6WZicNolC8urbgRkQPhFKUMv8K25Yr0Hz40/P78m1T/XL5Af2bAkh1BTXncRvgWCRPH+ysG8
i2rEozME6WA5FgHEE1u0BEj6Jm3Km3GnuEVBSjkwbg4FG7S9Z/xjLUYP06Ymcwhg6MGwLzCtdSl2
k1lH2dzv6QGCFYtTntaaEQsuy4vB/fEtlKtvVInqZu+a6o1aLM3a7cqMfWofq8lahuiHCpjMxaRy
ksqYVYmT9ddhjDSTfAzOMIKS9ImqhT/MQ7Pj1FE2DsOeeK4aXBXMFEyhx7kZ9zbEoDIQg54SEafw
38vo2iXPaJlV7iuj99abAJtmw/2JIjlPwG3SEhP5aeKL2w6Hw7bYiCptgUU2dCIroWOCO/Z19/uV
jVjyY/P4V8nfPdTlguC0I115Gfg/QC+vtP51FLBGqbDuRpmftMgCqdWtRUxdt8Q/lT6CvNfde9yi
5/GIwSIZnffCM6XBHbfi9HyCm4tNsIRnF27YIVG1TvuMd4x7/ygr+/pc1jw/PffUAWBJAHNxMINf
XHtnWXg6PzeRVUTQvFC8tP9uMU909FncEh9c52F1qddPs2pZcvNBFjloZEASWwmtln4LND52PFuQ
KtNx2Aaae15aFA4bFRIBLHJI0sNaVZvrQLCJ56nlBA/vb3W8ECwNXYjYWKM/bjaNhUsmqv6+9OlT
Eoh+BO2ycu2wW8fnMpxVM6t0d4BAUryInakyg9P7+79BnW9YaaeAR4g/HeMQsIpl0++6SheQfA5r
rG/TLUkuB2QkMKoSCxbnMINtx7c4F7nID1rX9d224UieZ6Z2qas8dpgGGsMGEDUHDkOpV8RD4AOW
+P7+CQ9V83eZ53UAZln2h/CcVwuYrA1nu+PGgSzZJ9aUOvkcbwkOfctbPOC22zTwhUH5zqWJA7lH
25DtYyqWuqhltyH/Y6TX8o4wWvUBpeB8m87j/7pUAv7zjLQqyY0jULTi3u8rsIkpknpxSV14uhYN
oKwSzNNCpoWcRhK7n+5pnLJ4sjKSO/dKhFk/DcDT70arluR6IoRuCLLUFfjQHTC9rrhIpbhpjZsL
GPiGZzDbddCWLcZFo9wYxMHOtpcqGq5f24lWiH8oc8Zsb1pW6AiK1KHCR2d79lk+GIxb0EHoMvJL
i868zcGWfwQrj4VvpR4sgysff1E6tVqDjPqkkhFnBZxFC6N/i82j09dUwhLMbdRCDBq0CYMwrFUB
4elRk9B1yqoYNGbaEUOAontUUpeR8fw6yN863wcYfsn1OMPMGqEiYoJ9qlNLbM3Zc03xYU70Tuhj
uL1OG1CmFGOOKDFiWNcKrD+ylqpTQadq1A20aEz+8IxHXfxEF3O1MxeRpO1F2xV8vKbpywQDT2bO
gFrTFT+CqWy8q8cuOH9AIJq2orFfbpoN/ba8RkXk97W9/sfPocMTjJ6Saptmd9Ct4I91KtDMHv1I
S8woI/AOZNW292LUpuDMJL2cOBTJyxXcz4J2yCoyRxWeGOHsbeKHl1fZ3rnXu3XxAPNl7Js9tTxh
t1l/6zBiq6u7b9pSPRfBpBQzjvaKFJW0jwgUJkBOaaVdIt+bUdNnV0XvINlw5qvPSCZ27Ausiwwh
ZUakedpxyT8cli65gc7F/yrUbH0LZ42qzhBvUY2Qq/dmOtKZP5j5WefNd38efSrEMxePQeB44rX5
Zb827XsGLmmzssg3415ehjHNTBSWCGbyxG80wjCgCNOmuh8FEjkaZhNB2dPOm9We1WIfAFLIe7Ki
DrlM4IHaXBFiuFxPPVPgg1UOjbs4R76sHbhdZwQbkc5dVjlbEbCL6/dX9ZvGRRs/91OhSMPNIMd7
KPsi33c3GVe9o9U6UA1yqbEjE17XjIRlbDnmzJ+efJTXAK7hVDcWo4N4tRRg30+5eAIrXNcxT68s
F6DVzaHU1zmQNbK+AazAcOariroOuNNN4WbyLjXzrFPMhO8HrI6bpaUu2Ie+v9Jo5KDVbw6slQk3
ns5nZFOEzPu8lovqSwHGeYS0aiPn2NbfuBxKHtwz4/cu+EI8EaWCc+odrwNiFNe/HXSx7yvEzui0
DezgXled/fJCv+UV0WCFBSwJHvLJ+N25r9rCH/ejIcHpxnVfvGr8IABcfEf3Cyuk0CcBJW0uQAtY
6nh6oTL3aXmavt+tO5QhOVAI7mOi/SSC6Ri+SR2Qv3DyqjaJcElfTJqsnTWMxv+3RM+ZflFajU4T
i6LgEiVX7BX/elpFr/l4913nZciWbYPDCGE0BPi14K2Fj06zK/VdTIQJTem1GgVV8/MndPIDsM4R
RiaLSa/8Q9MwoVG/Y7KkHyr9kXkjnuZrIScFJOMiUDx7FWI05PGJ8MuV0gZ2wE1ySWjlIKaSbKhA
CuWhmr9lVqrS7D0DcXGI9kHU5gjdBD68vHyNtr4418X+9PN/69bUi53+F1joxgMkkjiu+rJcrj0c
BfTNmrTkYlzbOrWqSjPSMKQKTfm/0l2+H5amKKfDhPTuQ11ZqcOP8NoYU6Kmo6P/5A9+mrt+BL4K
DHJNg7cjP0xdb9YOWbrDHeV3le0u695sYU6BOrlD/WESRfqKzQd3XjkD0RsZEct5+uVQXCt1aSVB
4vStjO1+yuD6uvkZo1ZtPO9tXFEvzg925o5iZYugdNXSJ5azVg5tu1ahM025vWz6bCrNByyVAiX+
ExTZbpUO/wR9AtptJm1ajy5v8gLruZkWPFk2QXxGey73a+qgOPBRZ5XrXhR9e2fHPJ32FnboYHoS
wPcqvUKqLbauzcuBzEtNzyDz08XOVbVBn0pv7UAm1cM9LryKvvUOlsKDDGPBJ/NJ041EPwoz9NyI
hnXcId3nNwZeGuZZ70WK8eYi4MTy/6BIGPbtb8tA5dwxLd/808D3TNc52aO7IQjO71FpLMCU/o5p
Gy2qwz3pQvpFFXtdq9h0IpcRfWYzdKWRH8voBRsfNNMEELyJpt0dEkpuJgZbG3gyS45FQbxqH4R5
Pj8kQTifpE37I2DHIDTYzeQ7Vs8wBTv3VC4GVgx4KPmMS3PjYdazqGUPpwPnpswRV1ifeEtTeFeX
tTzwLnL4NMM0FMjfjtO3fbh+xtgUK4tXRN37sG/HOBKKZlB7VnIPZU/rIEvlF08tKAvVrlIsCnGE
cMuucy5R0mbW6JqYFgdUVAf96fy4zbmAuEIjfiZOukBJRgj6h6s3pYgX4grvUaWv9K5P4mqZ3Tgy
gPXw0gdJoAFY1Tn22MkBP/KrOLwMvtrvEhZANaiVcQhXn1PR3STWjTXms3LUpL/GXtn7jh5FaVCX
JytXapBgLj28oET4SkrYME2c4856oWfJsb7tf63BILeUtEw7IfyDh5w8QG8QOUd0WhKdxJJOCozf
SuJ22P12WZqRC/b+7OXYnw+1j0lhX+CNzc6TPmVdf/BwqpRhme9HoaOVHTVmhoe7WC7GRVVMVzEc
kIK0Hzn3ypy/HtAt9caKZVUU6g3XfgfmWtyZuZBGIuPra9VZ3Df2WbLD6qSGuMymNNhomRGRSgQR
+rjOkWz2wiTM/MdeDbHkCFsnHmOhF0lhMgCJQB6o60eZxZmAd1VPud2jDtIr+9+eEzKOF65YaqfW
WDG+kD4c5aeleaGKT5WPWZOGhGL38FknBDSkvJCBsI0jdDWxboI7KYcSB/kKnXnPY0iwJhLtiHdA
RSa7XQV+a2PtuMIKNYrvpHBcWyQnA5XPXm8MD9t4tcLOhWGaZP3Gt3ElKhY11GRH6W0nuaoQUX9U
27qGWwjjGBRUK+RyXifVidArnEWrw9pmCbMjOFkfm9XzC10T1nQ9Q+V0IoTo5mtO8zF73kZthfLe
9sXKyloktYN/8JS8jo/anvQ3WDOleLUi3GBu9tjZ6o7VzbyJztk5j1cIgMgUF8I6gQEyVMGbeqtZ
S5KkJkfy965oRmaqtoBAiXfvkyg+OmMkdyQeQrslT6v87ZrQAtp0UN5Uo6t9Sjbkyic+0c4JAdnX
0gtkw5zJ1A0KiQfYjUFsdOxdx7L6cpIBlYoWUKmAHt/NR0JOuh9bWVNGoJyOvuBqZ1K4OIbzCFiH
z60/7aXjY+ysJ8yYsc+kq8DU0PVdfPtC/EeyCoYNvh8N6CY//XbF9pVRe59beIXOjQ+xjEhv7Bfh
mPzLDymjp8wVxImcVf5R89ry7ipDOhsIANzn40wRdZweHdNwh5i/XtxlVkLAOJ1M2/iYZ3acropr
JyHbFWO36SZYBjftaqyY6shdplmy4YkfH1ZVaE8L5boX+yAMMP7+O4lxN17K3ZzpKC55WhrlDXLX
A4C2VretkvSbefCP805i0r8He6GVn97JW0TnR0wEeAd4WM4Wd6DWJBGP9GyDy+V03mKpwoz8zvJA
Khh8KK9VmvO9jW589w15X/455QhuokzgrOHyRDClaZaXhC/3br2VcXGGxDz5Da8Pm8EDVaYqvkUN
wieGUu7twdYbBJdiOZBLOXxhXHFkA6Oh4hnTcGRfTrD1jLhoRargBC8ec0f7voqxGGIWAZSKFw12
Yx6/+yhjzI0hBng9DB13OaqnuJF6YYh6XjOdP6ZLPitqK32Z+h1j8+ZYOdKJSC3uZhItESVisnY6
tZLO7avOodGZcDArxMO24h/V1EotiDuVc5FQ9aRilEAm7+rL+XIWMsN9Z4GnvOrL6aJ+CHgf1dMM
IYqtKNpXyBj4rASl11jvZPNMhu7/fbYod4S3JLDIn7tLfHO6WgQKsRboBjY7cu4WH+6+IPZlOA3n
GkkJfTnnQuSTNf0HOuBtztfgPBF5TR+aUeB46U8R1OYj1nM/n8S9UjpV7GRkuCgMoLaNU5WhrhpC
3KrnZK7jWqoxzL/tH4d68DRLZbTWAHnd2CzwCY+3FjMP3e9BdvG3duQJuq0MLDx3lIADEIpb5XL9
tn7UV9fxsy7lQGMPsLVEVhjewFWwr1bE72QlpBqcblJ+jAtjr03TcBO5hFzh0saPScAjLyeM6tCo
YsROjCf1Q4L3tp+pglMpeIZtIOfZdfbaBwUgCOkNVBl8ippZMwtyu9qW6yxlx2BbCs3tS+bIekH9
D8IbPZ9dwc/Z7MBl4HuY3UI746Zuuq564nnaNPZGblXahj/MLiE8VvEZHEbB4J1f52Ls+Ps5b3hf
zYEWm0iW+kPGN/c54PM0A8Gf1hf7RqxE2fAYbaSM7rUss40cA8/1xw7tpCgByXouIY/Iheb3W3RA
muXM2V3pD+RAZW3kZjIfR+eZqwN48U6EVnmuGZcphuO9GEsXRo85zQ1edJTthPSc33u9c5o1hraw
OsgYjvysp90+xLx26oGVg0Pjn3OArLVMNtk37018rc5SQFmX50Ndusm2Sqg+tXOndodBGGuFPQOZ
nNicPYpFxkTeOIXJM0Qr+srg96bqM9PS4aRX7oVP9ZJedppIFeFJ5Zecq5auzwXPVjChm4nEC7X6
uJV7RHPG1rrLML04qekA8wmnllSj7soONre4yDVmVGIdqBMe8eQZkijef4gJ1+qzQHSozU8uBWDW
f1AF8eF97cxbAu81YVs2xcjJgfgVSU414FsY5dZ3WOjBhE8zQAcNJpo2fkv4PnXuYjOOtX2hJypM
pfnba9VEf4AfdD1KUSIWbncTgSdTib4UTnygcs5aBBfDAJcJ30E2eLBQ+RkvuhO7ENEnn0Fv8n5p
mL38W9nW3wRWkv9VjqfBDKVDKlcZ/x+pLAANRbtuxRHI0cvdM8FB4eW1CGyI1ca2Ic3vg7kIYtVd
ZMZhI2/RT4NPJb2W0UWndph9eXDhKnlKNEQdYgdtRhsAmVU3tg7VGka1kJ1IfK1e+PV7hNJC2nCe
d/GCExOEVRPf/zn0lPqg0JCV5m1VK91pLgQNCXaaCrKu3DlaLUBYusMIUUoZukPLPPZSW2tRnY7B
9vXkhz8tdriBOqrVJlBap+P0NDwZr7Wz45EGM365Cx5OfEHa97XSIe2ne7PasPk3gd/FP2mUzCWI
y02HAXntEHzLzUJCl2PnUO/zYaF0SK9ddG7/5/SErPo8w15na0QheQRPyjFMlEGkKKH8lWUehWOp
AChjz8DqlHK1o5n0+DiojSBrI9R3Y4NgJYdKWs0Lr8b+zp+Fta7pLRk5mQ4BmbB8ASqdHRAd+Mdl
hzwBFcthyrU8zWkvy4/Xmzs2AyAzeA7fQ0/x1qhRZ9+gvFtuCLeqj7wq5zSrTXm8fHeNd1oICKJX
XHjA538zIS+VZrCOt3AzdI4pdx9Fb4zVAeEQSyaJIJsgZeNg7wHFD+AWr8G0VlMWNH8FtYuIAfWw
2BwllSTAcdFM7cMZMQziLtcEyGGg0Et3ENe/aF93SMZrF6tQECJ2xOMrmaroT9jyzTjXRAZ9NvOs
N57ySimJAhqW7jrLbGtIkTEG7eScRGXMoWYWwSvBHPSh2iBu1UR0R1zg53rQloD84FQzi1CKhw7b
8S+EG/ozyDCOF9t/rnR1liWXF/rqQ4aQmSjms6VZOppK1mruKT0hHET2vayaNxaGkAgASP6ZFC1g
ADIUA6isY/hYvEc3EZ5QDOXBJ+6MKrHONhC+ECRVBs6Qtw1zYaa24ddtGdTXW421GebvaVL/av08
eENXW/9xiPmVVgIJerkunnjhjekivLtQ4cvafK+bg1Mgq1V+HC+fOd4bKn4VQpbyWqpK1+U3jD5M
3BSksG39PMumxd6mlopJ4XD3bYSxGIk4zkO+LeRczmIRpCDM35mMCzdzRZyhzHvbRXOte/WMA9kp
SrpWWqmERPSkk9+etS5FkIXnfafiBzhfsrn09T/0/KHMtLkMJhF51RtRZ2XlT/sKXbEXxbWoPXHm
6hTT76UiGxQX7PZvnUDVlxZMENsSaYHQMBkarlZikQf92C9eat1PT9/Iw8q/ctlx40GAVmLph7Jh
XJdqHUTa1duzgpqyyvdG8ZOcwQtO/eKlRQT22uh93A1SX1upH60tQOQ5w4FsdFeW3srRZq+4E7Yn
1xpMoWQFZsHZAG4BVO+SCqH4cYJjZYEDGShwpleeX+cRZwvjYTOpatORrMnqvdW73Ph4jaXfw5KD
RuANziB0UFq+lIWZ5B1z+Rn9rplWdHIjLTA/69lwA7olEpEekuoN15+3+7w+7iLW7/xm7dhliC23
/rjWg0AlRoDV2HUUp/eMQSM2ADpqFFhm56hAhALAchzlC4IPwYxSfSJCRDA3Iu05ak4WgHBa9BS2
BBK18Dium7VvILYV2fPSy7mDa5tQlXdHxjVVBar873e0Sfb5uhKH20x7lHhbfwass0rVatW0D6jG
7SBKrvHSP8nfizUegbLAIqWv5RJf+cfb/1kO4tye/IvjyXE4CfLtr5BHIe1CUyOyaIZfW0VJYDSQ
UfOHpNCnAYyr1CJkpzVvueDhOMS4Krgc8fCB0bMcWYei7ok9AZ4um9YbA1hStCHkgXXyYU+QjyNt
oTC+W5O1g8SSXc+bRdtllEqrHenQjghTnDp9ExFToegr0IQhzd99qd5rIZwcoUZBoUaeWyCpUotf
uGQ33fpznOiAqSE8Tzn6I/pHL8XaPojgGlxR7jy1dq2gOn7fAYAK+8FzzJZTucfG1mHRTVhF/EPw
hyvVRlKarAkO2NCx2udIG3SxFo4zFJqLRjIKperKoxn1D8PUJQb8tlWm+hTazNDMFlpRtfoynd1e
YLhFLIRCoMwA5LQi/WRyC8JNSdMNnnd99qYyYWH0WROGbU2oq+ApqtoUl1AXg/1/n7wVbhfZlhXh
BQMyQoRkq2T5iQUY2XV0BLtNpeRBU1uC2n2xbtofA0jZ52oMLGAquU/7Z6mG7qtKY1jI+0ZGwJi7
Kl77vLtuEbe0V5fEJ/KEXsIjaesgOEcNsjtyVEKEoxKw5LDCrcq8OXjNOo6Kj7vz1mMVQvwzfDz6
JJ9TTZmCP0w9e3r6EVLhj49v+vXRWnwgCIcNcy7s6IdbEBd0k7OTcWGqvhBcKJk2KqgOw3qNWXux
1m+raTcQRQL/RFouHStZfnW1z5Vrbqs5h+yO15S2SZe2BOuybhznEvPhsn8xF300TJd6lw7eoxLf
9yKTpgCXmXkAjPYIADj2sYDsmd5qj6N6dt7TatD+8LZx9RcghlOAdOz0TPz6SqgDXA4qh9OX0hdu
o+xUzk4UM/8N8aLl4p1BIYspNl2NGtp2uzX/7dhYAIg/cHEqIlelnTHL6+lfvuDwASVzEfj9DLD6
M6VNwThjQ/r9seqgz2urZIEGRsyRy6wo451Im+dyMyg4Pq2bHBl4Kr0dtLQ/tGvR/zfEjGIvsJ7v
+7RwH8VVWXVWojkHMS/vOt1IzzZYffsDY3torj2JPyz1xwbyUPQs2C3KnLnT5s5XdnU1DT24J1wT
JL8p4ByMIl6qyNLIvHZcB/HVUBWEo9g8KfRJ4GPwfmZIuHnpAoMFs+rXPXw5aUUmDqvdinLLwsn5
/3OcYtxW/Cs5flQSRzCu7HihFFwIKDQzpH1so+xwWjNJjuHRgyFYhlJbSOXsgPOosqTkT44O57gR
qIDkQD8QFOgtItPtpMzqq/sOWArU0nxupU7M9afedCs/EbssUrzC5Q5rr6SONnezvXSxm6X/knwR
F0rq1GtZD897Og+NT1C3OSuGgq0J+Tf9rskAftB/byza0o1aDelI3Vw/bITkJaEsMCLtSlrAjPl8
l2TUJ1dz5d94+8wjChR+GvhbK9wpLbwhe9/ZJTLg5NrnqNhlIvcUU/absznw6EM99YqmVeWop15y
TlKX6YKar6/YuS998sk0YlTtbHy8+wa8prcH2GX5ndIsfzSgnlfIpWLXJzhtu9fzdKalAlkyYT8s
UGM2e5Nu6d6pKhWiBP6/IfMxVUoGfrISd/8tF3A8/VTAITZN1Klb2/sSQpBNUUoQPJhTbn8RiESU
8TtRYvX6SG/TUoNRC0dojI0fmlH4kHIjWev9eN4kh8yIipYjlphuBZbZ0LN5c9D5sxprZMjPO7sW
SXlwICkqyNfZsOfgK/OyTTRTnSGnHXdyZXRwfwH7c5qy9mVwTsKfw4dBSl/n6ihZXGQKOTRXjnTX
aZf7KpiOBZmzkUM8xba/1SlcggZkF9A9VRBt5qUzjEjACVhDMoATQz5IObxYsv0xXGwyUnbM2q1l
aTo94V23+pweGx9NVOvlGJJnUJqZoLbC5atAmgklAI4DztH7Hg+8sFZT8hjgbEO4pEK9IDhsfoPa
VgG7cRkjhc0FEbPwv5Oy0YWwgYUKwhuRWg5fzDf+iDh4C4tFnfAcBwSDHaDAQ36mGYfNxV22yC+B
n1l9Xlr0e5QQ+SDpnwrCZ0+BqgGGHCtsnorGFZCj20Pm38j80mZyOxJmwRjoBnqbCzT2YdD3MFns
BVinpU3SWOOSJz/nikkekpTXsxnXVTMzZ5yEcC4CGZLB7roGr11FR4x9nVarWvkvNGEX+JX7pSsy
4R0D7KIgOOCNh8b25sjhkhWgoYzygw6wIZiNi+4XI6Y4KFLgIXD1q0GY8fx1g9psMPal8nrZNxjV
mnexul8JAwExomGY52H0jwiw2bz7wX8xmKg5uHBiSrG6QGSiy9fRojJUTn87N0GwFxSbVoG8cbf0
G5M+S5ha49+zFZDlhbwKbQxmOCQzpgdnVXYiagppCdWUSmMXq2z0MCo5S3xIR26vHRvRQpqabKol
FPcaH6WJIHoPIwmefUSt6wx9ZB8jnop13QIc9GjHdKLVbf4Kc446znhfenS2g5FhRvCz5IkFH5Rc
8LQqv9Q2HidsxyRS4Zyp52eCnuHyhj6BgWIgAcWi/mk7tkOBc2+ourCrwGKWyumW2UClANJr3ySH
An0NWzzUZwq6Pj/BMlCN2ZOxXN6liWxb+MaMF3hkVXH7jZaXJJMr+ZWQpAO5w62F8SBdX6PAGJ7Y
/WlRvYGYmMkJ8Q9QdPkk/3H4YwCRBo7LqlBg5yZ6zSdKZrlQVcVxELOzm1BY3JB6h4cd+OFYJcMy
w9AwdeE72RU9YQYs8oDHQ3xdN+6Yq5bwfPVdfcg2q03+Txw/epagacib1J87X3sRmWfp3xrhVT95
1KXWHzE7buXarvKcbQ1o5r/8Yy1clizVO4kkD74wtovNPw3f2b+moy6UP6RxvWGJX0ffNiDctHPH
FXHdGhFG25DJlNH0Q1cugBN6Xhb0k+PpRuGAFgdREmQhlmoZXPpNYACcPs3LzsLlGOzYZk+ez1BZ
yaHHFemJrdl/KHeYpMkwGI9/9K9IgpzA661eEIv1WIwaBgTkum/7o1kkCJfNHb9MtSTJ82i/iAZU
Ta6eG8Cp1MC1G5vOLp8jV7U5IEQRX4iH23EfXiKs/m7FBD2IG78dztc4R+aQsRR1X9/5+mY8O4bM
AgCNecb8cQ9QY4zP9abUhbyX6zyL52ohhx+2FVY0nch/hhuqJHs22nhO4g/n4VZu7IqbSMYyqHW7
7zoKTxwgHC/yLdL1y/KyIorOBsG+zkv2R3Eue66lpI+1To3ec3a9mOqkrNc6frMR9E4FNPQRMDYn
q+fiL1Whr3n/DERq5xkbQGX+7IWZXUpo0YZYyTMOgM/1Zx8Gq+vG22eobyePgpLAJNnhD1pBDWAs
9nM5CkI5MEy7UzWnhGS/PMbfMM+k+bCgQMdSxdK5Ei1ZUu/qcFk1gC2Yj3ctzZA8Sw8dBx+d+fZn
q9fVBnnCRoIqkEVR7ItJY6hYL8S9xNsPRoqqOCRBHQ0lEy+J0IIQNfDtPvO2yMGSGKGQyRT5l/8k
fCc7qSn3MUBAFG7Y44JSE50Ue1/wr4encLg8tSzhzPoYbVJ0wJlLw5DlHDHuNefO0vbeqS+ssBbp
79+4pth3SaKK4LLZ3AZA5LCX41enZxnofi29LBFHbC0pOa4kSs0+YCRAou4mQ/idgosqoMwNb0dH
a/PfiyNf1w7tx0J04YvyQng9/AjtK0mtjNac0x0vymxC7IGesbkus2iBMMG3Avqwaz88rQiix2YG
xo7qlgbVBObq4+b/LQGurmRLEBitREvDNsgWxa9lbNcNOMfzQu9rVuOVzFIL5XPxLSqd5WrIK2ba
qv01k1l/YTYujbIEvTm9h9jjG7WIKCrI/U7G4PHUeWFtoBw6OvNn7Ezd/faN/8nIkK5572kCXjRz
JZoXXSvroW4T3Ur2/CL4iLS3+sSwdYTN4mHYS/KzhWkMHPNNckEv9YC9iRjXpmaApv4xf6jjiW8X
8v6QzTvZhmD0lzBsD73zM9wEmvYYzdPrrLdzwxZKLyGQcrthgVwoDfPk5QspWynPYDVI+F5ihrLr
ns5xWdqpRt2Cj6LuKXCN7VKfNqoSgWZZwUY9ReoaElTl5jp+GzvCijZcr1E6NXEpfDrkegsWGmnB
6taWLTl9qznkwEWQ57/e9IXMfUEPvCVt6tKD9ZiuCZLMiH7WXgQ1Vn8DTTD/D0BI8aKnh0L+PFrS
8s/pSd9ZKce4LvGeyo7QIpU0nZFm36vwEc1lnJk7vGcmA+H9UnTentFxr+JMkRGYbRQ3ZcHjZ8+k
1hlzyqd8qJED0Y9Bq1tH77oyIrpaHeXxov8V6PpB821QosO8AaBnEe7aJBR7hB6PrHmbV3hCtsjZ
8i53aot3qSf+ezj9WjEqgPJRpfRS0Pj3CVvz+9JAeTyvfgMULGMCuF3CnG/5FhUOh9euzWItM5jS
8/KPk5QnXFf6SSEE6dsd5GSne2BgQ92/muR3XPicZz4CmS+5klNVxcw+0d1HSav5qiIZEtY/fmHY
rkR1KUs+EeItL80ba0LS60oTDVn3/6bI+4OJqD/GwVGHR17uSIvRSR5IHzuAxVvXnNXQo38uWhUj
YpHgTuQmBHJ55tbb1uNqFV5ZWdvd+LxuXV0H0d2YyFtCr9PcA2IIkzAb303rcS15SaCm4V1raeQw
STC7qY4a4SW0hilerz0WdwNwj5CVAe5mQhh8teOxBNzjX7ZEvNY5kPj+gCLEzfilJH1Q1ieEep/o
OOM5wpU7gSmsqyd3CBk469zTBm/FR69BTRfLjD9jra5GC6yUipjR/GwpfLODiqzJBWeW9liMdU97
wvUpYzkpvi96sY9SkNCA6Gzip7b7+IlZRWVqZSG1MvanWRyx/4DLLzOfqN6ohRW/EmI+ktTLqNsn
ppkbLuOZQjXZIPR2l5GQd6Z06dxkGElT1PcbCAixwlEB8WdC3Tlqd3RDtN5AWbQsBJCi/MyxZWBi
OCIgbHOukxs5ZokpkZGYcZP2CkVqOfk5mgQrw1MvlofpR6z6TwSyGoYQk+uESMrzuB2/xLh7g1wv
h0bj2XELrdNx4L7d3f8+ZzQUj7ArAlE17IJr/yqUbLLgYtwLG8J3YBXAo0pYTwYKxrxzgGIaiBRg
SBk8WXzcwptbOg6ORWM3ZL7gpECkA24uiFwblxYbSZbBoia2n0qkCgyd8nsAYSHobL4IZ0HrwK4R
w6fUTj2BHVdgc2Nyqh36ZB1lk+tVslylPZ4XdmJYPM0UuvNEyr3Lf1AkD0v2DHrWSHRvZZFStuY2
CdWNZ4aCuZ/Lp3mS+DWkD9MC9cA6nWSJ/Np/TuzOTDVhptRZnb4euklIM6+Y1FbuCrEnod7AHv+R
97I5797j34m0MQPo9th5S71aA5yHqxAElvuoelhh42qlOIMOn57U8UEa794V8DF83EHJmO/AJYeN
nKCuuIn7d1y5srRhLB1EuBkKn14X6ulnOU+PDuAe8s9XimtrgF5sLCpzV8s4Iq82qhjz6gD5iKFP
nNfFL8Mbw9/QpI+/zf8j1E5bIaFKsr4U8+LRe335NXfpBIlYZp8oIcmqvdhwG4F+Jx+M5fB+LD4J
rn5eYM77dM9tYYOWlnF28E8FtWcLdV5ajVXYrn4ArD1S3GC3O+p+EVmSkq7EV2fI/XV95y9ueItV
QWm9OHuJjNLGDmRiboKO70qHV3zVlrFL7guy54CQVFsXqtQCbQzrPuxtwmyDBInIctec90t1iIhH
SR1OK13sU5KnefaRzKutGsCeHMFmKrIIeB0twpdQfACFixsjr26OUj7tAZzaE7K9AgX+OlQQX1+6
IoYdhEvRQaIU0zj/prYCyDLDf/IjqMUoQMav21ZfAmf82L+3oUAXHp0GU6GY2hOGlXFUmwH79CAz
wkaetToSBKtr2egS41pCjSGGYUfWhvmHf7yhZvFwtQycu8FJLJBxZfsZS+od/EN88Yc8jrGYSaad
wNGuxGaWhgD0U/ubRnAepoX66M65cPMzuiCGyu6wY3Hv7ui1AgOmLXNOl74/3CmE+4r5LKKnmeVr
V6SpM3wVFqpR/p5OQoSVuAv8p/r0d+QZmmgdLZoynqjWm2uoLuO32zKvZqBf9fTfK5w+MJM6YbA0
U9/7C8ga4r9x9wcLpxa4KEjRuTq26nS8Qd4d0gGJMTKYXzQ5e4AynFTHL/vEWxGCYYQ6RjVY38h9
hV8mGH6utwg6jTyNLbviVxGvWHZgWi2wxOzWvJueAxKy6jMVkIjHl/NVSofkJl8HO7TcHP6tyKKx
Djkyo/LtMrOesFNbUNUeOiqlWf7Fd+LYDS9AOhi7UkeLxyDNSaEXTchuWsINQAbpL63ycyHfQvhs
GcN4A55ydaF+CEktHblsxDQN4tQNMdfYEzyODPXcenAZunmDjn9s8Uwe50G1AGMaeV+9jH3XGSqV
ZrZwsGlQr5sqh3CGbqqiNEFjUePz6azxeky70Eg9W1nx1+hZoMDFSdENSJl8AoqfxrJwcaMtkhG6
Ui+60FhXVk0ZUeeYC+vSXJsD6Zar4I50ouMR1AaA02b1smAYvFw75FggmdyLX4xoS6ejd31GxJAJ
XmgbDnzv3p6dvi3Y2H/j9LqnEg1tjjmolhT3B42CHsnltOM+c+P0O8neipKxv+iHttVQDYrV6225
OkxNwApvQZNig7QdENlYjEdy0kI/kQXAh35wqv+2TBS6MUFWYvnoLtV7+zThVDXnRSZAYs8pf1De
fdXhMNgjzRbXDUQBriLqzg1ScLbhXMLbHvhJJOcCzvm9HVC6Ol28Fk4pTnKnhiefmOeVJ97lHO8G
OHbfeyl/N6zIeMQqkXNveVwwiuAHILi5tpe+xmxWh9I5IiiSWxVYFcXPgSKojO+gNyEjvEm35NmP
AxF+jDTI0PmK+Iruu6SjhXs7rJiNBxggHDH2+z5wlR/cxhMJ9EB7xR7d8fvcTMbLxf/sMtc0cv4P
9mbMVfP5KgdEz6MW7+IO/mRVnMym9cPxYA0ZMwKE2IB+3bIbGvDCqJ90Z+2YzVj0sScwry8fiNfF
x2sp4ilVLviQB7MbRuoUoqdixfqLL66o1BdtjpJTWuu+D1RFJ+jHUdg7971lpMfW62s81y8jPWrL
pZmgSWdCbEe0a/l+K0lac0HtqCgWCyzk9pOz6cNBGoFk/DS/uvYluLOa6ia3DP0EhZa2cLVNsPPF
sFxq0ZcylQp3GG0fe3U780UV7TvPVrKwiC5dwnbRs3nSdnKCsCmIskxKqN4bgIQQ2X4mJIodNWWl
rzKs1/OhxqZ8mpPraPzEpnISrwrMRAfw3M9C3Y1GLK9LGTQk0+q6/YkXfvKVkI8jhcQAniWr9Gam
drTA68WsK+klb4sXlhihfbpetYCs6s6jHncezmcwjDwFxhRFAuh1yt2uHgznHYo3xannWN6Nc0Dt
qYc9gjf2a5PJ2UBODXKgln3gAEZ+n8GLkm1WprULA+BEN681y/KtK+NXbIxhEyewRwi/I2upNC6m
RhH8qsqbMa5jHvdkOBypZqEW0mQ3Snylrj139MOs3hSjNP8P83V8luDpgdpym9mDWLbvbWPuMoNQ
3aJbHegU6v5auSW63EdZ2vus0jtwohlRDMmCOV2SwRf4txp09cA0jX8IuXpwDNcZcSbjPhS+8OF3
w7iOpw486e6JvOGqB34+bZChhX852oVYrpEf8qV5zPKIq6N1K9h1zgtDpSq9q/DY0wJm1Lh72f8O
l19H8MwML+uXZl1gy2NLPcEo7FP5MdYnCbjP6QlMdf8EOebaMKTVg4ds7PTxFbyxGONbrbgC6jjX
T79rsRSX9ULK73Mj7RJOxsw9hHosUirH+xzKfgI85MNuixVHphmR9jQWvWRiBizpSJ47Pl+1zrQA
xb2lBsV7eAifcPtIEWFJblp5h9Q/dPHCrBxu8p3ynzGCD5nTOGWpHGyx2+/aKg012X6RImeCeacH
D/Emrqw7e0wdcegn/4mchq2X5Y/qIqhl1Q3qVe9+LuRILZbj73B7Avt2+a8PTRHpqrcVexobkCKv
4KjojSAFFzNmP5WyLgqoUpsiFrtCEH3+mMgezEn+9wRWEWp25lZ9Txupgj7oj7HwIXffr+DuFxvR
YsBakVYVQJ8RoRHdsShwT8gFNig5emZqc+rWWoJ4lqnYLal5xdEfDOKNpUhsaGSdidXIaMOUrq6i
WxcojAQ4P3I1WbSrmt3NqoXUsOLiyBQ7cH0Dfrmvlcju1i24JxcqzSbrZB1U4SozbwqFSh5+Gyq6
gE1JMk9JdyDaaUTIS7POHupZ7ZTkH47N2vjJTMLZYyzrV8SB4TaPFlDMO/sqV57FHTZctdxrCBG0
wwIO8kVJCmgtynhzU4GnPGALciqCwaVbRIZ87nQ5jv29SZqqZWdShKrfAAD0yJfQZoadjT8QTMtz
+80NzsXrcKYbQCi0nzpl9TaNBJ6TlQiKVPzC0A7z9fFhon/tWS4gGtWlt5M0uatVabLORloYGd/U
kAxa+YgVUxeMtP3fUvOwloWWpj4Asy0vLS4MmoHCIQK/kbTbtmvIQyt5gQmnmm1dS0R4uz5myRa8
P0K1j+M64vul8ibKIUH7C/Lv0f+RwvaYUgG6WNNhvQZfNlKWYKk6jyV7gDNCFh79/qiHLympIEXe
6OanAE+dx+ldvnNVQ4fxMX9PoZtFo5+R6mBMQpoSprtzJidAGZTaIo0mX4bpS82oOXqjQ19vIk+G
Q74JiyQc1ea+T+cgwqA2AQQxVrdMXch8GQnP+tN6dzrlUKs0kGHGPt6HJRoZw5rUxHsL5sJzQjF6
fhDW97ShY0MmCAQUkuQ/22H5htKBwbNeE8999s/FEbJjz7j1fdqN9YYSNxQcF+1rE6PXsqu16jbk
gXd2i+WtQlfzx2BFnwejzm+eMkBNYMiIeG/oAHr0eMLd5ljNeY8nVGTeOfZTPlVe/8mfrwhLxkTq
wKPWr9n8FJtzi/qEZuzSRSyi5fRfZz3gGyJaByLgwqZ8o1wumlTbnISX4OLq1vty1rCdmbFILxJA
93BgJJmgU32LywWOzPCwapr7zQc/iBizOuEIjBmydZWQEA7LgRvImvrBndtYwMV/gnRFiw6FLY50
jpcktprdqc8SDYISYQMmTq5mu49Pon8HyMOBMx17Q/0uglkWIC+xBrgxLP+Y+z9UCsMXsLblThA1
bmwK6VZ47iPqKugrEiWBViZsr0oOuZgYfjFH5zJPVBqRxyN/qiExh4oB7dmGDGpuOeOw57oWF7Zc
YjZ36UNBrIlqGJ+gECZFLrFeWOVg6XBtWFIPtwvrdfuiorGFCI6AhkOSEQhQ/l4i02zB3uRcOIBz
4FwFuMeRMTp5szBqQYxLhBWOKYheAYafkTqwthNz+uLRL/cYDHoFpa8vSbv0QSYyb5U08fJ3/OAQ
fgDw87wI9N8JszOBKeRxg6NbIdZfz3SyrjyEfGRvoRG5ih07jWiVQcx7eiCFBvAzzuxbHouxKeif
QPhd74XVxIbXxmYv5ianogVepQxPjylRx27aTqHVb7orsqQBAN+9gQp2MJJBuxW8X22U4akUqJIE
IGmWy+f/4m5BLufF4eJJvtxp12p8BxZbf5NDmS+B0JKlx6/PnmJp0LKdfRRy5jKCM0oWWzne1Cjc
TB7JXsEDyWdk6J8ASgq3ETMu3TSltjRY8tBKcAVOPahdgG5nQNui9uUwI5Z+td3Wzlm+QEQfgGBk
RH2cG6DjNdBqP1JMU2wVpf82y5jTVqz17wuIXvSYFhM8Rq4VIGMroyjwTCD74fF757wW5B9bQqm3
7/sAZUXCtgRGoaWjzON0jS11mxkFcPlOxyHlpVkw4p69Ae7pMVPA9B8/euNB2onzGAnqVpEm/gFp
oA5PyX74tR8rZ2UKwGKxY2YcfkJVABAgk2qXYbwJkDKUQSJK7uEF3SQsi1/EmqZibPtEDZ+OJHYP
PNAcwj/bu5p2xRWUErfA01rIYC0I+srOomAIo9KuUFMi+TqrVvXLFg9Ia2J5KzCHgfb/O5mfePeQ
1IOQWoGKxw8FZHXYDkr4YPsMSnTgdNCcBUs1b3bs+GqYYCg3oSp7EWG1f+urxPP0QeuEeP70Cx2K
2bipAnKmubscpKGIQOFACAzzsxEPE4F9dFf0bQU6JVlbfpqae3LkBgHYb0oJk47imW5bz7Ax8PKh
L+JoG1KJWQOFNQUQhTA/4TSKAufQJ5ozZmuNy25xH+RcnQwtlLtTflNz7Xb6ow4iKXfNZuxe5HSQ
UWSO4DJOgBZjNA4uEmRqpGzb9uSDyOjuZTHzm3Q9pNHWFgjetUxs2EaKzy2EhrwlOC+qVWgx5jpz
xVIASFlkOW7Z/cj2cZ3RsN0/Srvikyv9k1FnPPj258HGmKCVMh2ogmlUHJsFmSioAZSlOVIUB2kH
STGs63eLtDqEahYUFRdGjxSNKoNUHNNHIvZtU5zDxJWjlHuYljZo58N3r9K01kEko2frPFwHfU1r
FsbALUb7xLDBbL423kp8xNntbT6oIcElezzP6Lp7dYjj+YPpAnTfT8RtVYyvi6mX4Ygd9n3PUbvZ
aa0OfPIhf0UyLe0K9gpaKnoDpDom2uEO6d5K1XDnisbXlkjD67pDSji8AoCVvV0xsb0mNum+ZXBc
VA4Ubwhe+NO5UQBRy1Q1m6mgkzKepfZTwKT2fA/9+3Tl5UUoGRIzPwdDjDZ9iHQhjLe3ssce6iML
aUsJFQSGblEk6Ao/V89MxFnh7knhvBztXcw93ZbpfqQ7sjfr6Tmd4LVSIWwDJS6UVNwR5GcxRGue
4Gv6r5U23QqdHgP4xgDqAWzZvsmAXx16pYJK3+aWDdkQwUvfQo1Zi3adm0k6xn6j/rdKo3LU8ycZ
8Opo+x2MMd1n3BXnjN2zi1PSMgxNse44RYLfwR0Xlrvebvg7E5GKE8qWUhnTkMUehzRx1Nq6PQmh
qgK41H7nIcn5h2t2EKmZGjRn2X2XLhPynINpzxPej4lkIjylKwyiM4EYmw4lLF2pTzjApbQ8Vh1D
YJTcJDgRItpm+HhVRgRbwEjOmSQihcTlgiNVMXD1AklmUGOj3LT1u+r/MQPZg7pofoD5n+V70ae5
4TJVVSBbgyY/5uZAKCjJWZCsp0hCQL9NTOBQNFHJ20k3dPg4JxzXD12Fgf3US3xBepI36ZnBjF7W
4TFyXkN7q1uJBaW9+9xg8wVxVgsAZhmCpZ7XzMwjLrUY9losSmgPo0bbxrr+oWBxlhpOz9xPFEox
BLnkhy9kLDYYfM9tCT51NN0tiSrNh8sFrjK2lichX5mW7kMyHP2aweuaXKasRAFS3EbaidmSXL1c
oc//MZGhbVKiz/ycSuqiW4fy7zK7LDx0yZQB2WwKC/HXa/T/IXCrgUF1abodvFShG//Z55PnWq2u
7hgHDpncgTKweulpYrgmwWoY/D+0MLbtmHrbrN4XA0FWH6TL2+4aj/FOJddHE8D9jkFulL/6yl3s
EWpFipEOqgjJv3nQSPGSxDhNzhuF1wxOkbJyN2S7TZy07ryCw5D4825wiMwCkMraQdl8fcxg7QjM
/q5zVn7sDvrnCHiI2yiOLn3aMErmYW+ZiAbVUcLms6eVwD2UkIe65HBUJsoAec+jiilc+GXwq9Z0
K20qAeP3aSBmxnWSkmGskJ04kBPFfFggd0SuInJH/o4QPL52eFgADHuTOzZytgRSw3Ydo9afQnPm
b0OPzHEy6RBbnA4mYvUDSCKXRzpzi4BhPo7amf4FUb5LaUuxPCFA7hrvLVLvGnC+Y85zEAks7xyR
eE00AcY2KA4PBO3njWqEURgJBISEuyMlkLbolUdk2+eM3qaSaivDMChJN6jp4mrzayig5mNdIAUk
7sqKzPiZCntoXazWid0xufr22rslh62U1o02x/2S+3L4Wzm4CNCQ4vpbF88R8BgZZ4coXs4qcr6y
QcU7g5PLEwKLfcbnR9bzY8Z0GTI/JUIdYUrd4pNE8F/QdUqqpyULVAeDFjLHNcn+DUG3errwYNiv
e71lJzWuz7yqKTJgT0DpdRDcwzlzvlkld1/M7IaDWrBVKhBKBNM1f0tNW/BInSY6kCkXETjCEw3d
Z/MoE6/wApqRpLJ1ZyZseXi8TaBwr2aq10+YRLInkMqfdtHANdpXCt+6QIsNre8FYNM6NLNfwiXY
AdJ5GuQKYvvrsjANrNrO1dzK5x4vmjPcp6bGAnUP4KCj2VuLlC6S/JRZK+l0ur8gPSJdrU51ZLFl
Y4HhxkmE4lxrR6duwsEx2QNNsx181QPVpxGby06P5X8O6DEmo1izg/L7FsMvJ5Q6ke6ApEjnr9X7
+VLuKu3euv1vfeC+p07DN1I3zwivhxsw7roDQ0S3i+pX6rRDBG2vhNMPsPY8niNd1odQtB3xre43
wifwsFqq2KRL2ZzqvL9L7HX1zq2tXTHDrHm0YvRIcpoQwON0SCh83IEFuuxYTTIgr5kRPryjsC45
OCpR8vyB8HT8SEF1dEIVsvHzBX4XgVz28USwyKR7c8PLE86V0JhlxekOQZkgEGUYg0SudozgzVaU
6ohxO0rHttDq93tUnTEsowxaQGtzyGf+DKwaqeO5zI5tW97Y1tZ+i3e9gxNN26NuIeY4sfdDZw7e
J4RRTZRm527FhRexXIeoni/DaBVV0fZ8KpD6n7JVXPnMTeffIGJacdssR1tsO4aF/gjV2TE7cujW
Fg5eeaK40wSFHQGwFI4gmwHQUwYYxiBjaYy/osCmX3XDpAivOAesvdur8NXvI8YtAmSXvYvlzdct
EJv+oaHpQav31Vs+pOxH4rOMXQHxT6F5Zv7ZjZ3giH5nnHcprxvVt5a0IboamI9OyxDikscXcElI
GYfZdLr8xRnO0lOw8QJ5ETXxxqjG9uqyUE4u8iC7KGN2016+O4smk6+BHcGH5PV2z7X3JaUk1mc2
RaURh3LZgfMwinNM3umDfir1UAB1JMlEAHVXJO9AbZNU5ql07aV3lCzyLQCVigXRj/ImoDfHMCBg
iZT1MF/KCUv6S4g4dpWXwbo2VKxZ4aqs25GyFoWV+UerzPJWkOmwsbPCGATz15POeR5yA5zYQ5wx
mEpbhC5SQbqdVfQGo2LkYXHm7Atm0BD7ncCJj2VQJhwHj9x2Fe9nTPdXjNfRnX6YqBaHwjqNqVWE
NlUkumsmSSgxKcLnMVG4pfn1nubp67o6jfiIAJbDmfKCMqN+byT9Zv7YjzmgedtfVlF5LMHmJlvV
SEQ7PjtjIrSKY9TFxAV6gfDtzSR0DHF5Ktr6iS1u8LXbN9FeUBCEfINdAB4urwz/YHmlbvsqOBsM
+oGHHpVB8/aWiBf4aLgqIeyeVKIXOL7ocP671Mj2l5fU9xI057EYeAaD6XnDmsq2tJyMMwG2LGMW
gFX64XXDpQp3jLoOi7sq7cQuMru53CriXNGOHSedHU5ampQGIcrL+DozL1gp2DMuqWdmb4UcsfWJ
iDYvmT058Aa4px3hv6sv/frY7rJLPyUHqDNyEVOgKtGhdvApD6hlfmaiBdniPRhEqJXNGxm4szdS
xJnwAkWXThU08vlzU0ISlXPSVRcl232UR0tQE/x5BUYnS3LK78JXBsn0TWa+RHJgWmliEj8Z6Z6D
TPmzMnCJYbJV1ypyaZrhyKfQhHBiyQ3AH98yiP2GUX9mQDNcdd0JGvyfPJkB2cugkh0Dg2Y0YlBk
cTyCNmJxeCvVqn5TeIT139jI3wdJDj0SkA5DToUjPaUoql+VeI+d6NdHmjNzVCQpyN4UnzWssOkq
p9gaBDw4rlGiEr4iqp9mMpbLPi9vk32FltPDeYtHBROLm9uTn3LKYKBnOQvEPL9eR/RUpU/buggC
GCoHWdcEGld+9ynOE19KIw4BIX8Q/wuDYbyoU7gDu9Sl1c8kJ7JxlPkqzmUK1xtqKNqq0sPJA1wf
W0l+SMn6FhhmLQyn9ne6B1oGBDSaxgS8Oe5l5G3wkFVxXSZ2N8sEIvzoZxrOq9xdnjKydzVbzGpS
5TecF4QnVrz6l6iTnpfgl+LmI7QEseOnLVfrScAdPaVs4h9B3wBpnyS/Aogm+Y7mUNUTD0rrqI34
evqC7uKVhn10CA77e17Q5Ptjf+LCJebaO33GzJs82sMRtVNJz4EtRw8HOWohtvCzV206Ye12DPtk
NslC1sNQLf7hZd3DD4MaGCDABcrPWgBIgo5POqsKpV5ZC6c6ldxifOVIMFC6ItKfN005A1SlUWQr
YhWILD1smBPafcfI8xpmo3FeS9cpJqo4jXbo+oySATXe6G8QB9ipSaWBA/ns5KE8S7sPEQi93sz3
zojYkF8yRb/hZ4/s5hXQD0VpwT1KPjuY5KkvqvWzrwYaLyLFfEtWT8ongF1UevLTwy6fPweQMaeU
DOrTBbBhnuNLAaHuBYjNTTJUNUhuQ7brEvXabs6YHjyuWod6axk3imqzlL7hXH64/uxq5sjsXRgW
z3ZEOEZ4UcIwsAfTTFqKjO4PZZUWDJZPaEknxWm3PA4hbfZVlNsnNU3FR2/3ZOaAFmGiPy+ga5ya
PMHEy8zhSN5Orifw7B+oCHbZPiLu8TpQ+J6QYCuCybR8aFIYuTm2+ZdCRqw18Cwh7HjgT2BWfAks
x35UE3+tPsbILHmoE6vP9whaSQCnczpsM9ViCOhGF7e5keqDW2/sX3XXlGi2l2K68WIJOxIVV1mw
iy9tvaYh+SUz0weetqQJrABtDBtYYH3xC/01dn28U4onZGxdwOD2IbRu1MR3PfOASrunfjnOyI30
+DqlaJpIwFJA+LF+jVsj5OmThLsftSerHe456oK6XdAO2ECiJLRuBuw2tRYH8SKUqe7qi+XNC1Lu
XgzGQZUW50qpHWZQA63DJSjUhtss2hJuo6ScybLHU2c9jK66innE/X+eOTJwZsVK+Ge3bhD/K7qg
hBQyUAPzfwZgQ+n/hFkH/9FBlamjcvgWP0R3EQbHpd4oNtCPOOsZq5Onkouk6jNX5wMtAEt3ZrYM
NU02YQ/8K6TrjP7netU+/pGlBaoR89V0AoCsrFRm4dwYOiBwe2FOAMX0HKtSzXNTqfsLBYY7zA+e
pY2e60iy8ogskNL6/W3ghG3L3SFJgvj29TYSVlxFQ3LprDgqqn/2ev92YFcVrmk37KBW0Gio1ZgK
kC7fcGb8j6DXcCc5VWHxo2MFGvT6lQCiU55JMr0hEIC2rQjB6sNMZEL49PtrQyJ8YF0FDZHMQg9f
u0GQW8yPUks1fkav59EVMN2aDPfP7Ipc3DV8i8B4Ua84H5U+v6i7cYKa9JTasVm6nnqKL22BTNgk
dsQlblh9u49L99AU9LjDOmU3EWhXXAwTot3JTC1TDGLZn+s+v2CxFXvtnouUwiITCS3l4mKQbm9M
epZWJ+ybSkJ45bfwWFND6XZMp+JRZbB/EU3/umfAY3Ep8IiN1Iq3SEV3CvqEQsC9R4W1ovcIuhfU
P2oDknOhqlYMgxgIOBGbT6R03NJNSj3SfkcPWLr/kc3dJrEP4T7q5tDcxCGM9UmNKRlH+8sHYn6B
RkIaUYlKGfRqfhhj0cIX7fsjmk8aQg6V//wd5gc2soISVi2oQ/yv+4qlHAiUyIAwtRLBiGCsVWFl
iYIj8WwjmylCmEu6+ICausikwyU7cWIwpXRM/WMAJa5nB8ffbhjfvmMjoMhxCb0/9hrQDQwOmpxH
oZj78mJ5LRbu6SbCWq8D0laGpMn0B9a6X25Pay8ITMS2/tPclu5SgmYsaaDhNrqBCnGmb+S1vOfZ
qAtu1oioL64+cAgHOgQl7Qfk+zlGum718A1D1kJMmZJoq7hSKL4AJeEqsi9iogz37tF0JfHuYp6i
NOrSac0mW04rzblKp2HxcDiP4nPkG6NoJH8jjysrVxgyEeC1r3vJWr7Si7STSSt35el2pqQ7F7/Y
8Ktvk/YcHnoy5s9LBLT7DwXYjAxDy5yYDcCri6Qra8g5jnD7en9xn7xHvk74DQ8clB9KV4mYlxtA
R5LeU7r0n0kUTFgNq/SsEAfWAGbvekmUG15xhYZlyA/KuwgCdECoF0mz8515itza1RpdV0vvmqbL
LlBeKo83raAIH/aUNu5NYO+EZk/1ffCTjSC7Qe+rmolBUoAoJVfZBcF6FaELNS+30ErPlUUQO8Xt
WgeebH9UIXjYCIoUgdtwjtQK7Idof4/oOprjGlMhBTHEojmcSMtIcN9IeUrblhJTxTUYU+sKz+jY
JCVVMQFv6RU2xarQvaH+74e6WPBNTQzmk74HOwDI/XzT7AQAulKRMTiEY8Jr7+aJoNiPqRtdJdJG
UjlrsnQqcX20hDPAdYZypk0cmFRsWfs5DdR+fo7L0KRWrBvYc0vCxtGf1SESSrpx3UbYn3mXPojO
ObPmvA8iFgVHM/ta0MqpC1Ahv4Up+Cdz5m4yXoZkPOPwpD+u8gLvwQMdUNYsfO0mvQNdVSJ0KLd2
YS5miLR6y5vv4b1IOVqNFCN8eb3P6fLEEE/oQJPRLuFmCWBIRzLYcdnARwKqI4S2Fyzp567Htqtb
xFMXSKJjPNBRgty8iHRyADPkncvcgt+WX2remVK7fnH1Riqq3S4zsbH5dp4Z2Lo2VEXH0SEzBkCy
G3TrhuGIy6W5Dp8BB9bhtrmc1ePKwzq1sdUWQcuYrbKcyMpcwz5Jw3qIrAXAAjPJzbc9Ky1XVzOQ
ys9+uzsto+mAzN5u4RFzxWm/Wf7m5vIVdb4kgHj2/Re4vfr0Bf2R3c1qzC5Cxpol09Q0HZSActZN
YDEOsERxgFWAmDmEWKvKHfRDgnk2cpycKPGg7IBzYvGcUwv5oVI5nukw1w/5s3+HftBK3I/PHI16
ADiyPEwJZClOp1AnuHhKVYX6vdxlV8QhvtJ6ohg9+7dHgcTMZRcrKrj5jpvoKgV4o+aKhOM8vj/d
7IzehBvorc8k12SMtMLrHgGy8Ae78uMGPbE0whXcxB5LO6tZK2fy2LiOBnEZ8Hmr1GXB+5nmCBjc
WYZsv1pMX3HqfkFJoL99JNZNU1MCza1JXmMuOPoKUhKeZgLWZHkYS9uDchYdETjoDANYvFZgj0YL
YXxLPNNthCephXuZRA1Y4+N1KCrJvMbgR88NLF5eF6frVWnLtFtZ1V6Ti/AJeJ5ggj938lG3kgHm
rIo5uQAZo8dXeMKLxLALTTYUEyVJu0+Jm7K91bExr8rtuyJWKIQ9oMwklC+z/26MDIw6XKOyTyMy
3PAOX87ggdYhyvR2YQoofZtaj3rnIUU1ywPTvn9nAB9Xh4SqNod8NuLVRKLzA4oFE6JAb5ukO6hQ
U6wFLyRhl7e0sPRz7z4QaoYNwjDWSoHbUd8pIhNC7DKxxwOUPhn6X7rwmAHeCW/ChtfqUDVqxp5O
pijRqQP02wRjHIjChc8NXdScAQRXVdR9zBUhwdrT+pGDq7Bhfw6cctYuYOSCV4tbBp0kdu4vj1px
LO/4Sk1gzOjipdssgaY3zo+0sB9R+SWP4ES+yN8w15xEakyD0IBvg8Fo1IYh8rDMqosTrJH1HWFF
s50qrHv9+GzwUxboPM1FWF5x0GymLWyywSwlxJY/4gPf+odegI2nUeT697wIYBmeuz3R/3L0X8VX
4bLrP99+bT2VGnRDae0f2+5QbqYd/c3vsU7208iw1wfHCVsp4zsLKcTD9avd15zwq660AkXikLx9
+8f6BPNeGj/TYqmC6E79xDtN5v9OvXcO0NQnN/f6QP10Qk5i4HYxg7ZyMk75Y+KVW6WtqeJeZmPw
BBujSbVc6bLL7q3HQ01fYD7hGe29iA7uWSEBbnHl6XaTQjxfaVGpcm56Zl6xCTBEZq2w0OJyGR3L
Ee1UTUbiOUYFClDewCOWStydxgfc4d8Idv66UhE7+jc3DHh6zrLwCtrPhuIeEFEqh7Wwizc5aZPU
W4gebWiGjH7LEi76pjlmF7Ug/k7PqMaFaV1eKXEMctVwxYqcFq0dFk4Vg41vGpft1qKxkZUAVSMZ
qDDoVZl85ncP1lPQ583krj6wF2FaxhogvanSjcjx07BF+aSuFcow9QUTR0gJj79Gw4nHDJqMlbiS
T+d2BK/dZC7ysHGFGg5DjU6ojKibop6br6LN54aFcR41jyQLPHpjVZfuLaUMqP9wA9CiaGKzuDiM
k0F7pcMSQxOGLf6yoREzYMCmAHFqLJGAX9p6TG7CS4W/3euULmc3vQHGfgK9DrLXjf8AILYYf92W
Um+e/C4SCk0KI44KwYKhJWfQgp/4sFDrakxKPwG2Xwk3Ycnd/uQ/K8bAYgAbIs/XBIlH6M+j188V
/yqtUQUZJS9ZDJlDquoFgdL1hLZrwA4kQkcGy6JmdVsiZKxvtjDmFsOuDQ/JRLZ3H6hSD4BsgvqV
EzhdDz7yDZ3ewL/M3Q3r85KzdcHmyCwHWkHxdtRFx7YWGD8HhI0ZS/DfvWqIXq0C/emEG1+XTq25
BnNiQ6yXH6MNxQW8EnXsj9IyTs3nWUtceI+cUQl+6T6KUghKvTKd82VIHeUqUvmkJgej/BTqYp0b
zTtMrNCFHd0yYVVUIbR7m/gnBbysrAMTSRpQ67GRENyoTWelqqqkjs+tswUQZLlwD6FRaZs5Njif
S5PMdPpbfBOqA6JLYJ/klLKnZoOcIxekfuauGZ3MLmwQ9hQYxbqmSziC162zW/rnzbwT+M+totMb
ZQXZNrIy5Ahx+CO8ji3YsywbpmJJ+jiJL7Kdff93xHhOwk0wO2Wzc3+2uUGnKiZZXZP2vVBDk+po
EuiPiYoIwTjEJfdguCo3Hzb7QOZ6ft/IZGsU8rv+bEqaJlss7qBhkmx5Z4JMllI7xzC7moeK555m
WdZ5dSQTRxye7yETpExE/QZQj4JT446Io6tuJSerFId03uofKJNDtHE2Sz7+f+2PunFTICfQZzYD
XuZubs99GTWDySjS76G5x+ROjnob6TElF8xoVDhwL5Bgg0MG8/SuOE2N9lX9BCpVcuooEiNjMpEb
ZmFxMv52sBn3vkYWs54UphiV4NG9TbGSeQl7Hx1XzYcDFki4fIzZS9xTBYQlAKEDmsO7u6ffS+Q7
l9NZBSPP8sBHAUKWuQi50E/Foafbni3dbmvYDIZiURhnHCXqPdNVvFXlGptyxT0etOONRSv/h/sJ
fyjgYMzOp7EePN3TrrH4leBzIhC0h3DOd6+K4/vLIN9pzbD8J68PnPhCdL4/lF/OQXBwM5rq7IDc
NWbCeQTSUGlQTeWIlArnLzRF15tWnbF+idcw8WRhalyjBL/Y4n0jHN7jFHRp1+SdRe67t5wymRZV
Jl55whROYut5HEyRyPEguMGdaHv3GkjjybKce/KqCfumD4aySPKBE2/8H3xO3y3Wh/RDhy5mURJu
HFL9ql/AjBh88J2o+RFf7AdQhAy3LuDVbTD6KmMZl0QK0e/o4Oa+n7qA2aT/+VMpS/IQpvrGyNi2
m4iCCRJYs0vjfWxeaJhIZxlX+exMwHmy2/df+6Wplg3QGXy0VbBLz8TGdes8TU/7QBHp+PpEA9E7
naRaDZ0PwOBIDBCw96j7ISuTxbPR8d/U7BL/kHkGQa5lEEgGOClj4D/a/W/fV/AAc598YyyjkbwL
HRkE1U3hNNS8nVq5Sm3Fv4zsKzvMhvV7k4o3q7SjqEWBneIKpDgKLEfeqEhnH/8mzJPrZgr8oG5h
OtcP9osqEixqBiRjShBrXZ3B0juOrCUzLn7VrgcQ5kg3hcyW4Wn7CCwGvE8WeIMGLGV0qjEJw8/p
Eyf5USTI0qenO3vAk4Vl37Vce1R0PK+GPkwIM8DfYYif5CWiPCofrjbPVwiFGn60AvaC11uuEcUX
dKNvRutTbbue7Kk3HrP0Z9mFYA8PqwWFrK6aSKqWyfX+lhv70K1H/awDRyHsCOKOVidjVUxsRUwD
kTBdnvU7ccuTUS7aOXYnzCVZrItRPv9wvQxw3UaKtx7mhNjq1r4gmtUzLucVJGJQYCkM/pvUBtjq
tnn5q1b6WtmXyZ2t27ZGTAFO9D95mzHd6r90NI0HEuAnm/5OZt9oRT7T+XEO5N9Ca9sc5Q2P4FE2
IW2twuon4KJ9gOnp44+riGgr6N8WbV2+yl7A0uXUS5daEGWo7KbnHvW1Q3cOdaPMOM1CQ81mHcze
pfv/fIM27qRYsH1CC3Z2K+bnHOSwCC6cSGmeA4yVcZbN+PRKPSEEKrbFwhDytF5YZadoqxDhQvm6
0migCrO44R71RqPsS/UrNSUFXoZx4NcO5bcwYkgeZft6BlKmvNYnEvCgYHFKEWwDVBrCHTZ2aJW9
FKkBJWE1VpXKGIR/EjTjpaeRZ0QAirld6UHIf2Kpvb5OPJ3OwGnRzUHdck6lwa0lD9/iYrmgvyCm
rgnBneCFWpnIuSH0EJkV7AZmmufoi7VBnY7A1UDdxJ8sgKr1jI1vEQ0Yzs+2w915+VNwT+UQtiTZ
P+Z+u9PMAPLIKkGUqfNol7Bm/XthyCoYwEm+ssp/9X2JksMN4hwKlGnrBJLl9AJgobBN4NieNV2R
vtNmDQMmy9gy7BTk+k72FQvnkIIYoikcEZwNoWDPbtczc7IgB5FT6IqPlzpwKwrcV3RO+ydppsQR
SC/1KlWmFy/1pkn8lxA+LA7ONBRuj5VuHK17B2HuFqF47H0kWmXebwXVNIssTRaZZUwerFIBMRKx
rFqfu21+vS8xt+uJLa+1drZG55B3R9GhzOHv/SqhN8Fosd5jtoEVwyzYSIBUFJFh6jm4A39q2xTb
ESu4V/zeSeOaqv+AOvtmeLPMR8n0hhDx9JK5RBwCNISmSa1erPIsh7QDW2eQjN/9i+0kXWWujPCR
8powuNK3JU6Hke+ngnXA8wMEKgAs+5dGsYzc05EdIs2e8w7RrRuF7mZN6asseFT7Ea/6qcfUpr0z
2Ba8jH116oo7AjHlR9n5opQSZh+KoHcG8vvCqdwSYYkGTDOcGmSJ1+hYl7MuOyG92zWr4csEqvsk
wT5/10Qc7B/OmtZuen/mF+AuU9q+W2HzM+IShmErakiUeJbrmiJLYlPaqH4H7CQcNyawxhoH8ytU
VzUfQlAXOf1a5zxTO09c3r/XoV3IjmeecFi+u1/rY0khnFKFWyJ9FEGqfdTvRyhZ0fxezdpdrmsk
JO/1EKxPe7tK62czfK99Yh7R2nwdZPOlg+PrAskTPkjReI7PCJ2aQlwb3aFUNBOCKYzOM30RuQgC
hEhO/xYSaZMY2fpNbDzT8n1qvLAttgAJ1SIazhInszTeEupDetOe0/frZmjIWdojM38/uTpuIXsz
d47Tb6Qnmt5IzNaef5GMNKsFSzBEsLPJQanpUmcVLEd9Hh74vk3TAA2hNyLJbMFyj6A+sNywtY0R
hjR1xTlZbdt2pEKAbyRxQA2OHXhiN43f7RUYWB38So1eQMahrLCTKMh4V8M1ltGfuQcz9u4gqkmv
CnlmvYjblOSkIm2LLCmH62hNVw+3g+AxZEZqTNP3+s/hIxvnOow/oMEFA/QxICiC+JHem3XmBuuO
d0Cmu1c6wvPsnKHhBka4S3dqn5ZBrrzoOpizCIqnvoZtcPvBK4KTx6+g3+A/V2scP4OWjXWD5hax
iz3VrjRe60oDKMyrvQkMMMjgL+M181BqFiqmgRI4PuYAzPXcLVQcOZRWnxde4bAOL+zjFUTkRVlV
uV3m9Z++Eh/d7D26wSUwuWzVdkYSDZ87aIpol8b2Dk7WTCEEpO67WO/h42Lf6yVvJ2dE92KQn1kM
a363WqjhLFDR3NgINFJWXU1BoaJ3w5z9kDMCZB7JVazfrF+COEQOXg9mSVAiLcIXEDLcOXzONIXb
zWcYtgUgMRgaZWHof7XkpMvvMNv7H8i7wDYRktEG4wm2tfYs6YYWINyKJVcLp/yux8eHmcBtqNTT
8gj8/X/YZRoDSnEe55T26GmC2okkV2UgzgxRmytoISr9iqZuBpuVXYjMULR/0PpsqoFt9F/+cfTm
UXpWddkv+HinhFLdXdndpWgNd51U56ydoI1bWMpyTn75nMlFUEgMiInFOY/eeRkG1jMbyiwTXGI+
uc+qFs643ZGrlaeoKyT1I3g+NDtGQ+sbQD/Y5UX9emzgVU15HOThIp4T9jm5sExLNCtHdcwC8Rom
Y8fB9cUrYB7fxMNhqf4kcq0pEyLJ6trLk6XlLuh6a9FXwVxBeI735E0yiUmjOwsKnLRMhHOIcEk7
d2ztfgPApIr/nfSIm1zd1MqXNdid9Ih9G0vHb1zOB9X8JFWlxmJ2AEMZLAJa/3WGEPyEFgo+QQxT
DPjA3FzN/uGtMRMZr1a0BP99y9jWglOUF0COdmK9hKxMHsJdlC0AbQfQ9QBx/8aR1BC33nFDzLGD
wYHowNaLYSsvdSYlpnc1QD076kx5VqdcJHGXPqfgHiq3wiTrgX94TMOoqmmJRFMuXFiM+Pdm9MNu
L9d8fnxxnJGAP8suQ+8X/73xMmOkPLvS0retAmp7uRtRCE+Kl81qsGbhOH3a7Ne1cWBOPXHGSzli
hq3tstlGgBHor+4i9zki9OXMbmyxKmKd0g9V9TBey+CDKXdjEsOnYOEy1xyvk8bUrfLcKijlIdP/
3Exd0+6hVJGSE1Utd5LrnmG/db+YHkAxXuUeSzZslREHX4XWqWhkfPUK4RXerOkAzjlWBFl9qhVF
T9AbXy4WEMegfqYDn5qUrY9jwMDIS4c9ddEFP828JXXXU4Pu+Pf8tMxEgSZMoJSvTEE9/2QoaJ8K
a5hmXlTAS8ritQgugb8+8+sylJvjsg3XFYoaWWsGcbhUYNRNAk+nczzpqeCxuPdEp0CfhhL9434e
iRVxUlYWsygIZcwhbExoS8umHGt40wVyrocbU1kmLNRmB/T2AlowpYmJaDisMt2KXEAOGR48JMRE
of132onrzjpm9ZitKL6v5mb2KR3XTLd2VI0M7jW3ZAFz0e3cXv6lHDGCcNAoXzEGHVUaH+uxCbNR
7LfRo8FNb395ZK96Weflbx/zCbJGIvQ0Z1YqGvRUjPdE65f8HrJKrBNk9RLNWrBrAm403HbfZbsO
nxLqllKxr53tnllBxsA3xGmPSgGyMFTt+NX26Bl1aZYCq8qYRXcoFDNG0n5xDpfvR8OWYexiZZ+3
NLBCZIwsJijZYKyg45TVZrove71a/gn2sjLUzbe3zbwl0lAf2xkBwnal5Lr7xDDeaIiRSQCV8YXo
AB78f6NCGPtAGBlf0k90o6xj9TiBB7EbZYvo5gNS2IhWvV7BSpYwpW5XQmP/BSMMEvUWk/7HuUND
pC87lg5JHV4jFLj6BPA4Qavrs55Uk1mSWEwVz2DwWQMknp55S4dir2R51j4yOSDr2IphgxVh+GOU
P2qJtsdWzaPzYzfTemQluDleEEg9v59UJrF08RyPQ/p2jebr5z1OZY+KkhbMd2ooXl9Il/f3vhYB
J8RRlZa2U5XTIM1ku0rC5GmqhQ+KNCSSXtpl/zpiXWfWeK1ZaFsUKBbqGXrsSgDuOoW8gnOq3c+W
zYxI/HJnjyOKehALQcrOtZIIA4RYFHMINBcqiEYCLCH9SJQ3DxgLy+PfWj78+lPKCTwP20Dr46GA
t7R8nHpGO+poY4UHdJIlclD4JC7BJscykht15vi8uIr8g6R24x6w/ajvyv3N4/26oVbD+4TY+rr2
PnwY1wiU5ZojkineDv9M8Og/XJ0qey0ab02krToXUykQ7hIi3LL9rILrvb+tMkXsQxBHAYBns/2C
g98T711+sC8G1JLheQGKCpFTSnLRq162VptgQGDxsl+vAxqgk/E9ZxqrDSZhOILnBv0ohmRRAUtT
Z1KmE+dt3LVnL3GuZEV+jE1+IZdyTAeROZzNPDbQJY97bNKME+5n1ZdwqQF+79ew3D0aPzhWi2Vs
ZfnJ8CtRR7L49OkcbbUwpAcoHb4/CjdHvpoWQ+jV+GFeeZeyt1lpncvZoqx6JRA6QhnGC0M3gduC
IAu0DAQ6nCUCrzHkPBf+dfd+BuK5V2REzeZUJo84YOJGtiSvHV/cmYzlSaSG6A3zoShhUkKKMMZp
TAHiVBHYys5sLAMkrRfA3FFl32Ql16UDVaE8KyBk6QoSseV/r85GH56uprBIFM2quki9C8pB+i66
xXcDeoqZ7IF6IfGOv3KnMth9UNcg2B+lsHuXXYqFn0bQTov5yxsl1E7Xz4zL3RDHRBz1EgnbhGqC
aqSx1VjFY5BNEXSpWAUIl4tA8rFwv/6pYdROQ+NX9ZwT/nTFBBoG9aTaSuBSDIepcpP3FrUL8ZpK
BhIeA10RUQmAAhtfkUv/JAoUuUkPClvLn3dexX41NzIV5PqywdvfRS978gO0LFTQ+4h/sHroS25g
IhChhJdJZWIahnU6AMr53o9EHnkIwlWtUGmaFJW5XL8bbA3AeCLzIqY+t+vItBxzjEDnyIsWr7YF
92IOoQLPHEsrzEvTHLiKPbk56dKqudELUHW9WfGosmdSW9sSG54z2a9ap6mhbemTexYIZEiHW8AC
wwUttCDw0GBbbxBHGCO8v7DPcOKNpYr9Xa0C1mGYTBJmgS9jBUrAdlncmWEmyvWjgwdf/eD2r7YW
vn3/uUIWarEeykmV+zPv75+gTsjP67Noke79u5A1tok1lse9IeZhWnSzZWID9ulxozIW+9Lamrln
tBWZsEI45wIbE6nDflC4aFFW4lBIRKa66JPGz0KCEVpJD+VAbpFITp2LndOZfa1cccWoEfz18Rtf
OVmJgqFb8jBIcyPo9BM60PzvFRek/s7EIELrdyUwfOBfSLXgd1uB72c6Sc/wZ8p3QoiPPTNBJQcv
TxaqjCE2CaxrqE+Yxizl1q14qPMiiVJPS70O5EcXSk/WCGzIVnYfEU5YrYg5frXWzJmN4ewa9z0G
hsodfoGl3sKUOXdVvR7sHV+RQU7XOmqhuKSy1qeEaSRr/uS22Ox8t8ZAfT3B8k7nsI5sPjm/0SJg
LazyzrbrqDRSGq3bAgnAJ+X6gJk2UQM/Deq1O5I8AO6/1YGbMIuF62uUiUNt5qxCxT1qSiIa8sDr
ySF1jYCaKisjfphN+Ee0mzNY7e9olcUBk8FKIsm7hg75rs0vGrO5qkRsPPUEipZvMPniJ0g0U7Fu
cWNtgKaUMoz3JVbrU89FBVs8lCNhxyxxdhnz8zACQZWs6JRrTH5AUgOBuRn3lty/DKJB98xhXjRF
Ks2VTBsqOStPBTXTbcWEYS0ub8jsGhRLubXEtK0wi3AZe2kzD/Z5jIXOAXJjPAwwSZ63J9JenMGD
zXBa80dtO2XqPyagHTCrnwHvNXOBwhNzsvw9BoiMM5+kVbG73UTqCs8dMdi/Qg2S3ifrz0IzZvfU
NLJ+pjVlR8/b+L6YEaO9eirOVXPNv6IZ02wAB5+fNQu/c1wWeBz+1SS8GTk2kS4/mxtPTngkjU/j
IcklgXkEXgWnDu+cmBlp2f7009JbNEivh5c910w/OS3na7jK69eKta/tT+Sy89eOCwpTOKv2kjNu
hkYa6L85SLOA8V2seqZxhs1mceMJ0S1yqlRzX8WBDsJVUQuSltn+xyTOMI1vYMSlpZYSLaMr9yT4
rX9okDzDu6z2xBFZD+muVe3q8AC0WaEFXuV1Klf4iwy9OBn2u9qDenSdLvhLixTg0kKdFhgMT22w
0hIMhtbxdfZOq1GffO8lOAlsF8gNKsXOgaXwYgSiGN7XDl3uQrNhjcNZZ03tyOMkUmzmSsNpYG0q
1pUY0RbHBRnx9c+fvwhduEiGHnYhK+xrnJ0D9ecDoGabp6QUZNiAd/T575Exz0Qddb+UheAhlvFD
J3gSNuomrPfbne8wwO+1zyTtZmjARzYzA3QDlRgu69Wv9LWAwscea6XSoCReasF7PfAr+OZA2dOE
P8g8F6BSj5bl9Nco9ACta8wtFCoke0i5ps+WC4zeTvATC8jj1j+vOXkmJq9rvbLBCisp3D4yR7HW
z+lNiI4U8daANuIyh4nVLSbDmbzQTIrmOl8bYyCrVRWFLuXqBISW+9z5XAWfKrTVhxLqRs7gaSuk
QSnbj6dcS2wmITxWBCp8py69ChYEg/M+cIrDw5hJdwoei/3cB3aCwOGvhfigiBh6eqJxDZuo+ZRS
WryVvTd42wZuNqsPU9pYzdCbeaOi/5vwFhpRlPexVxSxGjxV2Lvd1CSviD2mEBn2te5wKo0F77YV
s7E7FY/oQULou7J3C8foqJ4lCMLq5jN/LTBnImLSagyIlFmomc/3WYge1L8ds5Yp7RBdRWAWpE+M
HjtGSUu/v8Z9Ha6iQT3erpxX0beIGShkPVydITuzkXOnCrl1egRc59rVzk2Pu3VNA2bxKTHrbsLm
c7OTx4KJtxhZqJj0uVzhNX4CWBnVg+xO4TvPUs2g5WnaymZRbcbT8H/Ujj3pWY12CD8Y4RvfUA0e
MFliYSkrdkIbbnwBSqhG5ukXGib/3NiMSzDCX8OU7eY8JABqtEMKk6pDl4CmsOyg9JBT0W9O4wSf
cZ6BOVkHzlne1hiJ9eripJ9+9EJVY31vls8Duij9uWZ9zp6woXgo/ooFoubuuf6bXAAI/bwPEZul
eeRQO5AsSNTku92A2rwj28NPRbuGguNfSwV8EnhBzjQ/2pgGUCjpx2OLUKOtQ1fJnb8jJsShUVPh
+zqN+GaXzBskji2CytqPzXd9cX/WMI8tnRvXh765TU3484Yii7APfiJz0N4RYRbBYSwKwivLJtmm
lw6Rh//anyKLzS4iO3Pzk1ZxgprAy4pasYhZaruZRDRpK0ToJ3JyKcijsYvatpU+s3WOBj9HDbHo
zgGNwjSpjQ3C+STI+GmPbOQcZPAIy0474Y9Blmc4DSODAiP7EpF5IyrnLUeHVMlJjvBmonyvpXl0
VbfqdoNY1NOw6E1DkkXyHEArdFaLqIjxWG9JcC6PKIOj52VuKIUgWOI+108zkxjedZWAwJzSYkDt
XhHdp9kDl74D+QN4ZAsOVJFJGhFvo0822NS+lpPmhu2bcBapubBmpABHvxKf5e2mF6YEtyzRaRr+
BkCGBAZmgatt2Bfxa/LYMAQKS28ZtMx/AlX9hFy/ecv2Mfis7njCslGpPN0QW/420kJxhmVA0jQF
TlJuyJdSPCOJJDQ7zJP+neZ2dfmEMkNqhfQLSihLB0p76pErMgS7qvHL1otGaCcmIhBd3jltjbRY
Zeu3arEftc5XmhK5HJPuV/TbEyfjPLt3nSON8erzNj69YwRdllyiWbNRvbKQGg0+ugyCQmMcoC1t
xe4GxaGWzdqfQaN70UIoCqw0or7Ytr/u27VzXWi+dt3W40SNLdkHbnw7lhgfzLZlxYa3lD7qNLcg
7SyUIuSup8AyTiN7bl6u5xiXfPgGJ0dF7OvA51O/0mhVhxa4kqsRIe9rmNGtNLn8c6MBBvTZUgSi
9x7HzLnlwry8kCpyoy2vn++PYUYL62iRtqA8Eovp0tEdImjMC605nGP762JMZdnvAAEtmTgLssyb
j7XWest0pZ8pNOnWO7Pz7cbw98aR3sR54EUghnh4YCPYhtitr8BYbgtOgveKMQnR2I1NdJL8yrgC
SFr+JgUx6G9qEHVCWqDYutKaKX/ZPkMi6i+Gj0TMOGEgcfWzbWBWi+Bf7EPQejQR8X13qZIhcCQy
Mf2r7/+vipCYaRCewCePHpnV7bgqcAaDkEiiPgDs3IrgE8P4hkg+T7sV204HmPRSSdou5Ct1HPR9
oWfY84R92CYbi57J6anww7pIJdTofs4BdSq+HfzHmciMkSfksZVANst42jaKKMYK0UG8EnRFMi7N
+/pb/o3wLhwpDIVCDvx452fP6JDeSFHElZdDYpsO4FVzq4Bf5AO+x9VB6E+085FSytHAyUEjHj6d
8rqCU4OgJNaj6Ccft08ugPXSnuLqfH6ey8MX+VsukIFnUj7v04qJvE5ci2mXmJ1fL88cpbyzmZZG
kommIP1I1ww7qPKC0B5FlojJJupVDn+TQXER/abGI0kxGJ7rBHwVCspaBgZdPfe/FU57gOUjSYXn
ES7G4icsCj8i2u+OSX/rg8fkR3ATCrfKumU6Wu9LP2lF8HZoQlNGDYxc0nfhiOVmLYoGDapOUT8g
CZy9iBZnHr6YI+VjDpycgbLXQYu0FhHC/+PB8wQHKJXbPzCuSPWexH+EtKHY29i43C/e+NcRyT9p
mGN0+zqEO1e9+FWzK2P3Q9OxO7Zl8HHSRkC/0MZpXb1DIIWhSH0UjFiICQT5MNkr8I0I02JMuasT
ZpR4N6O0PUX8m5smRwOJHwaUdO5PgwM2jPelUq5C9hUYz1pQp+/Ifyg5MnDRlk0Cco9cV5KOsNUK
xGJMTMMNjx5/GuCpYB2QLuILtxjwYU2ICHMEMP9jPCs04qlI+wYBNuJ/aiVZZmmcMYo6vwZcg+a6
D1mEEvOCtbXIatSlPIzFGCwnT0Wj+zC5eABAfOCVNY61MEBRmnczPnWXDqcHShDq/rMqOv5PQXpM
4mzUUPXsq65BbFgsgh3uZ5OkROBsFUyC46aHzCGuuLA2ODnUsHPWg8Ehtx0xnRyRNhlS7b3Vb4f6
wyIkhsT+1RSUGJ7xol6ZzUO8jQ8kYHLvK088iRxczopwaS3r/vTjbPTJ7v3ouHyKIAjWx/ke0mT9
ImlQ9106wq3PO0/iMpr5YHYAj2HE54YVIavgyIY+4gA4rqfAQhUo3jUvWC/RPJhZDWdrmJumYvBl
f4IjQpdPQ+q/OV440t64+o7YKrcZa0TTOuoekReCRI91qDnmE96w9J/kveVeC4kBYEc4SPIHT6L1
awWMuxpEHfeaJ5sRa41+WiGSoQHIRdkN3FAkqssxw0T8Oz26y38DonC8dpABjrU3rV6N1zf6kzu/
H1Lj+jzODsOpfmQO6pUzzXjIqSNfHhtZwmjWUOqyJfw1IyZpt1usa5lkxfbLr4qruC40plU15X6U
iF4DJ+af6dS/wfl9NNhj2ImAGvqiMeGJY40nj93XGqMfeh7XzQmBGTcYdaNA3p7J4b/b6M22RKhJ
3KUk2/Gv8hndH6+cqaqR0+3SHWLIDLfU53SOcvDbvWKK6QBFkdamxGV2ojN1+m2zlOryz16sB2Er
k/s589bvKN6li3lJAirFu0B/Oi9V51bJo5bPkYGjLJI5MHaehCar8MYiKrqBz+kIPMBBsHRWW8KV
khp27SolGD+dFrfon3nIGhe7ofy6LyaWWKhOaVWenNA8lZfSrsyBpISMzBWQiPVsGh+56iniJSdr
M4HXM0zQ1nDUdCgs/kd9TGvCvSUaUFMRTK8vRr7nFQ6QqB13CwiDdFGSLl5FilwZcjp3uQSWW4mF
RccLZQej/x5yXz58Tfw7EYRmnCjd373Vdg4nobGeMiP0p4+jewDHn3orSzT3mgzJqiUCmmApTLu9
7zQiBBnaP7uthueiyq0jJxdXiZdQ8xmSOufoidhjsCY7umIVZihoVfS0qOwTfini54vw6cuLcE2p
+jtelKtiJDnKvvhsKn2jCuen1WCgcM05tnJFsqLi82aWgoQpXCIIfdNYyasig54/OAWDeDXTj/Wy
5bBAaMVNKE9uPQ2YAkq6+aj3Ocb21Biv37hc/6mKrn+UOW0zFd/YGlPCYlFcuWnRQfYd4Z/FeKAp
E+0FzpjyPyQ0VNQaI2o6tf3c+yTIWxtWmlrVzX1aTIMcJlM5NJ63v6ddcB3AGHNrv7olObqnGr23
JV5BiQte+mFu/mqtCVPwh0oEuqka0EdZCEQw8Gc6icHy8ZMLzdeSd15a672nlhrZ8QWuKzJVljFk
JB78EA3UXiXuf2kgLk4jlbqHL4/dKZX2MFLyIWuI8uBQRDU3dlsJBvOR/nEa8uDXQcNcftGcgI8W
8190g6LirvqTMQuCeAP07AUkhLlALdyVctfLaGY4qeZiWJp1587OmpDaAQuEJm7bHkanQsi3Darp
w9v35fJof4R+/61qusEEZjtGKoWLzJOlnxo8L6NfpGMQHsJhz/D8FXbrkscc55mmNtWM3V+dOPkn
K+0+lap5YNmowJCzoCry6fsx4YGfIXWvKpyyxM6yUQ+vJhgTYVhbOgwX6dTeWiymKpXjP4Z67/+M
qxlQR9PbfP3c3bKfeYBGiIk8XxBaqXK5CaWMJmEG17WNtIwXE+uYsXuFNcUhR8xOY2w8ciL3d9pU
YkmgeUzCH5fhV0R4A1gC5xOB0p8nxGPzd+BJWpnnVUpfuw4D2ZIxzbapB8jZjfak37tf2n4rxI0P
rumyikxnPu9Q8hdZZJAZHHSB/3yMVd4LEXyX6QloV95IbZ3a6J6eo2hnTmlQIIrTHmt2f8dFf2h8
XiWtyVH+titKPQBngjJne+mJHDwLftg0OtCOAFw8o2eAV14Ckid34sOCVJRT3LApZPSKYU8LLlGt
ei2bqaYTaiOIvAo83KjWbr4x4QOv54lFM6nC7oPyeCu9RXzqx5SommBW9HuEW+BktfxJeSH5Kfup
7koCf9O51b8ONejZ8ieE3bHobwDkRBmExmNMOLRuy7de1+HKNDQF/aDP58oKFRr4bVkBs3jfgyJz
OtC7EodLmEnNblAkbZy5iT+yyCzqaQYJTZxL+EFKlBQapvFtUPpAQifaxsM/BDXKjGzeIn9yhXqa
YKLaH4hBOCucy7+NivUDsmMzhi5YBAdHXlBD9QH8DnHD7vTCUTjHBdCynQuWvWEESy+s7suLbFKC
Kk2GHYb2rR+tMC1WEa/mK2EoyOr9he5fnTmE0k7FgiFKZCMj9tJDEe8MGAuzlgcqCQhYVEeQBj1/
xHdJu3qfmnwQVUmRGOuIyahKO+5IgWsik72V9k0svAz4yUYNx1XVsTB09jIHG3EWOR7G59yFQhab
0ILFWwUvI+DEpd1/14AyNmfG0DyJfS4vw9aPtwyaqd/Rix3ujKUB18xgfEzwPvlb8lOhWlcqNUE7
zJe1ENRrDF9vyjqQ8GrM9gTqxhrqXT+AFGPWEYWJl9WLx3QJYupzdLMLtyWJPttCQT5yFSAsOXe/
GcOuZDwh0MuGAHkh2DaILN/OQos5lal4+PdkAbaVshc9nSH6T7oLr0CIbEISQujHTfiTCNEQF6XR
u/Uxl9GKVbABh6HTGJwvE3/5aAJr8C6v6B6C9OgZpX2/FMdyv3dhkF0yo6XsH4RWQ2/Th/0eY5NQ
vwBXA8zgkIBZ4s2nXFPHwbZFC0+RI+zBVypdSqhwhOT8ckBX0XY2jehSRN/YTkOTSpjslsmHEX/3
3TiAhH4xNv3iXV+xyzXrJRnZj56zcPJxRuLmUVyMQbqX7A2yR7SJf1oR3IAd76Hxhkg4N29QmlTG
7wRTH7+PEWOyhxuHkcgs7Tznpr0kedVFo90t9Qx8TGCSxhn7o0RUul+DVN03jxZogAKToW4kdkRN
ymzypf2Axr+UhFmyDooqJMJwG63qkc7OBMfGe5EFFHlD9Cwit270RGuTNbzMfSd8v46dbmoE42gD
9MfWL/f0A/6zDKMK4dDJEXUtqGdPZz7/31P7VVjyXQXCuPE2x4PqoxHjdjuJx5uZb8iLrQlPiA6v
owsgJe0KaOC1EWYZxYYWbVJwPEh3mHYzyEKbQzDe0cdRcO80SWI7G43drqKsH0/Srmzc0jCYXvxH
gcGwvmh7qOykNiz/hmOdhN0dlIsiYMcErUcb5AqiNvgTE+2fTI8jYTvEBma67MAUZXUXbmE3ryMx
tqtfuiAbzLmRAbilNYCRfwdLeLpR5XP1rj2a1wMhYAA3j9YiF5Dj/IjUafZ7ETEj/be5xohIVXcS
iRPSAlKt1BM0OYSIjS/cCOQRB6z1rTLFWhOB6cqA085fgVYh8m8Q0wm0UqB/PAsMixWZCHl6HS+4
uGMgiEhfpwr8EYUPxIluZk58etQf2q6oWbdrdQnLYcnptmxGFShC/LuNVtLelH87Kq2ZadvDkcfh
WmbvVR5i+gsNKprpYfr0Tg4We/yHDVSIOeVWbwDhw1BujuS+wXGLW0EOmezrpDd7PcWwRdlxasAo
k1vBSnwxkfKAce7IL0vW3yQRSrohxZhCOSAI5ReCez+aR5FH2RF60ew7cj5AklKF6zlQPQxASt9w
V/7k+C66xr5R0F+uWTofGM4dKKf6nK+GD2yw4YvNhK1ZsZoHiQElqZ39xJHlfjlPTY2maLNY9NjF
KKoqRe6N3YZaP1H7+/vUw74fWL7VBHaiM5gSt3nsGYLWltaS04MUO6CNED47Ozpn/urXpAatPhJ1
Ry9fcV9FGUM32abou8m1aeND6yt9f1Y8wDq7DJu+Qd50sCl7B+WqcphwU0O4LqKjzfdmUVpxQOYp
WgKi7P3BlT9/fxf2mPOdkgZxFidPFTv46rNcyS8LwCI7PE9gwoPhHlWoRgriTZbNjoU2ItmLY+Df
hoW8/GRJvNnVgmCvxFnktrXRcr10tUNgtSMQYth2wZ3pSq8lRYd4U1iK6sTLiDdWklYnoikQGivT
HE4CTzfb6gpRy5Yy/aNr+Pqew164dpjmMopBfT2gKJJ/qafxK3/HYtrO1A5pA2RBEOUjAs+taQRq
bCufhFBoEvAp2kgk0wb5EB5dHUbWEQUevtX7oTa+FbFd00tqaFD5WnpB1r1NkZuhCHt+YiqaoJf5
vMFW/m7ZcuUiP4NiHvL4q11YhdSHKiz+TWSf8Blc4HTyPL5x2kHdHYtvsfl6o3KGVC1MhL58PM4H
xCRgjVOGPdI5vaAYQmL1gJQqD/Lg0junrK/Q/6IEnFQFhA6xOV3Zvnc7Bp/VBVw+rIdht0Tdpqnt
SvgV3gGdVeqNIW8iDmxCgnO/f+t9ywdrRGrow8on+bP/cDUawU3sCvWRir21WAZrBugE1Q3+aijh
tNGPlg0ddRBNul7+Ggc+mklzjWD1nyqzl61ZSQuZrdUooB2fIUbcInNFfyPeFQI6iXt/sIKrxVv5
zAbrfABRNJAZu62G5jfv0usZHp8cAoeJv09IBH+58N9v6PhwJBQbn6I8Ae1Ow+OVFHvV4vccUgTd
YCIjidHXWcDn3oVxi9oM73iWkOj93HKHLgAtKVO8+H9rH+mIPgLhDdiwf2u1UmVHa9mOrMO355pL
Gq4vX396Cttj6L/ZW3HzKwCuC1MvItppxtS+auYJkYOJp+8nMRuuN85b+gApHa+/FnjvUb71sM8B
Ne6X3q+wIL2jPqJGPybjnSrSNzj73Som8079MngWe7Zj9gjc/fZ8iC8e7LFqWYRds1UsaPEflT9C
vyuf9GsgeY8N7KmledOW/k1WuWMOgspGvZqlviAOkoLyYlWPhTsmcZPaBKtSUDxv4b4GwRsBv7OD
wr3CxBLsTlQbsjZYgZfdkihIu1xq4BtPCtEGPToheTfGAXFuWBjZ81v8atgYc2kzwOsX1JWyXP8r
g8rdCfc2+b3yLpEZmVQkHC/62O9QA8dimYHRc9qrRAiO70t7z9dlm7SFT5RAYsEHEEZY77hHCrHK
hAd/RZHPR0feZkHkE7UtG92EvMnEVwMAW02NOQ9YQjdCF2i/guzAzvKrtXmTn5qCqKDhat3iv2bB
XlqJYN0DFg60tP2cGobHSSiVNwRRFbDZLh9TDRMbJLsyiD8M7KOu3bSa9Yt6Fx4PGdNRyyH/gCgM
uG925U5ZFH/8bNUnEjaE4Ii/jzaKkzuxOcx/op3pVRMuLmwaJzEvbhcBZIEmgnxJhjM69PN4NAIk
lesqgdHky9xfNDWXu+IPhnwZIlseTdJbfsq6SEoDx314LZBu8HFo3HJPAYUGJoVttvQ3WZqZJ0yF
PuPu3v4Xr4hyXp2M6uleyiFJjL88PLNnuKuy8cG3HzjeqZQKRUSHdw9O899dQMhsX0GAE252hXik
8XyPhqHo+GWYb4ZIPfnJMeS+9T0pMVsEn2rNfJexC+rxTPbOe+RivHXEL5NWQT/eI14vOK5s6+fE
ed/DtxGaZp+56gDeynQ0lIEA5fbl6b6SsM/UkUTyvnwrypXP0vQzHYuOFhe/nwoCyIj6TLswuri7
WIvLnRKki0OsWKI3PtZOe69gCQY8AHb6336uX9G0V5a5qSs/tSu5++WCJ/jRHoRi5AxRzWNgaKFA
bc2QG3rO4MR9zEkwgGAtxP+sGCQJ+aXifV3HuHnadqvJ75Ugusl7iWmR6bJVfZzg93gbGHLJBlQD
/rd1T0p+lpzquTkigd3iJNlc99A8dCj+cwUtFD5q054D+D0n+BNg1yiuglQByzVSQnSjlpCj8wUS
j48V4G/SZYvb3K1KaM3zvfrt3y/bz6+RZdiX+UHnQ3byTv8tuiJxzViextwT5zOhJRunRbnQSTtR
r6FZ1V3s4t07tIa5lcqYsdG1Aovr5nNkjYga9RXZb3bKfbEsgdC7gxcenmaHSxEBZocfGb/kiQAi
jeUWeL9N1tkWhl6/oHxupBS06o2IaJYh/rMD8wyX7SAUxZZGRcYfCLAQ4QBSsBjatrNa6mzuLhtV
618SMzNtHzNvqeRMB1phmGQIXUDbT3sligZjmA1/Q4YBpv15LXWpy9OKCmVZK3vMjLmUqTiduYLn
Aj0sNkuw8vBTcp5jc1F3so4xwEB+17t6ykp4yNEImZDNNITpBvUVC3fLYtOH65hWZDHhXw5fuV5Z
pBai6I5o87J7q8UAjbLj3v8Qku8moPBuOIHh8EYBeji/NjxwXqsYCA56pYM6wJEbD//mfWy7rrAW
U54vItsffa8q9TLHaM/pP436WHF13inpHTJKbMaRwTm55O56WIHy0cikqr80jt9oA/liTo3fdkGH
QAHk8w8FX7RXbU3RstTImWWSPLCr7zhxDjYZ4Zbs9t24g9PO2r5TbjgmwRjhk6OMl2HDhK5LDT5r
/eIL6K70C1AIPf1sKXUezz8nXEJx9hUnCIkxl4lsPLdDpkiq3Oxeia0E7zPSDBSmNuMM3sV0AA+r
WgBL6Y+NxNLHLtKwfq4H4Z/NTI1V01TAbjcVmcwlVsYtTCDYTIyM58r597VP/M/MmOW9WSkakPkb
JPkAD4yS6URNI9JRFpbE9DHEQrqT1PRsZ3+kVcg+dpENCr8rQAG8kQW5ipd8LkqZdvVZ0bD7nYZi
RQCLl/mieLA7JnjKrIQFj6wuG0u7Z+4Wv/5T56H/TXEdk2/hgfOyVLTbq5ixiRDs+qnc0IH3g1P3
zzCqn3mMdWWTXz+bdKyzaGdU3yusWZpM8WViikUi26eLxQ0boOF42o8/vbNridg7+CLS1saYz1Gw
Knv+y513B+4IIc5AV2DkYFZPZ6aFu+2YyVP5CCzxY6h7v+MJ/LJI51vdxnQhAqV5iJyP7BkDQGET
/z/wBgBqCyhBBHmnS3M+9RtCqFTim/rex/WR6Uaqe5xW88mIT2iLf0OEBTsWzHbkVmG6wYRh/SbL
DdtxvXuw9bx2qJjvCzSWsHOYKhivC+osVpwQVzaQbs7s+oS6HJRsgY0NAjamitjXntmPoV50ahtw
j4mIpQVBHXSl2NJImETHqi+qgkgg9eH0GRQbAMFuvLuRpCT70WIHnEIe4BubJ/Zy1L913QsqJ4uY
OPu9JEkyIpk+5DxkFB7M8VTIK9QS80NnWW4pYVWJTNcJ3IBnW+w1ZxUPpDIUgGI3K4LZjpc/MlfR
a0fNqdfJ8rTPbQQeXEp3/5tEBxHvtBSr1Oq/uwzrUvFrZ2VVFAiVP4EQP96tD5nkChL4QoMMWP4o
ZXJeuNe303QLKyzXjV3TKqNXoyv2hKiY/VP2qeDzznC1ldfpFjFO5dqn4qK0bKSzJU8jS3xK5W5t
1lVPbisg/iAxcpTA1k42CFHpvYWscYO9WXz2INQtLDSgWEmlquxAxTGTxNNTMMTWEa00Xi+Wihbn
AFUn+RyB+DOpWYHIMNBVABkoepB9GZp4ILceYD9wIMnRKwJCpQHgb9rSulIBs9ztgSPNzygExfXa
z2TTmo+9U2jZnnraZJczD87af0DKb53MB6MXwOSEzc0BLXJzl7rYCWCmNtVWZ17/eMo9gJfAZbVd
p1d/Hh4o5Q5QpkpeHRPcZrCF7lsIM7npLDMxykDZ35BYSAO40GHszDOFKwXUF7eKQUaeaXCMD97v
VvsRmEedh4Tin2fddj5dprP2DlnTv6qm32aRzmeYMMgsLFMwLbvzLACo4Uw90BZ0ozTrZVQyO42/
CAwu76K4/VcVHI0LJ8uBjKdMlQLok61DNi4zz1FeuPNXNenXLKul2dXnCuvepN39dlzj7irQKvY3
CAWXyQwLfidpIPMsOFXD7lXZJMt6pDHIoRfOj851JMdAiWVI5tARxyX9ILFFnaKLwwIaxQ8868xp
x/KSbkgAqMrymLCTWKhVuPOQUMAZE26R6Ak03oKNaRvngmviAOx7/wNclkQCMIw/57I8BbTbvq12
/7uOnK0ZwxPdOCmo4H0chW9z62frQkdaoXUxW1dS/1HHJUx9trj7xGYKgMfXksU508Asas8BF5nf
fGRhNp8w06MwWkMkC5eu6zcN82V86twdDqbcYncp+qic4bziYi8CjYrH7Ekp8rtR16OtJkDMqGc8
oy2lxDmoyaSlS2QqKpz0mbaSOOigVnrH/NYZzoVUCwAdC5NSn3T5haRsowZ0wL7whJw7Re/ONG8k
lQiwB8Cnn6VQts/EuYT/Az3oJKGldJYXAnJju165+J9ngmixIZOlmbghvWh0aRBBsPb1a1stDC2J
DNZnKubL5BE78SwYSStoPNm6bofgXXmFffAA2jmCIcSnVRef6Iv50TQM8HloJbX5znrnEDJXbsXd
c9jKLjhfocuYWiHl/dCBMIXOudAVGqC1Sbl88qIMPsM5FlmoYLfsXOT/ljg8oC7gxM+ak0pDwrT9
YOptZrxjR19fSAGUWSlzrS1lrz5qrV4mVdjweNshIdAEsliW6s8ehI+Ncc98aZVQzNh/ZxX5K03Z
NXMTOEF0S7xwXsc+ZpJe+Ihlj1b2UTuvrtEpbR1qe2kyqRXCOlEs6xsLsszeSpa7Udb9ahUzFkBu
DVSf7/LoUKWzIm74LZ7awQtxFhK1Rl3G+xXhE4OG3DUe+bJR2nWdyoqLDNJOjYvxcJLendv4yds8
/nviWcQai+VseuOe4ct18JOluQkjvYm1tIdgnX8jln4htwWTpIoifIGgzQp66ux3zWLgokcyOxCo
9jVWZ5BicxyXgjL0rXH0PW7Vyh9Fm2l+dWMlRx3jDRLcSp80yJdmKf+Ejcl7h67rbCSNO0syfT5D
r/Zl0IJ2MHfQDoLEvxg9Cs77h65IhzIjwBV8jcqF3N7akgc5YzwL/aaOUeaUrEh5jcLxntjt/D1/
IWJ1IpbJG/KOswQOeEk+CSM/WvWXwm6lWvxHZ4oHDQTX0583aColeWM2GsZUaSeVBe51XlbxXnMV
55J2YtBmf0DaIu7b1sUD1mFsp1anX1Jzsq8MQoiIG7xQcf6pY8o747QCqsdw2gs5G3qvg0mjZWmm
bJgSJYI2sJLKLC1JveW4EZ1vDL6klak0HL+rVc8lEw3z5YziMgGn/i9FkdoKMxPRtXJTLQ9RYh5/
N1f5CbYqtkXgPZ1eesp2Es4Nm3aG79VvAkJM/Vvt8/MvedS4kxZSEo1EUxyu7uqEpzI6i4vCyGhS
DdS/dPZJyxj2x4eK5tOBSVAEmVtgNCikohGBuhUtIwTD/qdF2z9BH0y7xagYoDRsJf6QR5/8rTsE
aoyNGBL+7wnATOcMTU97S5KLD9TXA82dZAFkx3ZoEqw9LwWDhVuURU4fzEfpXzc8VZ+6MsCpxm2w
VFmlHee+0XXIq5txQhvRHItIYcvmXOHjlXJLqoVLYgTfjBH2aMWWiUzDpINiPvcPl1XmVzBnitkq
ox8FiDHZM5p4UY4E/QMy4QxZ34ZXAJLbfQC4MIWZ/juds0PrxYnbiuwrTEhx5bYlE2drn0ugofNJ
RXtBZQCCTHvX26XGhWvdIly+xPe7sCNQiNpgb50tFQPP5XJTFUIxxzL6AO13IrYo2x/8f8Oe3XZI
vZP1EQYqcNaOm6xlWIwxppOXSP9J9FkxdjnbqZM71lLiJIxN7W0mZu9VPui8q8obuUvazZGqKVzi
4RwUUZO7WrZvA5AujKC/6qXN7OMwHMxCT/bGvwu6+F5BOUie6yn4urBZLw23seaO3JHAMbJLPDKj
evZxlkDpxaOGyon6HacdIAb8JX+k0xbH3+DqaBlrSROvGEudGEk2wcyxfmqV5r2kWVoJheD3kwR2
EPZoX79U1zeLXTnH+qNPGcrBh82Dxxt5zDaX6z84n09ktppTy5JiI6mIfDGr1yzRlBtIZ3EW4ENU
zU9FvV4phWrfY/XIOi3b7WR7xq1qNIoeR7X7n1gB1LCqDdQdp9iXxoM1UiNXHVC0ExpuJSgusCob
wHgzZDKUJyZc9CQ2MurAUgexMzTHTdKCw0lFGtfaUSY0DCDz39VZiWJADtmPY9v6H78pjXZZr/mQ
Ntb0YrUlLR21624XPZSXH4lWqZuP0QDDj/HeESMuB2WgSBq+AEPSo4OndbYEBla/gI8lEmQcfJiu
Wk2CuT9QRU1ba4I3cxO+/dL/mMGQuK/1P5uqjH8Y+XHEZwtp1MplV85uyTzaxpq/Klh1Rgz45ihP
pDq2T76/NVJtZ1iyNN3+tF1SkAbIinswVJp14IFSCp8S6dNPf4uS2S4aPERVFxMm6WLaoe+/A1Fw
10iOwrwb8LQ8lCVaz4395BZN+sSM8rrZU49WlkGyKMAs4GTk3h0tpTg7DIsmM9zR7u5wvRx8A6o0
VnhSy6TaruZXGWDiuAOpo4Sgh2RZOaH8ivghq4oOhieRx4SZGuwKgNCKWomlHiUjRy9/2TOIo90F
PL7bDPYn0ACz/eaywov7CUDSOwuRQxXpRPHVuxGPUE4stbORW7FCJmoJEKAsuy/vJ85jFCSvmKkj
SeDIC5cpWxiWZpLn+sM6iJM96yp7ThdzTsLytp0Vg8DBqzp3fHvkgtXeEULo/cZ6Rudg9o07kvoH
+0zV82nWYEYZYzSFm4YTgJLs1SBMCN2xFS/6oaYz33+YkQZiDQCBW/KqBkxw6pXWnZfHJQvJIYIa
24VaOQOdpVbD0i5Wxw7fXJYsXvK+j/5hfyi75uS2p6vWwFbD2iJ/yG4IPa7IspghRZvBLpH6X6Cx
B9fiDfDqhDjRwAg2FHGOLUqzQX8x63nFzrVkC2Q/ZasBkMhgpCTTLa99X1yiobUIquApnFYclVYq
ObaUxndB4C3w40n1ewF7lBXVUKZn9r2JMzE1ajdXCuT0oVw/bxUwsqzuYQklV3tdkwptoAcjK48y
O3/mldHC1nwXfpTNILq32CkHAwe6x+K4XJV3ZzgLEvXPYG6H9iNlV5HDcqDpBAkb5oIH6Yb/FWKV
eYaLlhUFNx1SWTzwlB7li1jott6acEIXorlNtSOV+iVOxb0y27a8KA4UndrjweE4MsH0g0TG5Ay7
jyezrr1yPr0eTB1K8z1ILRA6fgGGoz2VNhJXf2C3PA9gXRnHwFT9///v+c2XaZrEzwIX+rKy0Bxb
XGqxSuZglqWQpItJpuZniCWHudsvQWlz3A0br21TYy660G351cjyZ9eB/47iAqrxNsBOXcQnC5a+
l3MvRAogXclBaln7n713EbaBUxvPC+4AOMXQ9ljo3Txp9talTuDiveyuB0t0IpW5KyGDeOObDbz6
NIDNIv5PjCusmhrUAoQWvd7ILe4rtpoiW0b8QQEzExV8y4gasoYaa2slrJfeU/6W6KklgAQCPCq7
q/78S5RcjYRODzxhJgd3THmnfJBoum/5AA0Cr6nIsjzQ8o5k7yvurHcOwf/X3jJsQqRQcHZk6A79
e2zE7FRpxtosBfelMjYPyBhmPYBP9HC4z/TvqmHimoH8QOjuhNgqezK5TeD+YlRvOc+WFmQ/4j+V
/rtp0tdFCPuRXBlgmTG74G0cD0M4GC2OeNrUnmRvM3WlduYTAJS4Wm3tycB60xEtpxdrdkaCQ5FW
BVk09/yN5BCHqvImXNgXtuMv98aY6+um/suBGcTbegDmZZ9qV7QBPITGnxnINBVn3nOCq812C90x
p4ToF7HLAK2C3GlwUSc2S9cRoDjauSm1vSkbjJ8/CE1QGjpQNsN31uJokQw61B27DYLO2axyR4za
mwO8xVurZTrDZJM8u7oHmXJ8zhY9hdo8et5elrTqfGBD68XcN8ATpL063Cp+7LC6OEFEC4SgjGhq
e/66FuzHVOWuHnQq6bliHzg5YhWwWRvNCyYM75gvo3uUF/2WZf67MKbEfflQPtvge28W0s+qSzgb
i6o93btkLEkHja4I2P2zz67QsDFKxPAmyP0T5DNX1mALqi99OSi0rmOJGosaQ2Jj9JtHs4nCymrW
6EnJwKmtyE+slRYJ6RS4BCBjMc/Z+LjOkRds6e25+eqqHAnZOUpteWLnlfPTHwfUk/PvlAvossii
4kYyQB8eY3x60sMo3hJtUO2lKZe4zzOREP22mI+jN1tFOLFUW60xH9PHFHJBJECFpo+tlNPP6zQ3
pBroVu7bRzwRgQZ3LvdavAdJFnoMEYg8Xd5ZtO8gJdGBZe9/xeLmSUrGxjBqLFUFsnHvUvsBuJiU
1FdKeNbrFR0AWIA5Sc98gcIhrjqA2k0qvloC4hUxco4v7pqxt8kOXhzZUjoyUjiPAn90vU5L0PBH
sL6PL1NBYnEMDw2GcRZ98mkmohXf0ZlIDIUDH55++vNNP09GmhsvEMl5YcDCaNDU82GO433tMlKL
SxkTEaHmc1hCp9s9U0jVOroijTXZNEnHNDCt9lQtz2nMDppXy38hW6SQqsKGWMoo/CRb9jPRmK9C
C3UsaT7YPFig3PN9YhLhuS4T5V8ShZZ7NuuSZFlyQazAeWeuGIdHuKzljOk/Oo2t8wUxjLD4BCX/
9++C7ASrDGtIGWSGLiJcQ/LDNQvjaS9ZxmxNoHhee3ZDAm+t9T4z/ypKKAkffzlxKA4GJqi6eRes
iLrd0IyegwWMgmsNRrMf1iS35xrgDAlHcfCQBy3LVipycKv0Yvl4U3hBjUeNvA3huJfEpwJ+sWIE
Ie09sD/BV+ETYy7/diTMVlPBRKJs2INeT/IsWpWmst1v81gDDsGRD0FAqlHWKuv2ohNMVJeOd4lv
x1rBMdFIKLYW/5y2V9KjotpAWpVgRjYOr3DA9HXjCfnYFwxedcPpYyoG7G/bFSFjh/bpXg7gQOUN
uqmtgGzps74MrW9Gn104N9jV+ieUE+GF5SRu5VYuMnUQfiWRae7h+PTljkddWs2M+IFXMr7PIl9G
4Q0YcwxkQIx41bwdKQCFI36r5vN3eNhsLqeb5R86HbiDON49jXvc8kux5SbQTbmIsQ3+OWz9eQrP
WKrVfNXAr43NzuVyiKtMGl9chnF2XvGKy5WWmSmx+0fec3zmiAj8n4gzwmBOgv+JcCWiEPknV8lj
2XYAtoDhW19kA4rABFhsaJECYA7hfV53DSYaEX9RWZh/Mr2ilu/bLgCWINtzKai1Nyect6Pf/j3J
203CRfAYU6IGpPh3fl6oWJYNQux5X795v5RzPsskzKQTj0z5CPSYgi2qXG+v+JlIud4WPcWw71/w
2dBBomK1EKUb8e1BU3rk910mIFKweb1OaVZw2ID3hcVnpqtYF6Cm7r5E4UmFX8abQeAevPlSkdal
vwzUye0ja7ztyWV1znTBlqANMFzEp0w5BYtFbStaiSj5f4zsGIotJWm3PL+99zIHdEpILTWDNE0Z
5C4vSC/7WbbAsbBGdAsuHsWXSnqlTWnH0sHiUG6LkB5dR59tVMAKUdNLpnS4oYDfjVtUvq0iVcP0
RR+d4RXIIMCHD3MPRY2qiUNiLGsT7E/F60m8hFNTf3VhHw+ppDhSV+erx8zsM5xZ5SRd6WSoK+lz
ob7EP9D76u8HRN4RRKUjgXiirtfFyjsq3bCbOJK2VzLrWF9q1smzPzsj9x9EU7YGn8c1lbuUwm70
o/1btu9SNVYp3EE0u5d+7TOEddYZ+f0crpw91OaMiiWGPwQJjB7G9JVpwBh5C4Wdl9KSERI1Gkd5
Cd3In48c82WcxAWq+YEPIlM/jLjSYYSf08Jzak83e+wKMvtOKIwgAz4sWS/bpJSv194KhaxCjVqn
eQ1n/z4YbCs14YzhCU9KNzxfeosw1Qcd+EtuNHbjc8jFBh+1YxEAa7yo0TNs9FW85KBlW1IQAPhs
qwiJQfaeTLPEsvuBWLDbe0RrIKrnny4aQQs57GVdd5J3npUnTSD8zQactSiWW7N4E1JQdR6ESdv0
KDxhpTYX92FSIt4tN2KCvmmJvE7OzB+4XPyikbJ31tUqmm11U9dnCAVHU/Ylr510AHpY71UDzgLj
An5i3WXTugbletPRPMi0/PHBca5twbmZTgDjnbEbjcoXsufcmdNiNwJuijjGBhacDSpwamuKCV1J
jZk5OtbVlaTTfBcaEWXEBCEdTtD9XSu6wTh49bPaTnC2w1U8x+I3Aq3N2FuM8KXRqaqEVlHxtStS
QJkPJx5jAImSu1y1xdR4SbgXg90jut9m7LGn4UYUG/SX2qX8teNWRo2sHPccaQbMzrRksohwujru
2bv4tA/f7cURfWDv0gB8iV63z43BVmRmENp0MBnB+J0i+fPDMF94SySwcN2gAEvRGykba0MLTgna
MlAkilRxTGeLqBZrHQKlzrse8Dmd1Huhd59U30PffIsZyKcaYp6ZTN7Lhzj4Og32nCC74CmHoJbN
E6uGHZv9js2XyYtrQ6TGoshQmVgxQVno+ZjR9l44k/Uma6brm+PcvhLZ+RsLL4cIipmV7lIj0BPC
vfysoTcBwXYpxuxwY5FQ3IwO5r4d+pQEW+/XFVkaX5oJ/u3lfHQgggRi4NM9nJIYgYQAn+zJjg50
jBwuN+RD6a1cTYe4OX/DSk2UIVx62sguEtd0ZPmP8Mtiks7Hhnu6sCn9DxHN2VAj7xY76DyAjMyI
Xv0Yy5fddXREwjgq4e5JS7CgWEVLyLyfT6JzXei3EQGG1I0MblReQdlOFcgbfJDT5/cSo2cmlKbY
kqKxJLlvn3/Zqs9rePqw84ukjezPhfNUP/9r6m3kX5KFm8iGUfirdIxsB1CJ+1JQLTGG5E0CO/4G
ztJqWmXfkE5rb/oLm+fzoKoOOzgYHfRwUli81MVpoj9v/91isiO5L/DVtsGrJYcHnqCexgjy2937
sOFq0tWa7dy96KYAggZ/tL2MP3wNx1JgS8aWh5MgHJ0yIYDraIXbp1LIgtFQycefPtZWC6XO3vQc
zqX040A70FpwhbP/q5/pfGBHwiVPSnIxpm79MMCFCKp6hOldO6hhMWpuUA2MBz7yVMIgidIZ8FBz
AQG9LKrEXmKDRdz3GvH9l9aAugv1kGOrA8q9kDQYiq5lU88MHkGgeNIhwvQHZtPXOvhC1B0qJJrP
klxuOM6X+1qRgyVvcF0kdlkoqbN/XVoxcaq/mHico9rz1QKvShLJqulQdoBKFKvB/lUaFkONrnXy
xPhyYsTu+WHykkhDg4BLIsn+Oz006VCPgk3u8p2CkU5bXhXOsj8JehYuloavcv1RfPMNVCdq1+1n
DIiScELivvuJl8KaU7vPyLPX17Kj75KyGJu3xP5nVyDPghRhGRvgg+YgeK/u2D/wa9BR3+VwsN2g
AOs00DdV+/Zirr20eiSoDLcuClVFNiT4Y5uqvBgn8Ke1fL12lrroCMo5eVHZ/KidQ0Y0GI9y++Kn
uvLGH5UBfK7KIz/TtAg17gc57x7MTLJXtRItHLKwyEXpbQiu/qvlLoQZaUIVTaTtISC3CsdXjn2h
4OGQ7TMZXX6f4HJHzhOfqkDQFzqOonNtVjB6jQdaZqbk4LMAzn46zF79ymNsRn8Org7Pfifz6HqP
9bh7IeZkrDL8kVc6Tlq87Xl+zgTKd0NUiIAanRYl8B3nno8u3SNJwuc4g6xAJKrlRhFVZXVooKhg
A3ewf7mnDLZk4iflz7mNuBEvXBs3FzqSLujBwq72aNU8XNndDKtJXzvBv8p9fAw6y5GcaH7mqzmF
NnNM6epWeskEMQ3xph9MhOoJ6ULz3GqNj49uTytugsgjiOuEDWWuZoa+47HkO54eRZ+g/nSNcTth
tFWmcp3LT1U1IcCAdwDNd99PjIABORASLXK3dWDCunrj+82dUuKsK0coQZT0MWH6k0mPYUPpdEW1
NbkR/rXHpuOvxRle53RU/2+RMr5P23z5qM6bY84PNvpgoyXrmQH46kFCfUSY8D1BQsbCO0L6Q+Q5
JBICHb97gz9oxn4Me+OiZ7YUvBZ4JJy66qjaWY29waJrJM9DeSv2NZOFjrIugurfXVG21L8YFbjv
5V2kkW3BqMw5YxHUKyY01T0dj88Cm9ad2kK+0zwK9ukInM6smyCdTE3zvdPLI2SQ4s6z05WYjjGW
79Xr/k+rMZ4C7Dh0UqEH/oiYVdcs+2vMkq5uVS7iDJ6xE7VAxsWSaSHtrGa19bDf4j5N5aC4L9z0
44g0UCrTQrkyTeeK7fGJQcnBjblXAyKEqGEZiJwIiNunzCqUinAeoArShrJwWjQxwy13ERv5D9/U
nqyzHC9HPnQEEQoYdwK2n8ZoUDx04ohVPmvL8sY3v9VUYPszxjnToW+Ew08UO4tLwFc9GpFzjWd8
z9IAAnm1U+d+SeykWEixth3N3NOonolN1HYBuCdP860OFWqLpzr9+4xA+4xulJZi9HsuLFg80X8h
ZZLxf4EUI9nCfckvfRpd19ohPHugg2w3+F8Iohxl3Uteoe3IVEg8EeXVKVy8RBrP3bFewN1wRUaU
BU7DR7qeW+n0j0GWlaMlvyxXrlWsaxDWB2ug/RH9yKOQPPZjwVn3pqkH9AIL5N2auGrohg6WV3Z5
jSVbDYvJsikME7KMj5qrxEXB219DLwJ7dju2mrTOnYS6Dqz3tkQpOgY01TUAbWbOf2X8FCfQ680K
DxUuYapSZV/tVFD8xb+ZE5zJQY/Usv2qxt7wX2pCSoMrXeCw8UOha8/DyqI9yK+HkqGeJzH9lpTC
tYyO4TRX8MNeqUtGURDbu9kawabKoZZQVRPHQLtrWjuvuLL69KvDm1MjVpn8NKQlYqoATpyYPidr
KM1Q9R8P4WkJ9QhkaD/TvE1XIdEe0nNXqYg8AY7bhWOMNvHylp5f6+oJVTuzIlJANQd1n1p5Bz4J
4AwpyocCJWCw0exJ31HgzXB1qcsHXB9MeWT0Z2Yr2tx6rNrfflZecbck9JaRDCOsu+8gRUc9eKxu
SrOlk+T+N+9xoXiGrjYCN0Wyor2xuqlWGDmbNd9+V5F898Ys7NInS1qHmixRAVYUZkVZk35ayDrz
+8UnInIdIqsvjy1Qw4OA/dNxp5GKl0U4nf3vzFQQy+PUjRW5cvXIdQsaABoXcz1GFJa/EFdcJDz5
cjE5WQggxBI/XFRohFB+r/4AAQo4XbRc+HebBMoMFGQXMKuuFlwBvfBcXEXGsdQbJ85tjg3ETOtk
ZRTyeiRAO9MOZPuQ5MaGdWm+a6AhINIg3DqhYk2wbb9rFolxW2q2fe4cjgRwQX0KC539fvDrM7mB
eLWp0DijvtDEk6n6XCgOd98DvagR46QxDFb2ech+se+HELydjAZ2qWR//z1GI+2SHr7dXZpadGVl
t0htp+qc1t8Yja+7kOy0lDwUJy2FidNaLwgldmqUlE4Xolqqluf9tvPAYnVsbh/oeMSUvzuD2uGt
zhgkiuhAbYRbWm9I7NUqcuGnFz/nuf5VNiIf8AtshmoAP5ghnzER3pj/hg9mjFCdj/lW2tbghhqR
x/qWchBwBOFw/r8I6tbFiPPVmXVi4q38ysic6DQUwhWDwY+XZe/6Yw6CFSAeYuE8KUaygpNO/woN
3FxBxxNL52xhf6Zt+dWJnG9gsSlF9F3Fb5UWhq8RatOfwTMFYzetrJvad+fBrvFLCoNNUUkhF6lV
wBl6IMtoQssccHtBmIHQlVTcs7urS178ilTLiRTHlsqcjtgc5iu9iWsjsNcllJP0gdxXkMLrtwFP
asc4vh8b2bMYhDfQAFbr0BDoS6pSSN4xENO0/xLzpTYn9gcvdzRzMHwBDGM/Nok1AzUZC8RyZj7l
Rd5pk0SEd1XYZrZQcr5u9DSbt/XqMH36JVNG0YLpsPtCNIKduiHOlqYsxpXapoZ14ueQFX2h8kUV
ctjAZT/LoWpOADYDR42RwIoF7p1txgqzrUGwPdI8cqiscagGQF35fixKVjfJ9v5o2xqqIEr7he0n
mjI7IX2N1JMfi8JgK1yPjDggD7JyDSUw7PmaxkObUJBzR/BfhSV4yJZC+lqdLa+rqvcJUJkeWPy0
i3akQieiqNPymYc/Vo1eYR3H37mJZk1AFa/KHiA3VDYImwnb21iGS5iW3kWGSBzP17Yf5zqB9AEv
yITPcfw1NfoihdLOfqQT+1hZUIISSmQ1gKF6xLiya5vZ9ht3lPNCNEnxOyhm+ZgBwwCXOT41ruER
kJVpEcKN84CE1Hcx10muW7hOxYl6eTp2uUPVsllMWHPQIVMtO+K589wX3FXfcpwCjkEV9ElonXpF
r4uumD3I79SpS9Tw4sHmlzmHDhO1P+v23JBQCsz/CfHTFkSetaNTHqVVs1O72F8M/FJT/B16XJRa
DoxZvX8H8wNdUgVCc+t/B3lYOytn8xIb/NwEUaEFnCUspsRZdbBleJvkY/yFo6Hx6xSarfjrjhk9
j56MLNR9UORSrv9MJU3vLnS/T6Po3PoPj1VVyTbgUFJv/7gzlVdn5ULu00JHTZvQ6JsvdPBma9R9
sa0Rxez7o3f3B/6iiMVR8G19iMmmi7WrF00iV266DqKZJXjzh54OGHENdTtRGc+2ePGQ3pss0w5N
7ZqfO6sIqspBmLnlzlamlv1vKorNmCyvXqstkkiPc1nF/Ht9g+P9MkkSQ+JuQG6KUF/6lgGB4ShJ
EgsWFBQ2bH5PW0nhVdh38+djAfObUHPU0gbVJb0CAorx54pbiTpYhLKKfScENShfwBilncMMWf/q
GQHRqwmcR7xY+ir36TNi2LRmxRbctwvhEgfVwQvfw4IWc1AGl1NWW65lZfdPZQisQQO3xGyF9lF4
JL6kRfIM5ZEkZQmcvfPNqj2NhcFV8hmQTRLFICEQQeq88HDJJXwvLadBL7YKh8JAU9oVT9xPhFWL
d9YsIQUIfsNNuZldOl6yLD8/SsoZvlcwu4/abJnY+KJ6k0PhfEBAohMyKeTsJBodCPcb29wcLFZS
VlRx+UuUZ48wMveQoacZSvLvdHE0Y+0PAcewSBAdH+eoeQOlhRI+JhSeBDKJBfzl5aHif97KWoTJ
R1GhiBpm4YwY+G8xAtm3cuvUuydq9v/gfCUZC/p9AHhvGRSw9XJEdggaZbqjghWf5PtTEoEEn7jL
k9lL4Rk8tyV4V31X1FWcPn0lOytRefdQj0QQCm3KZv+TpvkgQ6N7Ptn3BrxJ4mA+AdlG/oa3dltq
+pbzOisk2ALf6r0Maohf8Xw5svayckiVjBOFzkjSLgJ3fcfeMLauRaMeERM/OT/4VnEKQYcTNXrn
UdarxlVGIZj6Wu7XEGnwHROPn7c9yVkIoKuVHpJRBiCRZ74SXTfUzs8qWPT+76Y31kRxps1Flyh6
OFjalMJe3oBoaoyt+jTE84oomeejrB90k+/tiqc+ior4NKiBfwiI5KS9gnLAgN7DgGMmZ4AmRprt
6ItldEbrazJTIkn6PjOQI9YP0+Kwu9cMdKOWzbXKDCPIvHiGYortZNasOeprrqTRSLgb1botV/+Z
anf3opOdhvqCkldNPaRDG9TudehpBCwrl8Obu3L7Xt7QiFMSYtD+l0I/BpMdNgzY4xXQ9WUxwrds
wGGK35GySIbJB/+vAzqw4koJro1B4fsYbdJ+LuRrUQJ6OTqBUGP/u3/UC2KETbEpg7W81wxchPDW
HYAyW2dZPQRjwpkurIE4ri3jXKNUReElpKGCCIkgYU8r0LJEzss/a4qli4QPGRw2D9GXkj3AHH5s
tpVUe5i259m0rgnN6g7nRPp9mDuGwocJWPdfBA4EP+nbdsmlp+NdPGJPSN4y2rTJppLRh8VfRn01
ldUU8MPBk9KShRI7nViwkmFJqaZlwoj26dCHmP4I7ncxkN36DbkiaQaYS5GAHD/4TqavmbF7/Bvt
hh9wuHlTCDqOoWgREcCvTIjXnuxTGdJYuWFWAkbRgPZHgAA6dGkVGrniLY5K7s0+NZbgjWCRjffL
+9TMHdrSMHihjV5ndOpg4BlapFW5jmmrHcTewUZNhMiZV1TYW9YwfZIUZMfjPqLzM14g6gImiQ6a
/SQUCP+gX/4wkh4wsxfQ1wS81c3e0Vdb4WFg90WLPrGll23jKaicimieYzrpV6Jp2me+smQf1n8x
HaImxmR4IZLarzZnLReo1Bl+VFOTJzfs4Li9dZ8h5ZpfCrOrQwvG18uGKNvG4t2WGAeZtvPqRlH9
uTN17XAfxVwMf26+cvVoFk/eqAfOJPXUkFmEjGfDDwUEEePI5uv3pAkML3TvbzpJRdrvfOhiF2Se
y5i51GIbKy0K3P8/9Jeb6gOa2Eg91Fz42SxrD2uUBA77NLsULKH44nSN9jmLQxN1jy/cPmTctzaB
iKhuvU6Q8Bfl+BbQ9x98ATbYknsGb0iqlfXs97Rz1F8mwJUXNmBaXiOXiAtkm8rpChoRL7HRUDYf
BsSnPjP8byxjr+/w4NNdC8p1uBTq/MKCOuL3oV+jP8RlxsNop/PGmaVAtDeuNGU5gY5i9oZJPT/q
rCZjA6LRGkJBHkw/AyEuVrkEWGk91lYpxXle3eqQN0PdI+1iZPXMaFMt34WEKWrUai9i494AN35D
P8CsYDCWb4Ni1se3c2mnlIrvj7RR6cTae1Amq2IFKdpSdpmdmPj8aD9X8bCKzBOxMZ4jJfaQam/o
xJaFNDKM8jFXm6OUuXK8r9S+suNwsYe55KRg0jeQPwBFiihi60m//4AUfbnq1J6Clj5YiBX/pszL
J2eMtP5VLFQPX5i8tWc0usw9Vw8/wn/BhvSC87dW4BvUt+lTvuo82JxJRLYatTH7/EK/ztyAM9G2
8jesshuivTUGQupmmz2YaqkBQOqXfErHtm9/ngN4eltxVAUAJL3IuQMP1WFW8OCkvpyVLuh/hv0M
YBn9DyGPkeWhqJ6VCxAuA6xDGT4ObVDHfRnSjqY+A8z11Ic42FUdxZGq9qdOf6pIySFtf1VytaA4
22ZtrR1qheDPxwSvwPRRJYOfeGARHimRDVDPpb/HXwJ5Fl8YanW2S7kf7iiLOOjyplIPWek59qQk
eiZJ/wOxnLdE7ci/JycgNyg6taCQwynuX8ybz5z39h0lpk5RAzvobcAcWEvWsyNwrKGrbhJmsFdr
V/NsJBsSu67nlrfirInBlR+peJ4tJM0U/7tMCAaNTMGzDGIhCQ5DalrCYcB/xFQDeiZ4wl/dwJwB
qqBr5zMxGfpy7laqqJRYvs0V6ktz3TLE3580marzKQgyO+LROJSQVUVT6fPc4SERjACzIhvOH/cp
h4i3cYyla8G+Y+WbqCc8XAPQHC9TgFYYQQwV0nb2Ixc18EsS74ulPqdLV8RwBxQqewY6PGH0RNiH
/W8Fw1giUGNcchuKQcDSYiPclZYfKQnUnA77nTHNVYXBkYoPLcEcuMrevC5MyPhW4s1sBkfFpxGC
iLYYF/K9JwaarSRhFVDatlXABzdD0mvFp2Z1Ojn9PzErLe40BrVlNKpxUBRRaUdgb1R0+Mfk2LHO
317CmMmH/Y3doKvmwwvlqyrB4MBzVK/VtK4g7lbCYntL94WRvb5G037+0Z09Uvbci9LNH6UbfsBu
twSXf7iZCwbQZFEpkOBPg5BKOPxt4a5VK3zEvdTriG4aRGIZKCj8IJ3UsIC7Kru473kqaqI75M4I
q/ubM/Op6F/dVkugaakX99yeV2JsmWN7AAmRrF5W7JiFgUDiTPgVpmxOeIilV7PxWMHa8HPmeVST
fH015CB4UHcblEM51p0dzRmAVbfATpUgIzBSgqgibhCUppQwPa/TrraW9eSfPMyRcNUfegq3dS27
9YrvHdU2aoAvLuUpXrbOwewxaCztcypP1SpCvEk4dAFomeX6DAXUpP73wrp9rKSLS+IYw7+72T/e
cBhLbcYDXbbf26eZx3sTRQTJM5sVfJW8fnrHm7C1QEggaHn08wZ+wnDlPWwLUCIZXL0Htz8qWXqh
WB2EkmOvJWTUiNzsDS8/95fFKWaCzFkresOLvkyYTOuQVx12H265QnWXrOwZrnDjxYLRGzAWElQH
qnzU9zWnvkTgaP7VDxUUqFBDZ3/+esternjc+VUziAUGwc8nHDTcYWe+dIEpO6vHrz8hQFmK9HUQ
U5Et3kueTtviGiVx8pIploGW4iGQgz7ovx1xZLbF0NfbLGK3Ca9Wd7hQ93tgCyvqdf+yCBzz4D7w
DTAEYGUbdrjNzfwpIQN4lROvSs9ONnIP3ZrH9PUZ2NWoB+kY2sV4Zny2/KxF9SKi8BpR664XUkje
TFHQJ4QHtlxqg3qnydCVD8OAsZpTUwW2ndgLT80KEpN4acYPWOrUUii07mtH/ASBZsnNSm0paULV
nz09tkt7msuzXsAlOsEO+owelXjZwiHV+svPmtjRfp9Fzk6gpDSLz99GWqHIXp/yGHT2sRNul/X8
CsSEDPdQ7hAJqfuVuiHnmc6gA/0FaVc/PzGT5Q9yjeNGKtAaS8pRuinY3jci5fBXan4No9Y8JW5w
2MU7f/NBfonInQRVXjK6jnnow5I01WflugBr7d2QiGmW+R4xU9PzENfrjx/iUOgvenHC7042uOW/
drQVBvuHJWUO3OeJxExUhoRZYUWvNVmvLTR2cvLTy/MGNNMUGV/9hUFDi2MLIQqx1Q4Hm76EwMbS
EuIQAIvIup/LqQLUtp5ke8bya7Z/rsfnEYWckzE4AxHcIchp/7K8t3+HyGxLbzYaOenf7jDm20Kc
+ZUt/A6F03lhwRyD+Cz023lvmfuPfmIxplmyi9QUyKL5MlMOZaKqBhuafR34ZOqR78GE7WN+o3am
XxZUXrqcU3B8hhcclxn69Fr0KfB08wNXOzV5ecZLGfNjuclrrY56y7kmhG405dhR502wp/IBr0Vm
ZfCxCEUr34Otrf9zkbfoQzAV+vggIuM/Die/Vm8hyNKcudRkCRLnhiFwp9YQ86Quw3/BTWjRP/VZ
iJqW2oG+rNcX+lbpY17nrDEpQqbArs2tKfFS4DG6tF2KGZRnv0t8l9tmIgyMByCzoanx4KfMUzAE
7UH7/3d46w5uzVL6Sgo7yuQDFZMUM6yoYxsvV7dYINwQ/zPsOQG/aF/ra9vmhbaHFZ+UWtvUS4Zi
LQUGXSVVeNZpo7E+SeZrKHKZQovvXxWUqi3jsq96/Ppboo7Upt3i+TIUxcuM0dPSeiwTJlVf9XtU
zeYoihsxqq+VlriKBV9rt8KYx5MX9zAQxWDJ7JDGz/pOuEXh8T381NJd8os7drg4Oooupf3R9uG6
mgAicR9Kvuqt514mAUBnstYInChss6V8fYjlgReaCaMcKYiPoOiKvfDOgZ/EP8RjHk1BKrl1J6JP
bI0uxWV9C5g16UFjxtP2WyKtLM5BaXdcTEEd4LDEhwbLcI3ItYWit1LYR1BQPw1K77mQyvrBJui2
y2VyURXDuB+aeXqpOTLFrS+JcKv2NETZIK7hTh1YH2zI2YR/EaDwwukDtlACr6PlxNaXyjFRzbjh
16zKjxZs6uUFeNpLmedv/wBsD5+paqL8V5CD1eLiZS9BPZxSRpPTiZl4U6WjXJTk+97Wc7x6lTYa
zAyVZY0+8PWnxfiGLHcNPzXQ13I0G09iGpkyHrByIGsrafva+U+Bot2fYLGThNUpk8xjet/2A0lP
xFk20PxeG26mEHtWdUO5vpgUaBdF16O9qU/ZA7xmdEJWP3Y1xM33jkG8mx1OYLC4JL4QMRT4czdM
Ojdlt8USIPr8+kS4s1OwzUosyzleCDCkydAVjeIvDXeTlw6m1MKN7/WEtHc64nSdiq4BgRC0z960
myjnOsTXzufo6UwdvqG19z3QXljUHSEiDmOmOmO8mqKrg09+BRgcDm3aIQrQ7q+LIpdOVsm8Vxop
XWW7DaHzChZn3p4+1hzBm7cXABwP2W2rPB/CSukWBY35PEKidAm0aFpPIcdDW1rReex/3MJCL219
SyCm9to5r+MgYQL9R4DYrYbKnv8/bAuy1vJ76R1JE06OUcwQekY+yQPa89MGipnfi4joiz81/6y0
2yrA+LHCOljZt4PGv/kUus1s3HztRdLxyPXG4QAYP+EtcR6QaFWarmtjayQ+hxWL4ee19atkP31b
MAWO3Z2ApIAU297iqrZtao/Uxb80pag0sdWNIG9dcARJjKJrHEb9jnFNagNfBf7YBrYmgvBY6603
mSqIhLd5j7yCrEJjQBFe+OrmnmMaY+2Nd62Sr+wKN0wn7h90ly97tKtZSPWD61mH0OYlw+cStGVf
py7Wsinh1PIMduJwhgs/btJtFJT+DGHpJYuzrCGTWKAvuydrybtO/lOgJ/vY0ES2RMw3Vxh7W3Rv
zqK8tuE2CWIZPExFqEez0zOkL2kQiQsZP3NSH39jiVi0qQ1GnzlD9J/ri5yC/Y3acYHpEMhPxjN2
g91HqtbXB1dwfZQOP052V6VmO5vp8gUvBoxAYgY6EkxqfwH7LVOuY+ixGl/KrWaFx5zSeBOBNAdl
OmiFPdhNpdK/2yEgW7ItlEUsQrDCRq8wYMcezKqPMZpyfLwRiNy1eH4ggtGXPmCz4TubDluxDVNA
GYeylexvognoJUKI1Dqsz4HuTEChcBdZphW3C0901nRfX4slU13Gun8z49knI8VrzhQz8vLKSOcW
8v/2BrWGzSRFTjHAORDt2Ew4CHPaRaucfXp2NOLb1SaLJhYguQykp5BWQk52DeyA+8WYtLEMbXxT
g6xQfXt5QZ6ZBFyYu83yJcIgMb8GnPW3dy4HepCx5uBXpMX0GeERpttFfpTblJtv0wmMGfJlkUIP
m7/ypKXtRD6L8FztESyvFs97FjHoKiwIiqtDAjlUWWfF4Gb62Itm6rjj581d2MSwEdaKvLuvvCv+
ACmIMDpDHF0OrWYGaFMAbOnWxbzaCCr/24hJk73OiABVsSaGIziRY7xsegdGvJdZZjgKuOqiqkGF
0mdGI736FE+k5o+5oxRKFhv3POoeuGJJwVlGdVbQQdcAp1Jo0/AEAvcCMY7c5j/ezBoY4b1r8NQt
SJyc8UL7NmkfmJHq2V9sYbKNdyJFGOnXwH9TgEiRLVO2EHp3OOOgYzbg8EBNgizA9a7vSRimLbit
Fk6+3K+cQW/3kCZY4EcGVarUqMeNXtcmjlLVGPWVbxPXwky/rKJqh6pzugbsoi3cbBrVrN6c7Bab
Td3H3hunxRnaa79WK/BMgXF9QwnWxu+dgEeiYVP6w0YVd2G9jARDsueJmUhIloJpT3HvgRV4O2X+
uvLQVN25A+sMVqcz9RB0qEAa2OIOpQ4+FPtQfwyG/W9/Xj6XtfYMhHQ3lbZ2p24z4LDqgcY+3ctr
RC/mZtDmsvZ3/AQRyMnfVU2Yh2E1zsH5V2TEEean38gCvBtXwTT003ZOk8/tufuPb76KvM+dRwfq
6cUOjM8KYYmPdmuSpSooYR4dy3v3FggdrU1PSro0G7tl99hiHIWp3Q64O8Dzank4oTLt0JyHQtFd
VJjwo71SnY5ZnUSWA+WG69V37Qm6GcE0b0hb9gSkqrnhszP5yystnk5UqXFNWI11mvrKhpmQrhI+
292Y2GuUBgzRGDUqyeWt4Gg2UIFgKpP3+SEgLqv49vS+uxesj5YpZM4bBAef1hqOL0VaHAN50JkQ
BIJ45xmy0KzVakiyUgZR/NjdT5EY9jy2E6lB9uL9sjo6r+TxSh1rag+WdY3A5T2/Yd7ocwold8Sg
YpA2bf8w1dZAjmooPCo9RXG23uOBTgJWuzIJKQnuPb2Sr9EFI9jSzzvEeXOzEokTtrYOCXHhSw8q
ezGPfHjbCRYPpA4GQwZpLxZa0rzKJUCE+tN3MoBQn59yRClH8DYRJmLlApwk4DUYFxY7pJBMyFhj
1CRB4Q0uzhw+sZyIozwsUGnsSoWUiRHHgZQOG5fjn/C3Tmv8o4KdDnl1kuI8Xa4dlv2Q0d0NsC4Y
lhllZ+p3YTv0pD/4ObgOq87epUBYEurzht9J2Pu6ThGq8WjwbsEtcpC7824chG1QoyzDCcA80JQv
xHILwAV/I8W7uOw9wGkucMS1WpjBvKY/9FJAXTtmucV+JEnbKwBiKLrzG3EeHG0yRq1Ds7HVIAcB
PV3qNMC2vJP+d6lFoYjUJI732nB4IHxPtY9WSOxzDDP6U6vVckrzu0mEcZY3SjfFpmuGlbaPlCe1
hBGu21n1ToWEh0+mavl9OpsMaFeW6KrVoI/PxJHoNsR+vJtTUDfJD9Gz0c9Gw5wXai83qUEbgzhn
+AzIISkXf8vxTUIhwjAudgH9qqxYH7odNCdllizZ4LubwuSXnawDZBQhs+K3ILsRp7ZwgKqEXBr5
7euNF2S9s3BG7pn59vCPZI+/T3OzHF6mgUxZIs9AIJISTLI76d6I9dbYC9JOQfhUpKj2aANVLDk+
tucwyYtKYlVmIXTXncV4coIWZhHsw5372vtl8hik388Ys6vcr+jVB3MgVBv3xSsKZEQqC9FwawYu
ShnZbb+mAzrDn4WjtnSJuxB3RL1K62Zb/EvDNVRyWJlAvRmh5YoidD5upD2+C7ZfVoLqJFqgGjT0
N5U4zqnUZGnYdlgkT7T6EHqPZSDkEcrG6+D8iPrfOdOHyU0XHItcwyhUQViqQ1R228FX3DpinGu+
cpaSman67ufBvQ9QLOE2vgM/5bYjRYrgpiwxCZN4sX14LTaVwvjoRYYW8iR+7TMkD0XZpybP5AFX
tP458sUC0qDWRg113+oPLieCrjABE5G1b7ncINNQBKJA8trfOWrld9zfyCRfRV8yRxD8f0s0sQGI
kEuT1kAeUWwHTWmUnF5ZWCN1WETUO40q2ET8t+cqe0OztTz8SxD8zloTUvOnwBVWqt2xYn5I1TuM
4Lyo3vUDbXNkZU981wF1I/7nSto5Q21N3AvK8UnBea2b0KRA3lS2Ejtj7Ct4gNz4wmuEyQSMKp+E
6thVDq6s8nB/7rWYGj/ZdZx4zl1Vqwd4ycPq/yRhBdGIMl+cKfKbUT+6SFQcnvEs3cka4szeb2SK
axDRiGKc0AQ5SN10KENHjW7ySng3ni0/cJBx5hoGywZF0u7vTEknkBDifNuhofxYymrqXfYxnxvE
p3cstxYJWelD1ioafYzFPBGGWVWWF6Ry4JynjSN1hQ9nrrz7TjNWAp6ASya+beWbnvydNEShSjTk
ZRLhp6/esPbE2WFi7U09gh5+p8ebu6rN2bDSZKgCv9b2GYKsoLUMbZ/Cp/3RSblmjFuqcdD0Chxw
ehnTIvTRMAE4gCj0ZUryAX2+/o4cqaKJLrpuxQKT2J61A4/L8XSTl+Luk6J4QLPPAhsjNNgPj2sJ
OJFJJJST829FCB0M/U0HEQG8DgJKCc1H5ut0rTVn0/OItUWSqilDDqBvIPGttxbuRW6YSkHVZCAu
uuJDaHUC4PL78Im5h8wfOSIknn9kmCU+kttFtiVBkaYqzgkylqGG71CXvbp/KQnxownfRCRR6wJo
ydcI1LxcsxCRBmZOkpmzXwtzXX51dHgBscOCIeLb2fvYu4wuAb8xOK8850T4flmABJkjTVVNS3wG
++lBqdFqQ5+9NZsKtFeSmAd26kxNPysW5rQXSn82bs/4FoshDRo0QvI8tKyydZg/vS8n28wYOHAL
PxQAi2vAZiVUOxVArw/n/dGbjAqCLCjZafwGcJ0JY96Nee1pPcrD+Q0bxxLqYYZD7fAoCPNboM0u
PnQF3np/jx9I4RlA5Vcqbr2rvhjslaEnOaJds0xeZ0SDnuw0ZLJnC5Y7OiqWi7vLhbn3UGfU6Vuk
aqyDolg/CeYvIAjKHwKAC3yqNQQQ2mLwaeqwzWq6W3vhV0EWcUItM28zw8p61lflxBV70DFtoRU1
mZN4sfKK8Nzev3xmpIJHDvcrmd9Vi/iZzaAwTEldxK6R33xkIHae/ZagEmO5jHVgjEvbulTRyjuQ
5BwnnsaxSCZv0VdHpUH8RmVkzWJOzzffgaQeY3xZbW+y40M6g+9MOO5TEpAPiyYDCJusAL4qoCu+
gprGy01pZaKPgjoEVRYiva4uzH00Kosky+7RbqHMUru4hmUBNBNtCNpf57Isr0R9cji28DDXKRzl
E+F+azofJFCRiFEDZC5iw//bvNXp/OriOaF4rXHgbNe1spXjQa4kPmDaC3TgWwa/AEUNussz11MI
kwyk0vpukAwy549XPlv/khw2IvP8Tir2tZZBEfE5O/M7KJIMY4w/lzOqD49owxNqwGq8dthv12Vl
iPwTdVDFgOm2nfOMSIrMyE/YhhXzubGQDp0an6HhLcMurxJP1PxI/FplqBXdUdoMgZVFsTWJixnL
LupcIFQ2EWcdEO2OhXE5f6f5pp0ZNCP5YHoHtLWZkkhdPLY2MU8LhXJvqgukQd9Lhj0GEg8OIgi8
OhaSOrA6WJcdVWrRDaUfF2iClUKDUHpwh1CFcE/aU3/QH3aWmhqwTedHewpBhLtEoGiMNqDuaieL
zLgwSwlKeTHOgcyQoAgomoVvmCeu2InydvwNpFw5ZaSUQ7rbHa8mHB6MzolUhzfSaK8xGNKkZ9I4
d91YyqNa2wym9g5xbFi6/Q64Y600g6V+qIz3rw+xuA3MJD8gU+q3cwbi7UxLoydaWbQnmlovC8ar
+UWqBF0mMcZxWKXZYGBph0+3gcOvCS5/DF/QQ26WCPgDMLqRZutw1DAvSz3N697PP6zKr3Mb0oBP
QrAYawGwzuMD6ESYuSkBsRuGe0zbFWCNfLyG7TXs48fma/PX9zxslzvvD1VRZC0Qiytr63sVAKeK
0FB5rAn0+paqtJwal2BL7gXXE9exqbb4T2RYn4EttHyIErU6gZl/yqDqG26DOIY1OXuTOxJHo0jJ
79vATxipPx/BOwIBBSgb9WN0IVTGQXG897E+rtxolJm+aVMBLXeIC27LvLxz9APIvOv3anBomHng
c5ESDnaJXuCOXMATlloK3boWsDETHAJFn/04mtdKO9/o2+hxsuAldu8Wu5UPZzMYBq7K06dlJ6nY
3KISW7Bh5iDiySsOATh/fDCNglJDIbXpt7NX6HYOAaOKq+Z9NMDTfzKpJcmNHyvO7UMczBnUXxZh
SWFgCcQPhuLEVFTgBM27785v+FI4XRKzCal6vPNzxB4mJJgZITxJQS/1UOjKdr/FBOciiIYFQWBR
7wBVE74mI73GbsUOOSx5l+W/XymjUP6sYQkLv+VwZghlMj2RX1LPT7FA/KHXPuLmQQiKjrNHnf6k
Pp0iJfem7Wc0I5AwVkzywMGD1qm4gKSGnV8Mr2N6mcti25eNlxnnVgAeBLm/TaXB8yfvU6Sxa2/g
WDQWoYPlvFzr6D7OoAfGqUw23wS4RsZzbdJcdVebwK+QZ7yXbTIM4pQoyg7jdYvkJLuxD+vgJHbt
pIxcvd+NBFNsufS5+wIKW44AaojaN0pufUP998CcHLHFDGcaMx+EYFuxgJcPrdiNWcaW+ap0/UXc
/k3PwsvxbNo7yrMjm7Eo8Ztuie3kv/ub0V14K6uCRZHK4deuoPmYQ1V3mTV+QpHDzEQEeNQnmZkN
7R7ZNRn1GCiJdpyAsBOffO8321GdBuIGnOMVpAMGqBS+dbvd/Vr6cHiLWIDtoD88kJ6TERQiB2qU
143jP0ZUpiaSdPpTPWMm59l+Rw3gekSJanbnT2zJAU4Zlp09PJ5faSlZ8uC1skL3hKfBlyq2Br5H
EV30ddKwf7S1cOXLx2UuiLDWaHL/myOkN6UBu55c7Fcqre3optwL3Lq2OqwLfzY0+6vyVDcgvTE6
s2FvswG+xffW8HnPlrpUYJApMgHsAssRX8TY8B8NZr7gWfaN1+tH53Mf2B/II95LqM5USRj0wjlm
//CtYuf5yfSrWQDi9YQeIr3AuHyuDBFNZ7CYuzQsJLVslHv2tZFXfuJFgdBeXN3k1PGx6RHT8sx7
1hH3W410ijpkRlNbnUsJTCnSLqpc8PLLETI88Ajvi6slOonhmoPEJjDa2QuJnHb3hdSSuH3FD0X7
JlgUynOmWNdkYCzpZj7vDiDeygGp5f1cWSbbZA76ZP2DOZowUA2WhQv/H+ybJL3nxj4r3ZGTbJ3R
i2Q9d3pQfSRqsNGXxV2I7z3iJkfgDxSOmrQ7hH4ZjCkLs+hfW8qtRYQE0pzfaM9VV0eO+Vqre2M5
zwAMvUrvu53IUnunBmDc5W11VdLR5Zx4KB23Bo2M32SyGjw9vosz+qKP60oXBxLeSxo51qxwJBcH
8tGuXAhNtD9mqCQVqAT1X6RF/cN7r50vdJ0K+thK7QDxYnAD9iJBsfBq93pZjQrf2qo9N+CxHTtU
B0Enhs861dOMHmmBIFN2PFp2Z4tvZ9jySo8XJYoMae5qUtPJHPRgvOBcEGlT4VgInFW//52iofSJ
UTJ3IFsFMCl0l1jdblUs1VhMaAGR0BzwFjJWsuK+Yh+jazTG6iX33HaQ+adQ1kWILnCVZ8BNpLda
AP7hSF5LNITa8HttoN8bH8vGPV3va9+b0s4jtKKO//N3vOO0M+2JM+lvZjQuT8gThmm3vs2C0rcg
mpIK8ISygOTkU7kl+6vXcmT0ISK2sQ5s3oDhKUDfKdD6ZUNEE2u7KH1f/HJUH1nrYv523Sfe1Bv8
xzLfVBWaHOAMlfNPu0DFBj7l559LJTZHRPJ8euKkkvXSWSqJSohmdbTSJC+JvD2qAUTcrhc85MNg
kaUiLSnSv1WB4XeTqbrIpcOR2hHh+ncoMi6cMHuu/ST5GTKqR2LheAJmdlCQxtcF2p7HGjZP3qkH
YotYiGJe/TyFnYHIxj+VPirzO3knPbBxUYrcKnAeJRdw1iEWg9cTYVTkUCJ6E1Y0SfQhZOtloBj3
Bwvurk6CZBAjUmijDm7b7KpzlWePCjHCgpPCKrzBy1XHXXtMPJ2DKzvZf+y8Mx7qt/JBdXh6bpBr
IRWdujVywt6TSBgH0kaXM3ngCey4La94/jMVzBDvfHaysXGXE6DrCFaXYIlGidFkMlnKhdX69Zm7
xHy9mPkichSbDiCEwRBvrcTz/U+Y5P0Zt84b7HP1cHvJ0k2O6EGwPaMmcOw6cnQwtMmSNbjjdDBJ
+E5IRuzIRi6YSOKOof3lQB6hSZDYjeOudiGR82WFjuQ+AhZLxNhXWoBPlBLU/PX921dLupyJrejW
Z5wcq92la6BFYZyIeTnanBzb0axBVP9X7Lg+S8qX1jm3poSUYCBSkoTTCQ6dCulFb/NDA0W+IFa/
Kg3IEqPnYYoGBfAwT63b9MNQlIaADQJV6ND3hGU4tZ8j63x5tb0wWLvbj/y7Nx9daHBMpYyzm37Q
qNj+5QvGuZlwkd0JAGeEX1CfsE1M78+MWGm8Mftc2zroH361M0zryuU2oXuNb3Sgg9ZHKGs6BLsm
CxlcD4ME5rI943mRbPE0UZqwW/fFmnU5BiFAs3oiMlrKlsuik739WqayO2SH9Tg9JRUPjvYNyJKZ
YFe2xLQe2q8+/+qeAIEhCjmgnFrNs54YxHcOZZmjBwlQ5QIuLK4q4zUQuKcAR4FM0xyijSTlgull
Fs+kvBOlgMjEj/gkX5raR0aZg9SzEFECrLqO23ICvuCO2zqjWEcIJHcoUcQmzYEpXMSLCkd7jXfW
DFZ/UXA2yo1OJznvGm5HEp/8XrP+Z+02P3UFn/zuv4ULBEafPI6cIAwLfRBz0MAWkIy8iOGEJv6Z
0WVItUX2uVinOWG26tCW0jN6tXRi8R+YDmSvAyokEqiMt0v0HNgmpWiM8+padyOwBeXHdAs/Qfnh
qj0TQciepeHvL4sbxYATJxQFLFKTYyn+SSwv9oiTDIb09Wd2Mzvwc2htif+3xu8c/LYI78AVqqyT
fBgJSLUEHXHapwKK+H14PnKlDn0/h/be8H9sZgvlbnjWXUP8V/u+gfRzziC6hHX7beBiVodiCVEF
j31P7y3rCHfFoKmp/BGr4RenSNCO15rEXOBHIybF18/nmSCDSabkOgqmIjDzbLmen65uYYjN/dQ5
KIumKnlzyYsSScyfC3cxA9RW89yccmMQTtyuYm8mYxPt9122dT97bOWE/3QZ3uRFQXb/UJ47Uk5O
jPpzhINwfc7cKcS5yN1RfXnv7tmV4bVpjH8Y3+9UxjcQ/sX5sRo+2PIKYuCjqHRWMbkg1fIVaIwN
RjEEh8NVqglHaTNRFteptd1/hn4pIORP00QRZI6KlzBiOosLYiYtH0zRERSoTTbvvQFjX6eEO5tt
vvzF2uFff2a57+tlcdcSFSyBtWlvFzkOo1q/PZzCa5+0JH5JwoMVMSjX69JXvLFK+VYVzz4aAQ72
JnIldlu+3ls46Ya31aUjEPZxun3dSxxWSKxmCvsxpgfmcEWAuxN6SGIvd2PDbeBNrZpuJjmfEpZu
VUShK9D0x9ncAa+07R84yMMWtet7P3ssAxpGZYycUnZ7eksu+FNooqYUACH7BAkp3Ge3O1d73Ajm
CUpUzNv9tiR1kcBXvDXHRbcZ+aRDCYNW++44gU/AuX5AlXwmd4J2xlgIXFtLfsSeulMqBvBMZhQL
Uc9HfudrY1xTPAaG44ZbdzW1wPZtTS36XVxjJp14jJjgmjJaabRC8pwwNpQueh7gTpu4owqaqV2c
Tk0uBJ87mANbCPjT8muBLIaFLJ967BEqeV3Xf+SKxyQGP6EH9u+HM1AxlfkCbqAhMAqa/vIl9qKd
+ckLVCoTpvN2lCVeQe+e/Av57QRRjQQV9NFvgILFGgd4jdIQs+frM2X0Lc90gJz51NqBeXk3frp1
pl00qEV99o9hUia1xqx8UuDvI3iU0L/19L3hrjDTz4hHrn6bsoQYiooDGjYcQ26Nn3zsEZL+98sz
Xm9qt14omPeZw6VZP/2DWK2kYvC9KoVWNQU0h3xuDLMjr7ftOuu4V79zKTb0L6ffDQIBiPfJT4gG
rKUZ3dLOp69tF1NB0+M+yDsbec8wSAYruHtReNBQnvjUGqckDewlF8jynwRBikYq1+91lLKeCm0U
ZgfBAXaJRHYvAI3V9NVUODb5hB3HJYtYfgq0iLm5dMZ3ki9pG2htLQFegpxoiCRk9dXVNSr70OZd
e25N5x+/AYlhAZmraC8Rm3BxIbu32+zzCfCvbVdmvV4BVOifGkYcvS+/RRgl+SCoKKcZVuJ6iYHs
sttsfRbRvffUVDZ5Vs7IwyoPCuPdrx5njnmjKNult5ha7/vStGm3KOiMHUCl0GhzfT+3jIW9X5fR
dUAF3SLoEEhtwCwVKcvhxRQY11yr2/JecNX9lfsw9C/uLxMD4t3ARr4yOlNockZyH2XEjrnF63qf
B02ifVmP3mDZ4R6gT20qKo1Hm5PvOSvL1GC4uBmGbSr01MYpcMB2J3LL+YW2YKd14oUrHdgUgGDA
Dyquf/H/U2pk2+FbU44ECCXoOJqCTQ8oftgdi7/BBV8D3G9qax+7y8rCAi/1tFjkZltwB3HEOOX1
jqLyLjcJQZTdwcccBsg9PEGAYvowacgXDTrVuaHVIuDQNGFb+lU8VMCMq4EFbKIgma104QybcKmN
i4pb2RxZ3qr1Xwa71VWK2r5oMkqK2/inDEZLrHr/fGsJUWxc91iTSgC1UsIM+1Gf+GZShnC5FfoJ
RGjwBK4VdbtmRRYgxtq+Peen8lIvbgK4fOu0bSbBzTzrkNyQFk2SO/fSXSHKaIvSz5VrIHc6FX/m
rBRSTbO3MQc2xgvkJw2zQm0uJbuvaoIlXPlr6rPQmEeP6PeN8Z+08E7+UnwCf/Ci2syslKCAq8oZ
MfYcibIEh/5vhokJkgIBGYid2VcOHipxkFv6Xux35d5x6hncmxPFkKm5D4ny+W9WLlFp6tn/TfTL
VqqDwSxoWvcqUZKMFvOBqdgmz6t+xSbm1LvDkrXtb6BH3zFFiUThn9r3Cn3Qpg0b1nwfnvM6ihQ+
27ZHVakJ2vGILQCVUSxQTNJDyRPwJmdAM9KxB+opI3+OYOMe6eb4ZTm2fbaS0PO8A9Ncq4Ask75t
4aXQ4oNX44KPpGSXoDO4wLqKCA9d9r1XPb+sqsjZ1d3/wxsAsLPwuCMDtj17PyZvdeOs6vxegVZe
dPY5nbd0/EIrihyj73m++e89UURw0FQogaFb0nOAcHzKYhQ5pGU4UUm+ypslKU+Jyx5GAPZgs773
AGcdFm6cIA25jchRt4SKir1jHOunb7SdeOdHRAATgIbmL2QCILtiIgRsiUECd/f+aqqbLl5sNr39
RiXhggsNWgTuS3pzeUlbWcaq6lDYIr8UnJSpwPmkNx68tPCJ9E8gGbamKZR49uBHVpTWg2fwCL/S
veKjxDr95nxsKgNlN/qc27BEL2MawRUw8qKhKQYXY0uwGqAdhmcUJSqibIgezK1zigvNrsC6th/h
1lgrmZirdCP284hH+VKDZuux7soIl8VVkNdqxsxNZbKQ2+XVM4qKsve1ey3YBY/qeB1Xnf17aD8/
QCjAFs+qE/itwQmzUtjyZQlEaq3EIpxz7HQpIF6oM1G+CjaL5I7PlkkggZ6aybLFjfvW+yJWhQ+G
q30d/9p+omxtUOaXvrZaEFc8KL/yJEfhrU4xGFr9t+no/Ro7OzSWzo/EKpGK3UlRxwAtqMRT0iqt
RKY7DTwA+AxlAvZqWzssTWOErTYg+BX0gQkTlr3GDsp+zHGgL4yI3RYNJfqxXp+3DOKsd6VmqQ9M
CjEjuMqKZPMEoQMFMteCTys6m4ptBucOEYUA97FEKp5XG7NZRaBVVDW3IOZacu39W53BiYOPEm0x
lMWWpDxC+Pwo/4yv8yTfMTPTmMAIfQsseEsz2vkUcNj57Wbv5Ke8oRhk0WcBygrGjLehpfHn/w0n
cDLvdg6G2p4nWxO0FZIb3X3cA+qqDxyXp9xq/loSEnzW6EgocdMpgwQAt4mkpdv0mcdon/VnSl5P
m5nHpmYykFiUFxolLKq3jgmuX1JZ088M5NuLPpaYyAxo3xqkyGvSf24PB4z2QMPeb/ILntOLmLUf
AVbcB5rrlNriEjT/Hra79r1u9HPpKSFKRGN+Zmym00NcFL6eGc9mtgLxkoswQRzn7+uubyq2eH+q
27BaA6tz3nRueixBWok0p9vLv8OBBn6BwUZtBLUVzHWjW2Dr47sZ6rU0JCzhS15C/RAwEvjZxSFt
o9vQnSK6vLr8NU3LxT8OJAAocEMd7zVVfjaGaUiX6uCe/jCw4cZhQFwx9xiSwSOflW7BI+F/ktbf
7Q0WFqYtniJHjQsL4yY2AZGzf9BOhI6tKkTRNF4L3SOlizNJ4CJ5YHrWPg04riNu08sCDWLVGBbZ
c2jirwEdVoR6uav3beAIwNXwlBIczRkzonP4HEiqQV6Sh9sp4bhUTDXK/7PQyF3cfhqWoIjS68Ad
ANglwQxJVzJf37coIwGYuXexZ5Gtw3pXf3ohpJSaWSlObhE6iMaAo9wpSjf8N64vpql9H2T2YQqf
vkRyanZRCXYNSoJU+YT+bnOsJ3bKxUjfndBqPpcyRPLRkSXXFPuKCzzBnJfbh37V+ZUQs4kGoAj1
PZbA+GoD67GVN3FYThXfFdUaD561NVKh5VtGqW/IU7ZZ9e0SeCk02tJM7BpvCngUINDm7LgXQQ+z
snCwtoOgrdRK2LF5SfoRdK0L2EdxiAJg9dUoB7bdZ2nqw2XwZq57WmgILLMFICaTIVGN40xuJHok
LlZAEzQpSGStk0Q+EctS/ssJqqEH5cL4jrvgq6V62Hr1Ny/gAbSagUzgt7WKBFAkzE+fUw2NstH+
nccJa46pSq6VeyOIMnOAynGLBZvajBF5izkDciHtoRWUIUO5RFUsJJ7nstJ1lEAaCVDIe3N3OBL/
agfyIKGtNq40X34u1ckEqBvQRkh/yI2bEvuiQpyTXTQYlSdKmZ0jS9tHhf4ZNCG/4h3MOOiOn0PZ
Px+HgSog2CZQf+OZZcZU1Ml5Nd2iS/mREPgGQHaOTpEcAORoniOlA5hFglL8ktCQP2pwjNMsLMV/
80M7FG/x8RAPbUKfFzMTHlSNGf5Mnrej0Wk7lVwJX7OWv5dpQ2TbEucchuqs0sX1je6JoDADefqS
Nelx99fGS9xj4BTKzRTKranFJBRgXq399HXsdznd3ndHFO/3arzskWrT6PGix3NcNwQ7L9ed/pgy
kggKGatBh5hezMAdZL3AdrwHKam0iojUJnIXZA3/VPmBuewYtiytQdOA3evxC8y6gYbZq7vdgZR0
GR7ziHntLyi7RHVh7RS/QWMlScbOq7LYLyVZZnB7bT42+30eikXngyxUeiGOJSeb9GhbO3qaftpC
iRauumAzEJiU+LckvwfS676YXzBdYdw5rzmk7zVJahJHsE7DGJvHNZK5BSVXYzkdO3e7s0FroM/q
TvFnZGz9jRH405RaYMxrvp4sulOFtSMgafjt4/2+/b8GB1POoeeZtfQqCB4JONdZh32S8hSPAI3c
Z7a0D7YB4pXYOhAqMpPlnNnfZJMvtpiDO8Lj+2IfOzkSaozh6ME81oY8qjW6bDS+ZaKVgjx3SQxv
//Q4rpxredXLl0FQTRDicg4GkN4tGnNtJI8OhQygbznxTQzOQ0IgQ7nlxlWRtm+4jr/BUL5qqflv
rdDOnmuXU5duWrRkkKafZvFgLuyBc+IssXlBNTFPVp0ouY99mpgzLLEuCirQp4pg3dqkdmma2UXH
sU4ZeFmftjL4xQ7mrpqiFnC6KxuXTcowoXxPz9EKnzijdpPabZGonwYBg8L4DXy67y2beSaXDADQ
mASvtM6XPJh4Osh1Zvr+pLhwB1+VGpZTbHfHqq47gDX4geptzISHONcsn3/juI8e58iZgkyw+yvx
ZPyGjJ8jhZPeTJn8l47HLH2E8RG5BIpSCp8tS1dubOZTznzMEs6JeovmdTchu0m+r8bzac/UtIbJ
cZ0CtAThQOc9zOdm8TpL9LxOQnI72AXrmIBAVih8LY7RkcCyqVeztzvlU00yEuxWXwSK9T1lK3mt
xkAQ+NQUKRCj15uRBOdN2FK1IclrLt9vsiWej2TRhK//SWPPwSQiUTW2Gu5S/GHHAKib1oO1Dtyf
Xh1/41zMAWSM+B86T+3OarP+BbuSOTFhptW/N96AKRk8ANNXtMcnyqmeyiw/rbPd0F/BT79fLe4J
HfBV68E5zs2rGEP2yeZ0lBZmED5QAEHFcuXAOi8M+xB17Y2C+k9w9BnPzTt0x3wtH4G3MHlRLHfr
LD0MWwfTS60y5OWp9PCM3RaSD7yZhvVDDQaXQFcGiBc2FC0kgObFDylPcnHDV1jg8A1yknv0FB5t
HF0zWE6jVMFJDJdcga9aGuzwuI+BgkW8Yp58FSnK4yDO2KRsu4u+xpGnSaoIXjpFBIxdF9Nmyqxn
hwmSJh5F7WkXPr2id+g1/tHn46Ev5aM88NmQRdwPQG2AEcN+DBLBeXMHPL3U+cVwmmQ9NKyTIN3E
iOjy7H749uav4fx67Fxl9QMvenqMSHHyZzayt2JghCJ5qU4GNNH6YRWuNA2bHkIf4tmb3G6wS99s
GNOpgh4Y6b/s9LhuqpWuzd1UiiLovyq9h6TQ9h9QwmWAyaDjrD96xqrfC3XnKAmyH9CYUbDObYf3
putqIEcaplzm9++Q5iTgeHyloyIGufP4HXYTWs1qmsAaDJ3uWt1CuPSspEkhVpI8e1XMa/FBb8SY
KUE2uBh8YFJoRQbECpUDWEFeFU1hkz3PEl2rT5dbpV8mo37lsCqUUXPKRD4EPDxybU7nUmo5agAf
QcTOSLt1YQD5LQ1/2ywNScGEnowIlWY3/Oit9FHdexqsbsHzfgTkHPnajQ7n9OSe7oGmkeEWbjZM
XE50XTFvNOSHj5VWdigqzPZU5isZsYrtPkELvlKhLDvUAaAj5SMDVReKkNozSCn1jRf5VFsBihzX
hzGWgCuF2V+9rlhblqil9YTw7UCY8KQu4yQLivoUcaFNUbmC+hCITvjjbmT46VStOfvwvNZLyxxR
qv4UL9Zh9LBGcib1yCLEnDszSkPkIjKZ1gaIbbJ4A2XCswmwW1jf74cYcWbOtKeDhbU2+FuKoxXV
v9fcdm9POhzIhe2EHs2LZdZUaSe1ezXwR1R5jMyG0Kf20Ka0KT7nvwWAFzQE8gsnDa41PeN/1zc0
ZmXE54ngT3ZbWP8cAJWjpiFAqKUg12BspZvupT555NUPOqidT7HWu0fafdzy/7v5eou8/A/fFD8b
w2wSkRrGm5+UCWp7VFOegrvnOSXOvNxF0qvWb4u0YrBHh10Fwuz7K0QiG4UDXk/EX2eZ/T0uF68i
r5R44ihmQc/TuhVmKQg9OEGGWGhIilWFJ3TGDzFzXWhvKnClOx+2ethXapBkjDObK/Dl6NSMyN/H
+MTsRo1wMquOpkgD642AK5BbMNdUk+y2692IL2BN5GeVebfjWlMKSJuzpLqft1mh3yKx5aGwTBzq
3yS1TznX1mY8mZEzI5oO7t9ax88vRyzDmVN2FPUK/8LE3yXQA/SERYpiBrP5Nq1FXu75BAGYMIkb
T0RwpPEhmUeyEAAD201Qlos0DqkgtYh85+8q4nIB4uqKo1vdIdTJ8Vm39F1hX8A/Jk3FP5Fcba5J
TWO4YIXVrRj9C16r7/Ohm9cjVR3onNR4wfw21Swzu6uWyt67zCUFtaAYfh0kqg0PdKVwA3PBm9kQ
usL1tZ7rmOduFYpcV9hPDmPpXPTxa2DMaEZ1wc5lo2R0uaOA0iK/FxJq8zbIWl8QE8w4XNbSBQpk
PPSsaRFjlujv3jjDSTkcSEemehvWQqCrKcXJGKzrCN1TK3rx3vtEgErsL1zwZwv0kQdiH12SSrgl
a13GO+Q+K4hI/i1Z1giZK4x6x8EgCjln5itNyI31oPi7RUwzzGmTlsvgcesy9aQZ9E1trvje2NwE
sz8k7I9ArYAbVyV28+97kkG3VLWkGKx5V00fDIVDIrFl+kXDOnXoyxx50iRlkREQyPhBpeBIOCGq
WneIVBTuxtrRL8NnAljB8Xu+NykNQgu+f8WcHeP6ivs1he2i8H9z67PI5VxvCM95tC5pDHaaxJC1
8eoAX8w+5Rd9XBBNYtJma2rMZMRvx8RBhmwAb5/9z1GY/581r+2kkhQlr4v4Jz6pQJ5yO/ZUbWxu
gll9cUXYj2liM/SK54CZxt6f3Yj4QIMQZ8vBq7gZ4JpFbc2ObOnbvU9LUum0qfMFeMQqsE0UI9t1
M80tgyLyQBsqEbtiJKNVQ6aZCxGNAvDzjg29lZamF1XVP6Y9Rmvn4pxfNISE/oVz5SCXz1EO/f73
kdJqHclOW47afy79b0OEb2osIphBu+9Xm1+Y0E5dhdqZ7le26ZjB9oGB6g3N82Ptd2ajG9293u0P
IVuiutq4ys+KBg1fqPrOutzWZHFaXZ+Zpzt5dT39xhIgksqlnI4BCpxlZ267u8g4WGsQuIrmz+IA
jrNDJmTcJpWHDm+qJ4Wb/XSb5NQR4YPTjCUj6XG5qSt5Wic9OYxFHWZRds0CoISb9sOmoEgKLLC2
IUa63K2wTeMW9Ab4cAjs2BS3CfKR+u7pYD7nF8pcA+8DD9YohOPZSQVNh2oy0LJs0gEVkErYHtjA
pfrMenKHM+igQXAouMfSVfbZsptLB1MAS+9A4qgALgWGAegitdP2W3P9m5drHPcj501p80pTQRPQ
Rt53yZhVMmIRElDFS9AzUU2+XuA4bHMhp2nU6uiie+rtbFVqaPQ7GByhrFxQJGUB0IJkB0LXsGWa
OEuRbBDWgJ829vU5Pf4fFdBCwnThuGc7MBZ9KOh9PHn0+2f04F6Rq3QUaKMJZjSMPGkhhsoSAz52
xXauyl6qdujq0BUnVCmvy1R93ziNSf8gLjKmjRtSNyHvxgYaNGh28+tgXKozEeU9jPdHs6deN2aO
aCsJOW1vHsV8FIQAPrlog/Jr5brQ9h5naZM+b+5ECGDZyXspJsBjKgHDYC/t+0Jx4RkZHtfSx7Fa
SYwJkfmPg3cN2tmpOnSR5tTJvFe9lojyDKqEULlVbDmjdafce3XIykywUfpjnFKtQfbIlGQ5gduf
XCVku7wo5EhY2Q/io/Cgqr9e50QmkYFbzBEWS0+cDTMrC/eoGezm9Xcubn12Xf+q4E0tGdFaepnP
credcnFVt7jdKexk/pemuX2ExPx7MjGwkyNugkmzq7OjR04kJePhEvzFAJp97UsKIGIZ2pZSjZbe
dux8bt7wdUHMSY1D7PNiTxwEuSLGt/97WGYTg8mdZvS9DUyh199sfYQtDZZK+rTVnZfY/x680fTg
iQc/Qhr0HZ6Jct7ohmS5p6QSBBWWCrJPTcgUq53Y+Lq4YLeWipd4f4wcgQhTvVprSh9O+jReKMDv
WYBUclG+zYTukYmMzqFGtvOvxRl1S+PBJh6yQpL4hC8Ha5G2lltH0l9stcDYfNi0l/Fkgtp0MRsK
PU1qbIU7mehrFWdU998u7CKeDL720RktbrAWyLfBDsRJdfHfvDDRWIxBRkxrq3sgVh+yuNMKEbrv
7KHV4bPHrW65cZ11EnnTdlDuaWgX/A4fLrEJhU+AfcpnNFbbLf/Hgr/L+p9MwxP1ehz/ccE5uU3Y
vy50Mje8UEkYjpRPDmC9Bkj9gcivJgP/rerkx3G/HqQOPfZbzGUb2QWbb4rk1MX44oT8PpD69G5z
kOVaZWl2HTRgKUwVHfALWvZ9xbgdcCw5CH5PMU4/QBQDFBaBxdTman91DThgJD3NYzsjDhDZXUtZ
lRrQGRZ3fc5zK8vhyaW1FwGOFbCKeok19bYh3nzD+r1u/DK7P12wvUMVAAHjcKTHmlaUQS8Iau5L
o9bskaKuDSuavWo+Hlr2Xw9FlajrswumeUSaQqQMV7h32PB6dObIh/onSMk+j9qpizRE0p1KeAL8
iYeIRJxqc9cFcjQMaLDFqMOF0YhNJX76/NOm6pcJNNxW/mRgJwkFqMl30tK12DeXy+Q6wY0f3mAA
vWm5hQqJsnE2OUXyuuUPnEXkqSdOzMUMlAJHVyvNaPpDv240tCMvoeQpbbO90PHaA2s4qkl9RN6F
Ccqion70LuPH9c28xWlsJ+i7HLkAMpA6EVFR8CLNvZPnnrFaohyZXGChbINEoYNsnspwFcpUr/26
M88iQV7f9cnUI9fvFBxBppmpHc6tan5f022xgta3sdCLTjL5zS5qYt0Ks17rFCJc63uFCRPk+Ec7
Ej6jwUOjLN/Yxf+Sas84cArdIZDIf9LYhGFrZALbFhrRkZAfnRoDuaZ+G3g7p4ea3H0nMQ+UeKic
CkohEFbRCRYEO8STZoSOdnLUsuDJaaJvpx34/HmwLS/Fwflu9ujVLCPpHa00XRsiY1Kg18HAmppb
TMYRxLXRHOdolVWqbzC3A+1DeUhZK4u3wndNfBiXjET/euP4zzMbIs6BynQq54dm+97O5d68vgcz
dD+HOHUZE6GE6JB+qGbYlKt2j7J/+0SeUxR4WKt30ruas/L312An8v/fXBpwSb7VVXKDEs+DGrrI
JojX8MaYrAEveAmQNqJT8XxtuR3bZeaXOWZmdgqIByzbGgtT0STMIDtLcGJSAAPrgS3aqSjhkzJC
QVz0nl6jjez5QTOlZHP9WvV+Ea7KZdwynp8zm/BP/MbuXarAeIsowrp+ZJ6kIJNCbj4t05922xS9
3Ly7qIEWv956a5nnthVQrOiS8V2raDtzGBJgwM8xpjxd/ItW0O8RiKMAz/58E2uUb71wnpk3TrtK
jg98iwXWipt08rqjS53qU06uaRxoEugLuJf0gyGUxT/HuwTPX5TD14xXKrIb8I4WtZe2H+tyqWZa
H5eUC1VICqYnG69LBTw7lcWsIUlVzeHAu1lOwTn84FdhW+BGpeD/AjuvSyqFy/nAneXKhZvfyRIk
dHcpDSyp321w+T5OZggeSt8OeDekhes0SEdfZg7P8zoAnubzccyCsA29YzVsoXdLsZXjQjCSyLCV
EqWiihJUD6TEKYnohCxEy/dHK3QJhDE5Jb/XByPeY8rkvNMRf1zcU5CSI1aY49abub1RYP6m6iMs
u2ZB6GKLV7HgWxhxyihyPJ5y5XnLMtmj//HYV27SO6pTerwsQTvWKFIGdpgTTl16tm1zO7dLIM67
X7XHpm0t5WPrVgH7pgCDv15H6zNpCadQWnhuJio9FiUvW2tuFDcUA/c3ik5luP6XnoqBD+mTaVxB
jwVrmcS3xXsOn1FmmUoeCT1OUAkJsearnPpGFxWR1ofc2e7HPxrLGzXS4U5mP0dxFXyVA6+eEGVe
OotE5bY+CEMebkkQnQJNQL4y5cS3MTDDQUFa3VShmcblvmc825uTGZiSe0uq3jSyAXkwUEtpbJ7o
3mbbnWl0k0Ua1f0eDYzrBWeYvbK+TBtLHvO39mDapobLL0fAurqwkNs9wskIJiPEVeLLaSO4Un6l
BmjlcGV5kf7E9hjBhEdwJ5RoXOfKL0q4vwuTmG5z9Sgx4vXSNtcvmW5XsQGp+E4LM7AL5aijQaAL
7asAgwHqL6PKeVQD6uKurdayWERIU9KDHc71/zerXIo68iaVsWCgy4NADW+r9VhKM6/Dsm1zReUQ
HUNmqEfLbgQTyUId5rsjoH9BVQ5ZnIMQlo0Ju8VGcCMKY31MVQAFaYmq54v3EgtLgJ5nABghbx5O
cDDFy5Ofv7GhciIE76ntDzKmSOBen/0iP4Hp2ZyqOuiop4WojE9gtycG/YQ72WWO/anzlqPwovkn
dsIJR5MXi9udrIcv/J33hZA/gL5b7+fl4seL02TsS2miOzxTmMYLmGa7wCxEtY2jwSevVBXLif5j
nTMpEOniAVHjukPp/6dFVJBjP7s4sykCjL8XQf5pS7Lh0DO9s6TKpmzP4QR4/SQZ7zrASkx8hYjP
Fo19qDjZiNl0vMpYv7cfp1AtT8HDcUZVWe/q2DQu1fOPH9m8AzvxyLuLQmGAq6Hz3t3OIU2ViHiC
zDegMuR152LEAqvHx/CA9ws672ei6NkIWEBqqGDCnWI4snrZdqMK4Jmilqa1zB0t9vV17pB+ESbS
HxGHqCIMWNaMCtF3rrVMJRQpoe8q4fFk/9r33IgaMybDs/8lJG+/8rucmyhdH+FJNS8tfUxkZzq0
mgWu/U9CfEeobkE5exYPzXV/oMUVp7M+sHwJK7MMUcJHvXsbO3G8h42RH7o5OH/G1PDqFtEaTW0x
nsZxeCgOzTqP6Evab+FfcP76WdECbHPaaqQM0gApFgPkyBlCvgNF0j1SfpUD7sDJQN2eurZdaKgC
iumya1SIAsqLtWtwZyG43i1mncDdC/rzWp6LtT5+R80iZ53A7a8hNLXMdLrdCQUN9ayQnDGtz4/V
iybLvwAbFNtuVJ87tdBJVdhJS+CrKpaih4bUTeXfoXgrB+0CYIz5zo8G6RWRlo3UY+DxVmOj3oPd
iLjh21ZE3bNdnmGf5/PiKAufxmslw6EufsNuDfNWnJzLrmYXia1F8R6sAyAQPs9qKF3Q6QO4hGdF
SgsDCT2yEqcpooQRyl9a6ORXvgEKGGr6Mkcql92fy8KuDrLaeMoiTie1GTlbCoBpDauM9I9MLvRo
TExjKkbZSgPCoxti55its7MyZyCzV4nvn2hgljNpOOTzXN2E53kmxASR0ZcBxT8CPRPIfwhIqfIy
R36hrkVpMZkiuBuswLYGj4dFHlADzmTSZv48BmJXkhAUd5tisa17laJZRv2taCABCumgL7dpFhiU
W47UEo3Sf1nzcJ7q6k1GQSCR3E89uKjJIVBDYoOhsDUZXfZ2mFmJ91uHbEO/M2uZ58nFtvIZqP9q
rNXySU0rbQosHHvkmmVBLhtsyfkGMGsQx9mK+ubitI8VilxUae/9UQoeAxbQVspc1yEQp70ePC25
Konds42efaWoGrXekA6vVbQs34AM7IhYrHWijv64dPyMBgfAYUCQ68owNpnKIQUlML72FeIlqdmq
zmiy82fBKl6+ClpbcSB1E+mkJpMT2bq5/YN2aFu8uIPFiw2D4Ab8iB0azWoOflkMOTJzR+MR27su
OQHAjFSNfeaFph3smfC1w7RWWVC3cxayNMoHKW/DLmbV2Ffz849EeDINvJFPRzb0TppdwcpQg0Xx
Av2UfEqVFmaaNHY4kMAAAq7zo6pfcS0a7sSDaQPEw3g1hPy7lDMNO2Y60lN+k8ppR+JR9BPTuszz
NqQ15VAUBYMA3fb9Lpg7pTg0Diu4J6fI82fvh+dlJWPXw4Ee0cf2xqdf6D7ghHUACUAS2KNxy3FI
gtr4mD4cI635LWzI9y4jlk7/z3BdzXXY87hDeD/C76R1vO7t1dvcYQALiIAilzYeckRBvTRPv0uD
Au6hyetzLqePKI22nx6xrwU4xvBHoWkMU9Mg/Z+6L5L7zvvUz8EpGpRkQ5iQD0NV5LoTNg4jRrpe
9hjEBmweHF7rzf3MQ+PoYnJDiZ+WmMLJ4MiiVq09c1i/ZA8maUCRkAKi+NDtFX61/4jXQUC7zvdO
zN65lT2fIVygUE2zGnrNyP8Qw6MZWSHwfZc2ZQwwJqW1OiKjffAp+n+dCR5GmbIBQNzt2YkeEdiF
vHsNMSKtVlGw8W5Up1r4Ioym6lTjJlCca/4adMBKcXZjPCGWPJQOuYf5f3hcVX2XvODgAjLNVm1E
yLKaWyunB4FJhgTpSSYi9qPv+qWBZfOq0j8JOx9B/uvBi/VvwvudeQvWRQmA3dJUS6FNiIdB3M8W
PRIdMdQrbFzbcGGVew80Kz/dmF2qhtTiLWA3HPsYF0ofQYtcdbEXkFo5xS9a5xAiLwqzzh1zw/kB
X8ZjJOvnl0zFpRGnG6x9UHBq//C+rq5S1k0HaG/zr4O87Yf2yFSGYgX8Pqh+8Ry50YEp8YE7eZaQ
FXPWbzSsvh2v40//Me8kSqF6s7gi/pwezezjCD0KVGehF0iuCCVynr1wMTiA9RjK1ZRBMLloJU1R
/Qhwd+jjjYTng7LPZJFFxXagKXmA72aGk7f9GJ15+7R2wcpni8hqkUBR4wy34KiG+7KE8jo7mkZ7
VeH6dZIpm3dO8rp3SdHIYM3Zhl9j5XOVupZgCt8SDvekdsfPhJr7Idnfi/DzExIhvyzln4aYh+pn
Y5N8EEz0+UodbJpq7GWuysETsO6n6moLmvZfSIwDpaR9LY3VxUOFBcEsVc081lEngbro9Ish6p2o
ddvOBUVmg5rjLMo0xTNZejBIXsyv8q5KSnNIQrTpk6UOTSSxB12U2JO7UL/ruTnRgBJgBFnOWCS+
KTAf7LacDuZIyJDdJBP5upEqW3HTLAzKp+vaJ0jfmKbwdcCXsPqDbzeEh2Qo0MPrHsr1uTwG9a59
3aIlevAlfMxJaBL4pqCMLxYC5AGNMJXk1hNxrmcKrc+zvWF9gh+53PQTR3/eES2bPIXQ1O9jzldz
PsFEkm4Ad2x6uRHVss1awVfC3To5YStA0oVBvfhLZqqVjELhh4a6x+FHW41AhRlcldcUSmh5KsM9
ZEi3cZaJJK93xSWJN147HbsEmwSj09MCNP0exvtBS4dfWnzuOZD0bfYyg0BVJfr3MS+OWicAHCKe
TPBmtj7cN2ZWcsRgekrA6CarLTG53tzjhw+VQVaZEi+vdZHfTQOTO0cdfmkLsr4tVcVi+puwCItn
O401J0GnRT3439kIZnndNpkydyZENrfrDqR1pg+uuklGOERbKJ1hGQj3Adulup79FfIrTvmEsUNz
Hf7unbtudeuHWOLLP+Q7BwO9DutffaOduvxR23/O4tAaUUpcqDglkFDndrp9tg3EDhgJJvlvTX/R
P4t8r8tVyXi5gdTR2nUUPFbaDLC5WE1Qlr7T+2eV4SFfJbcjJIYZKMdZ3Sv3KlYdqyud7gj/0cyX
PdObqMX2hTOJuYzn5zrVU4UJCr1Yf3KWA8MAguuiQZExBeVnKjRanPqFhwheN8eD3FAIKDRf5Ok2
gX3WohyxPGxnvCgT/xcWoET4/jWk0HOcJjd7Sb3UM/OhLeW2MWwMBMP5h+oACmCg2gqnSF8PsNrj
LaP0KgqVVVxzWUMYGCygq+NudgvP0+ePhNq4cFU4e0Ff1OBUyw7qkpP+QWVwDtL21ruZcNmxLXlZ
jrHDk6NEy6cZ8GPCQZJGZnm1QXGV4ln5WJXIfUGvBwOxQ8Osr0oJwha3ksZxha3S6v/vwByLnTkz
f4VoJcNQxuKiq3K/rIudKt7DeN93X5sZ0KVxyHa3AWRPIMrPcXg2ijx/0Xx06tFcOU8E9wSdTJo0
StRGaCIwSnuuK4+EK3FrbzHW3RqY0JrDqQLd0CHou9RD9EyLJqAngOB88nTf/3KlBvQj4FZEpLib
Irr8dd6yO7SCgVlKQIqxFHKXtE9kikkj488G+ZdP5SPCPWEFhw5+JKWRJMS2pLf03X2vCW4/Oj1B
fV5QQLQ9XXhZPXlWa9eiYLRkStHW6ZBUMZgbhtlLukWdIA7toZwNV8I5RvkZWCS91lW5NULwbH2l
NnF2WPR1xUiHL5+4byvLZ3nzytioejBV+bW7SH5jiQA5q+EGHQ+yIkSRw3W4h/jLwGflE1HskoQP
J4SRHnPAUqryHcVY93zzXBt81BvnjsRSGphM0d24o6KnPum2NJ/s1Z+ddzIeC5H93C2qaa2qqDla
Dc5z3kVIFahxU3/UwqfSbtkQcRmaEoGxny+8t0M53txHay0Zn5H0N49apeA1UQWXSf4wZJrOIIdo
oRQwus3awRJDHoO8CzB0sPN41TuYOyqpMEeFhejiwTer6kAUFrf+RyF4YH0QntEBsIaF4aV+dILE
1jY0KaReDJUZDwTBmbIa6h9aRuYo3qWqUUveqAfjBRkmd3N0Xa2Cs9KtANKr9nZpJgYKECJlejb1
kSnUko9G4oWnMoWKMvTf0W6aVX1zc2d/XdAxXrdbmQIxkCwErShnF7Pp9oTingUKqHoYJso6Oe4+
ThhaDsgOQdxWquV3zcqybfafDhHD25ftMnNtaCoa2Ej/sZxc1csJD96CF4F70SjWgpScx+fXRW7Q
gH6iCZxxGlX/W4gkc2Nerg5ANZtVAq7rM85UxmTfqBs4Y7wwXaqsJAnnJgyyqtI2xLkv9Chkj+5y
Y6qDFvReACNNzdlpof2wnNfHUiLK71246CecfZsvVPjOSNkbFJfLI+puzHD3b5/wWFQPhEBJ8mG7
oRf8b4BnilvlDi42lu1CXLZCGEGz6M8y/Dc0KPvKCa1IXJ2aMoSOhlog93YL2BfMvzb9YjDF+ipn
nRgQFMrD82L+lo7jJfzoLfXFQBIo0DOjmcUoUZG0M8Hr/rrronJQglzGongr1xP5IesBWlCAtuCL
5YRqAAbNLK50eLAPPGepls+hnL2gzKoJUDPQecafJJyqYCp1QFLoIF6ihBtcPIQtoyv9Nn3RKT9y
Ts7BD4pRWQjvFk1Ahn8SAMDk9UievB9Cg1TQYt6lgk2UiJVls+cGCjbvkNR0du9gQ+bv288Wi5HO
JDiiAQv560xL1aGg65qLDGwjqe7H/XuvgYMh8XXwXDJJMeThdKr0bYB9XJg6ZWEthJdngVKnzKcO
K8JHIlZDX7PIVcIK16YpgMRqWnMXj7+xY0+wor8Lnn9RtDdcPK26XgIM7ppCfFV2qzo18DVML3Ql
G6bm1J1WVJLfd4Hl7CBupif2LOLcuJPr1TXf3TPqb2jiflTs4sJqY3/JQ2iwqvKzRqeZ0AZdcB1T
AeJinrsjMV1UgG/rbir7fa6ScYKz3iwYHfzq0cVTi5P604lWBTCCueYlQZA1CnsbK+0aqAzSzn1y
sU5dUzrtNzYLQ7V72qVc08M17uuI4OHFdDoRQbVOS30Jb/1TF6Y1lM5do8znUTMF0g9qlQWYsQyQ
wUg1l8fnengLB8BhDOhg3Qecnmpccf/kj3zf+XlvbP60IT/aPQ44RI2ROm2tnx0KH6Pnk/QQrndi
gUbPwcXeDbhqMZGam434P2SBHHe46Sgo7RKbmSZLogD8VTMzztZlMw938V21psau7bYulSUjdUlf
kohpa44wq9j+B3JtcCCYC0S+5LKQSzqxnPhfc7qE4CWaZs9LX1JMw0x7pqbnNRNzHXEGADSouuUj
WjayUAaQoBBECavjZg2JGbSloEuEFoOC5Iq3OTXpOqtPe9P19IGt3lKmTBp2wiLmPpkvhhStnCna
hrJLpr1N1DM/gCYiDOVOVzRgPUYQmINBXpCU36KAntRFmZ4ZPyzrfS9P51YKsIe17ArlT0sR+840
1FxFRry0883Ybb2EPzDifD3aCP1gqUXGwEYHy8bdZ5LVRpjHv7f6vQKdrBp+PgzCC+LzMe6Wkjsp
sxtBH4QkJior7MxuHUXXKw7gM6Zx6P5yB+GucWLdfukqw5qLFXm2y1jutJNSCkJViYdIEpYyjrK5
QeXhHXlja8X4e+nE3WeaY+DW+uTpHNVNtcNbcDBBNTZDSdx83oIJlgDf2oBZPBiT8hzuXQJPUtlg
XgCYisGReki661nPTO9vpN0Puz7QxfnFuKHaNKTLWAvD+KigcvxXU6H1IO/+xKHOvg6nGlzGOmoC
gsnBQAyDxIAxtxfGQ3R0sBD4F4PbvLUxZw3/rzIN7hIHSJe2F1Wh14YDdIxLBQ3w8850ZcRp8eyI
p8MS11oFFLUHDhb+MnMLw5hNkspO7BnMacv1LilyVWKzbjBNIZVYP8YMuoK668xFpMoLtCvPKpf/
QN1OH3ysKnjK7pC9KFpMjOzJG0kQ/cvhQQ8mx8Ne9tnrO5R9YNt8eEjaQe42PryXsGscdKXDcRTX
BnY53dIVrDqPWpI51uHO9jP9c5p2NRwoQW53TudAl3BT56bzFX67P9otEhaHHrsFlxzg7OkGuRJI
0EplJFZp5HzhNN5vaq2kIhDYX50cH7DRRblgzjiCTAdAyMteAhRkviFNjvea2rI24Q2CcGmqCsxp
uvIPKy7dxRjxm+lEtnROz1O8tPjVZlCLyEIt8rAWzcVWTMi67aqn1jz8Mee+L4TkAXek4buaWdJ3
9aiGRXZFVP1tBdBaEYOT7kK5kjMe7t5F+dHE2BOYGSVRfF2yKn6JQJ3ybitEmjY6+YSJNtpxCtZ4
ebc9FYf+4Y498SCQkwipFxCjdW07zhp3CuLhRJVNlIeqYNCbqzOZODmlk9hzLdn/3E5SxJnWhSUw
JJqMDegDggLtTM/PdqnBT/kCEBEu+zKW/M5fslQ2eIGOcgj9G9TBSwb+3rHYwArndEDVkzQD/9O/
GuN2Bpn2bruDcMkDBp7wYYRkUUy49tA3EtcqwYlrpGHrswwwdKYn39dRB5YM//7A9eoBrTpb8sji
+ntK03VdvLQ8DtWc3eeEFDtWNctrwe65Ah4hnbgK8GZ58nkgLodoP10Y6yW3x5SUazQ1bBdD3b/b
ZsVIXRM+y8Q23B46wrNLqXPVVlTQUfZK44h+5j+ZmayqhFzTX+KFncisGyZcOahefo6vwBHVcNnG
g47L4wAEOq4iDBT1TzE5ELsng5I3Gs7O8aEKlTKM0uaU7qJouqLsYjEejUE13BbO6ZoIALpYKWQb
TEu9//fx2Yq5AZjOMrTVolut3pXCPVgbFfVoggXyzTkNEG116MLh3Uj1K7l+xSrjX7WUeBT1gvAw
X95LDNjB6iLM3ecmiX0Ya8SQs7VcY1vXXKPF5gh5o35gnOQHmUGkYIbm+6472XAnGzDPnBmUTN1c
rknq6YIYpfYW26q/WxG+WQGTSCjAKO5iKxfshHfNAybzPTY4ryzocjXZkWop1Uuxbz1j6hpsAWgy
GJ2ErTP0eAwHhd6ZtyM8DZFmkCcX7+TZGUQSjXsCRzxOv1AcrAIK4bUkLZVAJ4Em3CKVbVLnQuL0
8zVBvFKkafBeTRRY65X26tUP9wPnRnFeVaF4Q7enckqYGJx6xx0ot2KeK26aNJXow4EK91XBWCFD
3bdTDMJCIiM/WzdMe0vMsDUpxLjexFEZXfNctUAZwnGT0vQXAnxVToqn1cuVLnqtfNTqGda8mBfM
T1H/vnwezkOt6kLw215v1fDdnqPke6pgfe0dgno8ItC34/G5eRPQGvyQ4WZ74AAjplRGY/s9lMOo
L78gh77lcjNdjJCCGuN0fn+iNOloaiDYWsWAumpDo5jgh7rpVQAywVp5kpUB7Fsle8HgiVur9pwH
lTBr07n9gxVipmKOvyz2MYNF5EYykhz4Qz3U6hlAyJHWmAdGCdT0yMhWi2k4UTQZd/F8qlzs5p6p
Cab+z1ild2QenXsIdGyePz3+ewZsU7mEI4EWLJrcoGVu/yN7EarOi1v927Is5+gtxKrvUorGxo75
hSf2ZVpEKlodmOad1cKYrBvtgDkyOcype6lOnUSGdvyxN7Uq+kqCIt1qrVch/Hd/GdaRjS7hCrwM
4v6Em/d4HA/9eU+AUcrBHt/hTUnWzFp956EFx2CzUEgZkeMHCNAMB1GFRZ1PQLct6QUJx0IjGu+X
YfNn5zgDdkkBwfVhBQKZr30mpRTkNYUug3HnJ2cMV2z5T2s5JFSbXFNLUB4FKlnGu3vbRH58uZJy
2VJLCH/RbHYRB6wypUxoF20VlxN5gseOt/9ITBoYPCPfAg1UH8S3XrGe/rHQqyXcLzZ9hXXkQMTV
5PxAISqa+4ZgGPPFkGw/2ZQ7oU7dMi8VnNPROhjZWYbwFH2/KYVzoRi6w2vOFtPBsqfklEA6y2RI
CTBoJ4pqY4cQfiFb2MXRX8KAttvrhvr22kfUJC54OJRXG0sGZeauthEFQzFkvzV+G6kDRhZFUZT0
74eCZ1t92jTUyYACks09p2uFKBm27GW9OGH5j2gvjblU36LFkXgGHtBFwqPZxVIoGC8BJ8a0xwW+
UDsHK6hyZLj470W49vKxSXK/7Prjndn3RxsNZNMpdlq2qH9kPpitplEyaOufnteeWn4s3Z75+JME
ifedJ6AQ1/k4/4Whp/tNlzsfKlJZO7v5Y/dtehuOlOyonvvUxqzePf2T9devih5wZWQl1d9x9TUF
0aK3ljZ9jAMKJkvxyxrOJdN4u+kchs2xVM7ewG6klhmPeV7av+Xquk7Luvw6TKfMwNKsEPM7FOC3
BZ+2PrnTIZ60k5RGKFYu3DUOf2e3X322TmRGQGF5v9BOPeDTyA/BNaOyvBCCtWTwqG6TynrHyz4V
cfjoWWOjwdgp9EygcWuj5t6fC2hFOrK59lL5sebXiQw8ISAPxuOPIIaJcP5KZ3g4Yqdy32dzLZ+L
lE7aNP5lloJpa3ZIwZCGpxFORHLpKMv+zEgwHDGQJ9i24LPLPUqYCiJ5NWE2kY+h+D6qs6n6Lh8Z
2jO27eTJMI52HRMevkxtmIBZW9G5DSa2jF12AfFG42hxs6Tu4oGQ6EagvtKRJVkhctCiiLCb91DC
wSFDEY28d9LZ8ilJbHxdVrq18YfGeOhxSYtElf3Kk8tM1VtZEmYqGDteYdHLAise/XCNOhlh37Ie
goyQDfVosHVMWvoj7HPTUv4kYoCvcHboy9V+e3xNdq82lgD7cSNkD/GqHsFlNCWOLlsRwm+NPDyf
ikRQj5x2OUC4lin3qot0J5rled3IM7Su6xmGQytTOPJs1LtJN3J8iQ4HpMhcu+WIyuNuvd6MoXLH
zzI/pUwv+wXZYPDnGBlts+KcuKgqjJK1hj+zByFu7afudxtjHTglYsrwLqAUrGU9fnMNYqKEO5Nn
OtKbhYdWRoefwzrYUuJXNO7+58wu48Z4uFyoEoIZ5Acx+f5ES8EVoLhhYi/431Sfx5Qpy/7qFe/+
RNnR2kpRGiR4OkDQt8gT2PnP8SK73eXgZ7DYLPPH32tUdgjmF5L+UpA8kfYbZ9SqxIPbW0j/i7no
U33wG0dtoaLMJUa2uSnP9E55/1KAkZc4F4T7ONqcTRvI76HqV9/VVtjV7izZ/ZDty7MuYgdMf1Z5
To77n+4TsV69R/3w9JW3huCyQj3xm4IpgJWBu/C5nhdlqABATsLxm2f4hzO9nE+VzevZOOKQwOmw
WM6Yot7k2BWj1UkACPCmQ9U1sKbIKuAG7kx6ytBsBP59pmiblDTZUo8Ha8E/7nOh4A1yIEfv7ywo
FAjX+n9/6fiBPrPZUslnYWZaBx3p4Jw87Wskj8/Jh0TOO2iUyupMIjgt1AuhwuQMqHinWxfdI2+C
AOA9CfzZTHm0oeP9fFS0TASbLKTnKxFkXeSd7pGFWjhxBSfJM9pOXax0QxB2GEdjPDrlauG4tcDn
+BQYrgSJr3pSXHvLMuGcB4KLoVzMJaXsRdQvB5Q1CklOnvdyrB/jH3EmoARXgFNUTsqJw0f9YxlH
BLeaI7475ovXdsDPa5XSSWpGQfDy8S3BsVXBtLPRk/+Etv9xPFmiC52NNUQBysipzj05hht5ur5Z
tugn4tV7nzw47a7KBqH25hZjU/LlBr5AWNy9db/sz4makMYu+DwATrCVrAVk5QV6xNMVnmpJ7l6Q
QXKJjA9hdgyqj+nkyZvYe/HZ1Ci+Adp7+M+syp5aC6pnWAtqT7pjoRBx76+k8c9EBZRnSa05ON0R
w2Tbqq0egtFax2UeLChb9EbWt1bfnU14nY1xO2+kYaKNaEwEDRmAJQlwV9fPOcuJouq/GpK3geHH
YveQo3ntO6GA/luXlTaIAX+kLthEOhNSpVxH9kQ1PQ7jxHTv8J1bNMnAQpltYnDVeAgy1PnLk/Sw
hNoKjmymFjeKIhp/uDCcy1IFe3OksMagH+E/J9bdymsl3zRg8jNs+K/n3yzvVt0WbbV2vSfUEcBX
0yR0A4+3fqMyz+4/hJeWXGNYNoGp/P2pu+BccECNjiDUVZtCBswQYtbODCfiTtqx40EH+rbn3wV+
Z63HBSZA6HsKeIRlJuHHFcLdKzm4BbZ8tyXLKFamgtqV8Kfc5300pXsNJMojp9tZVYtftOGb1yFo
jw36hVXWlLzWDgNBEjNsXgIYV7G/iK+/rU4P7FPlCdt67fMCZHbj8PCaI2gA2iQiWr+lC0MBzjR3
jAcW7Xu08ktb5q4FXSCNCn2moF8HbrloyYetYw0wAgcaT0LBqR1c78joAGbj6Mfw4YyetXK+zqNN
DWfp0U/p8j3zRswNly8XU65HQCRB4Yrk1yLf0cmXEKyqntFSFZ6jsCLTwSAt6HqTIoKEwtQivTN9
ChlyEp6OUDgBwd0hfxPjiptOWqA2mH1PD5OGkGrb4hjZoDJtLB8LUllOuBbvp6o0yMwrBioXrWz8
YT0H23jGy0bYNqYIDM1QDway+k9l/VoD7vGqNRlx3sSJMXfYJb5wei/CGHAMdsSCctHTCcKVhl2F
VFit2c/w/lRgfM39Nni+03p4XhIQ9qW8P6vVN6F4mjk3r15NePHvzGUYZjlxzvaSjegqbUr7w8/p
KAZkcS9xnazjhzp0zvgFRJHd098GM3tO9qjwlgBPndRZ2qApyPRugBWJrp5i9udRZ0l3vyrt2idj
/4Z/042WiuaAZrvS4FJyjn6F3D3OaKGvB1RBAessboLPFoQ8rIRwKwx4Wklq9XxMEOtmvgTf7Gcs
ylF9z6Cp9MFoThr/8jjRT6XaVRhoxGL6OIqwcIzvcUp4IcZCWPbEGpLf2fIO44pqmhKWD0GpeEtA
AJFWmEy8YePnYmNMfWIjtdC99/zQxXtbrwQPIHjmC+V5Xx5BizR92SDvUWq7fFuqUyntzbgM8Skw
kG5pcGD6ajkTIXUclFSWorQ2e6X/yWwPY2fWJ+hwCYJHDfTaKu14Mov+oLfV7z+rL+nkMxkI0UcO
OflwrHlD+1C1WJYvywnACNYQ3DjciOXz8t146FJKZZQYvAAQVZjQSM4ksP8bP17ZvLE+Y2+aU5XC
3zyRwUHbtRIXrZ6Kqr2SzAJt6Y7t8c9MlH34nEKNqQ5v7Fa8W2l5Ah4DSiUPXzpKxPdUC8ZiOhWB
S+2Sc9yP4hhtZRIBtF0pYlQTx2dehQDaeowDn1DQC4l1X4AQ9i+/Z7dB6C7gr/jDNbQYhY8H5A0M
TTJKj8HYswqya4cnNnechK9VJJt8sQoLeKpr8p7WFSVpNyO0e9Lhpjxy4s2Y/ZmX7zjbcd7y3agq
n2CKY3rSyaKMx1MuZI2lfoVEBapWW9QNkQTx7HrsdyJg2kPohl5NvqK2YcjVj9AQs9mdZK64RUnW
Di1LqmbK90O6qpD/YFwMVfnIAYs1vrcHAzg5s8FH1qPUUHEBrNnqJWJ1nJM287MhhiR+EuxO9gf5
BWcAlp/9++p7ga+P02xjWPKJqwh/kPsegm0YFF8yPfej9kRxm0eR+tllkF50oKG0D7GiAu1K5xnd
83cXp0M74ODuBGXP5Fm7+hUKkDwOZQ1eNSGquP+jKvIwDEw+hfBaDkVsHTJvxK2MimVBV92M+8RF
MSpiwxTNsS2dngNB5/1JZJLnuEcEMxXzNGiyOfHpyFmyxzZ398wuOlixFauF9hIYFh8APrZri1hS
GlYt0abpeke2qF0mprdYo4B8QpfYB4l3k9tLQ/mNJH1lIcxNe4PFBDz3ghREhpwPQEo1xTkCAwPK
DVDkSfrE0OkfWj8Yc2W6yAo+GP6uDtCoKw8d5k3UnCuto/T19Oy8K1u/Yrq5NjBuQc+taF4wVzwN
txiQUFa9ERKWfZGkhKaLS/wrCnKuDPU01eU7mx4Bi4PRDM78q5r8Xu8h5+Bbh7VdTqScE51t74h0
AE4nbRsyu7KsUXSzBpxzyF/nvMWFdT65jowNv3GTCbfNwW8WX8C76TP1tvEDG0NXTMbGZV1hZMWE
A6IUzHYmv/tTMQ3rs9agVm6we5vj7IY0BXgKPXSxlms2BjL/DD9Y7vZjpoquRwEOt2i6QvY6Z7gC
bsT3fq7rHS90sl0w43r2lORRFKJGpB250JUAzhCG0jd+sBJd/ILszlBx/RmQ6LtAcCic2VeHJp9e
66wlRGn94FjyipliGwmz2FK/39+yE5HQyzzNSi5pjmJzR1QWPhWtYl8eQyR/xmz4k4u2S/uCTPW2
kx5/liE+NO9F8PphWxfACV+uKMWG2EZrzDguKRWglTpLgkceQFUx2kiVwxaCkMY3r63Yyoj1WSsV
zbMiojfGAm7h2ghEUkd7+QU1SGl816R+G7DQMISF5w4dJpB2G4lpZqFOXcg+vw0nC+p8SkDW3nTX
BOC1DxgpWXkW+N5bB6Eq76nQwdLWOyssbG7s3HqcLC+gfaQHPKnHYpx34KTTZ8Qbxr56NiJvXPe7
OFmG2OSt/vYTjKBkGc8SVJe9yyUxEG/WIaYj0t89MkI+QtYOkGTosgqcrIvtZzCcH3mEl2IgtOrs
KeIGqp+YZMkOzZx/7Z73T+vCGQwUCJk44aKr/sPUqk9Z/+44kLOSFDxIDPi9uGhm/Iu2EdpMNQuR
vQzSrbZmlL1y3e70U//MIKiYBDFcx1LidrcLwpvRlPTbD9n7xuc3sBT/OF501Gbp/C/gPRDRP6wo
Wt9FOKozdqKWabevNjMSrnGYBAkIZgmFPrveOoV5ihtkTm2bN6LsD3iP9onBEcOZLqGedFDGflI5
XW2I+7zN385wb9BhZ+6vZxoRgox3uhk8/kWx6CWSn2Jrqto7EwyYJgaxzXhYJpQnlEovAMZnagSp
FxhDsPr10I5FG0yvU9JvLzJlUo3cghdQDIfF/Mja2ESUihf5lC1E/fKKFJi+NcQYyS6Sfwp33Q0h
DsZZcD3B08ui2oIUyuTzJBGqr5R5XcWpjUT4mPJQGRCa75gmX7e79JkyqxMBr3IcF8Hbq9UGZHgs
5sWWbOQ8HGjhyeu6hBBstlz+3B5u5O8KezN0kIdRDtF2md/2vDU9jajQuP3mpuN6aNwXe+yFc4m5
+3Ur1YxoPXHqB3DKovFFVLDn4I36VhzqJUjaxVXiOj3FQy9VPfuhS+gRRsvwSKXga5/ePdmlFb9s
4k2ZNbkJtrNRt25JqBA3p2oE1rfseKTG5RsIsVfILsVSCxlNa2jf7otOTWvqCIvHPUdAUkoGY7Vi
np0qZ5PLCAxQlUO9xn+BZ2kQG0J2UX2PU918LrK0LeoH57gWh41CC7IbAOcxs6YRRmgZH5D6Eanm
RYQsSHFnINfXt3jE3kRe9SMsHAonZwK6Mr6fHExmroskyrcPylxIE1XnAE/l/rfhUcZBkoTQOCJr
8sHGkbAmTGp1n7pzYLdNr+a9D0aGLI60wjwK2U5+lLdIM+757Vcc8F39GFLiDHq9pFF2Dea3IC//
p5L2pECY8ckXMQuNZAZdAoXDvkyxNgWjU87HEhYZM8lZLJR4G2/qUrJI7MAzVVT1GiKzkN/20kZ0
FKJsKT4GyRGNZV3itmF40mkB0+tcE+GcuVZ56QS+m1FovkJExViZ+h0eMhljhaF8uIVtnKNsQ0xi
4ZJpZkGAxZLZbB7ndSVJR3Q7n79xuN5doef6nhhJyLLNbCZFjVGyiAQwXu5sjAKv6K4S8xu1YM6C
EAfohafg0LrhpVUn7G1SRlpS9xv7nl23YCAPlfvyt3nrTb027Nl45uGA/o8jlR96T6fM5c/2dQC1
9hxsJ2ih+MUhNMRuqcpuepHgg2UxwMoLBbh7NLc/ECMMtMu4trqQJ10NW5PSuA5EFOhhfsP8s7BI
sb6+f2AaWrkRT9nuoEz5Lv+loVm9OlpZoQ9lFpm8pE1MPTA2nucus8QmCXBcANTW5gqrt7uPxr/V
ihlJMMlL8XbQR0KVEdXI5BF81XypyMCbi9jqxZxffdl3MTGQthMXPRnVzDdKK3Ccmu+dNkh6dz2i
ECeoQi/SQeTfZXne2NvYKutazF+zm9UfmYQ9RL6bijEVJILdR2/b30z2yoJygTdPE9caLuuEZJf/
bo3t3xOHR7PnpDjbGeZ7SJ53+ktLcdoQcLBZm2L/QAb45hIsD8d0iavYngL/xKLFym/TN102Qo6L
+HPHioZWm1jR6SqopdLrGZPdMxsdnUG9UkiKNvGjx43HOrK7U/QbxVk5l6+flLPoWuDo7LJgZfVB
jEgx96TUac1Syve0mbe/t0pcC5vUtYdmAnHkSeYWrspdSAXCgCW2Ug4xRYfG0Fd5eTZ8QNpzlmHW
7s0yAwLopyGNvKmQ74yz2YWoKPCmpQdc0Cs/RFAPQ3E0N+3AtnA2/U0xYJV+hbjF3JES+bufs2UT
cTlPSgo9+y8hfOPbvDNxuBLr2T1Lpkl4khz+b98Db1Qa6DlIJu+d1fzHrTnA8FIvHyd5sMw7dfnZ
b6CCiq6aaH4QHrq3ArZR9tI4pnHH8EAGLZhcFH1V9rcMMDjstcHTjX8sD56z9gL7LU9Q86DAv1BC
+/1Q0TLb+BgvTRzzF7GY2abMkb2ee1B4ymTCr4sYXS5Vxkx9KqkR9RzQWQMWNqzVtCpsV2T3FLxH
ihhRQNezAxFXn+r9iDHKkYcgaUitnaAkq4XXudkx23h3XYofZBoKBFDmeoga2nac91sQkIEuaspW
fsC7wSsThAfj0iSvtuexhm6y+5uHAVEn8/Gv67Ojyy6El2f7fp4lJ+9PedvQ5irE6piIjj1E7H5P
gG+FXZCt/tPWknrlTbhIoeQS+NCUEphMH8GHUl0YLfS6J6taAxWrZr2EFdy8klzamubJr23Ta2wT
1ERNS8rPfTsvcvoIVzwKpwYfX3q02FgpUwgRAjimWszvf2efn5SodBn7It/jPrleXc5VPS01DbOq
moR7+pM+qjppXvR8v8QeEfVc4zGf7JonzR3XVvBL9bNqJIfTrHDC8pCDSaoNYTtXi7Y7z2nzLq0H
pay6eQ2tMuT9hIsZfgiT7XNb7req7TMvV6EHah7O6o2jgpG+mbaATRwzKKzqXCHHcQhsH4SM8msj
9k2DsV40SarNk3565715G8zF2nLXvhedAt7tZNDRDo7t3CaMHE3O3tNTKerFxnEUmCU6U0wi73Y8
9XvveEm9Zrh9a8s2/eYWS7LfxLQSxcHOWUgJFE1d7zcFTRuACV7+Qd11xEvKNkBShfgtZSNlVHlg
OQGbbw00+sSXGxD4hu+8uiT3JLJCe13wbY3EuPL8FWq3MM6gvmYwtjNcOZjGSeZQGqKub066FUYI
PucsR36k94wkiIG/jL78G9bCrz4TbuxUK7601R+atEUlKaMQJGFneHhC+ygIz64DzsPWndHuUMYD
zSCl2MFU1PGt72IgDFkf6/YhjdkNoctXAGfFljsDMdGYG88iEB1oa++JREBfN+sYh2yZfuKcMqC6
ZNNRvv0HBeGZ2M8bn5OgvhntHsWsJVvdbYaaIs/uHpK2fX8G2wrxvaeAAM9+iQrALEksZOgjllSg
JgaLmzqVuJGBGViUB/V8D+AM4FbpgJ38fEpM8UAUdnGv9G38vaH8C3abbxtM9lwHgU4ejO4cykZy
h1RMzX9+z5b+/SfR6CFyKwPwYA6T/QKg22FZ1KyGGe8DLZXGyFbghGXeDbRCQMyblQKD017mavV5
dpH0YXCrWm3YJOj0dxVinM46De+SWItkWF9fPukgG1PfrL2Kb/WyXTwsIxab5hOR7d/pxv8Eacu9
6JJnYx3jdUL/5NeERVNvr6a4aOgCNTXhPBYdo7BuQ+eO043HAylzrBpAGwrJ4HBYaiuyhgI92p29
EKQCRA5zRdiRHw0Voi8uime4IEaxZHhkzlt8Amp9ABTL0jc6FnY/OK4SbpUxHde4U3H+jS9l/xkZ
iqjz9zfCA/5BDAoLb9aR1ko65isjoLaJ3bGRalRWE0On0YIW8e0+jl4UotDxdDLQ9bEO7D7AKVVl
20igp6iXwrirFLCH+2jP5W5EHTUiZ9pFt+UApSqrgI23opjufmMK8yYdz1H61NkfHWXgYjCwnrqV
vYhkfNNkvfZHv4nHlHYluD4Xb1MUlZA0NXwqksnC9NoGPwEMie8v87nOw9yFSaonIqIiiN8v3NOX
jM7cXfMVrq5OfVq/Q26jDOMMmjHHBAxd6acVhZTpmauf3LDW329vOzldLZYdMhZ0LYbomQPVjy5r
p7SYrHPrW6kox5xGYqp3I7X2qlaG1KZAzV9wQCuQoSeXJAvbDaWh9vnCdy5S9kyQvuWFEmzgxXsj
4E/AxjI2XLTd13ule2GKV/YV/jAS89N+NH9/LGdyueOlLnSFXqmfS2p5gLohJSS02i0/OItZb3s0
irV34ohsMM75npABOp3o+Hr4VwRyicQ8ip0EBaaIS+mnK8KQhgk5xNJV7EOKKL54UZBZfdxjKlc2
WWy72yq67n6P5RZNQvryUGF5lYWbh0FafaV9t0g6iLexQupIjYEHLKbyL3ZOQn4nIdON6FeqUtnU
cRC7opX3P1RhQBbf/fCmK1RVOU9iOZx5PByRi3YSn0AGZZN+UlXf+W09XVpH5Lin1wvFTvoQQq7o
dOAOPg3DBW3CmdXWx1F4U/Pr2+rH/Kv0MKWZchkO3wBcloepVkiL17pj81FaEjpaQFb7s7aCN1yA
zrhsG/i/Wr2nGAjRt2tJF52lwncWaIzdpJea37e8iLSHLSNbjpOfKXfyg76kZ5ib1XZAi/BBFySF
jMFNiXgn26bPCq5OGzoX5D73GjYe/FjzH3kLXipnGYpmIvqb0YtUheqx5RFFhtj0fTP1kMz7kvyC
ltB3l9D0P4p83cvJEdCF3LOYLo90tXFAmm/QhVM72/zPnuBIzDDFE/huVwY8wodwEIPHlqhc/XId
iJ3Wx9L9v9Kqk8SoPIzAhgI1LebSuVAKFi8qmy+TXmc/EatnoTu3UFdC28tQHOD/6a9V04Z91nmj
NZ3LxB2BLzbXiO77GOvTR6u1FDcIeCPGXMTSh13uW4KdOBsCNTxAAIrP4jE3Fg0lzD+di32uFPam
Rq+u3xw6YXZGMWNGQ41h2jfa+5th9cHRuyxOWZB0ectxDMzC3U/DXbvRCe1PppSsMSOQqea+QJvI
R5C2eHb5xi631eDHzLPSN0Ef9C9yQVAbyvI+deK788H29SwU0fpIj5gHBb5i/BfnGni12fSNO9CM
9fSGLblsrV91YS8qPa43jQ2SMfzVogYps+ppj1xDhzDovkM3Z2ielQlNwVtP3krfo3ppC2Z1cgNy
QfQS5tgtwnXi9TfgdX1ppNnBiI5ARxtrQT+E67G871Dp6CUJ2LEjtYQOeA5gvdb3IH6k7Cdz+YNO
ko0IhlklEphQBRP4vur3hXQfBD6YqSOyW1n+DN4Hz6ftdxP+b2U/QuWdYavbLvhTSmk6WiovEeft
7h0s8+pSrhrVDftCwk+25KIGUAtqeChcH6LZBXCjwCE0ofZa3okyfGxM26ZUPENYWEZiRUd0v7rh
fZsv1Jk6NgGEvAWDkGDv2SoztQ/FL7pmwFO3F+2w6Oobb1+ody91NFXEHLk6LmgvagqD3zX8w2dl
+f+57FeugBdht0IFPCBT5+P+lQ/nMGTq10jJZtKREEGE512603/eAOotDphn09w0/fP5UzQbZx6M
ePVYpscybLcjI+ao7f7QrNnQpwlA9sE1aYFk74DtXYyFL3y5K6QblbSJfluOdjsr2QZYzbxwhDZu
ftjY18Xn3Q2NrMuQDaSwogZpZv8P6PHhO+IxVEC0x2A61aOXxmjcV4zyiL+bHdroXWS3bxXApsTn
0sIfKfmSyUZdoAXuuaNAyYGu8634VopHvm2lMyjY+ldFU5u8dph7fpN1Xrz9rRAq7wKRfT/KmHva
N3Z/ufSOKXTS1Cge/Aktbv0yq2R2f6qvLND7DaMABTq+yk4vUP7Ks8Vdtdkdokw2nV9M939cMbbl
2Q8rbK/pkd0flYaY/f+Da+QY5yd9Nj0cI8yyGvqRJ/+wHfPQB9IM9ad/SVhcQ1eL6y0mc9wbRhnY
KADWnrtRU+pkWlB72nrXGHFLAImaLbGsorRuBr8nMy0+sWBrbcPly5NXjs2FzXI8aYnjsNLCeK9N
kzCMTeqVdPksP0Fjb5h/053Qt5FyniQQNVFgZFVK2TIhT8k3fMPe/ZGQQudhQ/Biv2JjeygpmAs5
2U2ZQmZEBCy363u2IwiaXLdpKStSRGOiXIdc9+12a2UsyO8TXplC9S5RDa55ydcQvF+GvYzmiRMX
xckTlFyQUWpQpKh8pc5YrH5THismsuqyDcGWWD7dJWCX+JlxXJ/wWne/57hwYRKuPFE6JagO5Jba
6VnOwzEUQjtQT4vlnnnJ4HirfZBzlIe6ZJZbLkd23Y+YjXhAQgBSZx57qyUWOCxH1Z3pt3OR3ph9
EecfCNynHvphmOgHjrun6WZNeDf3RnBGpyl4KmzmtXt70HY1r02lV8ulTrsYKJi95sqa4p9eiEwp
K9yfJEagfbUZQGPEq5wkPK5rHyy6RicXa9Qo+BqMEOaN9XEbDhBq2borddQdyk9EAEcK7U8Sxwtc
u45jUMexXmb/DDyoUJplLMpmtSv0RqhcP36jcaA6Da0aoancKuq/uIelnh0Scuq5vlMr/HzKDNVm
VMvxv4+P2ZRAWreTKlib518nVs6KXEQy5h58ixQQ7GCAP0hFtDpv7oGseOcqBmgJ0CxWjNq2Vucb
rE8yLcWoPKVhpK+6H5JnyXDD4M2gCTHJ2ndoWWKPr8NGF28ZEf9UZZXoI4xoKKXLCf3HW0HK8+2G
NFVvbXIoNnEbT4j2eyL/ucg1ysDEUqUbUvjpvzPppONBz1XEHhwrrR9gyDD90b4BfQ4Dq1dlffZC
uxb0d/aSbj1Obvf/DA8Cz6Fxf4K5O2wAI+706jVq1JXSSheYpKY4/aVgfQ5hyVE681dKMc6TFcVI
MD+45GrLCPaF8CAftDt7m2XzFcEBZeuNFebdgzOXsBVyzjVSgvrYXa7PaXQpHdXvTyPWgjbG5Dxq
zyVhj0uxkSp+7Kh0JUB9LVoyMZJunbRc+pHP3xKvYHNk0wwqQQl9ARyDLJb7tHlqhR5ACoaBIf/7
HLjMmNMd1wQk/Ibg+bgwkb4hFON2HwC91b1w/XRMkV4w59tnAh3vjzelfZdWJ3ho8daG7rhqjTP3
a4CurHxfNRZJ14Fs51ZAqhMDpWUMS2+siNPrp9ST3tzf/umUU7ILYfcJhx0zXYWbyICM2c4rOzaW
zOHa5UTCRTyICcPdq2AD9+FTAJvooKIoKtgrNW4dcv0kUXhvXZ0t+LeGZyEB3X1IKxGmr1gR20YY
2fwpA7h6XrgrcDYwFSAvHxFn5CoijnWsEs6YvFxa44hWwrxc7dO2Ex2y4F3EwWkvslAW1/H88EU1
ykgZxAdo2psTi0oXEdU5E9Wg6NEPNInVQBjOd0gp1aOlojxk2whTlEJS74BT/MfRDjWqcfOJTC9b
/lk9pWU3n7lyRmVcox4dPnqUzUsj5pKbZ2bclmgcRnSk2acsUkmkdcrtLihMhmHguc/iGZNlWuf6
f3RIsUQfN8cGNircWRfYlVU+Jlt38VGY+zYzCS8obNdqSKJzJ4pwRenaDGNvdq31TdacZ02Bnir/
nVcWgFClXJ+TzPNoi62C4jssvYgq0rB7ixE8E4O7VGkqLD5xQPBg71UGjGpawZGP8hzxp2dqVIVA
BwKs/sSsKcChe+60ycUem+ZvjTOYWGu0JsgG7NYgtWFBbnCOf3fplCNFEH/dQyhxZwzQ73ZIRQ6d
hbv+a52IZ1ts+6zoYTl+x1bY6lB+ax4w4vhWOJU0p7GfBsmOMwhhiYHgtf9QDl5rPJRKVH6z7T3M
C4/9+wmoGv4Iq4Py6TXYehNC7QflKQb0ltv3Ux2wspJb8iX3aFeFlTM+FKp2m8MvlxEEnK0XxPby
KDOlY4vyups+gEX5FgFivO0sRkcsa2KrM+O5WtCT3iP6vT18CdbN0jeexK9pw5hYWL3D/aQm8qRG
7lNjRCmkSqXavMgptPhTUMAN1OcZHO9tU4fsbmX3ab6LdN/VwFmolICT2RdZXFCL6hBqii+fRNUh
47gV6m2J5K3/0CRjGbU7j4DXP3eoYpAW/C5F4eUJ3Ht4cpoqJ37kSVmgSHu0Ezq0F+cV3/7a/DvK
a0KTJAKx5/VjrhKEWN+JpgETuiJ9FIGXDsuFVSxtkOPJwF6fXKbsoO/ZHB7Omvq4VFAy2CHZdTl3
z/hygZ/ys7+0SpOxgcI/At+o7wOF3D4RuaNh1mzDtd3Nhq69iBAy6tEZpPCKxNwLB3T452VqqhWb
fSJYJZrhPtvgecWxzBSGE4BLexI2umGygv0J7jT1A4tULc7C1m2Cn43zfrLq0PKCVembR08DfxdF
hE+thURXC645ak1KZyV5tPMRuJ6PLZKbTdaZPoBSKkm/BwVwiEheekw3jVOQQSPTSMPaEHEpJlS2
WcBpBujQQDhKf2rLGtXm9MHRzyeDnnLDsoBVsY5aNnqp4NBKwJESeMN0PfU1uDNRZLkmOWdQKm6y
wAU7wqq2Vh3JJKZtUp7oYEliIieB9WHVMEWi+CbTBBe6Ocx3DAi4nHMvYwXPePwhlGQ/eK9/b0v7
P0Avp7KSHgQCf8XSJAjRJv09aU2v0i65tNwzjqA59TbwA6CHMz2VcCf2VGGQbwvfBZkLBhbH4fg1
9VTMmV9cr+9c3fbYasu+2aMnweCSCkzPk56oyDWq8ImfHdkTRCYJBHBbK5IE+r2GZbYoayDREVJS
o45yAywuCvcTKNsV2q58oP3hgUNKBTA2mcup1GgnLqPqLAprNGUUP7Ibf+zXAbfEgFmUkK2y4iDS
gq/77/rFT66lcNxwcP0kOEESFFw3KR/1DqLNkxIAwPd2wA5qgbwsQ+14D9fR5H7zs4WseyYfdsRv
VYPghY/HGwpx68vFrVdfIuffIKXktsxMPFgCfUvsxkdvV6lva4kHbgI+drlif74qyklCXTAAnFNM
hIlQEkpDnSet+CjD3ukaSIC6EnNeTjl0a6OfKOdrzZFaSiwrOP3DZgTI71E57OD/KNunHsdvniMF
fR1Un57nV9xn3IFX/HD2+K4LrhZAS0xlOquEYiVTCjYfNC9tl/tGPldTw38SAL8xlKqRTw5aTX6Z
Ln7Z4hogmHdHUiYTMdb37Ms35WoGguXYxdWXqvJwf17X+Cs9rWifhwJBvpd/EmgKO/tLfhx5cdPC
qOoLy5dMpe3x+1THj90XMQlNsDpngQxTVdk+E4IWJEIEFOCq93rsz+A2P8JAEoZHR9JHXIR7Edtu
Qi1QAzB5ASZehy6X2NVIgLQXTmiew8BmvlP1AiHJgJkysoMVi6aDqhghVD13vWNODNpx+LrHmlif
+bhD9A7fe1KBoA6B5AwrFLsEToKT4ai10VQtgb2zsoEEYMCDSzzo7O9FpphE7mp+SNXVyiQTqmeg
S3mcdg54myECqNOzeEqIJfOaejBOizTf0bl6ll+aaDm+pYysjur8NTp87kCBx8YxvBGsTj8DJrSA
OOGV7KbAY2YSf8EMCimrb+btdfuH0xVu2Yfrby3iMK2AI3HXZwFyIcc3TfRiLilnTM5yHaYNiJM4
b3xgoNJnxYNK+r7/4T8Hd0zFU9Q8JJr+4U2ad2prXgHdFYTYYDjyai02qNp6zN7rlWab5RMHMMDP
jsAQ+NfDFmh1QZ5u0pz8w4Finom2/LI3mfEd+DOkwD9qXMHRAt2sEd3ImoWaamXqgqZ6NXzE0EMs
prrftmnap376pqFxocNUpDQDbMD8m6wWlet2qBl+fdOeHRdOjDJYRi5h7HYy6dBxrr8DVwTbu0BA
4f75px4YQz1N/AVjQIrc3rRh3G7IzqTgyPAq/Lm4EsrTup/C9iJZvFEmI44GcUIYTNYgBDaRaOHI
tf44SQOfAO4lB2sUDOMYbGt1+K/LAeyvyz2pmepki/6fnqXChXoDvUyFOkad8E0nyrg9n2RIrEIk
FL5xKasO5riGVxhT3VN6uX8OqLdHseX22rGaqMvPzpMHA3Et7WVfkHOJHfN4n5MFGQuAfUerk3DF
DGzmWJSK+Hdun6+JojNK7IZJiv9Dvs23SpxZtagzbSMFdrS6ClGT9BXbon6pi8vLVtKc+Vfb4uWC
A4etsRkAHqP19fXwbTBmz6dd61BDQ/2+CuIPO+mt6j3Uc73kBoCXB33ooMyEHFaOlX3zVMUoUYrk
PXraR/KdlZIXqdvPmq7RcbTt8FZrOAmfMeNemHShHoZu4x6Vlq4+kV5iZiCKMlXqRDX9iblNZwVE
5liDfTxgS2o2Rul4N5NfypkdauirO/4NFUXcj/DrFJb1if4U1pNmkw6OQeaXXnwjvXLbw1PpSx8i
TfXiKdsrBsQhXx8bvXqY2C1WA/HT2T17lhPzNi74BXVbzXybvH7y2nU0oy9qEKTs80re2ug3Wyfw
s1Fwb3LJEqwN89xO7ZRn+dkRcUSB+5+vE8OllahHVGL4KENcqZJgSf/5epkrz658zR0q5vud9xrH
2KtDSAlZ3G7P+C6zlX3F6cFYycJ8TUONVuBcSoEvrYlBhfY7Gh2SRW+KlpQajxkXAXxNc1ftJ3yi
0xUaI38ixyhdSmJwAqsWwlyQ1L231WxoF1bBuAf5c74rc9OMxGkWglkhkKdRG5ayyFk6x2UO39EX
hFk8zCNyQdpqGfDlsVjOtysN+y2G52mpG7WOgnBImZLCPMz399lDXVxGwBK4E/b5o+bI7N0dS6Ip
5u/lEhmf6XrvwLqgvWW01qgW1A8twnMHorim/2/y1c29sKFDE9VLggZTgNr1xUt0FDb8zVIW6Qo/
ihEXkYgbwFEbPrayJefryVZiIbLWwHT1xiPkhiFE9aycCAEfbjAsdqjOIbP54oXxPOP3o7xFlYt3
yKjrwKtJvl/TL0ARrKBXMZU/wD7xftKxBwCPAWjgXWw8UdiVdzvU7B57HYpG25EE1CbSsTp6NmGe
KFDKEHZ3D2xrIkSDruZ60SbtlxKfV/2NHiCQdEo/lzx2sFfrpi8iS6V4vnZ67tyZEMribfNr8B9p
ABLh1E5BEsJoLHOvwV6Iz96JbktYkNeJlxnZT6lzZFKPONKprk5irCL4xUvEH53qv+KFKDm7bGk3
yLbF0L5oWz+sFvSz0IE8XnuBSAUQglGOQeub5zOHVLKYWUyGwN2X3HBet3N+FL3Bmxp/mTr9k1Nw
pN67vgt1736onAerx+rLreIxVICEuLqFBXFrw4lYLDSQ1V3nF2BSZehnIUYo9ckKti5G56vLuZc9
1Gh0ydV123PKnQFobRK9BgzcmCqWB44KgOoKDQAxA0W2GMldK7uroyN6FnabpqbW4AEaHuG8rIHq
BYEH3uBj5jtbrDC0GLUuhHppumu7QIDgsm8N1a7s+0MdR1vbKuXGNngg+muOSbi0o1LD6ou25BWo
3zyNtAdIYD+Tfj6oDoE7fNbdwlRUMEQ8ETOa50lIY686kxaeLe7j1JGTPxMu+EFOySjIe1mYSCC6
Zd90t9npj6gRW5VauChrra3ulUfDEuhht3vp082RTX45ViQfZV53c9P1C9yAVeJko2O4gjPdtpwG
EFrjRcl2Wejh/sxuby1V0sbZoOKEdhwLVpx8g4au9Zmltl4nhHw2T+DcEUBnB204c19Pfg7a/Fpl
NxPUCz241VwKeff51mMoWSO1gU7I2mwqH658llU0jC9/UQiClcTyXwOfYIQqckHAYL8W808ybmbc
+4PWSVGPtEck14q3fZD9cBp2YuYf0KXu7pKyRLi5kSL/cmbINoHy2X40okDqCPn3OeinU3l1JgL2
VdSIdFtUpbF4jag6u/ZKh99Lw6WZYjA6SICtcMwGiYElkyeBvPxPavfzhl+g2l1Ht5jOoE84ebl9
vcgQLHQqfOaAASNqeOb6C+458fZ6X8ZtezheJPFsA1AcEPM9ILl6ZoE/CQNgUC5JmFJN854WVkyC
oGw7jnCI8f50Z/m0xe/ko3nBTG7l0P8ToP8uRUQGv+upvV2FfiPoA2FbCPRnK702F5Lxs4cgpK7j
JoRYZM8gtr4S3DBWhAG2OeAqzyaop8SPmeXxNYHMO1Q87eY3c8vpHeZGsMDssMG9/pG8Dp6JzWQ1
ODQ33PW+nnuFRuLSwgstrqNQIdZknDEi015EH/wirMwlflEVdQhuP+L7DAPE1GD16imil+GbaQ83
xjPyPLtm+/78wAb2q9gb/Gc9GN/LdmBfTKM1qIKu804GmyhW84nrHnjNCeWUyN49vzSS8P0kxQcZ
Z0fNKoNc+rHkvT0mnpmM53oPMAHUMaKLE6SUEtNqUESWr3/InzCTD/7ytb53nRF9SNVr9Hpyjsu4
Myi5McLC2Rp9LX97Rx9bvNyYtr+T65S4w76NL6siM6/oTNoDpKiPFyWKGGxe29j6LAvPLVTITykZ
IK3hFgxq6Bsprn0r2ul6oDz09XZqCuLGsIOFipdiXbWQh5OXtcZEWu3YGK9CgVJlHPXZvrmSq894
52ZFd0bmk4905jAMbAXdkSXsKq3zbABMaGHj2gv3l4bp7lCmIkR7surR70mc/Sn10uzHqd8Wlb3V
R1+/rr/Fj0IwQcN0R1YHtdSJ7TUYSBfICukuIXIFor2rqxoszm6Z+SykTrv9E5gyWIf5v6dHMro1
/uw1Yd6waoKUn3fAWtbTfrb+o7nhJ7LlUGA5ubuHFsb3LZdrwYzCAOKgPOJWAD5Lkk4bS/tnQDfO
6o6FBnoOZCovbrlLoHfBvi7Exm2YMG6ZgiOBcRKAX+HqTL8JB4TD5SPiC9u8kG5VM1nbnnpE2ncP
s+Oln2frsV9oISETnmJzjDePV5uKDWlGcnHWqz6xLWFdHRzC9mGnlV3EyUkyUUXg2x2NEBkQtRxb
mvLtNKAqAqOlv0Mw76KUlB6ZWSKsbzeFdNhrKbt2pICsydHTGh0oYNFph28Az5sh9z0JfLnbRZZ1
OIuIS2zqphol7bcMZ5hgS4sd0oIXr/b9K2eriEFQXiCwQsQsOoFNlr1CNXkX7zOZe0HtNgmGzSWk
t5gNI2GfXJLplz2r74egGTLG4F3xeT07oCJ83Q9eyUTw+btQ2R3oN7yAxHLEwtJ05kQ9eiCwjWXc
7pKzRj86fWUTw6ol9WYNRrf1rwewUH9U503udHB0VE5IsG9WnhZf7vivxk3uQM2hvKTnN+oQkaoh
TzIOzsvvfTKqM+2lvgfjrKqFgnHhzuL5tcQMq6t5NEZxc0m3vWvza30+1QjdZJmZTt06Koh1/2Go
ToaLTHsf4r5sUgm8OfRqtdA0nch5qTzCH1ebv5Ct48kuObWwFYe1nRj6UhRTEbSaWVTxjPnc6I6L
6U6WvR6qGq93nzpsfBYjJ0SeoCzxx442MYBiO3IelWl9eQqjNsgVTeX0BV2fdHqwsFdqPnp9ZxEV
LNpb6chjz5qeOKLJo3Ojt2mFlBuBn/X1trOb7nvR0mUfuWhRRQMa5UdkhQ91b09+D6iGqi7Ze+tW
4W39uF0MWziL7gsJybauMiIPdqa2EmYCX0BZX2iv4MmXErHpmyhP9/QPflgCH1HJeAKpzcOHZoBv
7Kj9Yskp/aSbn+yRhT3dqVJqEZHH9MWntcJ5ePva6FMq+zzrvOZm6+BHXka5G6UaGVWKugNb0MXn
F5gn0MGydWf1I2SxpiC99jYkv7G8U24AyjM/RyNS3QnElzat8+KEy/KfScRmgN15DgOPX7SANeD+
pLlfwme8J8NoAB5juCzBWA+aTnPqi31ZYGEUCs9JAA3MCklAmTc4TBFL+2+nQWlLgaWVZFpux+jq
e6TIYzr7s8Rq1TZLgFY0GmvlA2pAfQazezHVtrb3XOPhLDwu8tQYDIwFSDq50mQJv6zZvNOeLzFQ
oNO6/Wc/vErJISgnB13aomsAgq2IabMiLHoaeW+Cm3ivrRN/UE3jj2ZdMhrlyqSoiXNByLJZkK6w
FkowbPPNH/kyaFyn8IlN1vnYenZX7+I5zSa0YK36ODA9GQ7IoDq6o2PbXP1g7TPNJkL4vwyMhwoU
iIMBAvju20PWJ8+3Tn3tIJYHvS3DxBckDu2zzLtlw+wS/0AqW1B4XU8fI2D0O93xo7kSqQmj8kYB
Bol26HyZ+RAHFl4xe93xrOalvWlSygwhnL1cQ+omKle/WAB7MYtDdVSzbLCIXfdca8jSnzOItCDC
i+R8Tgcpo52lOfmqvFyV2pCuF0X6vDu/24A/dm/s+VC/0Zr2z2NMOQODSE2d+mZD1MGW2I/RtBjO
uvJBcvX2zx1BUaK3NUlKhYMTy3bBtL9/+BvGFqcYcyEQoUJdFLft/HXXs2l6ZjoqoPMe0M2xWYtF
MiY2s4ObWvg41xny+VwS2HRLdUvKSQr81Wr6Zbj2yBXqwoAcGzL/Bdecl2UU5E5LqBziBjmid1qI
Tn3+l7cogNdmCRcvAG8bDWWPgUcOZFAAcnlD63zlB/4npbvQyo0y4PmymMrCLcJTroj7+1ct3Ld/
5X7mb9Tr9r6iiIczsYgq9N4e9Pu5JqiyrVVEYNYi+kSPWXz5/MbX+3sCEyHjvyOGr0wcwFf94zlW
Om39zPGo3uMPC8YZG4N5QWp8aCxTfBE4y3r/iHPtX+D8eKq5BeFRAtZGh0mouoyKU/opYCKvUwfx
Vr0annjYkNOALDnnKvZEXpyUyyyECcdVYxMxX1kBRtWt21Ul6YxJoZWNwsq1L6HOflOXazWZgRUz
WZHIbrzQnHApBohWMa9fCRqFTiNoJIzTlD71GX2yrt6n2nn1I9qNCHi4qyMI0jB+BhkptRW36uXe
Rp8JFd2lzdsmHi6hXvivx7IZD3iB+ap2CH8aUfFvCvsQNhpVvQV0ANYK1UB4+dEbuHVQ12z+HcPq
qrItSsus7Dgn78Dkz0BCy2tGYDWczkGoooJ4lqMcUDDyDHNcLSZUJ9DfcHr4IOq9yFp4T31oYEp/
OqXmfTMw3jkBwcyvt5fEH7ZzQkeucPfV6uXeIPgpNC6ydNXFQACldJMsy8vxNLnF7PuD0W66tsNW
PGcMwKQGruIiUMpYWg9PspvitebCy/IDImkN/NdKqcSNK/76BPAeEyCcPgx22El6CgUPm6jrTh2H
uIEEoa2V05MpSOBSDv8DzKnAcntt9za/MkuM6EbvqVtjROzxBt1hZp2xdlFSiRpJE0CCSA5PzMTK
igZjdm8gsDOCJjNCXL1RJT1PI4YjsSAYiz1cjkIYmVFKdbFSHfImi9EQA0JP71aKIHpGk0micubw
Oc86exaPteiY4hfPC0TsaW7+9cuwUCCdolRsbEjDTQYzRrhPVdcqDgHSY4nD7o09KZo1AjA8mNst
FfuGTFtODvywyGljN8mNac5pi2tcv9QBZs7tAVA3cwmpovwAbirOPpx+hfhSk3uDzom2QvWPYSZj
SyET/9kLqWmyT9VN+iZQU4fJ3+Il3ruo9d4K6JkzOKSx9KJKGKZQasKsbkqFIHIqg3m+hUEG7Chk
Gl/NXKF5O8TxSNgXLfVIzp15yaVXlivRp9m9G17SyhZqx8TVLs2m7pphCR+QaKX9CBNCqPUcX8mU
u0FsvjR5k7bhW/ess7Z7kguz8GHcmYV654/44/RVTWKYgdokPucTFuQzZrIsclRbx/AhLsGuq3Ax
r8mBYR6Do+7/8gxgPuGBTITpr50fs+8xgmNmWouxoR3dDwKTGD/r4JzYKdBuIblgSIlH2rm5Hdnu
iZ3AkzFSHopa0o8r0fd6AYnsq7/CsEv0CWxbBMNWkSRZ70twVoSlpthEJ3ZGFk2VjjetSYYT57cc
jocLBYSQ5bd4AfPAfuHJHCMFeXgZxp+b7GcdZshJFYVcX1cm13TJnaRAuovqt3pzK/nGGgMCDx+p
GbRLIsBcj2ezt0dK/tzBH1+1/tYgXvp3xJWWcGhxZGZUQfxI7kjLS4eVR/OrYnK8SRoEnAjMlGRf
J0dSOmmWruW9D6Oust6ey0SuV/EVg1bqBslQylyPgARPEkkm7bhL5aRuztSjDo4fRtOHZy5I7weY
kPo6ZTqIUjKetD19Wb16v5ozqkhziBfWOHgbbZsqJfC1/3BuqbdTSBqIorfoJLRDFVq2OFP+HkmP
nBUuIgwnnydlZtHVUgRq9TwG9tuW3TPwGGOsot+w1a8GAj8xcx7p5SEajZWeLpZdU0Vd18li8/UM
uzPKUxZPsDMGEieZKYcdk6wcVMFrrFMJtCkzro3uUrfphzE8xv/iACB6e6d6+w4uvwIQwoFdIC0a
i3oyRLQivQ5ND5/tgC30ztCm0f9v7uLftm2KFWIK3gnKKGy1tKwRQFQdSC6S6nmqxTjuQYSnTYQD
SJ4MUFGSqk1bQ7Qft5YhCpzOM7+1ae9Le32P43zftQ94P8KqeicGPcZADezqgHkGx3p28QAttj86
4pEX3WVfGirwY0xgcZbRN/QZ2cQBMX7PjnhRvotUo3o+tJM/cAjCifpi0+eU0bTMaE2jjfCrBetr
TjCZeE1Yo+ui/3z7ExqRm6divvob1fehFgRDZ7TYE4/L7eZEbMhN9UnTJS9dLpsEU29w3cABJV4Z
rNubiQpxoUUL/++GvUAXVwC1K+hfjWmBItJ5YUuwQdOsmjJS/gaWSEnPECqk7aVpbPFsYNPfXj1L
inRqdWhF+OXbUdwZeJR5NdB85Y0Y7NIdLiOZrmLWnDazc99Uu6Y3xiqCZl57k2cRw35djjDxo8hU
+w4JJAbmRp2Y/akI17UU73fu2QjrgXx/zde9e0osbpVLIHmsoHDkZUGrmdG2TijhicPtTQlZCfV2
sZQmYRiZOIumJllEPEVch5dyDIH5OekX8LRsk7ZV/HMXvjRfkCI66bwi23I7rHrxg5Lfzy7Uk2ug
b9AOu02NkNgUBtkO40mwZ7Dga9J55m1PAW1wug+uIi+TOJ8CC1kHKVR9V7r1Y4mXg2SIzJsD3Gkk
dbpDyPZfD5hYWry0B+oWAVWLZnMxAr83Tj+HKi9/pb3E0z3rufpEArE7EQkicrokdiHU8qT6bnRj
d+/KL/Hg3lYTViQVUi/JbYfXGzTr0oVqukt4l2VykAck/1yHIVKpC4lLeE+S2HgbJkkB5+YcmGfU
FGq+IWvYRHXnwPl/ruHoD0u8jTXzu3vR9R3psW9AqKL6W0sKQ+43g97Na+goKc6TSRENI4wHU66V
UZdZp9oaycihk24WLUCA/bBFZMagLZ/ulr4lpdbVWyTUTChybJNCh1Y7H2e7K4QXT7W8BbzrVPMN
9GsBDxl713veWr2s34ftn/+okclL5WqFy72v5NSlEx3VOGjVxyHRqN8afRFtRYXXM9zuOqR/uF+p
rw/Ur94jhHbW6SAcCiHXM+JGTQ1INkRkUDKBKydUshNQ14XWIVJoVaTys0/TpHCcYbQNq5D1ooAl
aXRBjhDwQ07rOZMrXgxTccC4RqcD58Abu/cXHBdB31HoGHQ/1ERBBj0eH9J/a0Lh27BJPL412fr2
UxLIPqgaRyh2u3thbzTvEioJ1BxmHc1or1gk8wnxvEPowxEB4zwasC5mag3j9xlZZHfiIK/m6uO/
TWIB5LUqwMYocvCW2k4HjYwBDskNX6Y5YfNQF3F8Vq+BpsLzRDmhzOrtf3FIb5oGnW6huRWZo9Kw
yFlYOmrd2pO+Bip5sndosAiZ9lQz9FAChsaFdNADjndW5UaD66b2gJH9vme7bXXanrfEVCker/9D
hhCCGWadcJ5DvU/6QrBk7ERsjtDBqwjw30HEH58VrVjTX5LKaIYLlntQCImhnWpfbbJTb4z7FuSr
Z2tpoYnOO5znAtN+aQvoYcVf5JiB70+80qqgSj5OohkhSftN9RE6Fn40uj+gMBu8fzFF5xvvLbHa
xSLXVp/1VKc56PY1J/iX7o7leho+AFziOgV8yqTiEjmstqGspNHNdcu965juCgTPi4AFuKk/+hO3
7uZkSKUIwkmOzgYwglzF25GewC/V5SPn+SgoWAgTnS5h3xu3JauMOXE8mzn0C/xzkH9C61CuRgko
uSdKEcFEr5EXKiPr0dZ5NvQMz0BMqqVRIKHhkdlDrlL5rw//j4GDtoHsAjr0GwDtFFqJc99Gq8Fh
Ajd966Stme5v+PLFtMrluSmwKLZcokMJLEA0FTuzh3ydNVzNW8kQCy97k2K/YFWbpuYMHSU+GcMj
N41Fn/9gjRfjSnsDtGWjUtPfDRZYdn5LbNUP6UVtmI2QRiqTQrXNQqUTq7IldPOhTlSyRNtZvmdy
YbSGsnwEm7Mv+EqalpUQqE/vgjoOa1/c9MsfuxRjVHLHMN7dPY6zMcyruI8YeZRj0CaMAVC8UpNb
DPNnHBSDmP92KGZVMkyt+iI8G53KU/lXY2GoN8w27rU4FGUBPtrhKE/ikvelTMBdqURxnPaeB8EP
eIUd11knH6M9ddrL13wmTTHHXCKSa9s+0oVE2l8tvXTV6fCF354/Mh8huxyikOFgO55ePPNXV9A9
Qo27mx5Yuq50xiypcad57w0dqxQGhiBMQ+6EpRjwAO6/zI2N+g74xk9twiPki8QkxnpcsmbCQEHW
pgIyYyRiX4EdKz+zUpvaF6b2RCL30bYlr5HGv1qCGouw7mcy2sQpEi8AN4PpJd4ov0mW8G1tYrL/
iLTyvDmPJJKY82Jd3gBHOzvz9KKWM4AIJXMmTlk2/fNg91YiLPsCakbJ5br5WQTU54AkLZhyATmf
PmdKttxdiPp8hwhKM8xCtp8gZrjv+eTtjMDOw5hcKA6sCyOiJHNAGN87MMQkWASsLF9L/QP1+jc+
6Z18ve6TIVj08mR6oYBKfavmg79j709Ng3fZPzkPYsZOMF5VRHRbJu9tJaXKkVRQNM1YgxC8Wxpa
wai1t0/9SdBlYVMr6p0yrVDXGagHnIHBDvuN3N9A0M7dF/HTrGyR+ayBlm6//q6hGPtxwv2EDh3J
nW4hjRvwC7bR3p0y4EwZdaUomErmBxj/eD+07owNvTiuoBxwW+8RwMBnh8mpYF6dOZzsPeCvJDhl
Q0xXTMVobotxPr0tFl1Ld2qCKGyFnAnwn0vs3DwiWP4zovLDJCWaDezINt/cjiewUxhR9dnwG8Ma
0evgkGXT3GPcXW/VhfJmXxBIXq5xlDTa6sq3NzOqYbgyrdhRcTXsA3ct5omO33QONtyZSgC2CskD
XS4rzqfkAmQMXKVWyZ6NPFhuiFwQpJRTssPts/m6nsl/EX0pUZjJMAVvuFeduFbXJlWWqV4roODA
/DuCNqtRJYujoahynPgCSOjAu4NDgbTVH+am7iLGD2HGVoQzVoF+rqjHDkDXxxw6hpyJNi1En9EF
9Yv2QU1ggEj6XsblQWWsuO1mK978g2q1XnPqobQszU7UwBshpaZFVxOqJGACl0vQ8diTcZouJGSO
4kUC9EGVvagg2G2jWiFUWEWOv2CcUuuu9Y9AI/2j6UUNaZh0+6XhNsL59g8RonndU0vRQ+oGeTun
VIi87Ty8hiKpdiGbkYQeaDIT79k+euP+sMqOOHRKpVAGdo4ZPqD1s2KqGI6rx2JrKg0r3oNQpFOc
yM6N0gemTb+Q7i/POWqiV998RVVCqk3fnYvBpLPZhVHaYs+Gy1Ivgsz32Dwv71a2Jet4uaTcDNyG
HhCfYVOfX3A4/phTeqphelQ5apn9z950HITmJLPkH913TyzFbjKzKOvDb3e0J+8eUQKvO6pPM73q
zUUBl/4OmUb601QTsHEt7Wzqfu4tya/g8T/sutuf21kPXnfCkgnYsRuxspE6JyuuhnmkdNjU929h
EIR0KBFAzkYCkeeXcKOnY+UcKCpPU1nx9eIDIZo3AZQXie4fKT9gSN2bMd2n9DGcb1IJ6CExKMSQ
Zs0/hgPJEpYhWhv07sFcJ05BNEbqHu2r5viCj3ppJKDuX3tACv7dn3o04mVUIhH44FVpwkU2o0iL
BkWDXSwQYKNi57NG+PV8jkmvjQrvTztTh8k6nXeThJtCcOk1CgdfdKwDnvitCgwdBOphmTGqYED5
3SqBEkFtSgcE9ioUwSd/1dTYskd4+AjQQ9cbMJxIvYMNvU42zqyR6h9w5kh3Bq/LTo2OIcEYGgbv
0lzYGABCo6klvllhdBZ+eIC6URHl9eWCswV+vJFB4FB7sqalDFOp7vGbluwxNKy0DViYw6RnOQbv
dEsLmOqxu3WZJ88WKmT7vYcBXtF5tyPgxeVshxFupGabzSiw0J837Z7y90XCwbNiddr9DSoIMj9G
l8arSCsWBktIzweNLPLg4ziTRF2V8EkmHG8GbXSVlNMxTjVph1vvw/ujMU+ir/T53yCD+P9SvEEo
BjLbZZL08/Y44odVMBrzLsPPB5yjqp+0noPBmemuQoXnlRplgmChBlrMA0L261oii55+5e0/1mV8
o8IJ2d1uZ1XVUCkVQugDpjn8mXbocLY1SpxW1un7d7aJrdGZx/LK2pz/3rIG8dtu1GfaKNGXHgf3
TmSLPMC9/JiGwp//RUvXsbDCt8xYB42w+Mp8xzNzH7Rqopj7eiWF3Svl6WNpAghHGSdCegDJ8JN1
rXhCHSa19tiOErdrHOl6slKlQDHxkvcx7b5uqMD1qn/VvvETt3MG50S7HH5VAu5sqtDEIv1i7ytj
HJAPleNX0rosN9Vdj74PsPiiiYTlICLXejpC+aUM2qTMowcx0tC3m52vWAydmEOy/9CGQpqynbDc
MBXTBMZsoTH2fVBN4Qctwm8746o50hP9EnoW8M3HokwFuR6BCIoYZCuul6LXkXhKyX6YDZeR3uj1
MLZ8K2764f4WR+yVYGj9VmvSlh3Oyqmbb7zH/4he17hhRv/uBERoRSW8uLM4qy8T8M0LJ90Wk1sZ
MJKFK7s6Iv2E79q5eqMtC6mr3Q1RZBVmRGmVx2fYQNopEZzj1y6wEqjG+1/zADszHzCw83gPUtMD
0IQl1w1B8K4WZYEePEFPmaCn9I+5IqZdoJrrQrEZ6O/zyo4u9U64clAilQgFO6+UFG+fG+2vD6VQ
dixKqU8UmPnJTcKU7fqAhU0OLWQFAaxPTTUN82x++//CJ/lDDWt5Ff6LW+ohjHa50TXZ5V3QZCe5
+wsTTDkkgvnnjiSxfmilkjJ/bUrMG0+JIfNKO26FVsm4yzSj6Ahdk/9F3nE4XgIx4c14Q0LvsGNv
oFiNeXRG16xOISV9m5CwMvjAj5cfCDqj9DVbKFGH1wrR7aLPBue0nxopoCXQoprAXU72PZ6cdIhI
PKqzKV+xxRfCgF2TDVaLNftW/wui/FwI8mLqpJZdmyEDaabzEuqPgVVcfZhddCS8KBC3DnP04GWd
nvUcV5RPu5/lgjGjxAoEWCNewJ+yGit/ls4vWGWNfRPDe0YmJ/S37l5joHU/8+l07YxiKlXVFTRQ
J/uWbkPR5qIR5nQmRhV11Io1BGOolrwGqbHeLHd0L5iNRXf4OSYiOR1mXrwrMgi2GifyDEJNbmVv
wqkY3Ru+srqEHvzXMeT/+dzk2RoRIuq10E/jqq7Eeew2rk2Yvo0TLf/d+js4x6pPEe0irwz93gH1
EOdkXek/RS2YVNVbE2cZmIuaRvG/ZWZyOnEVpdxjN+kvqPz/1xLsDoXs7xsPzn5u2wpO7mcc8ktl
BfBFLBoURGgMOXDbiwAfvSx7B/Ice2VUMYa705nVEP70dW2JWBw4BRJeq7ilgbOm5uXoPF+XsR/S
r+LbkVYhQnRuBsNreAee2zGcV4ghdZ5+hJZCqKoj1n9Wk8xML3KTH+2LHnS5fUtUyiZQUtLRuHCo
249J72ssh5QTufSAQJ+JphpbYT3ZS4a6KtDL+fZ4mJVpq/d6CzpMSr1/J+Nivd5XWMwNAs7bJO2X
vpx0QvTbVry/zlcRBolQB9WgxP1xiXr3a79gg/m6pefjTzu8GnVC9qg5XIrQL1cAih5UZ0zrBdxx
nyvdKMjnBWkFoYcF7lBmVStIQxtcHDERf9gJ58dovXodNAio/P28GEJLjL9lTWYANf1IC8CFG+Mc
YHVHINmaciogce0AvIpksXXjFl0jqy1Dcj5MPeIb7wqHkh8KErecpFbO/VNNfbwY7Rur2Qr61FpZ
AAy51tjvoKf3iux6TeZrmwz6QOusxQ/XNGZa5CYH+k5kUpaeNAHqE1UDGmUDdVpizStPRv4y7GRu
lBo/rwJjDeo8cUq7+1XoxwK1h/ZlLOMy9Hy+mkjXoxmA/ka8kv0iMO15x5eVHecMfDsTXWp8UaqX
Z38bf8OjM02iY3Dl/AT/Ac1NmgKpTtZzMbltsETYM4/D5Do6GC1zquOApi1XBmMMp6+mR3z1LUs9
YzvXl3Rl2vLv0Cq5ngKnFOjc/SAOxV2yAINbGZCesMCOoGxKsw+InikROjpOdXry7eEw+FYogrPm
Bv7L1KrIyG0YzOVQ0DRJ9Qba1Fpiw2VZ3pBBzBXfBWsegJ7kc3BKtupJPQihINE8uk3RVNOCISPE
Ad5VfZ3YWZIomaey4tlckxTo2NrhXZUKk4kYbZvNJlYbM41Mony9W90xc0A9Y1R+V/O14auDPsZa
B6+2VmSJFsDGFthtePFRi4t8T8rmpv7JsckpMKPAZ6euvPKt6k8wDL49CAMhxdhe0KY1ZhzCidq/
z/AtfE9JgHfs2UT31EAezqrN3FvXXCPBO71g+Z0SPfmKyXzkWJVZ2vNudoR1SC1IiOQ6x7Tn8rs/
C1JqLlryJjlFwJ2xBqaS59hA97D21wyF0z2HhbDDnNlIgoGt+aTOxak5BFo4TPBtgyzHWEyc1kti
9ocK3Ba+ILZLiuTCD7BDsD6XXRS09tPDA55FPgGymzlT/7jY/w33rwBIX9i+IGMGveiaZe+iZwlA
4iTkOOqCoZmL0K8lO+if7HrE1y5PPPHMyuCvjdGlZxZUSYSRiR3QdhBj796FggUeMHV2J+08U0ox
P8hj67h6Ql2kPb1RoYt1D9X96XHzfOJ+G8vGPlD2yMLvqHyZRAhNPTVl5Iin5EHujifO3eBeW9qB
iQL9T8fxwSDO0Czc/ZXw4HBNzM5cEIokgoTwbvPKdpCnkGb180SOAw9sEKqvW2oJQc0+pfrNF8YT
KAhSm6npLy0CKSs/LpUOnmOy+pGd3k3vqVZl0cFq7Al5ObYzV6qL8lVMVBWm857q86eo6gCCckkL
OkIoKcz80miQHSpKuohMNKUXUGHARiwZKspxqHutONjEwvZjZC3E2ljsS194iRzp3SgNEHSK0HS2
9v3fPwTMcdBX6M9WBHNldBJdgASZ2hGclSTYTYLnO1TUf7F8ce5wFA8XYh5lu6H+54PYibCdE+K1
MNBIq3T3/NSOxaPKkpG6BFk2l2nOpP/Yh75MzkOrQ72/rShmn7PRXsZlIoiY1p9UNmIu+zctxrcq
9CX4QjGG3LfqKqVeZT/atFoHD52z8YMcbrFNYcAKyra6YWnTQ1bKlVejT/2r/PCIQZuVkJxMaaLK
20s+4SsZiZcYbDGX6aCQ7CdcxOHbcx7rHp+slBDbuueQiBLn7/o7Qmk3WJEmGcGrpjB9dniG0VUw
S8blUt0j9FNuykMIZDsEgpvd/gWUQWhMbhGJ+Rh26LbNEHb9hsa+Pv61yu1ghjMzNZQZ+ISqgybB
48y06P0yBOcoTdIjyaXCEJglohlJ+1IgQeVGyoBGp9VTIBKv8but53qa1rQWrdPoku/oJR2sDLvV
DMdxynxZqAba3qRjagS2VNwYvf/YTX1+uKxf+sxlWhJ5e93IyR0TKpjr8ahmOJElHSVuel5yi7sM
JR7OT8AZpgmQwt2H0jIpKS/eNDubfm3qEAW27+lJgu1gvZdCPSrg2tYTYkLEYPoB+qZ+WYTt7XuW
4ehqk8PKd+5mpPMogBsEEe1QYh6vwP3/JEnW6iFVR+xNsBG8BJLwxk3SE7XHMbcjsMCuJGjKzB3p
tqJW97WLtDlcDj2H8ecmzk2c9fsGEymJxaJ3wUcsMaBZc7UriGkeVQz4kRWhu8LPlIWBj8A2ZKnU
TktAYgTMYFxjPrVKkexm7w3UvRvn7pkwlnJS4fML2QNrk8VF9fmhjjPNJthtkeep3lb3TtWq3LzC
ZfN65q2e95IdMBlN2jI3BrU5ZPpDZd2mJvJUy0zAG5S3YYMbz2APXLH5Q6fC9ZaoOzhyHhowAMJO
xpVfYUlUoImq6CgAD7Gyfs+6xFsT/O1LaoY671S8Du7D8D5oJeglPaLSXZiCz9W9Tn0xv1KOlyDo
kuZth8e9uD0+iAfvfBFeG6a/4mbX4U82oq7ZOoJo2xfA+ZpJuai5eaqpebhbSQ+v5D48p6M36C/t
pUYYFQEUYDXgxnHk7YhPTSbb6p4UNwnNNwjwW/ZZOJ9rbLb2RAHYEDaLMQ5z+Cg9cyu/eNrPebij
embc7seTW7+qVJlmVOIPLKM8b14x3ARanbWo6IvgxFYn7+6xoKFMyhaemzYpluh+rwM4mm6R8Izj
nva6yhu+DPiJOTDx9Lm69YV3mCZcoHFjjrsoLZDcV294m9fGWPWTO7QKXJ+PgDi1fYR6GSwms7j8
HUX405ASTA7a4IkbAlCyKW+/gr4jGYu033CraJdDTj97OtcPMhEO+el+LZ+GThNFbYF7oQ0FxftZ
UWM8yC/DY9Gg6Zd6wILyLx0/TEdyRKspvJ7DnqF5JS/zUu8DVGvgwW3xGxpRR0OcoiU2jfDHfWNu
kmUoxNv1wHEwTijNkYmbQFu1FdMUGZSgFtX/k+dlOvnKSdwsTK91u5hTHVhp4zrCoRRv4Y6SXbZF
gcs8sIyQuMkhV9uu/jfOu49HOSiLnFMFInjrhqd8lwMoIPze4zJYWiOsp4s5MU5Npv/qlYLmnCCL
HuYUosI9iDJPqhRd6SxwwtqvC7yPbXtNMGd8EgMKU5Pfz1KHg3CdE5VclfWK3GcmSKeEyfVPYYzn
fmg6mEgQbOeyjVH3kFkdYNRNmSSkn4OCrDW3yIIyRDq2A9rq7f4zmRB3XCDnwF0FAC+Jhlqmn4dI
9LKgTF60E6BFnbCGQiZgtKKFdCWfRNWzmEFi6SWDOBnvfhJxrbvx1zXEGcF6VYMI4ERwu3tvI8l4
zVP+4hFRRI+X2ZKRp0NgYS1JEGkh4dPNtuNrVGQo7c8Ixjxcl4zrPDSrg9F5ZP0zDr4OoeT91z2I
N9xdTZ/M1GhhPDf18vO7nCYDR5Nw/iligDp3wRPG1Q3SgL8+v1sG8ns5CdJ4lt2ijmDw0seDAGpp
4KrEHnGpEs5A5ghRZ4X6zXRjDh2ZyIdktKKFfftxAgE0QGfPYJsApP1jwjx/pW1+1c/k0bqFWaI5
SSF6KhG+ry6nHoyq4Nb/AGeFy1BDGj6tjShrMpP+JyhkUJGwpsjsEi6XNbGSpe7Za+0ZRDqniFmP
UUo28iUi8VNiE+wmkjI0hv3kPBL2tpUp5HZ9XDAceUe4Vl9sO/YqlxRic5l4izrwvmW2gFG8CwOK
s3InGk2QSgAj+fND8H7YBsui4qyMwqGk1qxmtjVG4C3czLwJYqjAIXhEAe4Nhi+rqPsukkUvnmvi
BRvAUavb802Xk5lafkcj5T7gxB9zRe3S7duJQSLHEX0tJBDBiAWyrZigtj9/zRANsDFXLYyqqC/O
0RZMExRZAB1n1umnkGf89a2f637FSjrICM78FlFe1qs3yBngiUgvDIiKUEx7YrtCaCBOavvbR9KR
OMFWcHoYgQ/DqVrr7P92CenRANdlYoXx7IbXFLLwM1OIppVemLPzI+ZIKbNst1QG4CMx0leRI96y
BJD3yMNc4nU7+/o6hfS4BTLbbQwZ6SlokghsVlvf0hbQFdxptF05qW5KKvTBizOFLdsb1vokvqCY
P6P1h/HHFY6Ib2TGPVL7v6P6U6MvUbC8UR5yEBiaimeN5i6mOZyWz8XTwyyV5DrivXnZwig4wvek
7PLIML07rrPJiHecoKW9ZyyZnCxLJClShah+L8O8AQq5SWLf5AR+rwBxQtnuAMEGI/t4dwZnDGjg
wf3CQXxMcu8YEon/Eax7HeDMJmdwy/UUfF3DX+6fDXc2Rau/CAx8IYAImp+DV9ulm6q9y20tiXWj
He4zbrpTPRqzE0tOAY4yLsP0xcg4214QV+wdO8p/RudO4eoGa14zQsRLOcD3fhyRra8T+/EznaXJ
yW4o720MJVngPCNca2xmck0AhuBN+vAR+2cETnytf79ClXrZ9WlD4Y8WSvRQZCzNOjYrLWz6VpFY
hA9dU5tJiTggocwsL4P/nk+Yq27J+esY0w4P8owfGTym0cDdIpuvek0Knk3FJvBWKfdBmpsUFRm4
QvXR7AcYvWBVs6/b6IpioSbbXnA/H0IuHU2YYiGv2w5j6OK8pF9TYgEp//Y84WmC5UxFxP5xe/Fk
2r3v7xOncgDVveRJxOl9jDEtkO95ocJ8tl0sGD2h7WjNnOi0e4t5QpbGO0tHeaqXL91XcdSgH/z8
fXH8YpaF9LBcj3NYHCDmiTKKfjndcVojeOYAoz8vcGPo35L4U97MjQA1e/2Pwd4ULbzv8aq1gQah
wji/L4HMSruR5vZWNYgrl30ZQntD2eID70WfjsQtEkvFJc1VnK09g+AqtAmzB1MxsOwMGaYld0SX
EOPJmn/WSdiQ168Uhr6tzkus2EWfO5OZuZDnFJmk0JzaLAgyUId2bFKtVnZzAyvycLxeKk0GnZ/+
HHif4J37Z69+DPqP+5V0TxPHtjI7q95a3Y0pWYdoLHdIujM7it4lspJKEvII7SBTB4L6xT0CoYb/
wAilH5eDsCXgH3WY2ojc/HwMJzpmJGskU1W/FY8n4/etZWDPmr0bvT6zSr50zKdFelqqpXW6jsn1
nqi9IrGSJ+xlXTgmmQlPAXsVb+cww0JLAIbxNp/KzguT3BciRcM5pEHUYM2dqI+/XfMkIgAKwM4J
CnnHuabpm3qpIJ+kUHdtVUSNiVPJeyEirDEGfBFLpEMPTCpJ/TwiiZjkLM+GOo/AKEgp7yZlCI7H
bRGPfx2aJXgN2qdLVWQcStMBVWtUW1tOtGIksCC9Qap/cektjuoYGYM3Frkrat8lP1PG7/ylV5w0
zXYyOX5eiVPQ1+k/bxwge8p4P6EDZ3BiPYthvkzjtkz6FQ/PvUeqXRPeqJNF2LIAZs11U5PY1NO0
2oKgkn/QnHXsi9QcWHzdOwqPe1fih5legWnXAo1ZuGWOz3mRtD+2fb0p8xq7ZEYXN66ZrQKtVDC1
NtIODvZ0WpY38tTAY0tiXyKeaN8enBYJH/zSr9iJY1Medk6/kQrv2+T2ez+zEjYIzWv0SctU2/cH
bNV/B3zBXHscJ6hjSK1UiyxUh6leyfnbjNrbh67jPk2DtXXrKQeJP9NLx5+uYE5WnpOBY3mhG6YE
W7e9Vf6v4OZhnW9kCz6oyI68GPDtmnXD/sGjHm6mRTqQfNvx4k/EDT4oP4KUhN+Tuu9xxy2qulo1
6T1OrI50/2Lmr2Dd89fHPSVPNrEVQK0qUS7kbUYluzXuwDgWxgGyyNe8Iu+MPEeI8ff5SAzSSyWo
SfKn6858XvXFx+At5jJFVKQRTTAapehJtnmbI2+Op4byUYaCrDFV5zzKganRsJy24NOWQlV0XmQi
dd4JDQqISSmTccFYzIVlYD7Mqdun2hGtPBXGo+1vQ6LlR3c2IntqlGVVzPTjp8/vYregZ5MAmhwX
WJ0Ot6dX8Yqvm1TXdQCZyyRr/t1MBsgyN4S79L7XVC2irmdi7uPYPiP74qOUq01uYQZI0ug24QSL
tv3+B037BmmfjmKw0LtJOHMQ4R/a2CjF2+ahGe0iyZusx6rTWuwoVAeVQo9c2bGDuJIB4RXbyEh0
pr0uhJ2iBxSKSt68THU0AYWQNinnu9P9P78RcvK1oiQmIc6hSjUTaQVkEQusTtcV8yHs0mgAwAfr
EvlEXjrOb7d2jF+puCVMaSPb/6DWic+CVmkearYiqas/yxUb4c6F+JHZZuPUmpG+kLYJjERedMEq
QLkRgXFR8r0ZLFiLCSZaVfjfbkn8RQ+3y3GIX/W7cpnZrBQXmZFbSnTyb0QcAoAj8IxcCtQ0EsC9
oBSXlyTQeH9iFXGSgvTH0sLrYnM9TWoOgWsicRhM/nME30cYvL9Qbuc+lttfVmfR1JLMkooT7/2Q
uevvgGzi67zBbhiz7hsuO1LnnMIbtpe9Cd3IMkNmhogQMW5T93+HpqvHCNcP+qCs2P1xZRfkEm0s
YYn75+zP3JvPl7u0AbmQeSMvV53Jp5ndNY9TfVdgWNZo8Cc5Oee6ZwTHkiLebtNZ0WZZSb3HzQDG
DSrnWQt0NeTUCEBkNdGe8cJLmby+c3hArq0IvsFTAS2DjlIsASFcl8kkyP6TVjB1JrQJnV7XGGPJ
HDJE+67lp5DAvo0YRyymz8pgqF8XQ3bSSzuXMImxKJJ2HKzR7F/tVEZOPRLxpvPna6gUagBzubtS
kcKKfGzMC8/5f2gWs4VRrwfJhgykTTnud1nnY8o5lHCwelTG8iDd8jR+SZfB2/kHNfmRXQ7QfVJT
POEyYGyBhEEX9LZtOTGt4WWkUiZdYW/to5s9H85UqqdbekooWBv2uLXpPGjEXK67K8p/Dl9xZAhG
/OwnBrRExyKNopyzsvdk8P94LtUvJslW0Z/a6x9V9KmrtiBoAuwiID/Uh1DedlHAArkxfJxLJYjK
gNytnvhunjmx1Y269POqmNHuSDP2lKr54ziCZdP6BoM0fuWIRarTZgQwQaqpbbLMabuID8yEMH/v
7gm/NcXNk5HQ/5YXYc7U44LyTtVx/gIpWaQ7bchdnIQtk/+d1falHWNU5iQRefFn8BslfErV1U3U
HNPGiP2QrMrFzxGsSYwTBYFxIDwveqnkyWrOtdA4MJ8czV72VCMWVeszqnuqDiqRdo6ZTJalGWOq
5qfd05sJgBEglonGCRYx4E2+k93AkxquR5Wuj4iYsNE9swZgbrsH1ICJQl23V/0/N8VkiEcYOKzD
0B/ctVvkejXvzOMZZXXEfnOtdhm3/0olEsZIlZXegotkR+IHYGR0yQKOedH/OzJ3HxlYfjeKQu3N
6XqgMe18oZZuNDhfx+7rQ48xJoG/Ba3X2Kc7z9HURFeDWAKtqbOS/Y285beTiMFBKW9lXuzXQVYW
9vYEnKO2DDkDzyJjyAcCY5xYA3+QcGgNE62u3dZ4siFms9lscT4ckbgcqTjtfPfY0is0HFm9RN5B
ntnunkBxRgD0wNr/QhRAaphZpsDgyYzA9wGkJLQvqAo+gnl3soqjk/MuoSiYGYxppEhB8ZooRpf5
c0hNVm25A3yl+jlABlZwj0bbbYivyELEzNKTqlBEGIx7zsW/3MAR3T6DP/NbyiFKjZniKIMnHi/E
XlKFC5QegLIqJuLutbzx/rLphoNsCEq+tuSeLs3Pj+erJ6WWSAH8bvBlMUdMkzLzcRkoHBcnP2i4
Ui1ycyFiE9BmH1OxEKgOsq63y8Cz6oSCOSFwkEFa2OvvlmsaVXGVbBxvtauZ9bll0+Kiy+d7fcGL
2lE4+ACX+J273FP1QDwL7/UkPqgS7cP34110hkI20j7eg6ygpejulQWIn8i920SS8yxQcrk9h8l4
U5W3mY79q46l0U3LrIyhBGPBwnyfghsTEazICuhpE8As+E50NoDSXbTFSArTFkrY75B0yQRabUnY
m0AAlp5g7mlNQAIlWUQUa4q9dsLXHnsZzsVNYLYXjf7Ga3mb8JPmfB1o0yXrE56BR4LaG5z9JTci
YUT+2gkuphlf/gCzv9LcG0yoXEoyVyx+o6pYueVRLwEpwx584pGj/9H+SjWLSEBe2tiOcz6Bv5Wa
dbEwL/veRtR/jXurxkY8kjhMet4AFa2SAKofPeIVehHhxsIBMckSQxakhf0PsulqKYupfAY8LHYo
FUNnS4f4wmOH9jeJcIWjKEHrVHPdjTMk9rKf6i9EhfR4nIAM4mIZ63B2kYvR/lvlq70T1L2Q2k/T
7+ie+mKZA3VcbITy2JmrpI3IO6riAdVwntmTiqySaYzd7IO+HODMXBbef/zROjldwp2SszuFFsmx
NROlK1UF0ZAIYu5X6uFZ+KzamjixLFTr2nL0xMcJ0Axr0Tw8ay+D6ypawqeasE0BgYOdrtF9GlGn
g+D4pQZDJra16MNsauujhSxBbRDRGl1awCSj3gv21CaBB/u99KUzcYW3Bu/Ak+QtKuK4fky4LKNW
RXDwFjuYuF6rz99++rCLnYHnJWgAHk/Fh67kg1zZyk4OiZKcFoyEDPWRIGQI/OWuLtp0kEWT1eq6
kph4Et9hfe6A4bVzyfz6qm3iS6hlfkKjBTeYMWbI/3BVqE+uJG7Bj2REx390VPeY7MjEEeAOiXI8
44Y/YQS/rWYWeHnfVdVLPcDiaxA5SCq3KiCSH7kw+zMBzRNragSXbUjVtCvoaHluj6IgFMfm3UKD
RCkeEDZQQB94dqGaWrniZUl2GtJBWrsgW6qdfPxTdTDwUUZpzyaksiRCruQYnwN68VNQtAtffwoJ
JvdSE4f1SQytYckDRUx4nIQLZh20nBvVi6wZdsOjnUtC2wepleKu8i6ICYLtPoo05SwICrgC91IC
0Hi0lIE1/hz8eYydirDYbWEB+bcVh4lOy0vAXudC7iI3jl3V2b7c0KuLLJu+ycVFKk5XJtJM5z/V
9YzYyM7jqHnaI/a+ZLXima+wa98pKifwCzOo/9r/heI5zShQgCP7SopMn//QMW7hhqoMXyqRTdKr
7NzHGpFad2EhqHi3e0aTk/2AOFs5R+SQQs4krsBWDd8/7BCym5bAb+R5pA1Lxgjx44n6bca8w99O
52jL0YWK5/v71R91FgH4s18NDHFyeqnMTMa98N9Wn28s1G3a5huHnL/fjQ4t3oayz+oMvSzc72HV
fsyTq4TJvwuorXemQ49aoU93uqhVmDsWg6dfrWgQ63qPyvAZ4qp0hYVFevGR61SB4Ar+jvgf8MkA
WjoHkyWdOKsvTgQ9CXKRoLfoSO0BDgERRoUJ3fLnb0pFZeXQnJWW0gm+FJesrIoWnHZy8yZCY0uT
jJ0bv6CHaKBCFkgfZQlF/vpq5mm9K7zxPbxQkJe5FtA70Uheuhwwo6W2hRFUZOm4AVvKRJ6x9QpY
c6/xOJWc0TAVtHQ/Mg5a2NvZQjFnNbbq008oLxT10WtJGyc+Ya9dtRgEuDaWhwY8+zP1obpF7/8H
La9k1XqhzwJFEQ8qV3C0oE2c4iPNtIx+XzLLyE5EVZZyzgZnmIIKhWG2SIM2ud+M5WFvZqdM3plY
KHvtlJn/ogJLf9Tnb/VNqaUqF7DhFCDP10zIg6tNPm7N6hwZzXiuXb+gzb8ZjmCWcBPEKc1UUaWN
mPQV1UMfiFYooN0YbjG0AzoABnEel/XUFhaEJPc/NVurs8JwPm5gGud0NNdVsssC8LpS1d7SI1jM
Eb5yza2Kfw+jJKZHlHBgkW9vHLraq9qfANDcwIfq9MMpnTqbmz0GwUwy7HkU92G4FK/ZJ58vvJrc
f20JnHV2PoVAJwiRRugq+DWY8B70tYCe2gpQYXseKNuZugrLJNNMKXIm5fNnat6QvKiI3ZGgPMfH
GuSLwhSz8o4nd7DofHYJjHESmu+dDFN+Bk9L8QAwLyY/VAz3th2kRXHNxhvJ6cPYMSVuR6xBzSS5
EE5xjwgU2YJrooY5+v8LbRW96oqsKpd76qp8417Iapqr7Vv+uWRvM+9Ab2tyAxKr6eZyQ5TZiY9x
4Mdfgqg+eca+p4G6tQK4By5B6VULx1bUNHsc36KDHBmKjd/NidHO9tgPEX8SL5bMc1vU3YfCYl/e
gh+hyoPdf0F4m09mG37eN1DLNsju8oPcE42LjIUMIjbYOml9CfcXe1amyn7O0BVs1GP400Wdf2dB
taIzRuDl5P8/s+ttCszI6rJd7FN88PNPnRKsq2y50f1aYwz3ZgKo+kxph3VsgsiYSxAgfV98Pa5w
KzOUWP28o+K+dVUT+mqQqfsla/0BaJ1BJPKK2Kj8iky5IGB60jJMSBiEmnc29eyuqaqQ1oxq3fX+
21YPxxyCuWHj3zWKDWvigQjgr/GkPkXnYPi8bYz6ko0luIIfJFK1IbUhrtkoLTtPHLtkPC77PWw2
MO8pbouWklUomxWkr+XuEh4cFIpwKkThg8jmlsZ0tWxv4MpA5rQQzdRo8FsK9H6DPUoZoTLETny2
X42uDAHwKEga5Kf5FsD/mGILvErIba6wh2HKO4qQfxtro/fnrPz/kHrIby2m3z0GVkhQkzdDucYk
rgESZw/HTTaJ+wWVvR7Rib7gIr1E4LmNkxPM2hp1KmC/J7MLTkC5JYJVHTHuwU0DXpznifc6g/h7
9MC8VgctTwVK8QIrQp9SGm7cog/oVLcdrRLWB3+KWi548t6/QBDzqMQ/jCbcvpQG+FzCtRltnCqk
Dg3QV/3WozorVfFlz+tqYwq/aaYs0kmIUM3YMzxCdy3PgZ8PKbhDDhuw+u8zex1Bv+dnGHxkRcIW
eebX/v9nHmDeZECbYvkc9HPo3xVreI/Sx5U2IdgTZmfqooghvUqgu9KT+L0i9Ijoi8YLIj9Q31Bx
AcWxmIcAK3UUogphrol5rqT8s2zrhsnLdiQHwk7fxqIWnJNWLNvXHGSxA1DPovCMNrBhdKVlLpBg
lEMpxZiCXLHOEDzJt43F7Cy/Vq0qY/ZBdd97PK5Fnc2qmblQgwuuwmbaa7hdh4kPx9SJ15dpXxFx
yxXPS82+bYBN3rUIG3IJdu6ziqSX/v1cfoKOnTBS9Kx6FA+iQXSDspG3ZXyaF9oC1GgUGMFxV1Z4
Dk+//n7ktpZiOLxKPhknLvdl7EUx9YEKhRWTlEK0gjG42t+7nJ/XW025h+B9r50XqNY3pmjXebax
vDtMy86QItKyZzhXOeBy6jLUQiZdqv4rGTu+LblvJb+Y0ALwV6Z/+chPDizFwxEvpLcL4YL9gzxz
aDt83svHNQRSS0unPXd5dpB8yir31QIHynDmm/7hg7YImqdDIuMT1fM1DFXJQ/Vp+Le042vJPy5g
K2Gd0SC+NHXFptVwKPR1gKowdnTBaj3aPVdKWzeDDwKPRfbC0zUTugmy/u+Jr5rJcPAxdDY8cFCF
Qgj/vyPBFYlg2opk6QsAxnWS0dUhFFAm1Vv+OCdDOrA7UIVyFLjDMQ2r5iaTdHfmSjljqeG+Yywr
HLItSWNj5MV/zbs2YjMjUCFsOajf90AcSszpEkvLKpwpWiqhVSGpbo+izCq60fl4C7VkseiwhzZK
xqRibJYNG+hjhqf0jfYGCzlfqmwuoeU30RUjmjvXcRT4yDejSf5K57Akmej5ZPtBtKzNnZh4mpIZ
joYskzvib0VJOLaAwTk+GTl2vDNXjLG2Wn+oBKJSFlyL9CxjCJoEa/wfa5q/LZwuGzBarjphiGq2
5A1TlFuc1VaIqUqifcwAoSS5sr09xeDkmjrqGnK9OSEVDTtR2cI+t1chddTrevryFNbbCzoZtT1z
yRP5s1P5/d4n1loc0W5RziTJr02pLlXrwodRL0FB/a84n2Yjyc+RQSI7eXSiaHH9MQKIk+P02A+d
Bj2irXA4QSx8i+pCkELTVIs/tuIwOox+6xg/OKGlJ3AJI28chg9TGa5y4TAPwMYaR8MdyxutSWcu
Aus5076g06A3S0riynM7uilqoFFlFycClLC/z94agtFI6eECgnUBvjbkxN8Pg33AuCuQ2i6nVgwH
xC7qrpXzx+QxtAzQE8wtB/go7cU1tiH1hkoT62Ye0L6NRXOX/4YAlf739oW//O+mKuLaQsMH15Yl
Gn82ZyPoSP2vW8kbQUFAs881u0TekfAfp7dzAjzaryUc7UKqA+Ud990RsAYtEa5Dez/6yhYslZlh
pMShGDEVO7xL+ZlEIKnSV2SQ265jhdSsUyjd201ZrdPqYvM4hW5/wkPNoMBWmxPelmWhSC1Rnkxl
QUFlHkoHgYG5sg/YHcwSkTB40/m3SiZEePpffPbu+rNNfkfayYcEbYW1kRUEavluzFYOkUjg7MzE
DlWK+PWeqRrtCtrqjGV2FcLsxYZC1KJudLkS/ydgghdwo8OmqspUpU1PEZilPfw24BXH7b1FjhcT
DqRKeGIhYgXsWeHW8ZvGmXZwoXW8jxjA4LaWjCUKtYZ1SE5i4vCj+0gvRnI6Ago7Ihp0XCLtSTcC
fKhsbaKXKmcEnm51tXBG0Kmy3iI/+SmID7RUQ1SWeKmT+HiAHL54uP1eyOtPNKAbwWGTnaYLmgRV
dvA8YEehZnSjahQDwl/Uc+5+YGZcwn6FQ4DFzSk8Zfn1f4AkGlGxtE8lG64dy2r7YSlqklVpJgP2
Se/xqwXiTIttIXqsn6tTMYUN5PNMNv35bCF915qka5F9XHqdXHZNCfdcf13NKOqMjI6rgV1jDOhO
b++lTwz2oaRtVLV2OF1GMyaL+IJuN8KgCxPzRkEi/BZKCWBEAeSv6oHVfAjFcLK3Q0R4EV7gqwb5
B3JllHLqwZD568nacOIu+cOsRnQIbjPmjkx45cPhEAcQn+MSd6mAQ5zKQIyX8oRaez8XHnh2v88y
/gAsUiK0wm7nWJSlJvCwqeKbD0GTcTpCMY+V2knNLSq+x59Jjt1Q+TP1V5uVz1NYCVXYvy3tUMTR
a+Qa7YmHFMwhUPZYQqXmMw81LwzI5tksmtdDFFGR4X3Fxa24pJwGDmCrJMAcAvsNDCKiMx9Hd3Rc
cJX7GIInj5iyk1ASgidDlerOFBna2q2R+ND1E3JeeC5F8ff8V9UrGCRH07aRRJrjNyc/Q8ADcURE
iyMJyW0nQNJC/G136pvSdOC3/6pOQJlToFEPvxB3RRiEzQfxbdejtGR1YbcLYATseLBJxAawpdSO
ZvCKwfZ8u6rGUbzE5lc/Qvq//E5xYnTQyeH+kew2qVfaGbj/S4RAhLGGFTr3kJmWc8fXoj+T+kZo
SIbFk78yuKPrR+ApmKUkbe+2jb2GZUJuUH3BOjmbtq8KEBUh6sIatLUeXjZlCaAUGRvnb6WGw95Q
wgHPR1L+qyPTcXG/tcAFmYJ+ot1zdzLAEsDDiqipsOXMJsgH3XKdFVy3P2KMDUFJyrZw7/9tMkxz
5GPiPVP5COvy50qFOUtiOUcdJSARib08GTBy6f4z1WPgGPEeuRgM4xqVQ6bajmJ1VWJhLkBZYRJz
6oabdY3425AZNSkqGznbEJmGIIJrX7fIgOO51hY8M/hEqmSdTSFAKOIaMISb6fBsUyNW9FHS6kyS
pbHWSOPG70ckeORtY/7Ds9DozJSweNvto7kfowdW1tCL1eH3RQdDaB5n2mVvKf+Zf4wFw6nQ8xGQ
2FZ6l+a49vOhen9JIbSvMyzoiNY5+9v7e7hXKDo4VbDm04UY6+bHBDQfRUFWOUOtUt3Zus/sZJ4/
Gy2bKnP5SkBqnfAWIIsfHrYM5uHcNaLNFJpS8UZI9hNPDOL1TthFG4zuHDJmQnszUH2pVmpGuvLo
a2g6JCWL2Mw72BHcKbwMLGNgjnVrgbd5jotyhdQwK/LA1fGiDcBa2/uUa2VQynd5Nrv2vPbrXevl
WB7hKf57feAwY960N6rrecdNt4QCKRjh0YhKvn0q3Sm4bJdxP+GO0TMWEqQ+y54LZsNnlP5eIad/
dEXqRv66jSzJNSS5TdHQNKuXJH+rp9RmDbh+QZY8AFt78xjz5eoGf2TGsDW2KwQNMm/R72lPHjCk
RrNp6aOEV9aLExjONCyNnRXGwNMkKUOIGv4mMJ3uIcCo28xS6rvedDAQBwhtfAcNRXO9wAAR9Ub+
HWOBVqxWYbsYuw2dbrT03whRKaS/p4ak0M4Hl4+4/693TjsrUWJVtNlrIqYW47kZLjEjy96kjHUa
f0OCunBoeBg1Lc2a7UWICcfB5vEzJz6BAg6BdMXDHsS7Rg9XpPFtQPJuPMnZl0AmMfkOyhw4U7uW
SpQAzfAUO2L85Xrs5Crd1V1hMvYDxheVOq8Vh0T01spiZ7odefQEdqf+gyKmDuFr6xX+AmXZ2lsO
n3iWmUruXxncYh2ZywceRIPmV8Va3xqlhQpUEuIhMAXueY/BEOoQ6at15iRl1MPpRFEymdn4MWBX
735IWVEXNg4OXHN7SF6lupGr/q24s5MmHoN8ZGdBtZmHK5c4/zbiccFNz7iWYAIxAmuxRIkA8reZ
qu5rirKnTkeic0Kp752BZCyj7/L4y29H8bTI+ST8NuiFfFCQ6j/jCagNCvnLdGjYIHXilmLCe8Bl
46k+ocFT36dk4chUUQCwa4GBh4vWDD1S5ndfMxwVwXfn+RnGIWam52Wjok1xEaf22e8M3SeNYEmC
rhQsM2DNBjt0ug1d8kgWy5aDl6pm67HGQcXx2x9c6++0zhV50C1ebg5NtVCIyIQgfwtdn8XgyZVz
gq68ZsMmpPkJZJBNFjM318iV2q7//5n3eETxVAY+NWUKU5SLJXtjdRY95ihpQRIr+GyJkfbkLGmV
74DWXuX2M+plJFkkKZ6v4aJdT7vwi0ZdROw73lPq/aQYM01L1S1R7fsGzY37DszevSUc27DBd1z7
lpxDz/ahwu7O9WUdmBgcLeZP26CM8u58nSP74L/MqYaOjSZS6BIefKb54qNy70cB1O9eCpnYiLEM
2/SlZomC6Q4Et/ZSQM1w1GQTG7vlajZd0/U1WKrPory10bzF/qbOsO2wIp30qYdNJnrM85aP9jxN
iQFzl7M3meaZy7DRJaqSKEFlMtgsfe56hrPxL+A+ko6+a9T9DDqqjO7mpkOwD3HsyfyPr+Kak+tb
9XVf8UbgZ96UxZz1PYXSnyYRKHOH4y0+V11hZWE2oN8SOy/d2Zcnn6Ra5vNUBAe3MBc4cUddHaU6
dw0+lrN6D8/itxJWkSwoJwgV0pVbrznZlmNbxxfY0X2rthJs+3jzCf37lkHwmW9CHTC8tFgJlGmc
v1sFUBDV1fxcfq8M4ghql+jUhHEWc1jIIW0rund3qBcap00EjDhIYPv2+UZJcMS1/Gnu4ky4s+a5
RYvpe2YYmhNkV2nF8xjbcI4bk9Hk42w2dkIIIvBGlVROU3X4m0ZvDnCJjZT6AIqPq0/2ljxpVpek
FoRp8LfPDWBkteSwS8xqiOrDwUpCDNP2gP8a0A4Q63W279whX004sW2iRbN0pTHZL/mlcUyrpaGR
wIFgtzE3egEP84z8CCCc8LnvoGLpUFWL+Mt6kbE+jPs0GwE6a5Tj9eSfVITPbpZVDXGjpnNdQOYn
v9SI+Hkf9HmAUjutCpGL0TkPLYK9ESt50yk8qSM7eTgAKThT/6Mg1C5qnO17LZsB5eKcorHVdN0/
jEuEEVDAW5tudzS45pS9i+ZA4+Q1N10wDFkcGPGhwC3d9roZmuJ8gXBWxBjn9+9xE/Pc8F+ov86z
3tCQ1CnB+g6HwHyJCCeZfkbJRfb/Z7Ksy4kqVhQR7OFlvTNL3+qR3rfuPa8PAKDv0L7uuv/iGXTu
1vRi1SycuVfr1lxldTpjciXps7MO8Ok5o37uTyGfew6L8eL3HJ2vGqChZAa5suxeymPUTR/Htugm
98oSwLxG8q+UfpigviFwsQpjYeV4h7wfyiPXZf3sQLe3jP+XvEcDN+v43XM+L2ySDFm++htnrH1s
BQyhmumi+/tg7dYGKgQJBR1mcRid9Zu20h1ryu/Ll22LXoVb8CYsu6cfUULNim8iUadF59c++o4T
s2mNXZUmuiSjKs7G5B36mBgoFvQacjWVC/W6MAmlGukT+5QPW1XSRpy4Gs5m2OfHv+mFElfF+62k
oVprfntfpgK4LE6gqn2unX7iAQ5xNTPmvl+du2ipcC48o2k4nQgWtZacbpZHCI4IqxmIr9APQE5F
bznbzIWiipgnKBRkDqgAgWHX8zaMGPFtSS5QhBmw1EJtaSVBodjWWJSiBIdbinBGiBdxLh9iO0Gr
OWQ2M/+3YcOJABKh/Sb5UdERdzoi/oXUEzdHazd/6llegcBsftMbRtN+JXKMC2cTm1wNjveaxsUi
FyJ5EWIxteshk00RYBMkzXoaX/V7UA4vRPpwuHxxeSsZAuHLEP8UVl3UeL2hGAb7EqDp41UC33Ac
9p5iBpNO1/0Lz9IBaFwM/vzY3EVgnP6YTRn8w1lPw+7RCsxtqHbcxTxg9eaCTMjby7wJwX5Rj3x3
dRiWYxCafC6MohD0kPXcvekIBktI7qOeQP3S3DYmcl/I1L2vCV5ddugOCEJqizxC79/wMfnXNfc9
2BVeMAzZwe5Xq8JRRJHykyhxAPb1lAQI4P+EEF47LW8da4TGiNXXbe1oiDAftLxkfWguc5RMd47f
CFAfnrjA7/scKjQZ+Fc3wAHAES2rdyIYfWKrEvLDiELIfOVd+lsYHcEO7HU3DR38APFERhnd89qz
k/nvgEmo7mgKDjUGHxVyk3MxTg1ZVMmeeFlaJJhMKfScJkqoom9+iQeYtIDl26kl+FacKnvqLRCX
etvNGA3Pq5h5yaMe0ajDOkaj44qshmUQyid5xKvDR331sn9lL+nNLev/ycazA1FF0Um4pwwyTqyU
4Xs829sIB7wKOgyRtZhLJcNHfbqotUKpzt4G5lEfzWACFsDYyyf/AI1yqXxMyUSaxzp/v8Q1gAh4
e4AK+JfYPhyX5Tr+DioSnPBqWCO/6j3j29ZvSsyUtB98ZynPwv3feIHKClEkUIBnpXWjoItGWoFO
rFAKc/H5Dts8sDZ9WLbIWp7TkNXoAEEIKCaCNtvAq7OHy8SHacSQ9kfw9SIneNp4GtaU9xqZexQK
i0aUkFSIxWNgby+L5D+hAt8OBtakFy19jRPe+d1wcTbQmM8R9ntyBWDA8KF6uIZ5zhfDcJbLcdrL
5sNsp+g2CIhk4QyVpmf5H4xaCTGb9fVLNVGaw/r7JSj4IDEcqV51xOEN4tHIFCR3BFXVX3zPDyvv
0XztxSgIgdGA+iD3azLf7ECRWK5neRTtQpANitrMVfX3fb7SLdDxriy9ggw6gBfWEhb53mKxNsok
xXK922kQXR9GowBFbFDkL4G9F/KMWPtDzXCah6TKRK17H0jkUW1zv6V0ViW6q/5gpgeF6Q0vnk8x
fJ6cuFk/yxYaCH55hdCxEx/xAL5r2wr6RjeZHzdkCRS2wujG38cvJ4PHXPqw20Z2U7XLH+IFg/FB
srTkmwDDaQZcrI267CVhurF0wtVg+3lysPRBtkejSvey+5TCg7xsMrwz71AOdhEkHz+fWW8l3n8o
TlmmUTx9PbVUR/yj/dwcZUf2ELO2Q70K7Xp48rgDQBWrSpb1Squ1o8eNc3IRl4mp5HLMq+P9zhWq
IxMqlECXHT9tq5Wv/3YKn4zE6WbHSYvOl9kHSLMfCpPAdXPC3WxR+Pa2lbtHO319Nh4y3/GihlEo
VOb69aoga+IXyvfpy8cpsGEjBDzgWEc6paKVP9XNpPWeH+VD2NY/NyAUjTOZXMdTVhrBmV1yWvBk
g9dkbkAfG2aIG8uZWxjioAsANQGsgQiAq42DhO526Go+A2XygJB+RrJypGRjjt/U9Km+Ft6BLA0h
cFnmh+CgkVgRSGsL1qhuTPUqEzx909T2qkwYC10/ezp9Bm9btM2309AohmRUL2UaLA59tiApAxZz
TZqZgJruJckObHZUgLblsSqt8jeIktI6fB4PQ/2vZMIPnqbBstjjr3N5rozu7BUw3x6Vawh0WIXG
2Jiwzvxmzuow+SM1XePZiKoGi9T9jGT/8uYoSF44/A1/a/v4/0UyFRj6tPfM7wJ3meuXyfgT0YRb
W3yBnCTQTOcaYSjrut9mH7jjH4BbF8fPi/pMxUCwqjWAoRXkMU0wlSmHQ0dTX2SWqjBVDMRsS0Px
IhX/8h1dWbDZaN+ZuGsFaT+9Iie0xQzBnG/5vrg3C+qAgD+VAc4WutAYxTW705AlFYhinc5ZV+ZA
HnK1hVP9JY2RRZw2xX7KFYDZIBPkU1+CuLd7JjHizgL9hpHaIk3KsrQQ1EzobeFMNpkU0s1vGFkG
r6N4Jj9w2F0cHl2iqN43AyoaOxMjGEDyRYpPgjlJBptdukd+UqKsAKY858pE+4jXc3i0R/4gZ2ci
HoTLt5qgR5EXtERUJNB4tg0S/vcCVXheWilWlM0e2kqfuUnRQ6w3hN5kpPo+X5jHrgbwNTa8TTIk
JwRYSZJ9/FUEywzjDqjIDN2zFei9hlP8bCuzp/dc0px81WjskLHDf3gNPHwkdf6qtcztSBrLf9tr
erA2VsYBy3ogNdrNWcDIbzuNTHSftMpozvLMJ8GPLZIlhet0pKnLzmvMz7wDLI9fMXbBcDN9ajR0
UhZIadMrit+SPB42/aXP3zoxrxVQNWJEm5Wv2QjTBAB6uvp6JqJNWl15JOxx11l0JFpY62ktE0aT
hT1FUA80iUgGSvmuCNJLKPnKVCAiar4YXwAmT0qKsuHtrSQqMV0C4x4oerg2y6eUzmuIHffgFwij
pdwZfINHEleWymVh9G4fY9OqKB2I5F6ce3RrPMoEYaQpZKjzNomlKijzXH9fPo8xwsby79xrK2us
6OanXf6H1g+iQ1FfU0zu106F3nYClhSZ36BGII6ZX+g9xNhMnS/JxZPdyKLUgpOqoAhAjDJBmo5v
SCvI3bKhKya7cAjCLqUwNQGTUvyYax7POqEzZNMHAo013BAAoa2S7mbXlI0HIL0++peMbhqpn4cy
yVOgM3/qTSHWNwm8wePMfn38wsQGWJRHAPzNA3hOjjhCw4shSo987V2+gxbC492JMNp2qNZvBtVR
+OKMhhB1OKUDVXqopS4Bxw6Uflnu2xaOeBWvvnlx7y7u8e8sCB02cU5Wbaxtum8Q0ESOkGTeBCpj
69E2J15uNcpfEUb3Pvl2RGeMNwtrIMfRIRxcTJbVcMQZiSFnF33bYRB1wbpvulQM/thhUPRosA0F
4KE4N/hgtcLdqvB1ZyhScC2unGOvGPIYizQ9E6pn5kZcSIS/G+CEXQI2k9WwhhYUojnR3fX3/S+r
F0mSAUS5rcCIXbnfn4nErGjLwr8KlTDMq4MqDcJljLIo3f9twNVVgW5+ATWI28e5t+TfuaT7kLEm
8iuxMpmgmm8oiXmlzAeqT5xPM0Do79eDx/Yk4uPl5NyXlXED0ivceVgoUe92NQutkYsGgdOhgDCD
ZaDRZPo+r1x/fV1AMKwk473AZq63ozCr5eOByJMeaoq/4Uil60ZFzMVecqWjnx4Yxz85c5/mIJB7
UhSlFkapgkqI/R61uhBg0yzehKuGBuqkgwSOBrKj/pMNnGtVNrdfR09EmNd4gP+C7A2bBEQuOHwn
RCSDzdmzI827yRiYHwTBSseX9S/ByMGnitlPlRMWqk2o7yScSWSh8AC2qhYiJLNJCOLYoN/Mojz2
3AOi1JSS58FnjyjAnP/YAdFUPwb/3JK6spDAczyGQvOP6dHUdTSTf4cHbwXruiRv3fiDMJAg+b7y
X9iygqYDIXAJxKLLFcxJGssyBUXYlbe54Y+z0YM40T8wGKIuo6pq7zb08yGXYyejbIqexgf7+MGF
9MUeKd/PbXaS0Fv0wg8tZsTC+9URAKiq9DU+iW/BhSaa03111xv6QE8kpP4/0/2aeIq970q7FPeP
Pqf8kl/Hw9YmZLadNGHq7XzrVeT1pc46UAlxPgvXfwscpVHFS60/+pC9ArlU3iUqmezJvKgXkOF9
TZcepAuc09ftc/fkNGcpMzmzFhtqS1LCl5+8ND2LK2cZazZ0bhZ1xMa/mNw6s92b3hiS/JYquvUs
Xrfyx7FLV+dyYg+GZ+JCxFHAGhLDFpt5dt8ygDTTJDnUkCcAgZCF1ES3COQ5tZkC0P7QDYKePA0W
Xvs0DdFY7Ks/I6UCB1jCudg869mnB9OUY/yC09aaUsyjETIaMyxHuP4iwve+2F+I6KfBBxF+KOPC
RM/HemCl00GCnJEbVIHL2Gh0DR66F6XYHM8dDPOV5y3/YNfSHjZ8QkFP5BCEhvdoUwYsMyt3gN96
O2xqzlyYXqrc6q9QBXUSP+D7K2bosSZRaei0FVESGYpETkwQO1NoJpx1uHCvjqtHiwcxnh1Y3Lx4
wMMmFLYQC62w2FqdDCDXyz3oHJfVYgLAgIZyMRzKR/gkt9FJWJN0J7cHDHaGiuUiarY7zEHtGQ8M
0okJxUe1FGzC3MGRWyKyd+c3OK34yiyOjKXctfL5uh4eOEoSM05YRXRMEfbPU3phUh3dua0U+56S
Qfph29ggR4rJu+Eg8dtQAHjElc+lH5pjFwjU3NdI2ZKYML1Q7iM3eAVYi9ZlH5L64a3rLozxpQT+
a2JRQxKR1FHxEl0XZtN9VvqlOUrJqJVHGsEHJAPkVdR0+t1taXXSVyOpHxDYvGdZ3kEeYpgI+xj8
P75EErO9TQd7quF8RKMTEqq/GG9brdAzeGxhgpcPVQ/hZZJfjYkZvbGHfmlWbA2trzfb+PQ1u1Y5
J11X7LP0ZmeIfLUxIfyEhG1jeKqkCz2uE+xRxikdoia+ZeKgp1ScEzl2xSq56qkdOTzK5RzPy3Rk
OJdZwwXnmPQUzwZcC99oqa3NDfoIOn8d1IfkHph1iIgxHTzeZZEGvNK64VWm2HI4YxEwd6XNEbLE
uKIcxAkdteSyEnWxi3PSYLiyGRojTBn3EYTflSFwWdPaIQn0ZyMhq7TJx+Ay8X+9Jp4XJOhqRJcm
dh2SAnwZE8at/6PvOVodMAzG4XToUmBIWW9FbPLo8V/oZ3FFAREclX31NCJtsglwWYc0wvYM8IET
ecmZKmofyFt9whrx2Vi2ylAoK2/1Y4vUm8ZJ0HG7U/eNLV3WDocb7Ngi3Y9ZdTVo7CcAmUhnwxxY
kE0H5owyXSSeV+8Ss//A8ZRJhhembw+QjMD9jNTuTJ/JleO/YKagNreACXSiD4H7yevElp/HgIv8
Ok4ADyb046mqJq22hu83V2jtjMJLWuZ3SWY7gNlAYXXAk7AWC+kz64bpPWPrOfEHBH2e00jwRw95
g3sfFz+xxymkXGa1iQ5cfMjBH07jIF78ZuHTRFe2X/UdT8AxvYInR8BCznkJMzs0icmyUlbLp/xS
9Paj06qv9dYJFX6HhWLFBbSEFnQIeRGvHcuLpmq67XWdy7dgOKpKOeXxMpwgAMSVLQ8DveBibE6Y
U1gPWkTRkJ4pXoG2RlS/VtXHG6ajxD2HyHz93irOY7Ek0plAZyyVpOAUDhYIwZj9+PLDwtmm9sKW
E0yP5RcgR9DhyYIZfcUOeYnfch1K41FhsdHHgr/JHJ/+oyFIUfpV4M82M8FOYTNQXGYTDSWNhpSY
s9On38YVNeVmZIlpsNBleWM5WHk1b5H+5jygjgUHBW8C8Kl1Ku08OkGZBOd8wBE7m9jgZiJjXWfQ
1QbY4r2jOuJnA/NyhQ78mSX/BNfF7B4tIyoAlu8iGWilkYpYyEbCJwDcrUiV81UiY8mfTk+SeDhY
8cq9/nddT5SArXL28V1tKppWBWuvAUis5YMxcJxCFcwy+ED4vi+rALujbQrvsApm8OqlUJeX3BQN
ANT1JtcKKwl+wHZZ52NFpqU955FKK8gloh3red5qBjb3igeCJIPxHpCqVGnoVIBlV8DGFH5rrlGH
e2lgSau1qvpx2pUMok5y13q5KFsR4IBByGk/VQjmckS/zr4Ad6yksYXH8Khpw6U2uKWAtpakFIQQ
5n2WkHqmwmV/AT06m54YFWJnKgaqesrGwLS3vUaeIkSreRkklOtLcei21f47wDHcl9V7hv9jaHGN
sEI6HEjyWVP1AYFnf5N1HxABLCS6vrMgSXdOCG+OjEb6ZA+3+9aXAJLtztl8+4ZZ8BYl+g/NVZW8
aT245uOkKHz76mL7rs5GyK0Cqrc8TYYoUaCZianyagpLV0nSkSBRW4lLWgbC7jiM5JXsqgXnQz/+
it7U7ASXzB9KaiFtTWesbktGtOjLLpWnfyqaiqxHogfssYRHztub/D7+hFkbxGcnBF66U8FOWUHp
SkPOazLMYoAc3qxG+MmDpT4TLbVUH/MpBooAYY8V7q5Iu2b9LGKarxKbLZgdN6lI7zm1yGZl42WU
O9KnAxhJ+Tizv3y0RYS+wapXkNVMFYB9A5rf0yOgKzs9/2qh9aPpZTuFKl5h+1mqu16oVGf2A8zy
WAWTtErESRU7q05dzLlrXwnj/bfXAKjXnzYIA8Rrp7lPzY7xl8wnQX2SDvSs18FbGVKTsXOcTwLA
Emm7J73Qmlx6T4CVUNysLTSUhrmo1N2OQ9Csiz9zQZTfC3w7nieWkCtN9dLdiR/ccWSATErNXr5w
28pj+tLQqydFFh0TEgCxrl+QdjOZ9qmf0sRQ+d9eFv3BnonWFabs6KJ0BVtzP6BUuoge/WooNy5X
NXqtFBufd9lwP00nhHHWjoUN4jOh7aUpsun/lfvnMp5xKLbh92v3waD2O1EYMNA4WtMOzbIu+gK+
J3vC6UlEtbDuz/rWfV1gjdhql5oBEfmTCbOEnfiChgGNGYLVVWeUx503By6yToyNrjsoxsmN2eOk
OfSxLxiD/1uJQ75818S6n8A2Jo+dTXEm26Na3o3VVEXSbuMgm4FpY9aDwX8MIflYg78rH8uMEDby
5o7UbVjjFG0Aq1ZN7bzCvNeD+1xzP7D8q8SADh8dh43DRoej3MvuxYTqRyIyGjfrmIlvIpCfaYMX
r+mUJYpdvoc4r2GXhaCjUQytnCuGeLAwnRjDAS5tJbMqz61WrJaht/vzwLDsQea2Arbx2v0512f2
LIuYRhmP4nLWx5c7/bdVhVnXXsW3zR1D8KVFpQ+gb4ReEPzhNkwVuL3oRLtWOp0lpBboJMbOugK9
grRP3fhU/Jgo7fVKSzx9HZyWlJtyJy3WcENhLksLBSwGK2Bcff0A+CMUkrVqJcTKxHdwxWr9wc1b
zoLr0rH/sriitVJfQ6bUCk1syixg4oMuogKEfHngE5JFHw7796ftYbjYM1x4c+bmnYlbyH9eVhrR
eUxlETaBTlirJnRc1ANTod4HazheltJUjZg9AARC44bFoNkWdpqe9kU4EDzoBT9HrOb5Tmr7aipU
bewWaJvdnQjnNY18XNtY4F+NvPrz4Gc0FCqcFgyB1pY0AQI0WM1aKd28OS8MBFH9l+iO59d4YXyB
6xKsjiRXnKTvMrCbA7MqINlTQPh8Jz+u4HyVwyGLWFEcf4b8XMBuTgj4kNDsMubbeTprI5zQGBEZ
GkYQZD65QA1iwswkq6aECLCsV5rUZgUjVJzJHLubp2GXzGpKUkC76pmFuGaxjOV3rqn73S8zF8HQ
RznPj9cUNzRK4NPD7bpvVg4wVRrbZvA4/aArDTXBAbujQKvbyP3ap5BtsLgzljyip6PuZ0YBIxBK
q2FAMDc2hiANsfpaW/L5bBCHXGzBYoS+WpdXSmMr5nfmtZkWuSQd1AObrVHbzMSfkxa4Xjl6Azg8
mpJV2OJquEBat09u4dDeqh6AMBxAB4B3j5Sns+ZFNh5sBvP6ZDmLPodjE4Y5ZWUJOW7zH3hGtESx
PVl0E5Pw82t3lIvSRSBld02dk1TCNH70DLs9hNpRgYvFTgb2bIRvuEkceJ3XkWuINUS4r1L8wZut
NzsqUPaLdyEMO8/N8+FzW4SRIqbWb9gHSxvsL1Fq/gjDcfROioCz+jnqBKljwtjVBK+aQw1ELXgo
eeVCa79NzhpWQHLY32kyu8ncF908TZ+jlhvN49paSGxCbruTSTICARTfEy6i0wt6SeGWBkjg7y8o
9yeX7DIoQvgJMPIeXjLPTtFA4QtFEpuH8I2A8nMneZxWmtJC8luVYpS7cfQyk3TfVxcuvHdtiiPK
nstt5B7Qa8tdrTQni8fibKGw+arxgvi3rqZAHomkZURULS49eL+T1v9y2r7iYsSYBI28XkHbhds3
Y+ew/Yu0zDk9jZUuUT4yVZplaNnwqtzTYJ3T+l3gz/am+1X6C2sOO0gt03Nwfthd8HvsQxSDoJtW
KFrRTeoo8Z3A9dpQxVe+36iT+L8q8ZuQ6iJPKKBvO9Z/gDl3JGxZMuwTKgmQZMXgiMWZbnIDNTXB
hoB1/ubg5qQznQmRz6xoZ3Jdp/gRJGhyBBxjfVAGOTo8137U1bHie8hrxqXVy9nY0lRXJ5T1WA7j
AQ/daljpN1QeewOKWfqPj3DS4Xl0lcutVJM7WY+PLIjb6ynoJ7XccRrcR6JMDlHSP8X8zoapYkC7
2XHjQL+ZBGrittTyV4HRyHf7kJ1cgzEenNY2IJJHjrReYVM9sc/YxUBHZPps9aRWMeHheCTNswrh
oeNCiER7fjO0X1B+a41hjiyaAmCMNcS11GtJNG1/RBC4Sfv3Z1mn2bZNMg8QKo2eQh1u4Nup287C
MALHQ4vDog5GYvMT52cWE2PGLTLOHwiXSF6/t+T98RAsJt1AaUj/jpHy4EUiCpy+qsYwtORJWAaI
K/4DHxhlS9z1Njs6i7trK/A1U3kSp6Iqm4/THenPCbdIbudh0UkDeVKKZOX0+PkuouxCoEQuzAKW
/dUDSJqn+aOHgHXmXDyYV7/Hpx16w9PHP4WWts+BArmAcTmIFapdk7G/Cd2v+lB0u/hYxS8AGxvE
VXJ3aPPPs+6bqJqFdCjNsESOvYEGYZ+DJLioQURPFeNfCeU1n26+4itMJK0OmIDjStNy4IIkRzrr
Y7t7cbgbzwGSWrrKVIJ19GoJTHThGObS5JgEN0xyJ309BIN2lyygVNF4VDdqu19UiAMI0w1r+FQ8
B9PKwuJ0FVBzwJcMZ4TE7oqBMqcxz0n4lRULd/LwfNpp+PTvffIIgG/fZJj7u/wujv2TZqmaECzQ
+qRePpJz18UUMkCujODguX2OOxz8Y4fLKx0mKJrMgz71sbwWCh0IcR4hdz385w5ICCiE69kg8oPG
GLfX8W+bO/3gPnhgiffvIW56+rFXOFPOOfWjznE9yQ61E8YNcpQDW1nd/0mAtkWrs6VAaolKMIOZ
BH8dvtYxyAvkwG7VUMtZ2HehaDgYNb7LQpUc/eFpvN6Ae1neBG2YB2uTNDUoHZnDHujQP9eN3MW+
aaT9hdcD057S+SLjgGUrPMtNDeK5v+MA35cs1lUR+q75s/pd8QlVI0c3uzw270UqOzmq54PiZfU7
Y09Q44rxhqRFVz2DRct0VHLmdJ1qBAdArD578FyZpa5wwey2Rs4HrGtgSugW6L2IoLosSQbq0Z37
JAiMW+n7lsQsmPlI8UP5mTWLobcP5cWBHi0bjLIR8QREg9uq+tizUyd4LFrYrgfNap96Fz06QtLy
mTYVvxc5b6VZAf7GYKA60lGmmF+NmTOldOXetOpP+R5egRr9zPLHFFk91uXqr5Vn2g7oDDJjMn+I
n7nobN5jZuxAn8vSfufZkkGybST7U9FwMNzsSMKJIYIYsdJq6O+kcBzHBkW9pa61ZmvzepHIGA9M
oG37JOMwJTpaLMcGA1N9wi0EAvW1xWn5E51xHd3aHqrwpkREFyvIoym+yr83l0WsEuOyXDnp6Iea
r7sJ0EDSeU4CQVUhWSbjmCcRGMJ3cMVxznvReMd4rVZqhrpasonXSuSAqH68ddYniFfvwBKzxY1M
7YyO3rTF4D2pBt9vXXRrEcV6YEJI6vN64IKClWBUn8iNvsBW4FzuWJBK9aqwBkS2BeloXgQLuwUw
LCtlVbTtgZLgGqhVFIeo/Vg2hRLf/ppnSoPGWwJeG+XuVgP0hX+dpiv4NJaaiByY3hMRQF/ItGl6
rpGKvvfhXC1wMFXBNP3gHMkjppc+W+kabBF9PMx7vqYVEkLVhY2A5OkWFWpTnD2CHQvfyDb18QnQ
QbMjg4rq24u+c5w36B6ncLtQLtspPHA2zdtJQlZWH1DWnDv/sHCXJNM7p1Vpigc65gA56aRahmnC
o/fJ7JZGjcElDOvLyDO+lr4LK8gUJCVLmYDmZJw3teXQIsP+AKx97K+EUl44MJ0cfK/kUosiZ/SS
s+yD7GeXPqOAvevNSgKisWa9Qh+mQiHUtggSzF9OX0tyqx/NX7WNgzKB7kaeJ1KOMEITGyRzFs6u
JPfkiPuVIA99UoNRYDplpBSvgj0IrMmv82HMqYnFEh5l9HyMiF1cGWIVvWUcm9e6FwyFCOosPR9Z
eHAnMDjJ1Aq0QTIlwWjBUAnml4Ejsi4aFptHca/HQM3qd35sKJHUpPeToGp6g0nJpRNzowEfKwX1
bUwqjnu4S4cQEb9HbwV8v5APybP7iGUQlLtma2WVBdA2VedO7rAc58CITZQLDCMaaIOsTgQG7uCZ
JzcLmqyNEVUrDVuOxGridh5j8c8BhrABEFBGRiHMACwWjrs4RLU/4m+MKMFbvSFr6dqUF2kEvvDF
K6EsFEEN5latCVoh57WF6BH16dd/yyJf1Ah8L1hOI5+zd8liNMEaZ9C3IYpPhuDiMiv/ivLk8otN
rkTSuG6QBTHWqyxfn1/j55shFBxiCsg1ZvBA5EUNhcByv3XcUDIF7pwFZkhHkOAt+smq1NBighQ/
iZzltV+85+54jEcI5xa28Zlo35xiV1XGL2rNswgiX8Jaj9136VbnEs4l5o+ZhmQtW3Bn6wuVXDiq
6NeSW06rR4Xe2DnXsUHPfs0iTzG20VlR35rETzP8s2ylMcsK/iqDo0Y3iKhgmDxxsz/gIe9dcP+l
tzAcOGhMxs9juRmuEiBQ9DELb5MUf3tl1wulzWOp2XNqJ5gAZ9Qsm6A1JChY7HBiUnta9fWf4sBz
c0sQy2bc3Ya+YE4Qo5N1wS/YIK5NB+gGiaDJIwqs0ZCO6Gsux2KUF1wOmtZ6lN4V1/Pl9uP5ZCHh
zb6MMHhDH5fg1N+Re06z+DyGiWfVeE8wV4khW8lTp9s6h+INWDU9bUaU5AKHU4eNPFdaGLSF6Vgo
dPnw3Ed5ddAaQ94XhBnGYJE38y6tJlngZvcWl0hcVEMkeEV3yzwjC+ZRVMGVCrXRDaMHsKYD0OS1
7VDzzwMp4WLIjx+C7HypxPiPojlDY//nc3yKtsqOokNeC3EYwUevlEJjBETEpUJkhTdvQepIz5OA
TmNbHE2Cf5jSanLEyZT5cfRD69/m3nTbR1KA2VelSIeqBxEfJim/UP08rFIK4198MsRvs0UfxXaA
2o83BWejc2mNVdo5C73aRO7YcD6r8O0+jElGFjFT9tW4up21oTXQ4TAP98KtUfb+474Wld6jp5vr
gDQuoTjGo+JOX5odUdf5rr/Qo678JhVMV7Uza9EL6Q1Zz3/K2t6DYg0J1tyx2rdkT5dMp5fkUI1c
wBQT1xM/t8UAOFGt/LjhbbW2aIYizMHOYLa/ZQUBGx35imRK35htfZOx6jEOLzNIMbrX4Qul5lO2
ETyRfq4qkqJjwM1Eemfc1DXF9nrYuKNCWe/NzfrryZlP77MyqfHAPWAQWsA4nn44SGAlj8H5nvRa
byu4qSgFLgVXEsnWjDHAJQnVZ5o3NMqf0bKGtpKDkLr4ms2znSSFabX53nhg+qHReFh6/hL784D3
52B/6RVWHtqkXi/C2TOt9x4lzgT/rbw5UPQegP2rPelP7orcBlObmTSfTUXTTVMOqfKRVkiLOTSP
nREGsecua5Ra8WnRXinnviyBPpNBY94uXofVqQiyssb7FP26pDUbMqRoGlVvApRZYpq0sfu1arM8
45JJUa2tDaKl3eUbHzCg+P+GeQwR+GPRMhckbWuVx1nalE+m4J79+Ew7Ks/4PJfJprMKDcTGrC9S
Qc4/WhzkmC6jnSiv65db6/zkoZAnOUXQmj6eUcxyqQoDfSAzFpNJZ++L8Nwj05tZnPgyMXWri3YV
EUAH2R+0mvSsgyj7NmbfJHrE3aQXl4PDnjKt6tzk+1If6PbMCpNw7r3I+a1vz5a6+QtxMXVlcHTE
jaIcl6bIpv6j0Xse50xVvdfnlNOG8Gz16So7uJ/j1KAkxWCnw1iQimerw0j2DUuHh/g41aRO5wyf
TUHsdj7yrEuzCLmNOdTm3hLgC/MeA32V8ZcvIO77U+ouFJUJxUxmZbVc4xuVw8MkExYSb3SZCevq
lqgPFxJAPo+kdZUkPEr4g8r51OnLGM8B/o2niRwu2CdHE0tzCDuY7VyKivHnXKmug3KTaX8kRrhw
cqc0DrUbHaIVH8NkzH7a8uKdp2ivZItpQkVjZBXH2G/tBDf8JcpAvG/Ae57npcL+QviBtT6bBrPS
7q2XukgqM4/5Jq3EfSAShovyQIlEgXamXVG+PJFVaYkuHHb/H97yMT7JX8j33v1RdazBmHcMnEbQ
vN1SICuGQ8QDSn8KYhYLzA3wRZSV7bub2xMvBFWYZ4d/dXv5ZbhkaDSEpI4ARpDUXBk6ntGeA+I3
0gtarIOYMYXnqCpgJnleV+bxohZlQlR3Mg0Fyr/R+xblRnc8/nxxJkT+2oby1tv4fl0GxUgE/7no
YBMg9H/boOQWQHRZFWF9hmucaHYI9t3s0cd+raHmw6SB2ys4qO7oVKPeTncGiimUnrBHgDdy96jg
UUZF1zZO8Hm+XIib8tRi+COYpx24p7OfvazFpnsys/ZtvPH2t3Fi3V/4OK0Hq70wekg4ZNUSAciQ
4IjVdA8WZHfiQnTFsV6VY8RxNRb3Q+RtOh2BU/yNnkcdQnA/iQwZLKzc5vl1DJZ9mPoPPtH4krK0
XP1E+cke1E6aUvw1Op6Z02/QkrQ8BvMmSCd6NA4Z/zSWrpBSh5mNbOUwHV+LeHYc1VFG/nMWPGrS
YmWhUqNee+ehrK3kIsgTWCAkG3EjndDFQLNsPVEio0iKVbIaEsqPZBlpmJD18lC2c1HwumBFKPq6
bBRH7vAJKyOFdRCjGI8sJA4ksQJXOWDFBpwcYinknZnYFm6hv0hT2CjSsuTW3UDUrEsE76+NEp5P
udY6OSlX0yJRNfhypVZL3n1s8p+4OAnV+BQhc1Wjz4zuHXjxBRmiAruQCqHsWpe58IE5HRwx3XfH
mdp4AN5nIZJIBCLjQEUJwqXoJIs8RwL3VoA6HC1pvjoJcWbEj7YJtDBNNGNcaRvjqdbPembDxL/9
FatnmfpPHN4Jivt7/yOm5RfJPjoCeiXXIpUKbykhwlfSg8pvcHr3+wf69fVxQMHreJe27RzEw0/V
Lik2U3Wck6GasEJzvo1uj+Gx0serh2KvF5U5jWJZq1Fo/qMmokZbmcsrXZQBxVTN6j1Q5p6mmrhz
5gSLE5b4VQ03tnx9j5o+Ht29yF5PwtMgVuVsxpjfOE5RijsVlksdklkVxDJzTNPnUuJFrAZaxQBq
NDqZ1Rp9lxnW7CCCvq4ylLcTt0LvbeWNJfpc91sHPaQeWoOdyTwytJI0Ssfr3BydxxTWIHWao1eO
jqU4bPlO7iAHVpJAsap7vCAS2RNJpbHstga+0CzectCHfzZiGAcVAt5sPIpsUQf+ugkYIZ04YTlL
G8GsIwq6Y8z5CJHU+JwWQHMerSeVg4xkCrVch7hK6s3oTzAK++dsi0R6KmptuTbULh/9upHlDliB
dPzHsl3FPVJ3fTO2NrBYf2/QoTm2l61GELK7Pe8JmlK/AspzansTNQsl3+S+86qmv2dvtaJbl+aS
D1snOPPfldajPwFsTkWYvJ7R7Led/MzEHBO8g8X4qe/y+kuRW7tUKcBuiTucV/ZQJnNwSlLCItQd
SDodoxtpnWhyo3nKslxktvI14GBDsKybgH+c1xRmWNsvtkFQn0iekebO3576SpsZNR/PkGi9TPwF
K5UJVKsJz7ZaTQEgWfdf1DwJxm1vhemQLybeFUIJ9bjP27N0E+Rf4L0p29NkaFDhp/+eJT6sXqy0
F4L0RZCxtDWxWFOTjL3DI/S31pzNX4/vwBIyHAX2OvoxQC85zhmepj2neyEZ6JJiX3szkh3wsnL5
EbFbL96uHZcGCJtUctmnLDHLW8ZduuzKWbvuCR5CQSegzbiCkgKxYYZ4YBXhJECbuNU8iGmIvG7t
fBKSmmYZr1d9MlMpAuD8JuVtzEfI/OlVPVZNDtFt3UFg5Socp5HL0Rb8FkxrCoP2X4odgHVVCD8H
87NyP3X9nSlNYpqwC8i4YTE0f4UqVh40Sh+Pg6MAtRAH0QjGhwBXKWft4/4UXJP/c+3qa1eV2Ot1
5CyKPdHDT2aqo8/dpM4ihjh2KJ7PbzyY6t6Bvxj553xVv9soJzy2bqAun4gZ1n8ydW+aC88pVyDX
lIuMNKh0Bk2LhNu8vwYQnpM82e9tFL/BlBKuOVbeHez7GOswa4Gpua/Ap8eRuZ03lyaXafBj1gJ6
1ePtS6dWqwqexONjTDLJKItmdoAKZ28Xuav3avMpgUaSq5ZKbazMUrzC/WtVJqNK18GRwI5qBfIf
OM3KB4TKSs4SjHHUWxusj087F42MdHcpwtoHQCsZpIr0/cDjPzEAPTw2FBRf1AuFBDPUO7vfR9mK
OTdJQHoEBF3idZ7CTKniI/8OM89ySSKcOxx/DAdCNkLI17eWh3CFV7I6apBhTIxmBp7znPO7NLkM
Irq/FPI1RopWd1mSBqt2u50+3YS5nYWJh9ZTejd4mnwFqrGPqjdeaI/OiqfzL6Q48D68SXHOS02P
ZEW9HLxQR/S1QBbskJJqQpDdo8uYHUG7rRd5jg6m0jgWLZyS5mCgKv9sw4vLp59PPrAnzdYwU375
a0iu3jwmh1SeztHyqw0NQmoA7of7Je2sO1rGQAFvOG0/h/Uvc4Wn3aVNmiZfcMxm4XltOc4fbR5/
Fyi3dkAtOyDqkH4hQ6PzR9qhuRm9grXlAdgPz0OF1D9y4OLyiHIYyd56qIfY70++sSAnJLHFRp3o
u4cfWXy2+e1yJyzrwlrRCxiviKeZugXKwqyobioYlQ/6rOGpOd0zxN+M3sJ8ipOlZTU0rpCm9CTc
Oo2Aj64NW1lYXA6pYJ8J5Vy6P/KUhDbcvZF0eLynAalwVlLSozIvs8TggXH9L/SCoUDqzgW5NozE
JT8oQY/DIigZdRVvNmqau5EYAJd4JsrZXspVh5hvko/ugdMDzRI4zycbhQLJJr10KP1prH9DTADV
KCNAL0Em/gJq6Yw8T90Wn93qbVW6zlcgAaEVcQTixFTx9RXD16VBkiphud1u1oWMO4q8hiFRmIxF
/4HV25g7z8so/cw3SaB10VIs+iCvotZb8ww8SUksCPSaNnAP2O0e+KP/AUYvLITMCwRGRfwlMXZD
SVzwp0yi4yEN7x+GYOr0rKgjkbIl0znUUi9J2CzhmYQKcfsFj7u5ghpLh+CnpAjkI3fi3IGu4zWy
XGXxzZo3pmhIzLbl1gYXF3Drnmi+tnrGYvgpeP/MlFrDNi8zlo02Ew3SidZSVa4rJ04gHNMMdkt6
wMl6CTv7DXGZJ1kDrh8iTvfpWI2R0ng9eUL3BjmajWb2Z0DpJC1udq4CGTiovyyjXuX6Sz2iUWg4
IEFYdtBr0+EVVSHm7o+YKwoyS1mw4H/SjVh/Cpur/SbaWGIlLsWxpGD9J7K4MYpBmTyePkO/o0A+
J48jZSSPmyd6wSBTbqs1ma0SJKeEpYbmsISVO88MaxB3MPqRIWqHXxBE/+9qIL9MI2+bukHJa1FH
6dgx5zdslbmThn/yg8nJ3wsEZ7Z74PNsrgxmfxR2dsdnCo2hKUEvCfUmJ+TL3MNQDzxOeqnx4bxw
fQEwYTLhcUUNPP+jMjzvdTNEkfPBz/SEfypRPixkIeOF7y6D+LEjtsCNS/O8YaTCXPquz9tfDtLH
fO4Sx8xbEsTUfsvLczd9JF45NmWlbMowlMz3B/JTreNzwj4PpqiIXsAE55T3wpO0iEZWH/krZVxI
C5ac53r2Cu7gR2gVxPRXDyl855xrCvVj2H0HWmLP8ItAFwbwbQBrvrO0VEl773uJEIMi58DiMrN6
PlwpJeFg6ZVf8q7dsvTaKm6FERInJVOAeIB7vAyQQb3W5pvi7kc8nWap8nxx5FInhaJJYUcI3Vk4
Ds0vIfOO0H14XlcvH/EGa+I/SXW7CULgl+nF80YbLFhAmId2CF80A/fIN7f/POB6DiISFNbJ3JUz
XC1VL1ehBTvf9pR0Ua0fO5OW6XKh976b0XXgr6xd1NhzZo4KcfHnWpzJGrc64K8fJc5OwjVBYHKU
XiLl+rdFDZEMxPsSLWZB1SBWa6Gd+Ut41DVvg5v0ES1HuJZ7A1VDBjNhrgAt8X5pO0EHrpA1E3mi
G8aO0K7eeIJrQjjyAiwiIcXcRJVOIFnlCPIyJE9I5+5+rfldeKh9MCQdIXcVKQ1IyLVEfIjqfDT/
79nfCDs1t3zUDzmnREpJWX13leBtO6R0p6DKUpQi0b1SvD19A/jlhode2fUER1g42p3vsHZX9ciO
yZlq89DqsvpPO5nXTRVGzXU6kioj9EM67/6O8Xbrek1jajoUUQaVEip4n4KATiXSCorzBXIweabI
6u5BhNXQNnGsug/hOba4O4mAYqkcZNDcPkR6oOLxlrHj4gvRJWktsoOoLIDEvjT5B/1BdkSjqSNv
hZoNeuq6a1glQXVHpgMoeojKQgrYUy2yZmeyfaeGxfLVQlp1LwMrh88NWDC9K8eGWSFFIkEL8eyU
l/DKKCkEjp5j0sUQkELR/kFlwr15kwEbVgzcACM6MGuUyAI/J8D/MbvHsByj7LDeoIYajyJqgXax
/23SI/hnZQUnjHdNE9529LpHzJhD01Lu/SmrLDNmlaMdGrtAW++jrDEoS4X9QhNkKFHsvfuwz6by
o9W7IU/FmAxnLYfnxQJjNEwjtakKZ3O0g6pDeIn15gcsW/ShAKCbLsXqk03iQLrrlnGIB8Dvn1on
ZRKM9gXHDUb+7lcwrdI7GCwUHFgd3QQJj3WkTy4CyzsSpIDjjYWS3mZBNK/u43eZs9+rXLZKObGd
RBekzTIGARhj9KavtPTVZWLpGfh9pgGz6xquydb5KXtCNN4SvS0RNe8pn4t6L0cJVWGVwX8MHFhT
KKRZW63XfHsPT3fjyYXOmasBnCzH3UIZ4kXDvdCKC5pihQCT6HiOCqgGtJiV/KYq+zrok/6gwrk1
vtNDUyjIQYtPfFEcSVVgyI3+pdhGhOnQo0iob/b1wMucHZM8V+3hSzSJFHLYPEHurOCp0BsMj+lg
JXNQXnqEJrjXfSzq4xYVAfxkJraTOnD6jWAr9nWIPHbDliOYAcpUQjl60XF6jBYNPHy+u/BzODpX
xtHlEqJM/j8LfrNvI17I4FbARr4FEhh4ySDbU/bp0LGC9yu0nJuYCADz8kAj+lLV3a5bxbRtOPCC
wDyPWEhXp/9S826MK4I6UnE8RJ+i6AAhZncQqK+8EZyOPHzR4uoC3XXXnzS6OSDbkntyf9C+qTp3
jAiqMkUgyyVWdmGPMJDmK+0hNAuL8B3o9rImVtVsZmnayxT9WeZBFOKw4UcV/ZoriMh6UfC/KUqV
Vcr2DX7wjNQ0sfbT0BUI/UVtE+Kw6IPDB48wwkeX9YpPd6oDpq0NpqmBBu1wnX+tZmhtWRJw3mOc
mQSTKL2bMMqGnIXDYh7hRqotHspUTlbpaf8piJjsvgmw2b5iqgL27c8Wlvn76+94jn3BZlH+W5+M
BpqNhtnm6ZTDiSVzeYVbM75JjcbO2XZeq0bsruBfvLBx1a9YvK+sbEk9anpscMNpkhAtZXLVmCR+
6ZQC3NwpiIdSva6HCPVoLFdWVX8awA2d/Gwq/2fMkcY+p9sG1A2bWhSnlG8xmTlYph2PjbTgrF16
2TLGLWV0VI2W2PAoiBW4LpgzljsECjGNI5JlnewGIX1fcshj3x7ZlTj240OF8viRmHA2e7aUZZJS
2Tv2NdNSHbK8Up79wDHbXJBbSqu0pClLP03C67ixRiXzBUn1wySGcHmuG1EANH3LIedNosT5z6A+
3O3SHVq8dc2aGVqsUua0RYQkIUBlICABAYCXKiNP3GlKfO2jS3vym2C0wU6tbM/mppEqEdi5eS7R
KvGHKO4Cf8ukpN4UEL9GTJOl8w5R/eaHdbP/pZ1K7sZa5QI4lrEMhL+3tzoVIcfgl6UTKsd6yfyA
PfMpyn3OkFWlF+ACjz4Wz0N6DtRJ5dUbwQt2m5L+gk3w6O23GfBLTaF4ABjf4Y8hzbFJJY3ae9nk
creTBedYI+F+89x9I0Cb1iQdSEezIWlFQ1/ksWIajDA3pb0s7ie8ftdaW0hDs01UHOVjoSHKauI7
MyBe8uvzWoi6dkHXAWqyrWA/3oGspIPLVIIfDkDyd4wItMGN2gAr/Ktvpw77w3xUOdmoGwldL6Sh
STtRrE8mn5O8mVealDpe03TDh6vm9gufHf7hPp2HqxHu1l4XConi/NmJjqAn9+lNiTB6G/zJNnkP
kGi5QJSe84RfNAltYg3Km4rbiyl17ssd7W6qic6blOM5ME/kKbilKfA2t23uzVAGo4445kBMhuyH
spLRQbX1iJQSR6Jyal+Ky8dem+CudDbZD6AsHGwLmw6eK9tDFXQRge0JYdlAUTIaztk3IQx2R9tF
F/R8FcDcf5GCY9EfQ4Z66Qat1++JJpPF4Vb0PRcZxM3ZcF0KeS4zkfnr5tRfm0vYbSXQZxrwMunC
GNeo3JuSemc/sRsRspoF0LIrhojLuckIEInhDxda3hATqv+wSagfqQO46bf3YYZKnO+kAgBPFXcS
x9vX15Wt8QZjmbMZvlgvUDbB1F8f+568D1x0YjbsKPQwUaZ4F51iiCWkZZXZzK2f3lLj0iT4eMaf
vY1VW85E7ANQ2mhPnnZEiHExpUO/WQPZm5pYlAAe0hEd5iKiHUTmawAgQEFIKyzB6stThdLLooca
0jnY2arg8u+mV335T0FdgMJfMMK0yvqhGGvRRBKke/FYcehdmsX1eF0HR4vdwJ/FQqBQ1eg3lmI8
QvnmBhSnuxxvvgWvM4H+jbQ2u4lKHUBcdWvcK5PC9rXgKyH0qGTQGmmUICaOv/24f5vUbIQpY4XU
SIsWcDiLeoH4hDPCQ+WguDD3h408+WhU3TleedpAuicqHQx3srUkQ+oiQU7XWIMk2Po+eq09Dy98
FcgRm4Ff3jDGYTOnFFkmVvhJb1PaUnfRgWl7xYIF+OEd1YiGhzLh+H+TpCzbhVkAZztWZxoI36nm
oLTu4L2Or/AnQrB3q+yGRdOy5A7uxhDjzMW2tg32GsXiEee++n/ZSv/mdzb6EHkAjGzI/Nn1j2u6
xFzLM4l7EoxKW2keAtb9NpqPilbJwEtm+oWZp6X6/ciyH3lmm6No6YA/+hr7IMiM+PGFdJ3ilfq0
nBuCup7URfv08t6vMNHPbYupKyCQVQS5WuxjI3jLqOJ8oi3ukBG+ye2azBsactiFf4i7EOjz3jfy
3vp1CbpHa17d9m2jjYuJjCHEKDtKyF5/d5YPi8UsZIReU8kB2/Drxl0X25vqg+ZeT5nQvLpTtPJF
4RCDwKh7u9KpfdNuKErdaUr0lA6t5m74UPQHxe2w1U1JeIhd61zYp7GTbc9MT7BCGvFmi+BBRwrN
TW+ib1EDwQRx9wsuI9+HxPaZKufered41OjoIaHgQnhRuHEpyKd3WbEtTSuKCMTljgT73ClrwYHy
dWVutaKB10t7byAwMZuSrlQ0x8OXCw0fYLHR78ce4SMJELo34T1qc7kv0N8dyQ7W7SaWzCL1ySVO
epAlOI/htaM6z9Jc+gwlax1mEpA9siNS10BzlB1ppK1mkP0Gk3MUPM0MFcuhEmi1Qc+zVROMp5D1
kEoBFAR5hY/vfUyftqJtOGc1/h09aqpWP9ZjKcG2gqglQnZTAJ6aGSwpOkFFFO2s5AV4ttdn0twe
cmcjN3b1sZmNUL1nnghDPhkCHbFj/k9gaXn+It8LxotJiIAz4cwl/psqnpqynaxiPT+MATYY3736
FQJBirRdcYJwFm1fpyFARqHndk+Klkqj3UH+q3Ql8W2XZnbJeEXGNSA+CGPNEKi04jGP1zDk3O2v
5uUnLIrdQ+k+DnfggtEVmCZDJU3xNCNkGyxXIqJy0yFQKoy/23O74seJAj3y5ohM++Rm3pX4FG0+
l7iSfEpD878T24DbuzlJ1MrAzVKcVEU6GR50FnscPgMCN/pX1mYBstXqaXytgIvnhRGM+wI/B0H7
Gqo8g75MCEDKZDXyjyulkKUFMJz1zQu+RxL+F7msAWdM1AM+E5TzAd00Z8AJ8r2UutlLm6kzUikP
Yo9M/mVRBlEnk0+6LFmGSQTFs0zMWar77Zz6ir4bJglqFSlCsMCcP2Th5/A3pd0lEfd3B33J0uDi
rmFQ9t9HJDZzWWi6FBtOf9G4pj3kOz4jOswlu72ZsN4B0QoBaBFE47ZJJJOa9N4BpoKGk2sTNE6G
ptNNsEvb1ZgkvwVXtqoeMMi8GvopSZ1geHJkjuwvJWdw4j2yJVZcreV4+K38U6Xml9NuiSc2k/Vw
6EDaB2UdgMe5f9xd3cOcGerYxxioxRZZDmCnhDTwIMVcpfmQOBvlfAtZ6FISaTx0qH0485yOpecs
1RRVRaIBziAapWl0DwhjijAeO8SwzveCV69ESawQ+jBHLCKDdNBZoxgcripJurR3+PccMxpobDXF
QTGoiiewVGU9C1DQ8iGp0+Tsx1fTLcpMmdQJ2SW8AcYIKexd7u+Z70vJTzh6I5Iy+O6t3K+K/741
Bdq3tOJYdmnHwGjV/Qj+XvyPqgEwevL0IWEtAFQ9uH16Kmyjx+JViqhHnOtX3A/MFkq6SSyjoIYA
9mvIbNuXoOrsKnNUFU4LBRx00u5AIGxJxrj1NsOvG4vNSzjn5KgVM5qZinxk+lcQ9YO2OrYiOBhG
+ugGKoO2OGpEZrVbM6TAEDCt/MkTOoL58pN23+JKaD1jBEOVBEexGTg9r/bKIEBF6BXmVaZUnyLw
XSSopZJPRTClffEsIdaUR3nxbZhfamba/s0t4m8ukjTptY8lUjWkgkEobQFePqdIDQbPAAUSNUQv
46dgki2rKNaEJWMlOgNWPbuPJtDspe2RMwd0jl0zZXAQiYcHDIK+kaydntK9PaDbcLpF+lWiWXLN
jiJW3Zk5Oun9DQQd6i33hP74CfujyMfLkXjEGsV3YO5hHS5o67E2r/eXyqeXEN6exWrqSK+A32gy
SlXJU2A6jkB+myiSytpzN1enCEjC9lrKtDfjiFQwcTw9/aBr9ib1fXpI4jJu8CdYJkjtstQL73O7
Mf5sJftO1a3C7V4bMuOS7hwVDjfO+5kO8jTgy7tYCKqd6UFNuCzRMs+jpNpDkgO12Hi+vCoBI0eL
hOGLuQLJi5Xqb4JFuRDpQxfCwdose+R+GuWcoHFpN6g9aHcoYmJMRKrTyRjpeUhkRrGCZVfXtkAY
hcxzpE2nQWyn1Z+iJj3HCG33sCKuxTy/s1GMm5u0tj+jlPgpPdOsgMTZ56Iy5LxesY9x3C7Ynb3u
ZvprqKjhiLIdctx/KxD3yZgIVR8WbtI2XLu5+ITRaM/Mbex4K8jtwmcv+3NkqIjqsps3YhPj+Sw6
LgdZ6r6PHxUDQMPI9/Yarfs4vH8XhOZ9Sp2nOLn8LdTmjAzGDVjci2nucJlCpaXb/d/TaHKxh0tH
SlTlUY4KvtIFLG8DLQL4svto8xl5DnoVRUSGJhBA1w20SS9BgllZQLmRbxtE4NuBMl9lT0FxdahW
YrEbd782baCAdzLntDj34vwKW3+vY+mgxObkUU9hSVJajJkYtkgyVf4MHytUjpF8mqsYCoqykJm9
7pXxx5jSNDTh139/XfGx7npuyiAfTG34hCslaL249dPjufVHpdKXQ3JwNYRxWLnafoaC1GHnwegf
BmrySb1ejMLiEGr+fHEFDvoEnNbctxJZpJtVjw4TXfLSmqOKFtMiWBkt7fvYmwG71AktjwT4Ek6L
iJVtG9/tTUA2+1ztrCMSyOqgY44qWbeT37mkhRtY9ofUToQYgm/XF1NRyfVllur/09B8arwiNvV+
K+lQVlW0VfP01WIoamxuhuMWjFPrqxQYi1T0idpErqoY/nALJY3vVQ5l9FdqexKRsKMeRh0DUvCZ
VZyM7Ivz/ad8a3t4K1zgc/fulRXTsqUCLahcYO5JFpb28N8NYKEdHmhIEnB/e6v0dLyrXVZHYnnp
3BpNcZD+xj9PBTB8oJbeHJLVPTYkbfUzxf/c/jf66ORMGmLkXItOATnPchB8gNlI/FJGlobMjeeD
BdI1zEjzp/7Q3zTy3T+6JSRsg/LKU4s9hG3B3XlgUfp3SHMzKhwSTYMNZvwnO+fJXrn7e86SlXg7
bIDB+Ubp8ASSAuaVLRQyb1HOB8w46SCToFUeiQgKCmE/Gbu+5LG6kw6DY74XcHvYcFzu/f1QOrln
72PO7wpPUD91cC+xM3QiGEXbjJWtREgwL86P7MDb/nla6IV+4HatDWBSH7QhNSB/TVE1WiMwIkU8
bmqwR2FZ+ZjU911ukYWjGOpcphU7xZYc2SchViYfVk4EL4UG8f4I7bHjS0qNeZLo2z19AhO5wIKY
22Gwg3KCR7ciaGQGvqCUVq0p3Ywscbn44kNzJVE1od80KQq1CfaIlLx+U6sRJwGqsSqjCXGgeb0u
w+W4emD95wQTP+mbEscZJTSlA8Dij/mlX82fwjM57PgeuOe2ubZ7wwPH3htW6QwAdB0M0bUqsXwZ
0zjqlAI8b2K4kglCixrhJhqYWsAng63DGf8lKji5ploeDSzSCPjNew4Vtg9q83bm00C4o3Gw+bYM
X+RfEwM6bHCW/DMp+EqjpJ+U56zhrKBepqgEnH15k0uf3c9zMFuW/wv/A7YUHMTmAfP4ZWDzid3M
WkpMpRV8JHrKsl6Nn7bt6bICrx7EyJ9fiI6TXa/Ip4VLNwmu1ktaPPgTDWJ7Wkt+3LzLe/TxIXmE
CI92LL3lK7+rUdS80X4UVT0XsUOqIkHXyC7DoCMAP3oz9aIyndP58k5FO19RPQTe7Lvxy6i8W8wp
OiX1wxK4uGWmXb0Qko3gdAYPkQVXOjpkj1K7F+oT8cDmHIyNa2k2txJYUcrf7WY5/JfYUVxFHEQ/
YAlbmcxqly3djBkuZtcuy1DZgEc3Pq1wS3QDs1ufXZl/2OFnnM61Peyhqc6sUne6GaN1wFGWwsdM
Ne2bB3fURUp5Qtii4DTtOOfySnEN+OS4O2t+Yg0ZvIOJYOarvbYJ6r88oUsuoSTuS6mkS2ms8H63
UoV02JrM3/GJhqdPGNZdM4ZJdYH36B+Md4c/Oq+lzJyNPS3p/EA+lvY1j1C3rF7DSLHFZIBEBC0+
1tQizdnMmisaZTMJPV7Mt8wAcLRTZJw7YAX3NO3Mr6od8ZsVI6clSPtydicHoT3JM2XD3HHyHxBj
GrpEOo+PCD0dhfi/K4g8zVNBsYn8Euf8ucJfwuub0jLX9RarBBpQlxNP8bDAN6Cr4gW78zG+7k2t
8XQgqzUFI6bJqQcNvSNo/KMDaiUgfUbBumMjpYhzS9Mu1NdRiJupBn6H90u+G5uUqNvg963Asuhg
7dFoL6wc+EfUxqYBTn5cmADu9Hk7encf8uJV5Itn0eECMIK1xERxywVCYyCBOx4kSVEuo/FMIb2r
+IL12a43s+RWfNNH4aZeJR7HcIyWPkpMNycUdhViPlltvVGnZRcX3zuD416BD1f4rNiL6lFiMjC0
HRcr3mvihvacDZyKQRM7mQzina4hwNbFA8V1QPY+6CXYfe7ZreWGsvu/JDUh7i11IbVywi+lZScs
Q4bsGqQ8qIgA4qfoKctylbhBrYetX//vATmtDQ/L5K56mcpLSvdv8erAuywqy+1wYTkQHPEIn+gG
fQNmqXwVvb9rEJLkLO/BJf523EpktJ1+qiJDepsG1hFjjJ89RlnjWL1M/WobjkNiho5T+40++wN9
zpSb0ozJpA9vRTSAhc2fVkQk+oIDQBtDPe9YI8U7ifNFOVsvfz9P45PZ/dUAeAbEfhL4hF0iJ89k
OxDzBrRblbrUCN9CLwnH2ARXhJpGNaI1JeNIVT3c2kLOqfk8S8W+BVTMmrRhHBX6MDltYDYqiZXe
CjjKs3WFpR8qm9Nn1QSC0DU4TM0LxD8rD4wt0t/0Wb6d8j1107ZVcj7wBXSnQYblwrijhOAM2qra
vOMt594CwDcuR5dnU02YzGkyiRfcUFb0sfv67sasCE/K0kYcXDN7XX+pLUP/GnpgxpvpOU8IZ520
X8CkhqaGuaX+qtmTytDjhF9IPgqGtkNX9Qr1w4A9TTMXgj+18wIZbRRvEmm8tjktuhMqYR7izrRb
TdNfbNzwQtlvGjGOFQO+jbHxPE2na4QMzb8a+AcNL4gRfmH4MKJ1tcNZIJq85e9zhV/Lr1VQdDgI
2VAKO+puqoDRC3aRZBRTmuLf4CYven13174Sf2YYkumCUMyKCE/LoER1oUX+SnZWcwRhbza+Dc26
tcGphGJ6DHQGD9L9KXuneUcV9dpKNbyXw9uoFkiha7gNTHnzoMTSjRlt60ovW0vMedKtmhsQimeA
jXPHrIl6xlVmZyTg6eok1I+eq3NB3J+SAIwgjzF0s6b6ztg9kx9Sc2UDLNR1TLw0R7e0A0XYWP7n
k+CmX5XZkjEBTQuHkMkaVHH3ud2zps9IeG5wA5eIPb7CF2G8V62qpICge3y66g0SfF3lzZkiMIjR
DfUwzin2hDjui9cr/l18fBhIXjsAySg0jwew0dnDSkaP/INmXXAidq9mZd2R6eAxvG8NiGgpwqMm
nFln1zcMTLa/TMV/RI4TomlSD7FIct61OAYSg/QT7N3iUdG6KapFLCt1IqCWYpnzAmj6br8P8z/X
wzZNvXFoVY7ddWkkE/vqOWpFBHG1fpOC9kJp4jWQElE8LendRW4L9SL8MMLN302O3usbwOTpQwkO
zWy98aoAzAPREANF2Gjpv/y5Vy9AxVREyfXk22wQn/Tok2f/ELqjLWISS6/vLpNsjKbLCZdmt6WR
HJnMZnlaJUUA1caSFClVtJNn6i65N+DpW72kKc0XC19RHdk1Ri1oOVkZwt2MIGWAZVJKaUAsF+dS
ZqHlgYhtvRxzDDgsIvHxc8OGuf2EOXgG96LsMpUOyGeYyWAZbQiRxltSygYPyOo59TzaAAKtVuUZ
4o2BiBuaUqHFaPynXOJ/Bevieqg8L3O98h6mq3Wh2tu8+7fmfykNRkiGzJGyeZ9jdXviIE2da044
zrAH51gJ7VASVQXn1Jgc5reUWae87Xwtx+dI3EL2QzfEqpEWNmw/E+cMpjhEC2rljz04tG/KY+lS
FKmInpsVkmnzMUS1KPcaZNsbNKPwWh7ksNalVkDLeyfL0rZawN9kAA4JixeROkH5ohqBQLnPzD1a
JFUSssT0FpR/PFSedIcxQY5xeYX+b/ZXtZLrAs8zFkPs9XKv0DQ7awWh+zC3jzimq4Ux5IXCen2g
ryhxtpegaE9CgAtXCfu2RrubFR6UdZjge/TVseaFcVBcNhPzUrU7/0NbVwuZ9P+VR74R5wBy2i8x
N/gbaEVpxFAW8Khr95ixorHvIgA+GFwTEGLUWSzs5ZJx0I/JP4h1pxKr7lxPtPmQs5t2/hTndgOM
5CFWR3LwerJ6Fdop4xOpgFDVbu95aW8+QruelGxNqtwMpM5C9zCVB3EjPu8JwdbhHlXUIDS/vBt2
gHdI7SnHySf6ILUwYo/CpdTDVceAe09gfBOiPDFTUe851ZJyILUE0LuiS863zvayLs7tYw69R/Qf
D4647U3DlPYVpY4sIxoftPqGw2V8fm5piz/HG4zqXD8x2w5ckRSVYba41Jq8Gh431e5O2o3doWjV
5YHewL1sICSTFukrG9eIWcRxexxxy0g0gXnrSVmYNkh6HJ1ZFerYU0gGmbJCkleZeMlIY7V6wZyO
WoOZbYJixH8Yza3hHrAs+dMFgeLa3uww8VWyHMdqJOIFOpgwiHLkDBgrJXzzr2V/RrQqR2VnBxP6
YTasNnw6bdRJqr7372UpwBlalsZ3q16wTyuxeo4OriXcOg/9UQ+m1tRXREaYFuMPYB9mE2InamaG
1Hf9Hz0N/JcyLqplOEUIdK1mvVXijXDBfILhM/8TJELcLGQ3Hfht2GyTlwfTSxwE+lquC+fSwYcz
FI29Ry2Vtk2HIiPEQ/YiBb/nwNq0CpGk0j2Fhm6THa7zx5ScPpYxXj51ElxGnXAGOmPpH0wli1Sb
uRE5M79QEBoBPKlMBHu2Md/mXxVk4PTS/OMydnK8ca38X2EgBaV+vWbTk+7bCQnXzcRnChmOxBx3
RJjx2mspTUyXRIrw8ALcMdfD/ghxAwMXgn2NMhNmkjOUoGerKpJ7vOrwHCg7DxBZkJ14faxDk1k6
B9rhfEjWYCCbiCvOWeXmVMogScesWh4VjkuBGOo5WcgE/I3ndeyqK1Obx1rD7Q3wYtAGlJ8iwdTz
NfrZMQdoY4aDmY9ENwIXHvHQxx8iPvgfVggHUMJVIAdEXzlk1S7kqoLKD19QknD+CDNNIQ3wT/1C
k2UaUt/5e9fmJwga57sfNiwuObQucZ+siBJx1OPKAMm6OmIobjQJFXmtpjK1Mcb5fofDWaQ7c34T
oWbSti4gj9TOBOhbizzRcCpuWIlcfEEXKgWoCxAdz53FolUv+kH8aOY9ZPq6rUyc9RAZIXqlNMWL
aNtqBBWdaTiDrV/8mpc8u56CoHWROBsXt4NIjrhm/dgSrKkb+juDRU0cZGbpfT58G0Stl8ldjCa8
/Q+1Yy1ulnOo90xv3aAUHq7GsRXbrj4aw4s38eWb7Iqm5LhgBTldIDLFCkMTDntUJELHsN2uLLhx
8X5MkiQWdX4448baxB5MvW9RMU9dcEL2LlPQlhzD43z98daWcGJySnRMKqS8aESOUFSijvwfbze+
mgiBZ6ERLn1tj+fEaZo2UhvR0vsnHkzpZoc7qj/txPxT4oG4V/ctuZtLf/23BFtsqBxgugBerHFl
ecQdFosxGOkzEpeFgQHHg/v2pagsJIg8fFsICvu5XrI7+sZjr/j6zFfMDL5ruK+HOrGTtVwe+WP9
JGL7jToJ68Yz74djDb4P3AbHVwps0jtcu/mVpZaZOgrciT/CZWdkhCBJ08qbPosa3sZi426jGGrS
zdR9rnwyXF5RIhVZNqKQXwNuZiTn8RA8dBqMrR8s+wWGxbs0CqCLRtY5eYwn0/i+wS1c3GEmqZ52
2FmKr2kvsmyEhS1AcVIROR54LLkcjYNSjlqp6nVTq9v8R7PXrDYx+dnIEqgj0T1jWVdY6UfaNEjZ
PsJ1dKqR6Rg6jJZjA+Ke7SLmhjWZDc6EtFANI6O81MmjS589C9A06AGQU0vNt6SsdqE/0zyT5sEl
XIA8/Kjq4lWVSBQmUL5Th3DJ4YuHPVtZuY2AhRebAs8EaOs/2wXPbXM/uz9DxZIhb0LuzM0jKiVC
turHQy8LzyQvTIjQsbaOalB3lB3Z3MrPJQepfAnCpvUCGbpgbaMmCxL77T/YjmUysfg2CrmfVcXb
jODX6O0c3uKgu8uOEwWB1MakooK/IkFyMJcrptT2wbgR7NwU1B3RUtgCzjTbhccBcEPJMQDH/l1T
jsI5dN+Jbhgz3w/f55wLFC//BssJRHGzHdKWPzBy16fPCpir7RNJSrkDgZRyA+H2L5cRNVmnaf04
A+Mb6UcWr9Sky0PP2Clhs0eEDB25g5Uj/fiK5LyAX1wcJ8PrGS7BPt1P6lKZyWun72zMsNOzCYln
3/u9IUSsZ/HbiqqtFbX8nOykBMEQ8yOpNpM/qrOBCk/I7aV66RiQOnF+Y7wqY2g4XleEoG4tjO+j
DnB3Yim09c8Ha1hu8wKDWk8w1ZFFJ8SHwzoQkIX3LwqLxzfwVkHgUMZ02Js1/GemT5IUcQzXMH6q
+N95TriOyXm8V/lJfIItQiTQWhxLiabBlbZY89JYlpvOkM+pnp1skvbsZfs8iR++yZzR+g9xK8aZ
I9ugKXehDhPf1Px8/wAii4k4ijLXGWAhpi8hbyTOwgfTAPjdmzDEcvvshITuxYNe+YiLXjcxt3sX
E8zlbIEnMZ1OclstxKCERzfkLvg39RtHccjOASjn7pjToOzh3UdzhhWLHHfNUSVWxXkDxk0OkLvi
fb6qqk6Ruhs6vHbwmn7iAM0fCH2TWrQc4pnenfDOAt1dq2UI97F5JuJdKA+f8sBBqsuw4bFeL+8R
cfTb4dzmtfVkZZFZP0tNnNuybS0DB6xDNuL1TjCW3A1EvQAlRCPsHT5p0E17jhV+hS2Nza7t3t0K
41sVNu2Evbiha2JJB+C7NGI0ZxRyl7kQd/by5pFmEHrt35Ya/d4q8DJr52Sujj2MnxgLnMDNkfPx
Wuto9IWwzharPpaXSJBp+3Zw7PKume4cavsKHwHrmoCNo6Pnc80BMjvIiIEG+0autYmZFjrTJ8Og
tHdGh6VdtA0zEVZVEslAH/Xu0OWzScGpdvOpHtZ5WqHsqP0ZmW0XDvW3Y4ZW9B99QYEnxu+RxmVZ
ssPS7vCalbDrr7D+4vMrDmjmjkDKtX0ESs+tZiRQOUcCdaDB2LP0w/Q5NHKDDT1qktMIZPr64UZd
tpgCFARZiv4SspwAw3oswpiEkAXYwRYkydhcNKd/t74h4f0p5RBYaCo3QT6fYs3q/5eRcWGDtZco
ilvWs2JIqyYokuogJkHw04PSP8KHrmBk7uJaKsvzhMogLKlEVZceOnxXAymPrCJ16KVoOkM1GZCF
cRNezpFGQOqCCF36HHX8drHPOWNkr/oGYOQnFzF2E4PJF2AgVqxUuU9RaNyo4jAWDg/JG6/1/Zcs
dtxOJTMb4r32ZmEngU3KNp8cxIIZCM4UMalOlYFxQCgaFP5YhGNp+Ks33uGOMyKZmfJYcr/kKKrU
Gd5d16ru5MDBgHigxZpTPhVrag0yYXozkUOkTI8CGL26mClXK4ae2Hsc2DQpDuNC3Ucm0I/tQODP
dGqGWEz4WGepaLfmNTtktgh1tVrKtaAZlcAi4Yckl88yx2kl93RLxwO4axRIfEKKoO5a0++QMpvj
IF8Ewnhk0bxFiMRpMcNgEqH7/iWVKQGnlDRZOPqSIqDKgmyQdtLC/LZRyVAMhIfxs4mnNq72rt0o
loq9OAtm0LCyHAI5TzXOD5Hh6y28+lWFdLhcrNHreeF4B3e+Hjy3aOFRBucS/8SZ/7sC+mkxRLH/
FOawVCWxYIcpIxxwVqZk8rv5H9+DKEnoDM/h03kk3U9/L2hRK+KAPbsm6L+sxNbUM1SCQLhJThso
u2Sgj0kfy4Tpjuv3g4rwjIyCoCST2DJAHVa/WV4zf3yb/iIQQ6GVMhnjo2WuFVNyhYz+9ervAb/m
2TA0BCrWvcWX7h83rw3SWlk7oWBclBzVK1nLndBXsTpcj7HRTnX6jXnSDeVKAFzA4K7FL1C13zoz
0qIW4JBed5bD2UowVD0hd8o1KkBMtWlWGQeH2/wNeezNBT6ZfWgnxUxMj+FaHGregPLurnka2uCh
LUgfYXnpAWSi+uEspHJZFVwNSYcIQlVoe8wbeSzGeSep9wVucsnHpivqCS44XNNDlWpvhl2pQ6eO
9sfNyXNBEp5M0bndJ/WqnthYk8qDT/ixJ4MA23fcQlBdwJira7iKvxeblie1A32heR0r/7ntblXK
obJLKWBLsSd8vCcSC7sPYnrT+RIbjf9Hl8QYLmGVM8ZcsfVg0fJog1QbxhDFER1dDWALJ6sQ1fOr
jH7GJbCXoEZADgzMEdES7nvDPyHFHYu/+dIwl2VC7Pm/25N5ex7O8XL1iv/Gm2VvcaaAvzUyxxIW
H9oiAOjzM1IMCfBFuEbIscu70yRMRXhuHMoerYc7BDrdcEucBFocahN96eKw78J6NqL9jlhxXQkH
SCQVZKtGp1HXEA/HHbRV3M+cbaPNQqs9wuhmYbV+8tYHqwuYrvSpLKohz+tPrMUIJuuAHw1pfW2c
5r7yY/4T/Om8AmVKR00JECrc8uTfA/y5BJ7VSIeNykqwNAmHwYhCdeWlQKTQK13Y9jlsH9IoCc84
dENOfhglrRDDbrW3Gk9MIoWpcjxkJFVjGsvAabjsZYJ2YVb43Zdp9/kptcJ9X9uKSzoQKNrY+TUS
M44fiFNrl8iF5UBSXC4vgvbXSlS6hTQSkFxb135iJQ1caxpa/RlLRjb/mdxEBLJRKKZL34QsbVL8
iEQlY0/P+32j4mVpHKtt7MvCBxE0Zncd8xqHs/UQqybrdbx83STeU100lmLfojvMuRhHPRlPscPN
J9jcRRw9uTPuqf9GZh4TplSLrk/ldBtdhHDQ084s1yZqsJm2iIiVUrHFrrfQgIF9feS0c/eI9WbK
7FqglVja9fJ2KPxkj/nQ7Xn6K5oqSV9fHr5QmyoqXYvi9ZSYLGPP0V9hIQGMHIqaw7GgpMeLbKtc
zOpbiCthqU6daMZF2h6BpQ8BhQmYzB3IXpudPAfXm9sXRHE/8FI1UdeHiUAUAeE3botqajg1/RUf
S/bl+eIMmhf+G55t59wgul+3ZxmPGhaMHtXhnmoK8gkDZ1UWGvQnt4KrtnNQHJ87NP7/pnYuFbzG
N93OM1I4DwdRBMWs7eO8J7gxHLo0Db6Ux29yJ90MafQCHud57kLR7ErK9Yt3uzqdlOLa7RYvqMfv
PAqG/ZF7Kp5xvdmdSI3cldpkDuuswq8DcbB09ddZwfqyqajfSYH76JNLX2K5Sbzdlvw3IPSHZ7pf
TByIYHcjW9BMFLebjNTsmvmBDGEwVbxs70BcUw8MfWshlHBPALTtHuh5sp81AsdHUp1C/fGd8L8Y
Iu22kkgy9MbR5iAPVLFEL1JRrTjOJPIG0gDyfsolM6vMTevLvtn+8m97rVfPeS7ae28a/F8ATZZu
kfzptQWtCSDQJemQBWeEcIGHfF5dYELsYaCzUBenFoW7yGOTZtxhDgisbqzup79kvpzn4jRIYDuj
2W46UUHc1F5pgEvVQNjtM6ZSq4UppY4mXgwSCCHJTEzo6n05MFjap2Q8XEOqbeLoE4955lIUTPIq
vA76smL9QNUZ2MOJ8et+0hBj8y+U2cDN5QXgn9ri7FkYeL2hWj2p/srf2UNL1wWWX1Y7caCPwVh9
TMGizej4Uzja2mF/ZHM66X5L1xqTsG4aeF1dOieYMvFpxSLGK08bMaxC+VEGAdoGx37/zKd1csAI
nAd5IKk5uTYY497anNZHJgJExuSqs0+dmaKXunif1sz0hgaV5eoqlsd0ASpjWyNOUuz6rh49cpda
W2SNF2WrrniAqCSVKIZQhY4UEvOY7i/XUAmH8cPJTkk3vbq0174uUNyuj8qgYNeBzBa4HLBOBvTt
krnqY0r8WyHc7hszBL6KSQeWuJpUB2PB5WtDKmcu2ZO3c1JPY27bgyupkUc3gXk3rn4tXlxdtT4N
kEcSm0Bab26JsBkdySeq/u533kiKOyYm/2ke03EIkrMt/Iorv3GZGeJTlHM4vronr8jCrmLV1P1x
hMBvoEqsM1FXHSTl6wNPM5SlrWIVNzx1bu/2Qtliju4Pjwg6cS6eMWNARE1nVOAFvhdsBIUFoqK+
pai/rEE6RiLBM67of4ifHVwFsaBgJ2W/jx4TLOhf1hX3pdNvwCmdEJSdkF+1oKCAXsUygJmWi8RI
45zqFGhKyom/yszofCT95kO89sE2JxnDSQOi12cL9JgF+WNVZa5Dt9wcdqCWSxQpxVivYrQZWa6H
+RFmnAlZb95jJMrwFCftORj9IMkbVZONvncBqXblw+MCjXl1xl4ajgOt0yCRK8TQYE7k34Z6sJFm
Rh9HuiIWrco2RgGf8IVLpOm9v/Y04WbFTYlwNME2pN4/WLDhaqhSIEmI8qO44jHfj8Ht+w7T4OJV
eU/grWigfAGyrKiv98Dcc4sU3FOA7/Ki6Z/3HYJLODRqsJYuGfjI2wC7psrwman6nwNM9p3mvvDz
YnmLgXhFAGNTStl9YJtxkt5Ou3UAi4xIYoNHRA8dmsIU9I9mJrUk7wSSvPHw0Y4jvpznviUsNbag
BoEfa7tsnCNiSb8OF22yaA3zCiXkV/Cnc5FLDacIgbyzOV38kpBBnhlTTVzgHnZSbIpBxKKRFdG8
ywE0MFyE4/iylc1MhqbjGKRFHJOpRPgchaLlHgqqXPaXXGYZ7XxtjpPmadQbMdkoXn9pbyHO+6iv
XmTMvqm9lvk3o8dMHjlmhHdej0i1Du7JfcVwoWZpDauqahQPsQNxXAGJVC/qBKPsE4T9DAWndmfy
00Hf3OMCkZHLb/iv4kxtP4LemqG0VzFLcS0kQbQmROxwsalhK5ribn+ru8hOyidGs1FYq5DT8NSI
e/+POby4HQELhsyin8SB4cHYPUTeU65Lwa6mL6RzPxiCI5/94knA4rDSw+1B278qQnm+noZXb/cv
SZMn6Dq6CIwfT2by67gP7i8IGVCAS1DuwWTz5vn3VBElSDJqS1HL19pzppEsERao3D8M8z8MxVEI
DCMIvX2SYzMjdvp8MRo/z1nnMqEVFuq+7BW3QgJgZlHIxIfcStUEwOa3qaVBzBHAtpt97/pxOZ9c
gQ8Hqu0xZxSxCpYMepYs7IBFhtjaxIIFzsJCvZQZhgxEB8kouD6AD4dJO0FI+CGYUAtJVcN9Ccdd
IgM7ERRoi/hdDkMjpvMNyNH9F7HzqTF8NZzbU+PabnGhhkZ5eyIyYtusXX6MD74ETglFMOvnmm7l
MPdNrc+qeAoaz2fIZiJ1hui+DXPowgunzeNn6FO5NTSmxlLv1+PBlZn7hqwlLVm4ljdzYJri9bZL
q7o4h1rM8//ApwVX/ZdVJNvBvI81LjTsQJzOLpLTmCjrg/QPZcO0Ggg8RNYO57zGXkdUbrBlMUD2
EYjScEuM4ERKaHhTGMEZWcr2eMyyLaA94Xiknpe/3JJUCGH1yIcwTX2S9bc0xBP3sdZrB/oOws80
efHrGM9ZYrsQqXhJb1Jr1X8dJ3avEjGioheRsXXBOCYcJX3oDrgj1imPLuEsAN4pTIwGnOC+c1bE
qgRnawcqhJQsZmqiVTYMXACIsoWL39gxZ/1XI/5lB9yafPAXEo1tPFOt2Z+KguH02uqWmRpKfkJK
dkBdjTKmb79ACdKe2lnAazMC4jcxYl2cH/2jmXV8QMy7Q3qDu/EsQV3rSu8wyDNNPH22QyB8amTc
izqcxy17jexMjt6wToK3vid+tM8IwcGYKHuIVmw61PxKvq9+YCrvACjgIiSwuHnwlvP1N7YG71VU
hyA7UUgzcZOfWdsiPq3DGP7P9YtDYQiV4neVkig+nt6nvTiMl1Oc9Sx9wyZfLnlQDPHn6K423V85
+2NBBVnFzYcEboGbQdpMBIOsPVd2J3Z4Wa8YmcfBvzw7SFB7sq0/5DjQJKJliptXWQ2Gf3Hmtd6U
tEqFaZh0PcjkAbeVVUh976ppOXH2ORMEs6sOJ+AzOKIM6y5ddIOINI5ZcHQCns0AqgOq+X1skTWS
EjDKLuwUIBIjY8rcZPNb/HNfBqZKev6YIHt/6wFYV43ogs/NC8z3n1HzjtjOK6Rgf61HaAQ13PSX
DMZk6DENlEUHDMTSt6HXlZ0F/M8RbEzoiOHknjSOJdH9nh8BlzNiU6O7xKTv4r/hBcguyptsAIgi
9qRl2uau5zw/ciwS3K5S4wdkKyZaWyzDgTYG7DBOrlRkdiNIBOzpLD0s5UexI7NDrz6yVThyBPXx
su5LeoQkVR2USIa1s1GKt1NanSnrGEVUFDupzukFhlEoB+Vtv45/GqJRF34RC98QHswdnz3NfbXu
abx1owz7Zo7+z/6V1VvL7ybCY3e5Dh5xKyKzwJpUaTIXLkbyTzc3VYXQyO+D982nau6uYBnFry06
NSFwK3G2wOZ7gMabax8A2TbzgHd/xEp4x9MMw8zGfC7LwisbTG0TXSggfXe3WeyaRl7L3B4p+d6b
mm4HOVwNfBUltm8ZiUlw0Vf1Bkh79Df961cT+rTnE0nUE9//uqb9Ra4BW/zsJA9nkQXqhFkNilkN
Ftzj2NBnjDaz+bXGhiDRQMVRlXyUFl/h5zcPNFIUJufgsKDi+B8/P0OeeRqYYMDKFjXJ8OpG2krO
XU6Iuyt2QQM12auGYkoP+X4r8Pla1VBmtWQpFz/1y6Tz6qjRQILzVfUp0jKv+/i6uNG19XPemLkr
c9wC0j4UK6D4+4uBrz8f2KT9TReeGFRFBLXEdipWek7NPagj036tC08AXUHAYcZDiCsJcJB1u9WN
oBFvP+s4sjOn3yvcwKSORwdiyH/DrRoRKDsMFogEZtdcYBW+xS9oNHaJPX+40PVpjQaYH6kHCgKL
TShgn6n7+qZyXoNHAl4jEiduhD2qpXDOzN6jNvn12eZ+03YWDZZaH6dkO2qxti9J1ZLdy3sMqE23
YJku1/3DJTL6UtC1+rMkqbZqy6EOPeUPOUyrCSPZ+8iMyzdXRxQXF8Xl1E6lbLRTMHnLWSfA7Lur
lVvF4Ocrz5VtMnFdXr/v7aOuAUYAmyDnqleGvCzxTkqUoC3ThfMbRDVV4HISjPp372F7HoQ1TQPt
OQWFQI1PVLu8WP+bXeemL/mrNj4nUFLBZVqWLYfwav0wAKFsXqDkPXuz4/TJELpAfLGCJ7YBQ6Wt
g/DcO6gufEyqPnhlSKPtEFAxTkGlxpZbXPN7L2gf7BaUg6Nigu1SAS5lZYCxJhO6cijMjPKkLlFA
LQq1ZZbrShIXW4kv9Ozg5/K96U4blGPJh47ALcYYqkWXJurK/l2Es/BhTc2Tf5Erqc99Wg/ZhDts
5NhaisF3KV77jtNeq2xNkl90vLAllQaAcsqgJl+Zu1t/nD3ZSPqqm7+1ExIq2qn6xKFQe3bTl208
/1Du9QBi2UAKtJCrIrZMMsEAikQc3kKV2MdxWBdZRDZw5Owx5/EM3cWyaAat47r6LHI4dX+d1o+F
36eonuMagIGrnvaqssutvQ9FJ7UPu2VLTQM4GdvIpvZ2CrGImgwHTTR+p/DkRh0R5tsiUf81BD0w
m3c9NlcCnkDrPGck7gtm8USc9kH9wf85TnhTD5Z7fKIhq2KIQnaIwZhK+MfSb5OZKDv+RgAKmmiC
cJzZMBJR7LxQjNJ1w2GPqPxsNeMp83IS98LTYMgngSjhj1apkrG2qj5aDqfJH/nYvkCgjSelNfge
z7hiboo1T/71u6sDtdl60BDA9WR+BI/VUrFi4+OMtjKbEKn7VeMJsK8D2ZD4Vn2dj9phcxwrMOuK
Wf1STj+IncmWrWYt+eGkin9V678jD+7fs1S8erRFCa5PhPKOA/IGAcB/MTD+eJLuIA0H8rzRq/49
qkXeOfZK3vpIDAHDHKk4uiVet2NAznqa4c/kbDwsV5wARCBs4CByKNmriF/LOKQ2kn3Ir0FyiDvV
LAHMwgG5J4kwReGBD4SwQT3aSmeEDBtP93nlS1iHN1UsZaIA5wam/o2m8fENZGMfYoyGHFaIxrDV
/MG5nfPaZoco7kmh9fhTZNsdY3wn7ZeCwumhTdYqkAb/GVVXzMXVPwy0MoB5jbgDZpWbqa75tNFH
NmTXbo2R9fCF+56KCqFN3THrBfVvX74q4Pc/7K0QS9eMYtdcy37oA2sqT1jEnXvwzigJaBqWdu4s
O2B9Xv/nDJYdriu+3v0eIpecQyqiQDY88DGJyU8ZSWLzrj0EZBLutqFVe4Ex2pQsKcGRBr1e13kX
6q7czANTqz5WEspJuQfRkYb0utvMu0MzyrsyV1lEbA6pLufPU3AbLEy7FK9S+Ghk4LZaD0vaUxPQ
mbofFP04VcuvCYtG38DJcbgxo8GHKUiw12sRPq7AJPMUCt8RRbD/F4mFONFvVxTPCRYGYqYpDsK3
oMDigRvZt17cWpTpovi30nbSB8QJ1ureGsVDKbaoDwB/RAuvV8GGE/JInMeM9eSt6vbIuZMoIvO3
mK6uvFijaPrGakYE3ju3IzXCtUrLq8JhoJFwlsJ2HKtO9jbpt800cUfm9ld4PXfr8uzmgr62J6o8
NLuiRDydbCsscxdzt+Sv6mLlJZEEJQwWrHEbMEfaUmd+nAnUyoX2t8NOnvFyTrn2/BWTwePrF/eR
4i5J74p49RbGnT0JFhGyqtV7lM9F+WH9+azQ9tFZ48McT96uRWforpeqWPyfj5m6tt9tNGZiUWhE
2a0odoc+tFaHHoaAvxHlfAiQ3VdtixmUW3TsAj2O9VumgO/+rettzTfToWfG1W9agQ5KZGzanrOX
mGXADFQZmpyC8j+CwHygtXZC2Xa1n/XARd/87OX2jwWBR6Ru419pgMdibjXO0yeM7Uf8KJSOvJ1R
uTrLaoANvl0CcSCm6ilWEq75rTJ/ifIKY2BhmMo3gv053vQvaARu0wRfOnRmu8KoWmmi5Ul2vH27
woVTd5S3sddtLGklhptEb5UW33tXLojli6WJUvHEwvEWnnXKfhT/WuAYnnz+mf71rAQfkDSsuWrf
0aR+Okk1SyXYFSK90giH8xNzg5/HF0faF4pattCWdlcIMv4g4LVw6ExMXunB7Eg+EIC4Pq/C4rm9
LpzZF7lzsUX8VfoLd4GThRT+JpMWcvr5DcH/iUyHBDGm+QwyOuOanx0Hxk3RCyCMUKbqhiRSGQjT
U1ll+RDSS1u7UADjrqYfOdl10sB6m0KNCfEVUnYhivtqSgKeG3ZESBzGS+ndPCodklKm0JGPLjyz
L0FKZA/zgK2MD2VyaeZm9/FL9heFNLXX35frHWmO90LvCwb5BXYa8/IkDZ4E8VVHl3+jELQUWAwc
6A/XeHMjxfSe4fKfW7kaOYniBqQi3BG8kveJaJc54eVidnQMfOy79bLXooakzehDIRZOhMQjqheT
KzKeEHAxqWdNH1lXI7QtzS1pHNvbHLzKlWcWhY2TSb6BCr8Cws7ZMSENJLHCO8rlFkN1EWd0ow9f
86JW9fCrn1uOWluwWqoExocAD+5M/zPe+DUElgh+RPhxXHBNHcVUFrZKZH1BSCvLam0qU4IgRF0i
eLu6zETx/8omdeZSubVd0lxojxwXQql8XniCiChAwt/QVXYcViKDpMbKe/G7nM2MqsSk4T8IrAF/
eUeEfKtmO4xJy+i55Ap5lz2I+D5Xz2zTvtt/6HkIe2lRSC8lEcMx7+n5rqHQLk296s/1+SB8OSE7
V2qy6hBRqni4tucTyPY0sscDTnOdM166kGQfNLIeTLy53sPOLFSR2rlsD5jy0UqeghfP3D90lDcE
UJDe0/3hM3I1HivjQZwbyT3lUBT1s3NobcP9rMfZenPmhRdqtTZJ0I78PNoEDxZ77qut3IcfYQDU
VYJGEI5MYKmeLyZ09QxAMGZQqXrefAz5LebM7zTcvPWu8qgpeZvUIzP4eNSPcLrsp8rQR9cNyI4e
ECikOUP/fFtxNC/hz9US8PVEunbtcKqOlYOjR6CQL8n7Egv0lcwar85KI08NfKqwTOpdgltPPAir
RkcesRUgm6a9xXoBfSNMXzbYDcZdFeyFEifRbical3//hfLhVTGT76GuBfTFsxzbW6dV/4Vzm01z
HS/eYcqn/BHCTndLBDrYjIXCIwbH3IuCvs4gmQbkwyH+8KL7SX/kKzCZ9rlS+pYKivPfxjNVu/+9
O3FD1lgFxlyMFXZj15p4h6FOSLuf5QGQifuHvLniZ529fjH3DBEMN8iFykTGRen97hTtUOyRNcQv
NU67U624dptVs2xB52Wmhpim7ApSaaNkMHkbWIlhTazmCmNvCByqUDUScSPq4goQsnMG8Aa2RlJN
VkPmB4kRgEJyQ7nEtvvTpI5FuJ5h9H3i7A02blmuFcuZO+I/dlL6PRkI3OaepF0JpUxV3CW0vit3
hDx/kxASf7ftCJdBug3npfFDgMEDOmz5t3Hwy45KaxgVzYqssYqICLxTP8QN6yWnxz84VamekRV/
qKrDDxgpUFaWBVHAHVfXz9jn9f8tIFGNaLCq//YFwriQ2LycB4kJB6A1Clywa/YPRizh88nhSrRa
DCAtkhgLgpvkF8S5Zb12fElsiL6RKbYQJA0Pydiv5AADRtKmvGYUJP2PK08W39efhVt4pav2Y7Kl
FFhlhdF1wOkPPQk/ummxi6eNS5CiRJHRUU4y2dhDvFWROVuP9N6sXKON+XxmkCCzOm5uvNORjnBo
o7Ekfeuqd3edIDdlpAbrgXEUBEJPmBAq9CCidUJWsUqzsdiOGkuGv656kbYTULrZX7dUcPSvZ1Ps
dmXSn8bQ4Eu50reQyjyofMvNjD1KqbxJkYXNVJhfCZmSO8qrySIDXLLl7E9F3FodqaiHK/JM2v8o
VSzhTR/Ba2fUc8HaKEfa1pM37se79F/hJoOrT8lEszlgGhE36EWmrYMcdbWl6Z0rVU+pVe00fHgT
pJg2laN0iQSru+y3S3HICGM7A3ypnkrNRr/LpKuh2zxRP7yluJJiqeeby2i0FJarrKd2i6PveoKl
BY/Yg2af3bymcmmMTqnZdz9Q88PRro/Euh+A+DGvv7aqyzBm+OevNd+UGGOXz/Zbwxv9V4p1DDmy
uDotWKwZ4GvQr0eB+hU7KtGg75Dq1ptT+zc5l9cjF9awY5JAhxJKOUazWCDYPGCHtRRSjS1tc2f6
YKdaa/XzUcatzbjM/5u3RzVnJLjrgehp75Sin9sPt2rK3+JSdRZva8j22D3AHJOjAjFMoA7HWEmW
8GiDDrjKNg8IOqTvfrqmIXpf+RSUG7lyzpr5/dXuAOs/FJdP+TGwD+7iJeIwfHjtBbin3khVITP5
If3ZE3PFEb1OD2NL9xWtT9HSJ5TqN0yutJRvH2o2EopogbyEQ5zQ9xhFCWQbp3E28Ck5L7d+ps9d
UPvbErMUUbWqqRs4amoVh/v6CAU1XJaPC3rRqtJUTT+bo+g1EcYgCgK5tFoyH93a6KMBpSUtuOd8
KLDfNFy0kVfcJ1Saz4gKdLAFJYrWVIFa2iFmVcIRJCUycUpScFuJCGFbNRtay5qSfTpPp3GF0oUO
NxlKbK/SzFbPLNnZBLlC+TZ0AUWoa5Su9JOfsx3FaB4vLmHgxFn4zMsq6tVePVtZ1dxq3PNi2qKk
G3Q9ehFtu47G81y2n5TVgVxoRz4pYxthCg/r4WTtiYcCUpCtvXEevDGbd6OTThxf+PrbdD4GT3V/
k3eMzBtcuJZdMq+DdmJVJZWP41dJH37wd+qYAxPmB93frhIDK3ZUkgR5vZRpfQh/bA1gCxsYBBfn
IcBWJPHIJ51hmek2xg3N7HdsDCePqrfYd8GnbiWXHYBIanEctnD1LAeh8Oqv59Hqa/cp+QonnMil
sBLjmA6h39WWsF2N1Zhg5hiCwPXxW5cG2fJf1pWYx/ZTYT5TzdYr/8KLRJhqV5sS9HEh3/VY7gXs
SSrN/JEGzkWP3HXGZRvew4HJqWtarznsXa1ISOww/teblEXhOMlLIP/U3AZctCj/EeYLftlOvpSm
sjUtjJfuTrmoOuYFi+H63w/DLtYDMmZoEHmI5rgg2LDSPC414mOl1PJTBUKep2aRM1Ul4vbSwJ8f
zYJLDRqFNDDGVStz/X6jP8gT6O0ZEECFAC3UvCmrUQZgOj3sBaRMY8kwZwy8s/YjRCw+HpynO0Jq
bZ7sXA/xLUbDqYrytYRFTgf5mm+qMS+buHet+2pNzDCZGtMxWIA8FYgLt456c/zSJ0aoAaIGUZG4
blwg7Nkxpy+0VMhyTqNGJXqcUNa1xOn8kL9qeurtzGSLNOn6J0ZMpv4v1RznUaIhep9FBKvMQcnG
A0Fhmku7wQQQpQ8cuRdi2JWmpn1G2Chx6pRmVdth+RhxT2CnWoSD+K7FxqAxibHepJW/850gP7et
wWar2Ll+vaISoBo4h0481F8Hyj11+8M7ZdE+58ThFVikd/ZhCAeH6S+5IY+Zjh5lFxE2cJiPhjxK
jiTVwMI4JgKx/iuTEtYVJToCE4G3aVB54uEdZ6KmgACvfhGVckltNV1vFUBXfcTQQMY/gBDgUWvR
3SZnOe4Lquke45NIYFiU2UQVBnDDgsllz1UKFz9Anaw5/Iah12ZAfX5ZgnqvUq+XyepVeuZ8VyjW
0BL80AwLaDze/qpAm0uorZyATeiz1JoGf7IaTzyNIcigEkUjFEi5qE3pn4VXzlMbWg3KMUtb25dw
UD1bpuEdnZNbyNXzNMYCVVDcIq7+7yS8rzBKxjks+6t1stWRouFSvcdQ8kxGi3I74xzEfU+gtsv/
3LwgkUebv+88vmSWJSlfNrUw2uLOX8tFNY/ZnIRKQxh4b6hcxNC+ADnTh1QQdhZzeqqYH9F+MMeY
sM4S8DQx4Da/zjrrqK4P7AlLeFX4dk3GEyZCpqgd1EPctUsmDiHkLiuIWbCpR7FJ5qYPlfNgFE/w
7nsFL3dTkVAjkKmCWGzCJyl7QoNYjkmNHctSJ3JTQiKX6yj1k4i60GVzxpHQMfg6KIdj/gJZSKKQ
GWZx2qONAEm4Lb9/uNliMAMOXOh1Rfl13FFEJcpP8+LAOMpH/POZD66JvghkNRkPLDQbLFWtNfLy
3Pql/cL99AlCUFkIVdTeaL/ZCM85yyCB2RVUmwwADJS6jt0tDcUfzWlCqa3+QRuTT9WBr4A0pJBO
6kPL6Bms5yUrFiP106XCS9YDzzRvR1rc6eAo5fJUe2Q18hET0uXZJhVEaG6FMg1QoZQijR/e0J/y
hRYvANoFnLNAWRoo82PJN1HDZ/NK8N6bVPsa54uzS5sjhkoWWDPVfP/vkNo7S3QvMSdlcF4+Sdjm
UbnvJgLDs2XIrk5kNBitN5Vwhx7nJVE01Kbd3+0Qs0luTXjuEQdS58BQdxvPOJD0TT6QFxA03o5/
H6Op3aUntMyzQgMGAIExyG5CPA4zUsjb3IQT+bHBxRZAfEdRD0oGMz/bbdL1lhcxaC17c2WODG4W
TLEQQgzIfGc/T0X+cSwvUArOY5M9TOMFa+1W5Xzrm5T2x0wtfqHts+D21AdXdlyD9OTAzV6SkEbY
JbuCwb5q1VaUQ2LtRCGa2nKXw3/48hHWUvEA7xt3Uo/qMzCvamzYAkXPXdm6EMgwYAmXi5XiYS7b
MwCF4Wiujs7lqWxf2g8zxKsrLkfa4y//ybwtCioptGqvT2fM95SbbXmETZdFOfedJ29qxhFBkF+3
NDiAWMZkbrp+9+6RVebIFZSlf4NyiWAdD5fyXnQdlwwsIALusk8NHp30iLjSVmufVQ/smUKwlqrh
8vma3GTls1qWwFsiiNSdn72caDFMOAWnJnzd5eISniNDrFkEpcO3/FGTWpF4Z7PG/jNtQj4t8lVu
Mts9tuE3WZ6KIYoaMsuqh6MiYOfdso2bn+KwsXf2SFJjIBVVGfKaBDduAzW90tBzqHyYymzCoODJ
hNpW/BjmeHwMEhhjuhUe1MGi0i1Odh+0o03GcgSGMQfPRiY4obXgkPH6VcBJzgNiLDXvcQvvMzAr
cQponyOAPyNohaqJ4aYnYklClTQXakC/LzCBaaskTgIIkSYBMDY0hp0fLLA8phKRnRpiUYSpmQ6s
OH4k/cbDT0+++OGt9CL4/6Gs0k0TysgChq/BWMdVoUhKI2B1bm/dEG/8wx17lqCfrmtQfeKs4ZCy
BvgYG57RyKSfHeKgsaJSkwOzu5vFFJD8WwaAhe6kd6hoCt/IB1MyWXYepHZ/WM3b7BwvIH9JfjTv
DNEuLAuQVmvPv2areibGpnlOaKFXqQuUOK+t6+Ge/6btZdZ97ensQF3UXNzE5q11w7U+BwbGF6c3
r9e+rufjTUHhm55pqbsH0EQCKHFvVttsShRtaOT+KCfFVpnj8Uj8Am5ui+3lgQMEWtGDb1mD5IaI
GgPOyV9jfKrkcwRWWxoaTg82B47KdNQrNRW2UUXXxN56EneRzl/1f1rLMK5reOF1okAIGY19zAt/
PsE05oJLVkriUtlf3noARnBlZszGNfpnkHrq6BPMAwTrYrAgc8hx+2hjNpV0jh6BDKekBt2NMLUu
TtWqMvp2xyOvuEZQCd6MQ2aoMvllul7AQxQyFr6xbso808gNVihATUeSr/gVXN3TIFAGK6iF7amg
FzrAhUPiF9Ap8SybI7Xt1L1wEPwUxrWfz7gzrpKssnqGK5wf5DoJOmdgn/qKBR7aB9ztisdzpF1V
kYGlSR61ByMWI6BNQf6Y2cKZMlBD6Vsn2qAZrI0ap1lE/tPgljK3/NDDiKHd/pjuqhvFs7X7Au8Z
1FJ/TPFUlkHB57mqG5+LmSrunrfbCEOh9vTFrJIL+RlxKQwIl0zzvug9d9M8hxn4p45MIcp6blST
dXPwMDVZ/DbTtChgMuoiAtzFZS4X2GYV6QlpY2Ckm7OolmUvMzYpYp/yr6JmegxXGEWJKZ2iZ6oa
myzcVwQmSQnbFfFBJMfOeOylZqh5DI5emEE6Tp3ZezH41/cmcsJbjG2uE6j87MNt6yU53OzSkS/e
N1cjz/qvY5MF0P8oHUq2OfzPDRAXzHWLqK4Pcp7ySGBRJoYSVo0U4+yy9gWm7uVpglKfcSnFfeB3
ohko/vGD6I6sYLhEJVMyfqUxnYw/IjY81jdBXAjiaY4/fJPf357Jn5Rk559VXOXk7QDfw38W+XKm
zFOGVhiJFUsymCzzuUFQY505XSQ6KOPCCPr8ShtHP86f+aAuQXrNAw+jmc2pVvqOKotBoGAEV3U7
yTDkNyQbSGM0/DYc2m6M1FoG2uWTtMN7Lz5oruH+r4NGPC6rz6ZcALWYbtMJqDAh8xZsOjoWPm7N
OVhihRa4WRw3QPJKcBhwy5toOzFD/7fiTbcHl8Xjhw3uLE6eaf5Texg/v2wga0kK1BbECg/rICaW
fg4NWS/xJhzFl2BitYKfWtjn35YWXb+s3UAWz8EUKD4/cO1Gk9U7tFb+UUbwp3kFtyNGJNuoBika
77kX2UDbjdZK93bjsqdHZywNisSr09VF4/JPGpai0nDGdREzhASoNyUSNAroxG1iIgiG9N0DBwvO
9yujM5kFio/NiljzmhhxP2a+M4WHSn7T5Wu6XFmjBR2ToB5UrklT4DVAx5/L64X2rXUebcaPKc4y
qzNOAY7nn/Vz6parkyZTAlg/1pD/1vlUjh5MzzppkG9DsKm6lnl9xqC7ZKKgMmjewZ8Jy3RXRRnj
KaqjOG2EzaXnKeXp+vgzrlTpPSQqj/z+X6RuCJLq7n0ZvwIzJrLxuvC+YlRcszaLRVTVK29dswlF
ShL1IAaxb4A6s5xOrUy03lN6gWt8HxFXdURylMZqMfBxnpFQ4EwyNOdpZ3HMsu77+Liz3oz632Wi
SwS6O7f+ncnd0A5BCC/26oKEpJB/XWXaIRMi41GWxBJu068Y6esWfo99nxuWfRMpTNqyB4RxHo99
H+dRGewAyyso9BxaWaMO6IFJbX0AuHvZXqt/a3upyghtLc8ncAJ3N1d6vYxk/RxUb5jD6mSJuyke
gSOCYAnjlgf0vkj7vVHzlYnfWycMW/1Ab1Dsk1sy2daLX9GiLiPLAg7wCr4aJTGLt30aUGKbcPsT
hPq6IjCQhWHGlkxEpIloxS/w4XJrSzhQzkUdHIFYPgApikkv94RI2kbMG7rkH4wY3NLuRAMkRlEo
4oRlj519uPnPRa02EiiSet2fDmFwQZehOXQXQbyVD1FEMzgj3iYEfZQwOKplqSsUdhQeO+KVtqje
Ze9jjPrfT8RaPhdOC+yr3NyY8e2UVPSsLMKFpbg9iudoyyf9jFbPGGrRTgxy8ZNFcMIpmTxPXrON
4YDDXmGOtMgpXw+b3ARIKa17n17Db9VPYXAdtMJjlvSwk2SwGak3Vyps/F9zKGhmn7yR7sI5O8CO
b3dS7czohstwA8FyqeaRWty4ZQeFHpkYK/aKzx0jI7aUJPejYe3c27JWPAJw/r1ICpIWP4gWZVW8
NZe4Hm2TckXr1btabrCJhcx7AHTKLaOjADK/lQyw5i3pluDn1NciDGjjy7259rAoozdsPKbHsq1d
XSsRZtdiVJ67EoILgHHbw6hEOX8ASQ7HPogh8mQ17HT9ETGpWXFMnOnmCgKtBqL6jD19vfN1YfIK
gKYnA5TJSFnhXUpAAQsV5KCcd/TMBPPn45691SosL3fi575mOC0NbTuoQrnHW/D7haMOduh5O0Zs
wj6Fep/rR333BbWohryWXbl6ssRdnV1cf2eZWayx2+0wNEqnnLmCYeup+tzMb6Y4bBZLMe45dR+L
dvgrl+lIlYAupI9q5z4DR3+N3JpYZNWC65BIZLV+s//Q7UsGsHKwCzbhXFXEL4Qt/0blrMQIEv56
xdSC8o5EZNp6BzZ2dse8uWQ0+PHFcmtrwQVkKoIbWGGnEWV0BPtfsCuhOoVULqZ49JONXDVp/NwS
MHRsEnQc/Fl4PQTuJdwKfW0I/TrVMHYIZX8DqJU6ap2o4Hi6DRnJI6241WjCpwRHa7HM/qInesp/
PH41RqPD266uWo3ZO4t4OwArVgB/a0EYEn2aaDARw0ukAQjTxFaMHwbd2ryRbmAexKSCRM5BtmV+
zqHRJnjEgj57giH5q5RFTryib2VXRfSm1wUaklxGRjGFMtKyzsVVWlvf8M1ydCahyCHfNoIFZjuZ
tOoqGqnczYRDyiW2fkIOCs2z+R0tK4LS1n9wffoOxgpadavFrhwdN7eFVl3t53Vp1j7v8+PjnmEJ
ILUh0np8NwPFf99v2Q5cb9UMfUthI/5TZ/RA4tcX8+ULrLEmuVjO5X06jw3wh/idE5A4f9oztEcV
UF8x6tDhWvKg8lbbHJ+H4dGWpIXVZjvEtG2vWVZ7iJGWgkqhXq+0B+xM8B9IRHqVTGL7AEhnX7Ur
u23CaFqcQaLiamI83wHgY+O5RWabVG4Aiki7deoaLrWe5TgVy8kKxImfLNCjCNmXilzjePgqQOjb
oQhEA5Y3L3/SHu1SaTS29d3ShG6TTfm8XJlsN0QavST19439WNenKInQQWo4Ge975kdx+wP9GSQ/
h/r7i0Be/rO8/YuFJk5zR4ix9rS8uu5+xKDBecKfT8quV+R49qjGu6oyPBJah0VyLD8jQLSUnCyA
Bcl43zYj2qbluQ04fKUYAUkPzQn3CHP/JpEjkSafVKx6IsbvkFrkQ2LXwMyotcWC+o1G0RoPpyfI
50EvIGN6CM9fx5N7hcWSenwtXQQvr08kDy9tljfG+bJ+Z39RnjkzfZjFzv4n0ZQMvbrFZhsfkvd+
/4haKuCbWE0LQmT1U9YZ0u+AOoKvEiAzuUuhVEcNSdtO9FbiTOOaMLo8FoPPLgdr1lzfQ0tu8Xqa
BhbBEbLWaZAEdSG/i4Uf1BUk7yG5xkhfvLRZlcM0NuddQsNFrXLP7giYEKPbbtyO3TZbg65AcCYU
KsQrphtnb5gXQZ+JmYCdDax1CFw0mQl2mmSFnngTynpW2xR3q5Gd5HfaIv2VyD/yCD4T+Xmy3oh4
1nbWwCBFIz78wx5aK0zETZUasVH3uM+DV4jUPCVwaRIJ8jIMORyvv8qaUxV7Kl/W7Mnh0hNM74fU
cZcvsVnQ6Sd8qjnc5R2Bcy5bEJqKX+PpnYTiEHFMk69cex7FPOUJoSNLz4/MDazmm1UBFEJIV4Se
cqmaiQumPZZ27pY1cGFqAg4ZZnT2gDLJm6k7JIY4OWXUQpdR/7GZ74KQcIDoP19DsuvgDI5YpwRr
Y06nS+h2MKNONKzSdqEpGIgSS3p6UYof4YsMkSdJBO60zUygqJDKM5fHUl3uPUjjo2blfV7FS6Sy
+VxQgLvo9BBwGeheIrhQGQDCivgzZ95vVHzeAiKtDgfQ3jzK4DcFXns5TRqUk7M0g4llP4jdW/YS
AH0bvsnBLd+h5Fy6kPBMMbOsfJ0p5vCsFAPeYH7oWmaUb93AgfrfNsa+3ZIyKO/drFUHNDK2SSbF
2C9DIB0QYlWLjLhk9NV/2tpcb0Kn8VX5+CXjpoQwnrWv9vV0c3IC6tNteRZ6yDkQXh6N1+PbFEE/
44WlTeRtCfvg483YVdDeucymA8b22MjabT4E44EpJV74m43ClKKgc3C7dWaHZUwE3ILQagbDkUYS
UImaVlWfUS/Fw7MMnPuYzL0GO0HZ2aSM/zlq2eTZhVEOhJSiHZg1JTnD1drkVBZMJBZ+RKAz/plt
k82xFHyAelTO3WthNLWRwDJbrXOX/6EyoP2IicveuNb7VXu+YlIMuMAIkb6qHC3o5ZpcpPY0rIZQ
Rwq6WKihQSYrFk+jZx0ejnrQ0rJr8OY/Im2aE2ebQfWgHN1u9yQoUmqIbQCrvLex9xGJ60dnI/1b
oisuUUy9zNfsD0SjhpV80vdP+Zi81Ixs7w50annRYR6whzsqpvSqI+6NvH0iX2ivqcN17DsxE0sg
2RwlbyD2/Q3qJQgHayjsiUtKqGSxnNzMCVmmhHmMZzWRwl9FnsmwDpGn6zxQRk2RyuJ+yhMpzO4X
bRSx/Gv5y83abf8bVKkGSdcviIdFun6P71rWCMXGhvUWV9ir8RK8b2XtV9dWcpzUg8ioHf3RGuYX
cm2gJP6eAfEFUcVNjQ645nWIzecsL2R0Zi7n//L6GXwzVPRilJpXI1PnhL3dxPFl70jHQ1aYUvhf
TZCPu1iJMIrBgnmFk40KsVyc/BR2bRGDFJh2IuBZ+qnQiL7ewbwrr1YP8DXp/eE5Kjd1oqbSctku
IqeotrrSzymTN5vFQYV6g//VAF5HX9RVpecVTjQxEDHSfI/2HLCs+6p5GYFaMHNKv8lm9MW5mB0Q
wD/+bJkM4HYtHaPlYC/DvLAiGBcReaneO6c6XCpYbXu0SKuI+/etbKZuRc5YkEaj5QtpV+TbQ+Zv
2Lp3TZja7liskF+EMK1PsAYTDrFk0PWwh5Ge1+JSjxCF7Xi3iwrWhKqxN9cy6/qj+gp4cw50ftQT
QtuD8aVR95Ty4F+bQ++W74BS+pBe5GEzc2W4A8ABh1HXxRoVbSUC2ZQr63DclygCytfP/jxBs0vk
s8iLWZL90c5J861pzUBuae0KLiP4qv5DzKgq1rFDpVPvJrxiVzX03dLGYjxYeiCy1ZlviXJo45C2
lW+0xL5wjwpKQ0kIEuREpTeEd8z6lBkLXDy4kf3VGOWertmu0KGsXiTTGYYZCIT02D71wrdecu3y
DVlPfS+KnwRsWUFSBGbkNy/TwkuO9oOD/1SlmdQ+tINXPtmuJEcg6o45Nd2AqZ5aqkCXtEtFbpMX
ZaI30uAghmepvOJ/8fYWUpgcenn+VmRoXt7cVvlqKp5ooPb3j8C/2pHc1sH/GWOaIFxI+6b3sQT/
xIJSNFyLlBX3UKWgMQCNaeW5BHcAbWlRRN0hHxXlf1ZOmlK0LCgPXE5YYj+EXJ5tGfSGcekQeY8d
f8Cm2JiieR9sJ9qbNNNeOCBuYVGbRkKAfUnfPl5Z8fRS5UhxrEi7HDVZAo60exBXwHQygt0zlxNN
mWiyUs2RX3BCMpiys5O4wTKIGXVudjAwcodsqBIcpx735CD8qeFYSmvpiteSo4cVcgKjcyGJst/3
i+cWRJd7zCG9J8xSs1SHc+PFGbmp5u/ufhm/B8wCVe88GONathRCOYglLVxNdJwTYvMZbmgnAusH
IOC+6g2fCgkvS5bmFLGctmcW+RgtHJePaIEGF/ArdBiwGt2ZEcX97XWE4Bpbq6T5+fMXzOB637r5
FevHc5NWcHpLPHMpGpeRm74a8rfglOl0ym7UICSiFkJQx9BmjSvmMN2rjlRsHsV5YZYV5ds0Xizy
E1QfJDRaPIhFTVYl+XRcM6xSRrg++G7+bZiYAXh+NSNoHu2/TEhCCy62raST19nU6NL/LfbGMnwe
KK6a7zFYM4W/jBmI6mavzSqpsgIS4wrPBn3b+2t6SpckjcrtecwLkmECVAyB5tBc1k8da5ImCweo
5JNvb+qVPps8xs2QRh5Xb68eyggGMyEItm+xu+3T9XABG4t8jP9KoIt6at7GF4ibQ2FdATexkZEL
zo5jq49UGb+h9DfQQrCCI73twMotsUhWjv4T905ZqmyEKLzGvHe7SNWhkyMxk0P3z5RfPMa5IhPm
8+G4dSiULzYHHvxUJcQig2AIEetqOAxCic4NiMyRqarRqRxdE79D8f+Ei7G26zK4mUhSbOvyhloU
vlrHQ1sI24Lm73DXar61GZmIxUru28siO6zQxb7oMCAcvhDMGQETA3vIRx0KpvcYegwzMY7xMV/G
HILA06DcbTvUzQUCKkPL0B4JX0IW5ArkGUYCCanYMDAYRCij2YnrBvkK2ghbHgggIOfH5Oju5fkX
Slk11M/pYLXduxCiCoEE6SqEK5q/5UZ4vWO7V4MD+xP4ZUYcUDkqDMCk/eZghxDtPesLGeYnVtcT
XYOxGjzcYvC996/dk+Cdi2JCwvhe6OsbM8fxWNqIuLwLrLKsf8zkipfdeIDcpVV2HPNQluq8DLWn
X0DawunNWr1oe+qU8/hXMdURiNfSroVFYDET6VUoruk0kZET+EEefTef853zW4hZpBTBUF1nZ6Et
0bLOJ1er5vThekKuQjJu4CrLy7XcopjVp89eCWHqiOnxQrp14p5mxp6aACA+NOo2bd9doj/5MmfE
iwSq4OPpX6rzvWHcX6uY+Mpk7LLnWxwD6+coI1ubkOPcKFZ9m2/clpw6zD8amI2MALaFEQd40VVa
LvCUiOLYQ+SQ7tXydRhSiVxTu6Cl87wsBEIGcFYMlKGl43hNNpVkLuqmGyQyJeqA1ncx3AszofKR
l/0N+opB4xudOUFLIaIIpQVnolxasIdWpQ+dcGZX8n9lErtPDd0/ionBcAPBy4uPFgVd9Tet5q44
S8Kiz6yna9B1BRw+lDH143qF32sZZvwQ2YSwPVRCWqgzgMVp0DgyVsz4Nq5ML6Ej6p/c7Sjo5pr3
2mNWGQdusHxxPll5ZTEUBFbWkBTndsqLzuJz6csTKLzK9zc4tO4ZwYHWR3RvVq9geyR0aLdZ/Qx6
omMxVz6tTjp2y8QwRK2m50Cn3RB5/rtrdpKOSYVHbZmo3BypKDNmDqtifFsw2iV3Sm/9CSOpj0Ui
M9N+AfJznWWHBlwgF720WVq8NwqBpKyA2Gq9iByUoH0ZPo4gAgaJLNhkuIB4w2/ja5TtQnTIWnKN
g54wxkgqJRZMqHsgZONxAtRTtk80AQpUVounsQH8dOenw/u6gtjsanObdrw6Tf0rP9hKYmSbsxEW
rOvV3hvJFXiUksm7Z5n1gl9Vz8NwnJr/ugBk3asVDrG1q7pox0sHhqzU3Ou92meZBZakwWGc30g6
AptNb189Xy0B1kx2XG/3tho8myDJaxD9+AqRG4pcr4FEyTZX3fwSb0bQQK3mE1kOgjEEd9CCVJ70
HlYh7taDc/onm6+kSb7ZTGDhbXHTepFyZH+QVIavRKz4+FlUjKSdaO8UvtU27zM7tX7CD72WTA29
Y8iK6NuJzT2SXMnGS4tSudBi/7B74IpKP76pyd9Uy3/pgAH9+8OeUUEI3FlHhxbiJ6RuIjWU333w
mT7S3WxMABzlG/8g5IgVX9LlF+nC6klTSutlW7R3QxZaWl0Nj3xFA5z2d6pFZu1nF1PhZ4niH5dh
3Xjcn352vsE9UWKR8J66TBq13P3/nmrt7te9MuAQNuBNKyVfe3iSaTf0IUAsM0LTPdELUFOtN7vh
pPEFWn6jmsSiOFFvzXXG/IbUsrn9xMu2WYtF6SwlJu6r9iHSboA9vssA0WX2kMxq80dll3jzA9iC
JL3s/SC/vwq87TbTIX0k10RrSWV5BgUWhCi44fAKIoGkWkE0WrHis3urcHfX24inXZ1wilSxT31Z
X5BtI1fvhhfNlN5Mn5d/cmdmwK1OzflTrKPXk1JwYG6iXLju4/ztTrcCK/VDwuOURrqSWrn14Pn5
XsSe41YSEbJr5PrIlgKRsHTHiOB6aYjR1XsXBY/CEbtvDkEigmKO3ov9ykOGlIrS7ELBYrpGjwgr
tj1l29pPYYOsESZWGcoGlmwPWhm0ZBLquGq1h0NE8sQExcFeYAYU0s6xShjaRdEpiXbnn2asUNwF
6C7i2+fYvctR6QBzgyf6zsbmwNSZnaPpdqbFgBZnlBt+TTxccXIONq5DQGs+fgVTNxXmGKP6w1zI
n4CcykFaG7D/cUVcjgG8O6iPT4+W9RsZe4LRoIn0my6zrBUm1lYF7+xeWQjsBQ3xTkuduYoJRxmf
RqHcBK6tI5RnWn/7HxTCSyLboNpNmCBJazQ1zXHyXehPqq1MPT1DD9/wKdMSI32sYOWYAIX20kvr
TC4AOEK3bQ1GgicNIUyD7T9amzPA5ksEQJdegErn2f+5Iv0UNFYA7S0EQwbavLLyQ+EnY8rhGLTC
LSUajSRIyRAHdp2dEPduwr8zrGi6Ni58cWkqB1Q4sniPWfkFvejmtZXGsGDWE8mvOvuYgRWleO/Z
9p7aNsQQBTIB72eAEeD0HQ6CgydhVmP2OHXpW5uICbTPtgNIvvGolJlMNfKjrA1YSZ4Eqj651Pyx
jR4SGiMDgt8ny8h9wkZlLw1laGEzFDBwx3aMmrnl0yKzPz8FT3ZMJRK6tYrouueMINR2UHrpI4sE
VUuZYCnyYZZcxAXyuGvimrLxXcQnS81GZg2zoaY8ptrrG8zfnz/NJ6cNsbFWcTaHrz/JNpEluTFP
zOt8Cs6e6ctfBhoUvzIBr+eQtjvFkqbNan+z/WYW4BeHVcidnwckFdulDqWFQG6CSdJoSgNPVXIO
Ao/o5FJAYUsK/hoae+GJWRloJgBjQQkx7Sdt7ICErbKCfXEEwjni42Gdvmhuu2DlriKhP8A3V4+X
psBOxmU5SkhXb3N7c+GlZ4pkDl91RfTDbJYeCSX5d2QEpvqVYyMDPy6PABprnK2IvenYXyHqFKLT
Uaw0y3GuG05Vewz2gr7ESetTPtRxY94tyfN+L1AXCKVdzYAeZlSkZJXkQcjFZeQK6zOIFiPWMzQJ
oFxl/sxNbuDkrQ3eFjCpiOyeXPZqjbz5UfDRx5EboTx8h4ra7LryH8oCEfgOwF4p+kDu4x5OXK6b
882NSnbwc2S8gHLawmx6VCLkXjao0T4tEcqmzad+kSOhIBndxuSh0PrsIbY8LA7trJUEIhwQi03R
qrM6p4x12sBSALE7PNEQLFDq1dbMYHiKwZiBGs1HD+l+rIewC8rcuHWY/K+JZKEOXJvX64xKLrrm
25car0+w4qpf3g74Al0iWp7mak6c/MjaUEkAefMDB3p3N+Dv1D2XRQG+f86N4tLALNJq9gX809MK
vbNki9mcwzvzdeKL43eGJLU9eopCftZAV8Vt6DDGT8xXC8NLyTTvfcOyfCvvb8eVf0YbxCN0o658
abm+d5dmMsHZ9ZPQcuCJ4NXyz/moc+PFcUCjOEkt1tkXqRQ12jEhy44h6Cflv2P6oyuBIlpQnXRf
HIGv9rIAFjYbTYrsA0kKJYknMZT5+havXoyMpD06P4FcnkeEwvBxCjohK46qSUL+zCT/YaN7qRqH
rnquE9V2Tj5xUMVXsJjcx1x/zm4tzdMLE0LycmSagfMlVYvPb+uzyCPpuA2QKxojpXE3GR+kgpL3
aY/XoYJqhFeK5cvfDD4Rg87L36b6oC/WqTOtepRil3z3Gkj+u9M5FhEF+x3dB0VKu8eDBfXntG3I
HqHZC2u8wr608HaPxYmpvivlYiw52EwdLD2UgDEuUJiCSenLvvqjLHIlAcg819ZUcz+ZB430UleA
5cB8edI+o0iotSWgdxdQqMm8f2SESEsCemiteu4aTSUlURAahNWXCQJpRpsszCqpaN7UBc/8XJ0K
6RM2+43Sr2ZDPDzec1cbM/8XygdR4e3hOaaMz/ZJlJrtfCAIrdto3Hm9Wi7DXr0pjgGYc0yQMyad
Nrn00nlYanytVk6FQ9HtNeaaSn1+S0UbI+O2j3pjZ/WMj8Swl3bjapO9o21hjLUmcIt9gwEugYTN
v0V2xIok8Xe7LtjHcJG8IJKPJv/6CXULEDEDL3po8jlgkFhP9bScVotU3uLVRsVXbp+t1tXkSSNq
n9XoXYtvsnLEbT+yaIn0zz3jkECNVPj0ICCGRmXsA95FfZRE2AqHksXsjD/13wZT/r9GCM+dcmBe
tJxq+1ltv17kFHyFKli5FarV4tiZX5jOzPiqMORhSWv96tQXgyp4edTYjiHZu8+bmfer1s6jmgYG
wc2jBXwC+mXiWKKP611DXwlZyF8AXAKQ4we3KuvmsseeMIAtJim8HCX6F33Lnexb/BDLPjm+KtL2
1TlZ9EtSV5Mwt+XBqzYKFVzv68nsCGx8t/WgnmsvEPPRRGkzyFqK9jGZmiiZSZR8I9NgVQbg7dQV
YAy6O0/HWp2wr+diYqNp9dQ0F1XXpwDg7W563AzS6q1XwGZchif1pKlNEycOw+MQLJ+1tBOjrFft
GgRRg6wJSUtwdV4YPasyqpb2UM14WhmHj2wxJCX8zSt1FT9RYmB85IBsskZL0GJQ6ovpWZZe1Qxs
76jJ2T/8OkVjjVD2Rphte6ah1PV5u2zmbzCu7WcFQ6Qbx7U4seEPz67NLjC4tcvSu2PfSpWiyX7V
Ds7rP/O13j22Q8D/jq4TWtUVZRd4pdpBMpK0UCaPux423rDHIDRLh+GDiJU2gUDkqFtcoYEfh2ID
wEy4b5z+xddJ+XIbGALKVdI3M/lmv8NcuhytVryqv3fCiiMxcAkr4pn29GanI/Or2w8vlTtv0fQt
pM3vsiIIx6wDqH9qitLmbs4vxXap7lvBTQlUYD48ktCbAtIEXBE3VGCE37PV3ZQtEAZmIu7Wn4GZ
QQYlb4qyrPIPP5L2QqpHuLsodXfzJmXVHYNia+76MeDyJW/IHrAq35RDJiq4NKl/8+m4MkQQT7VV
0K1J784zg0WKBswUGasWsM4TzHHyPpy6wLgHFnhN0zEOBeAEC+6RkeT0hyjM8VK2ZjYnNNFcnUPW
Ul4FlzSSQILuWMObHD6p3TxRZrn6jjrYkkwhJDPKi3IyJrgEj8ONkzeukYqurrMUqIRdKxaqGZBQ
pX+VupF5SXhtl/y5xBOuAaAL4nQsgoNKtM2PNDFsj5C6gPBn69RD8PmHA4SgsNdHaLkZCL+iSzoj
LleTiIRu7lSAGbGPXNrWERAgYLyMmh5x+vOy9fQXFNKu7s0Ny3ov5X8/fUrBvhRRBcYV2cjDMbOx
EMds5OYdmfjOtldZOeVsdoTHx31/44TQHJ08Zx5l/9Kt/TCifkCRguTn0pieMUWutZIn2uWwfm3u
AhIvxTFeOuuHp2QE6G3sMxMAHH9ucht8Nwsp0Q1ZoBimysLlmluwVbwvUizkdiJoUHZJzCPQDGJT
2J0TLdtTWxZQw0Ww68YmAFLi0EgXU5u2+HNPjOVDcK+BUH3XBwsbuhqYvRGasURGDsQgGDiR9Kip
fxKqxrXCQ8ZiIXWW95M0fLEUe3hAeajwpFXxkchhLbaGyLqiNbJ/OhAedB/XisjprAD56Gfo7Uf0
//BH8/h+PFh9ftaIx0Ea89Gw84ckggihi9O9u914/2uPCvkJkhZ//n3HMYI7zxsNoreD9vm+zmpj
LJM+e7jOj0AByPY9/3i+dDoSqox+Lpf7uU/StjVHle7v0Vg9XhsNvLfVf7rG6tCwsUVe9q0vyhEY
r4yqY8Z7Ta66xW8NpJJqCyhNjhOGCNkzZDZbYvS/PUhSysMRg0ZbPQRhCHivr6GxI2DSYkA3o/F3
Qxe2FokEGsooDLHw+Ux04WCteVV/EEyQ/AVxRt1pq4b/cXOyHv56bW9pNInqps8ahPfboe34bK13
sxvxh+oFNAjGLsKTz853C7ItxKhyLORy8TtnqgZRZbYTWhyNIlAHX1Pp6i60gwjaxxjDR5LYZVFw
Ncif3kuhQhPk6kytU1YUE78TM11/GXR2rpqLHclfctgFfzIIfXzuYZb78njeoE0Ehh/rRkLF7Nln
mSYVNesBh5TgCZ+Aje1EevTRjxvGUt8vZrttiuMNhQSpGzRJMG/Cs8VGclmJPPfVCQK3AUehp9T0
6Sg+RsWBTJdS3utU8qxreoGPLXIBAGLSzdG30GYQXmqGr5B0xzQJMLC9eGCjDDo1pBoDNFd2dJZB
u5v/5tkGf+bNEVvv7W7BCvoHUsCSrCvUn+jDqsuJnuh6J5y1IHqKM5wxnmS1Am9/el8AdIxG9OBV
FfKHE0P/02lhFYSYGJ1gOw+Cf62kCPmnuJwyXkiavBQOFmMAJsMlfxKe+MIs39qswNeJg2VcFeWG
ykok/FoNua8V4mV/9+p/w7mqV+hz3y6dRMsmWoB1GEXwgKL2mVHde4XD6BL9m1Bk/FdWpMJNK+uA
VMq2apd4bw/mRIiWrNiPclmcYdKraNr/whpwhsinosDxHxcDx1lCaCx+sNbPiIBsBTgz21OemFne
ss/3mziPzHzLzJvjdwKxH+7xXQ/hXyqc4GBfdqUInA4e+FZtpFRzrrv5uyXphnxoQDKYQKgHdXn9
0PEJZ8fEpwpysD2Fh0NZ1xi+EcKlJw2Zhl2AZ1tCdqd7Qrid8QwC5uzVbwjiffVgqbQLSONbgKCP
jeHbwu02vMN5uPY8/oHCBvVpp+j1K2CcRWWhpyyPg0B6deL2Nv3oZGbanoyTGejLkYg6Xf9yQnda
XRU71TVAHrw2klX9B5xjSTF2SEvABrrrjb0067q+Il3Qtv6nOGZk3B6Z2hbBamtBtY5pk5oBHzij
Sfroamu1wBLMtYDxDjtsUqiaWimLjOzqcUvDqCAC7GiRSPTt1MtxN4S4Vq1fYVSJeLn5DAz4Wwx8
JZ5fIOXNiozKC82m7R1gxN3K5BYYaHHc7v4YSzg6s+flN7HAOX+7Z697dKUFlUsyGk72mUcqqKt3
bcnBnEuSJchWyHV+5Hx+YilfOJBO/8HAChUA0su0oPyKZQ3l40E6dpjAWOLqrYoTIJokN3g9ulCv
dNgQV8dWh3dIo0yfOHPBsJrZ4wMF01kAYza/yNYb0sLeRmT8EvwaCy4Rw3L3kWqNcRp9/0JaNwrN
UIaLyo978A4DKmCl6qvadQ5aaNECoDDNLD87z43+0J+FdDMe64bOZ0+fDpehjhIEmtGSM1cmMd4w
nIwJcCvHAwEiE/wW0mdD+rlMdn5Nb4nyKpsTjfloELlWepe5tR+pngnmDCEYoHonw1GkK7yphFKU
X9bhNMjPdKySQGWwUSZkG8CfeEEoKJPERXM1PHuS9SYd79RHtqs7jM+hAGhwWr0AspDZ1CBzjp6g
eXqvcoNyL5FtV/+dZncfooXo3S9xH9Vgg+vcyuddxNK8WYJ9I9k+6Cj52CqEdVXhNoVirYXaFuAm
CAugt0Xjmu4ihkFbbQXmthcLA0s3Gmq7V2s+u55Gkhywt+y968jqtegku02YKcFxP8MXRVxprw3G
OiYNBcexIO8L4QIfNIxo5U+JgZr1pbjN6B8b0WtIwdS/vVZROTUAd98u/P6L19PqZi8uOAqtqe/w
FIlq0K+hyY/AkFEJLD161JxIZFp0VetpUIaTZk68mkhEZugDuQUb3IO+1fBkVaayhXlcIjck98aK
UDFJv/4zSsANDKNZqJ5KrWfDZ/2+jG0INwtZA0e358Vbpdi+zo/DwvglTYyOaD7KUj2S3GXTLIbx
W9n9qqBRN4jJkH5NXlFiY5lJi3dEDLcTLpqFgwpgQzGeqXBCM5LymKqsbHV7+dJV64XgsnYchhS0
vQLZHZOMp6Ll1L9pfATyy4KDUrJXUWAZaPACDiy0Si6CJ3QcgL2DB4/YHJJqNiBrMB03n9R3Kmmb
4Z670n7M86CQPlWNUuqBWgDtrRLcOjtrIU69j2KEXpIltO8EdaM9w6q2hhLTS8sAVl5hp+CKvdeS
Lbs2GR38A8KPoJh+d80ubx4mTjSjqFB47wFdx4xNy+QTSEQDP6A7pPkaLvv6LGBsMqbVAWtb6uRn
XF3yMbvu3xTSUUJxtJ5Iwr8jQ81sc7t2aK+jOLfYA8vPToeafHNf/S2ZZFo4xYx4m9OfLEBeBgER
Qdbr9GASZR4tJVmEqBfm6lfF+0icUE/G4AU1JeeKi2oSzwXkjMUv9qgflX0OhMcewGRltpaC1W6q
XgIM+sTlBw6WMIKcJ+03YuoOYhTD9m2v2QyVmHUSdCLx1UkUQTaL6qm4j1d/hCuk6IUw53p9F/aL
45I4l2uHvaQ3zZ2lMxiJFQXns5sSe56f5QhAI0XEvXMaBAJpyQypf60T5ASljqpZnGTs7oN+7oWr
cIGRVNvXRO9UeWjSdIZwMCexTm6YKOpyTmfyxXW5Xtx6cETXuvZI3cAq1Y7DRio+HXJXbS86c66L
Exuywp65LjodVq6wiYiY76ISyveWhFbAdu122nYp7kB+Chbi0sAa7059NMCe0fvafE7ck9Vmgb73
oSbyfEWE+CVDlAV0ZB+jAK3is0iElZ8IUnUN/YNDIm6rbgt4iz0yoHNiVWi1eo7wARXmQ/jH0oKd
0yPJ611IS3s4xsEiHKbjkfX5PYc/K7fuTzRvGeE0xSZq3ZPNoz2NAggpg5To2llLX0xn8peoH7T6
CerlxcbBFovubzasT8ql26OJHkyPtT2Xi63FajPNcKMFxuCZVlAaVa3d1z5sjILqYrUUeL6O8eEd
V5dJVj95MUo0sunFvSI6zJXiwnfFFwHM1juJGUki36bKHqvcvquOSSX33+BQTD8+MUoOTtX1E0mb
mYtsM8ibiw2Dp55H9hAOjNUdw+PEG8ICvNq+HpRFl+6sd04FXO4Cc9XNJwXMhEnRvkbyt95Xja5T
2s2xUVMJFAK+O4dPoqlqTEP+/p5x3hYpPw1yPkYQlT81t7qrMYgU44lRuBr+SWmggdG3SLnBOOGF
KwHV8PUbEw0AP2HtJmYsHBgBn1Sa/UHSghGYqECDvnfmNPWV92kG/BUkDAIErREn7KVjMzQ+HYoO
rCsPWVa7R6xveoBAkHZginQEgKTCUdQnMB2HBkNN6AFFXfL+VI+YEO4O4Xur5SetXEtYE8cm2UU9
eZ2gGXwrbafEqYcG5vACwuGo9nfV/SeR7KHuz/e9IvYQTUjMniS/lHEYhZTwanVoRLDUMLhhqr+7
ty52OJVvswhgaeZNWNbAVa/Jb4z/+ALv2nzqdQVlEoRxhV81JJv69wztHf8lZdyK6g+A74yahM6a
EYKfcjIJzRFoDHlOcB7/HTwIIIgfPbTNzGYKUNkNHiDLiv7iOCdygMa+T0dY6TR/9kJxEidi9qoR
bHk9QkYUXcJaddnRtUSvcXL1PsHyY4AweB78qK+e5G0ZGLzcNJkcuhiTo3hm9f1vO7tVo7Nxtc91
qz52ZkZJa9crb5l+F6EuXYt6EGh5GnxZ0VyTuJDxW+H1t8TeAyN0/+1NgerGBtCax0gjyop44vq1
wrK3Fb9GNHqJvQ1jQKkNjuBpltgMMD3/hDMPSDu7zTctYUmNmFuwi7I+IIsb+Ky5R3MRnJZtlhlX
qA2Pj1stCcACHT7s+SaypHSZoN+z7Mc3SLMCemSq58zJ/WN8/s5HxWgeXxYDDe6O3Hj6xdO3ucZz
RdvKADyC5X2kITLq8sOco7nVsrn4cLS6aM2xGqu5wLZ0J4GzLQGtnNiFW9gQOich/cYY+K72xlzH
nD0XPy5X+DWyySbKWmR7D/kFod6u+b6gvBmohHPHLR7sAeJHeqd+JXAC9IQPLW6e8SdgmB54Vv1D
ioELr5mDdjvmdF1SMD16nag679qaZ9/O+z9kF8Jjw9ep7i0jAmzjXchF5AOd6n+6mEFpj97rHsZx
nkMPDUQ2O0MQafnr7rMUw22gvKZySuiRsS0sKXrfkOgYE0EpJvkF+d+m3U+LRdnCuIb9Yitl/Xtm
bvi6D6p2+MASkv7Nj1bbeTqPgCLmZMTHA3B1c+nnpxH6zViHKcvlTL9BFE7XSyWv4V23l5GlO8Ax
qkqwsnuM03qUTeO4UY/DE5VHCU/UchrRCV4eKjU0cB4DXSCHQDUNZQpAAwdxfstxG4CLhkmmU4gQ
ooCDgzz64UqBU7Fe6/BRI6hAE8qJUPKwEPMmo5SY4B0bcmsj/9su8LKOVMuJD9yEAzB6K9p1Iv90
b5Pbj2AxHmIZzXHNdLat+6sGg+YbxGdtD4FKINGU914a7VRC2MYSA5K3nZkpEaOEPeKEKdkw1asb
aow2Dm2f3qJpr34/jz+0M6S5UOtMIRfP42dVUQtHIffCwpMhwbvU/AoTInd3W2rI+5pPv8FYe+j0
2r3W2ijDDe1d3b9IqigwPy07kVR94hfhzTm9Ep/78Y1Wcsc5Z1i3U+TSr3gcUOpWFktpucqu6zEO
JLle2lYVje4ixc0TPqLUxlQsmyeV5CRoMyd+yUAMkNnwZSvG+zXLpnCciFO3lucbGxJE38eoqSWR
YhMGmv6BFjGDbJsSmb9lRqPeCbVFySDZd8MTpfCp9/1NsQ6D/Lij/cZiex5uHCgy8vwgGILbdWmX
SZaBn1+7XrpLF1MSGiiebL5AB4aQhivc5Soethlk5EDNaAXBRigSJgh8Z601hjWLjoVegUqVB8KE
rs7ddEnwVZNKkM1aByvteD0psTWCBJFTeN8OAhnArLLvfePcQxBO20dGxw9TKsvxCkiZyTPsEOq6
bOC9EqjJsHo/fz344PbfvZhLrCZXCD5530sJlHhCEPI9t7FuHTHbMKylzaQBjG3LhKHN0Rd9HP0t
/SsOHLg4XNAIpYd8O6t6p/hGX/Xw0r3OAdUOmKWonzZBOo+g29MwD70rJKWd90XfJ//5tlvKBEFr
4YK4e8EZDDS4edNjNQYMe5f2XEB42qkwZUlFDbfuF440PVpQ5cP6XDYjYDwgVHP6PLEuR9/LJgjq
3BC/Ly999DFROaUo0XnkVdJebs78UnU7vT00wFbBYQpviXoZ/qE28tnIEfawbFequ9jYEkt4+bgZ
J/XXIBTKDGpjR+2TDkJnVlFL6w5noPq/0LEdTLvgPVvUsCjDoGJPwRo4XuLm1BANBEh5pbdww7Ss
Fn1uLZUTnDcZH2cQEMkJby/bZMa4jwnSd9YCjBtkKJ+VTB568qxOHmT273LCdLPY9ri17Tj5vYF3
AK4uSc0fv7DHp9tdgnjvgj/DLW1iqjkKtCSawxaU+Vb9qmnkIOtwc3LuwXP/iZgZuQ7PTYQR2yIV
8tTV1kHcVTGj0OPX+rCNnN0Z5lUUOnk+KiX6l6yZzN4tncWc4W+PujxNh7NNT3WNX2YxiI1Oe+Wj
lak1hNZVXwElqbrTX6ps1xitpuo784Z0QKdAI/MG2mOf9brmY9MDsMsq18uOiELwYbVtEGl/MfU5
n/iAc5f/v2MIR1T+znYZ2O2U68ObeBW478e7hR11eOzaVDVFhz2G25f2j/8lYE7Y6std7Xlj0ih5
0XfANAz44MiospnhiUl3rj8qzXu9tfPX5PaNoP9ZpYplQsKLHOHLocUt6ac5MJ+qmjwCCjgtNeA9
R5qY/Tey0t+1FML8dP2irHmgwv0e9/FBmAzAsl/E7bbS/KNGiaihbOTncSecja8Ycwte5qu3bQjX
JfsprNyv2eNITO9bkfIGLxI170+BPibMk1sPqcjt5wZxpUC/sEl0Nc+3Q1znDWzfdoLNqHS+fcYW
gW6NKBUPs5nj3gPcUJFYZg01GWZ3zho8jF26n8uAsWzl5Cenm6xN8RLXMnKEZMyN39IumiWoW0gg
fPo1BvtUQaWVofBFhsaUQZKK3Zw6JsM4t9XcefdEv+FjRvj8gBoth1enXVycv54EWPND1U1nCN6H
1AfnpY1jdqNDBaDvt6PjXY7QlcJLhgdw49owPXEbBuFH+hg2cPCwKTnkYQ2WA7laxqekhnYyqDvY
Azp9QABDiZLbL2KZ6XSt94+cUHx2A9KFVr6HP01vVgonqbXW3Eoecu23BLU7yjHQDNIHfuRKZi93
IeNW7U5hMLBZbQrWi0s3YBETK5jGc6EkH+vrz7xlsloVfs+h3SzGFEey0yJ8heTSSvRPRoXMnsrL
x7Skos6Qb52+n8ISgdZdH0ynq+nF21uUe5e4yEE+W0aEYQVDQXYsCQbLQwsC+0jE+UtO3h3c6SUL
SGNXcj9eipHuOV5NUmKCb5ibR9BVnfkkXtLn1b6pTxtO6sLJVutovhxuN4e5wivzKaYutJeOJSaW
kM1cjaXPaMjONIf80ddSgmoLNoDUqkAes9yOumhwH39iXmHH5Y/i7BK5QTJx10gnyjdWgq6X8X+D
6J6KmU4LNG0es9hXg1BiPe3JqBCHmQFW4JrgZNtEzM6Jp/D5AUGaXEGmuoa/9BYuiPwQ8XpJagYY
MLgWvFiPsYwOZFu1dfiyX9JtOkO4wWi2Gp3UyNGbUGfQaIxJeXCl0Skn26sBWqyIUPT1d/Aq4j7F
o00SH8OzjPtJmSB1T7vFHHsJA16kkRYeIcEFVKI+sm3c69MWzoWZ7llCpIt1CcVltPAzLdiasjKi
uekntF+3jIDXWggXoTtwYs0yPVouLpVVZPFaxJ+XMXQp0b9fIa9WSepM+SltTIlkICYNjDDBmmF2
or4hL1hBCtw4yd9ugWfLJRE4XJeL84+3uCpsk7VGnGDboqZOJ0VZ+1cN5K9JhUMkXrqklcdLy3UP
ldmptG5lxNHeqhwtOQX0hEoG48ctp3x1agUNuBPgvEPc83VptuMXybjL0muv4Gc1lkbRxPesT8zQ
SI6EcnuTctVXwkJKrjtp1/Jw5UH8k9QC8CO7/8CdfPAVNcolmfi2Tqc0JxBGJNZ45ZhPKqnHAAP3
CnYID+kznplvlKKJuegWGHlKBzvOn9mQ8Bp9EVgLjhmRXzkz4DbbK4m7Rans/1yzG3keFPgavCZb
hzbCzwZGdh7oP4OdtRW5yhn9XwDy3BIS1GRiHBDllTcXb0BhP8YQkGxqPXXRWEjBQKeZ4fSl53eG
2BL1ZuCky/rjgDUz9vAcOBVBvwXHQF3wtKvP6DbnhP73vWXvk4bQGc4FNTrpMV7NCwU5oCNq03E8
B6BWHNNoJE/wRsVDvlNjOGdpkpmDsEGm/o+Zw8xAhVautxv02PpgQQ/XexuY9naqnKoP1KdKgwFU
2I/YVvQaAfwCk4jE6AT+3HMkaQTlJBPf3UIfiYUliXrBs6otVn1OqdSpCaoNxsxYAGaiiuKaxNCh
5Vzjf+WE8ELsujnmdcSTkMRCg26ZM+SBobEDhbUb2MF7rmx2h6dxiE68mg9Q+VIWywpLaWZ0Y4b9
y/1O0y8eNPW2GXnWi+XYeMbnOQqIyeCjvZoU0uzSUeAo3loNqeQNPWaa4Dv6SM1zTRLiKgYeAvQS
QwHGjdJXww1TPs+pdhbVL8tj01ukx5tJZSnqT9zC0jME0G1TD+xvyrsONQ3RvH/e/E+Amj2sQ3U5
tIZPca++xaNTBfrNW6HvFjxVmGFoNimk8WvcDXA2W+1RY5evRnIFqz/RNcvNbiqFf7Dgo60JvOgW
90L0Z8f7JL2fmAfvzV+YpZuJQjtGcDLFoZRfF0Nug1A7zS2m0Hut68sr87sDm0nThNCVYmZsmhEv
Cef3xp+qBAro6OQ6zNJwwi9qeWwq1iGIAqFtRCx7SDy1YKoP95sSvSUZCUr1UrYY45g/RftWp0Rw
joKGQY+hYI7JcY1rq0PfVp3EEMJL2wMEVLqPU3c8HNSbH1T7j1jEY4HJXv9jKn/wblU1fKAPDWaz
cjsH65Rribrn1WSvQkj+XbpfWvGZ+P08h54fBDI4zrX5nTrrodwvE0ma+klvILEAhKkCXXNM5Zxh
uVZIapaR4SSCsqYUZi9CwmgcWON885ZmwD05GxOl9YI/EftPvFakCMDk6YjQllhC7akttvur/hVe
xIpk+n6VHQSoeRadGKdjBM+aaM1zwfSD+03VJpe2x6paaU8/GPIYavJD0lHfdEE3NIxTWvYxWoiO
YUWQ2+qLUT7Ld/CIsBTQACls8U6xAD5ASleVxAfoT/LmEFsI1BVZza554MpW6vk6jEe7uaq7n7pw
RZFhsUekDIfcMLIKXLjFZwnHYUWFEYi+ytTzngWT4hYvvTPfNGdEarFgA+fcmn7Xxxe0AnSgiWx7
he2vT3BACO85C/XuEUC14TzasP+3MAHYyH05hPl2V5MgihCEfDlIWA1M17JGw8uKg1K307aYFPbz
ymj+51be69Z9EkvJcisuyQxwZH+pz6mZLRyvEVH5rR/Sk32Cbmwfctb5m1BsbLwgP/j3wQTN7b4Q
iD3DQME/jcsX276XOwy2JGoqle3ocz8iv7QdBlbVO3qUNHxU+Fyjs1w0XD0EhP6ltjdQ40ckjvZb
GqHV03Awwr59uLghCYIbHufcc/uKsW/ZRM/gtDRHGOCk2xNH9/8UhC85BXAWQxi+p7JmrnhEjj6o
ZCCzVcUu2cbyUXl51yb0QlYZmiQjnRiAW1jC4Aili3DaRWegV79pB9du3iHP2aGvi6QdCZHq6Ecs
QijVfr4LNG1QYGUSSmcE2pWotRSzrPv4VxD6uoT5LbPFJOCwWB+gshLbcnp3LBCswfoMfnGb16An
UmyRzu4Xe6nh5ZrFUqXpTI3YIroYz+TisHE1VoRkzae+U1l+FLYH9HAvWS3T+bTaWFft6PfjV7R1
kxqFO6WrVSzcpGw3vjrK6Tks++ErWGVGE5GoHi5lYamiZEJe6Z7oPx5F/2e91/X0elsvIdkCPN+h
5q0jzHB69mavWr/e2lzTsBxMsw91nMGFETp8MAp/uRhGyc2flRUlKrPv99uhtln0JDhiLbbA66WX
YbhLUXl6gyweqwoIKSi40LyVc0siEXQB2oUItr6zO9Jeh8/D4ZkOqiMXHk8kr/fmwpoCTRYa4xvh
hl0bhVkJHWDLMKWwbuF8gDl++jNStBd2WA8EMi/SYMBohsKyXFhaRPsGU1OY2XuUOdtgnplKq7bk
harqZOy14+HrHazEExNOm18Fsx5SbL9g/Uyz98A7eaATM9z4ajcOnpD5cu3CCmWRBe2jxfmHvEYs
ULVFNl9Ht4DO0uBZWiFPKnM1d1VUX6F7q9DP+RjREbzixZcNyw/yXw0HRBfOirqJitbxjR1HUREU
ZI8KHpcpx0vnz2aG/yzdLxI5aCq+q/I0LGKUZlnPuEjPQJdiJtL3Oq4HK1MjBdn4mKvxmQFFVIG8
Bf54p0CkiAGbJ2PAqVdsdRZKU1Nc6+OBpEVeXGLBA6a4bvnEVXorPcIpNCVujtthElWUGImCHZR/
sNBSLF37wJP1K9M06QIFNOfonSzwkHrxkSo0u+aVFWkY/26XLq+qZ1gWEJlV9N+7SetGnzE1UJ1J
5kya+/OlvSpFXO9fgKLGlncojMuJHwPkBK99m+Ice8yjAeTEVuJ3uF3i4kIDUhLboNaLulsyWm4s
CtEQoU7bdeDT/yxWJud5FRDm9Gaew0TwOKYKbVWg6jFJeSR3FtqE/YLXnxZ2qfPLYWFPkZmOiaKa
WfgAinMpZKIHRg4qB7wri/L9IdeNV4BSXME5OiFT/cGCRdFt4J4ycgW48FWL+nDaHNbXi1oPiJf1
izkoiYyAcRVMU0lbgBQZBBoEe/E44BWzbUzqWJyuuCNy8cS+KD3x1qQ5MKAZ5xZk4c9kzCM6mjas
MkkJtudAtbCStoJUCQfbVjF0EMwReZApO7x2GnvG/QoxwPMN5Z3yKbvK5+0ebDoppFfWj2dUrjZm
vMBkJ8+IxmhwFvwYKuL7RnLEU7fSVGgtztQbG9YnH7tRrP1Z+iIaa+7YZU6GW2Xz0KoCFeBXdXMC
np0q+PpRRxTMW9PbwIGxGLmE4sOzsUNRlLc+jycaJHgSY9675l7WMxGhW4S9T4nQ5XNjkpbH7R1n
m3RD2GaLbrMCNhblco3obft5d81P5L1TTC2rCeNX5NuqCOvhMS/m7ExH5cfAMIN2zf1xy+weCtC3
kdKtDgEhWWK+Uwt6qn+OUg0E42BBDniO5w1MymbypacCvXC+iwIqxK5uaMXUG+ZthEN3P+GwxOUa
H1U9Kwr9qssgvi5Xn5s45wOjz0XdgDUb9NeKvT7GThjcKlIRdZJHNukYvVuiGZD86yx1ENxwCmYg
ExCDGWo84kxjon6AGBzlTbA49wMAxYo9LsytTrR5LMGZkC7rU4qGWYC6e1mR4mvgtHYiXjW5HXua
MJjl5uFf3ebuGaq/GU4HUX3A1QlBQcTzy3bDmjjUY8IZAwXofvvDqSACeDzfNgQdeKKIwX4SvIJ7
pOLIs2IH8i4knb0ZnqvZ/teEVTtXVTH5o1NJQUzWXfogDdhgYvtzOcvfqS5ILlhMh2/Y42dd8uhs
9d8gtGNALPgppoJEfryTxAMkvY03Ye/M9f5yesmGqzKzo9BRmVSk+uTkZSp7BXpjQzMaQD3afMJQ
DcuRJveMaqoNNKnS0ijefiV8dUeTDVQk0IVg5wPulGzCxgpSh0ioFAo9mW5/fVR5uJF0uC4V55sX
VHg4cq+x4qujwXcq2cfBQXClq2HFTTYYbBgn6d2tKCyR5T0kRHDzAkwvSMtRaYSC9YNjosTl1WgO
j7tMUtThQO6zM/jP5x/0yOVr1CC9AmKDTNTKwH0mZA3J/lVVjJgLuJ4kdujf3SG1/ijalSr5tQkJ
CPk8uwWI2udCe12eAsOAfOawFqdpqjzfqsHfpmpcH7KiXuquG5GQXcyZ1OVV3ymX21AsRQX1a8Vu
goGukUUPPkhrC3jst0MwDF4djOkDi/VG1CafUpzQXTI3d9LnXfGKXRIM5s2UVJ3mLrFsOk3W+BEz
kDJ0ayCJPeHo38y0sL74RFcOSabV0fcnFI3J90N1AheJ4wyOriFryxoKLRWDlQo+G4vSnPqs9jX7
0oRexB40UbAQideUohCR9u4KOiBtjOBSTT5AKsellwnV8eNKu+D9DQG9K6aSwnxt6LRBHTVL3lzV
PqxQYXBzRNiqMHDEBEfBJfj2+3bcPrCgDtMjppEtjsnYkchBhjtnkllPecGriSP9aJl73rKKqo/6
blw3/JZ4Po9G1lZVJEkJCQ/CNe2MVTiyv4PEH/3umnYnJukVmjOvzSNEIvpTlBtyudFwzdnwO3cK
clFq5doDtWtKxZgDeOkX938Rep6QWV/QfqqlBrxkTRS+/FEA5QWexQYtd06lDVx9SVsxipZYxBjb
zGSfWAR871ZxGO2zXoVYwUqg2MHvpZuDS8LRIyUng5GE7JPtPU4RA478XlksjvjycfXVBSYt1Pmr
MBcZGNTurxGCTdowR3pUbO8bWM1xEP0FxUT/gWsFIpjK9ME6kNwpW6EA+1Vjj9iqdDX8XGuH4SwQ
i2BFHYy4StyjdGyDawzilF6i2KS62rhZ/BKSJ1Z8UZnrvSK+QwfpWrw6CE7CQVJ2Jv3J3dc36e2S
d2X/f8eAZydfffa9+bole4DrDm5LHUcmiY+iVfQxzkkK+F7FzpUNWEGD7KgYgVamfLCF1vKdBv4R
ATkutxN0TtC1+P9UD/G1a+iu8MosHIrmV+Z/nd1vClHs9tki+zWkGrxwgcms3ow4FIFKLkcJwhuc
Jmy3yA+zQ18ZYbaqfi/POsnxuJ6zsCyA+4nlYxwOh2WOQGWcBZWcTCy/hpf/najMBTMDnPLHaiPx
AZ5I+2zcQSAsQdntcErULfzWm8vam9ZnG5gb5nRCtCAsSkSRCKAisTB3kklspmEmeQZkXG5kCQEi
phASStgYL+devxluJCF6lN8mDE9pix5CHMxUqisnxCqviYHMG6MXyl12zyELTDs9KO2m+yc6tLWL
N2Uqjlu7scmO8MJBdmCJHaGJbWXpYdP7rX853KRRfW3k0OQldO/zghNqrjz0Yv2+k6YNA/k/p0k1
0psL7SgRVJcp4uQguqgOxzwDP1EHLBltnC9eTkUjmEGHYWSsSbJJorJiVVSthEPj5FzmLmSgAPC/
txLjcf7N9Vo4zVTy81hCJiG3CS6Hz6naH/6vA5lxDSUeNgyFS/qwl2HVbIkIdARGuoNLY3rT8/P6
uQzgx6lGVpSbCeWq/hVkSR+lRi+J/LmhJvxSMiEKhunCGXyq97OzPC+OjJ4SfW6pZdJcuPN24LPb
BGqZr6JqrKR30TWVPgl2MuZGxvzTAq/xhNSKYxZ6J6/KAaywQxur6m6Od+JmfY31gUmhdpyxd5k7
F7ANPXvzVzXsehyB5s4VclqMzNCWlq7hAmbUjagAG7t9yNH3g1ot4jXD+7cZaXJsQDbeo5JXSREt
eebbYXmGm17m/BU3O2j2dcW9+xtr2Hvttw0K3OX4URTB9hwRllm+7GAicxrRaWrYBZQ2GDXK4Bel
G567HwzfAo0cML5w471rv76/3RvPnfZG6yCL3t4d27nZNupVXDeJzRw5C3cg9TvaFME59S/V3jH5
g4JkZyWoldKnWMTcZGK1b4tnTpSBQFtohdxB+w8zkzLHOEyw0pvKZrWKZIwT0D+ruOO1vmiKd6xm
cDveHOAA6ZTX0QkG1sFVDYPG6PXkrCLhSeW0a/adp0fZfrn9/GVjNNsZ27Sb2O/QK67cfRpLvRZ6
A7J9t/PFe5pYCUZqi9+W9zsj0eywoj+gzEjJwM5ziqsrM9/wfkD1ZBnI8Cyd1DHio/tRzHwz4/cg
d9I99D6b8Ylag9FZ5B/0a1f43bXv3brvfHZX581MOX0PWkQGz8sHERkwplZuiAWlDST7i96GkfSG
qD0K+bpcUBC1FVnETBrdrFtBk8U/pjmF58rCbGyFTUWJ/DCsO95ajGubD0YfXXX5KLz8YBdCAmEG
CnkE5oUIJRpwDcxM6cZQ6tL3PlAYpEO81HJ50S0/Wks1KQnpwOpgUthdUubnF6yZZrv3LSCQjldS
xumkENoTc2mC/1zTJmdSC+IuXzmb6NjXEQ5I2ageXcSft//8XaaaVpAKi9Ylhfd8ovJhj5ejzgxz
XhYfrK6P0r19Dq/lZP8TQppuhbP5ob41vYVF5clMcxocFwsVnNsxRh7g6J3AsjxUkW8Y3261uokF
ka79rHylbCCErQ7ZnURaCcT+JZY3ctumF+fzRl/DyvVldjs+01EY6qFa2Dl53kOAL5dHW5BLqW3C
PXR9v8dSwJj8zFiMN57wL8Y/8vcuBR0YP62kjNMNngsMfU9NgiVoPIdyaftKDaZSvbdlbGANRph+
OnPGrXfoUutnQ4dwpLN+XWWuavrezaldWaj+rmHlmhuTk2M6Nodi3csoY/H7o4Eb8p3apw/blDYv
LhWCcN7UqtyKEe4mfOt1Fbz8ya1Q+zJYtY9qDwDIrVce+/ERHW5IuqcuCzvv4VG3vXNXw1QSHWIg
2O1ws9sWyrpyZMIWWjsF/I1WLgV5vDK7CP/jyfj97cD7Jm+ruLJcOBCAdvbmUX8YMXftELedBekB
4vCNtzdTBM+Sde3s5zwFtUnOy7XslvUB01shSUDzXlix2ZTFdnkkFRZOmGspaFTOjb9ytH554CsG
Ao8gD4savFu9Oo5UluUBSJoqK5z1pJWy/cg04ppAitkyJbem0WLZndayO4rUsOebRwYqfvb0mOUq
rcm6A4B3Mrq+tyBKGdi2aUx6iWejUvh3oaaGOB6ZLE1ZoKHunBXHyRjCsmnabOQY8sLeHhJESRsS
WqidLmsaPt8fmh0ClG8mzKooq7rhVBz2mr2wGZ5+gd2nuRemoZ49D6TFDUfTf+goVmNrQcyjexHT
azY7CjigrdlRaYqhJxTckkhsPQLa69mikvufjIyvAKvMzCCE8k6wffWufODu08I45+zfInqtvIvD
1MXzVqH3zbN0ADAMjj9XaD95c1OA299lS9HDcAm32rWP1qwdGE7TYTgNleDfWr3A667amtr66VDH
RlpF0Kx82mOTFvRa/LYyDeUnlY7Xnl83Ee4wlAlQgoHdGyoPkj6npjsV5qBHIkGz6MKKqCquBr7e
aTxNlm/7SHllMPJpQQ+MF/bKuo13KUSfNE68Q5Oa4Fghbz/qAPFowc7sCcEhayYbm3dlTmhnXzOo
tjgoSkgdawuzI4WKIZgypR0WinRZV3yJQO9DlcUXZIBALAAFELiaWg1WaZvXYBQ1Bbun22iVXVCm
kqafOV+PbzPVmEVno2YVMCHbP6DReQ8s/p1idK6iB4uVdzGBUQC5vPCRRonnW6lLPnzwG2tM7CBj
XNd7fTkT5Nu/slF492tJxbSenug9pgjf7uW90t89MagKtw5+3PFA8hl4dc2hYVc00zk2+H67IFDT
mhWdY30B5GnvKNZZIfuxfU7Id+ykExDy1uMeP1G+9EhSdItN8ZjKBZEAhU5V2GAnJ8sRRn7d2fUO
ANeRSFMB3AeVkKF5SkspANJfIIQxYoWF0WcyYFUWMV4nATTGLvxliXxbPomLq+VCakvKAPBIyn/S
WPAXRFD8rgY6WwuwDSWiycfrq/PV7PaXeUngtKwFCcLN9JkOhoWh7FiZQoIO7BwNCFQEbBvKOcAT
/XLloUBIfrelZOUIvbbTt5WZGWIw/fGzjhdw94LXZxOenzlpbLvU4JANMG0l2WdkEdtHp4BN17sj
2r8IaxxHzzG0PktrLtBEdSY4DiMZGk4zf3YaoRz5MdCkl+isPU6bM93DAWqx698xoUe0g+MFZnVh
T2yDlyxLrrgPHY7w1400XAFk5Bi734Qdx19gdvxP6z4OtGsGjrwwCcavSiFM1Pv/J4SLaJIsiAnI
S2Vib1JxcD+m02vF7ZVz0TW1iTnfT1fzo/zkomOouCLzEA92Xe03iumTJgTLWvpItmru7kJfV0cY
FBLAjSZQkyrWWQ2ltY8umqyUGWsWZh3D8NebvdXoeckX8CzsIJnm/NwgOYArBadldgO9UEPoul7R
A1Fs3+2OPaYSzrHQYMIho4rwV2SMACtQ2WR3EefsqFCckxW1l2KPj2232+uFp9SJhM4ow05JCW0L
HBcMfOK4yANalGuN5KnfDouBspECpAYwdOy3QbEyG3wfH1Ph6LaLhlSIvF1XiYN51Ri9PHv9BFxM
3eMVIzM9j4g6vy4QtxEl4KqlcNP3XqEAcTCbUhYQUrTEXyho2+YHqWFf8oVam7dDqT3JDoX7eBeU
kaGGGO3hneteMva0v2AKeuo5D38jaauTdaLPRDfVLKPNe+zKFsq1yPFJj0TqM5hGFA+jSCf4qzWK
1uIxtxl0NlnNO1dRS+QA9V+hkdb5/ecIzE9xm4Nk9P2LplMQgogPwrl8ToL2wxC0wgY6l5QfVlFv
O8GzejNjdN8u1jTaioZK3IYuR4E6l/Fb96a80Pqxp2EXCQPMgqAqVOuQCr4XhayWRNPUtMH/kf4T
Fm3D/ficOklPWuPVe3BT6N2hm/yju45dL0Qoti6+Or3wPx+Cfx6WJIwhKYvkiCVnL/aJZkVbVI/V
hpifdF0HYLamxfZnBIkYd7W08TVyTJdaUAfL22snLrXU2//Hubsgf6C/k9GsfaJd3qGFjuVaaaQ1
jJ2eRb1YI3HaGqGcF1zHsd2gVJ23ZFe+zrMrowitlUmsJ+PYSJ86V6QSxk1WFqjU3P2EWHs+Qcb8
5l6/aWpOuNbxL7P3mHt9YiHUfkCkNnmi9Kw1QY1bBiAsMB4b41XgSCUhmTmVn/N16t3tNHH69Lj9
Jqj5IXpqAdJ/ncW3u17XMGNz0N9obDGy+NV2z55DbSH4zYu80Zm7F0nxzF8T4P2vZxPpMkKaCycR
Vo0pUvAoo4dYOw0StbAoXClwhymAi5KHdZF4DJgHtgsKkehm01LvnUhUqiSbmBhh4w3cqw3Mgw7H
6ZvaHaYLOzk/vUQ9/BHYUnWc+n0e2fW0iIbWEhc1szD3SLrEA5gE+GYrtpbD/+DfBCYcWxDIEdu9
DAzel3Atn3bv7fe5WpvI+NaJ0kgz8ANGzyGJAKnqwOu4poPmsvow/ixi/mmCURRpCVAA4+j9GvRV
IvdN+sL9Wgs1a9nmqLu5XosXv0tX40cR4+Z4VKb9DEabLrzic6AtuUYZn6OgNP0c8hRv96KY5RK2
SysLg3Z9E02SlMKAU6JkDFnm0PAfANc8nTsh/B74esQGxZ8PIOAMgSMnuztsnlpa3l7d0eiSUCg4
LyDexvY0+F+ZGlwSzbuEH5ETHTjLKRqS5CHXCZe0IfUvOF6UFAp2EsqawwKhU2JT3PAWMAGyEC9T
ca50HML5v5FcOG9zmV3Cx4pSlVVVEmodw6QwmRz1DUp/Uwk3o9tjx3ezDaSRtruUrqoRg4zNsisR
NfgNZgDdy7pJFSr1zNaNPuPXfSXo6006WN+e458ld8iUyPgrzSel0KYodY8CvgN6cUfGbs/jE8NL
gn68aoD9ioU/CBh5KcBuORF+8lnXkk0S8NyYl44QXhWbSwcy7HAKI2JNGwvtG36ZwdzjlWFgBuKO
FyZ6soGt+CIhyrRX8AnteK2rHGfgapujfAuzGTKY2jqOItWONteuv50ndWMxh4pTyHoeXiV8Yct/
mtj4E0cNV0K3tfzHIYmFBLn/08U00CFJe5xttwv/2ZI+zJXYWawXehugO7KdgbNG4/T0G43zOKZd
3ikbJJAKltiY/zMh6m7JJxFHpVM85Aa2ERaiMXvxZbQXbOFrckEkk5ifFXYgTmxGZA/GZhpLc73S
2Eh7BLdZCO/JeiQNtf8B/RemUjgGYgZWXuED+wzti1AAFsot/TUaeBDm+dOoAdK6U9hySY9KZtfD
mwF3B5dqslhylZNg03N92RoHNerUB64osapsC3EwAevygJZY50SbHscWEhePjMIHa8lmKn47TlRJ
I8M8KnDmAubabemtgDCxAqoaPwCFd+OVPO/88HxFX2f999SJxQzDSWnRYzynAtvxHCQH/CDdcirV
yoU9L06lCIL3D555q/KlxhcSBx7EWRE+SPJEnIFuHf5KE8hWqQ2uYdBo+pNNjjlZURkDC/eBcYHR
jHDRGDzED28wH040TuDReO7nnNuStoY+a0DtLntFDSp9oLKspmPBOxN9u6kfouwILHiyRiRRmLhy
XtZTe60sDI60NT1Xc4+B+DD4IzcK/dpc0P/wkzIJbIZYuFzgxar+DMd8/oRTmCmxl4oMXu2rqU+O
GI3dQ/1QFT08VPMbiAgDyMQnaz+v+6bG5vWnGBIl7E9kn/BZEuB8eZsNn+Uf+oc77XJQRSkq9Vhk
4fwmudgevznFIpqBptUSuRsnEmdhMld9acJFF+XBhgp/K/LJb1eG2NKiceflqoGLzFj6fqvVm8//
g+LNwY/3NuDKuD03x189GuF/6MqxohmkxbnP94QfRkhZ5LQN5OVNj+OvV5NB5YQ8GDaYGdR3jryy
E/A4Ir83SlGciZ0O0Y3XWg0wucHadU8+X10U2bmSGDyXncw1dX5v0MZNBTp5uslwME+a2CkUhLS5
LbdGWCm3T3Xpd9WqC7rzHI2TQh7W/x8RSyCWcv64CAdOA6GZ0bT1dD+4bHhyQYaQDMbwXk2vkuuO
gu1Ac5NqgAtftp9dWRY78Afu3XSLZ0lSsnVe7PboOKbx0d8TmSMJkVc6R4H52MYyziAnFDWGFOoC
QJOx4lwkWlkrI22L0pGhzMvoEV0YOyH8SS3Yj0Gbx6at+uQPqCJ+vOAdRuvyDqE5p6CmMuP6IgjD
wHoRpTasKG3KdXzEkMi/BDpbKHlxcrxbJfJkPJedAcVssOArA1JD81HwBWYes3stpxizzrJvXnPX
iCRn5Mq5QxS06AUGtZmq1mYzVB3HuTIxGNYWPa6aX9bpjrexTsKgIXMfzvbCCOULVw7LWlRkfsqY
AyWDr0RQryj43g25LoQcYkUO0ZbSLLz+6ZTtd9O+SNGjZEPhf2M3Cfw+IgnbwPUF3CY82CwK7ZwK
ouqnVD6me80H+P3Ny8EJneUTr0D/N1KJRb3JAig+Mfjn0DJ5qrZUaRSd0RNpYWjoOU6GCporBVRX
JbmIJWtq7LDHa6o1wEN1lfcR8IPvieF5WbKfDZoDvhrgbMs0e49cABZIYTwqTdBebDdveIjfTqsd
mcffG1nJeyFBdUl9tGE+NrWOHpxj1eYBWr8M+xRAQZVrhHqU54lR2mNyslEsLAxXRCexV8SNQGKE
jM4uQKBTu7qO0FAO5FDR6YHjHyDH2TWtzZg1HwcFrcJULvPeJkmx6Ssb8gWWFKV0YqAxHJbV5ah/
7ZOphDBccQPibO0vZongizJQYszzFxDszb+E+mJam3SDOBDyWhgjWXR3CUGRpx+raEvl8i86RvdC
vTQAO0baAJJyQ+sfUwwEPbpPTGr2Nuf5aqx0UICUlIUgeziAtPepA9UUIyh3Hz5SvkQC1Au6IZZo
EwtgUMLCE6BUcJMm8XIrFL3ujbqM9GfGPXNffJVoMVEU3Fpl0ezmH0j/goTUK8g9z9Q+/7JI6J0v
xfguyn1Wm9YPSFB4K0N8kFEzxZzaQkp4cla5wXD+BcVbRFCytVYXzMjfzIaL35CqaZ18MpjuhUYu
7ZCe6p5v+GublxsHdpx0skLB9KxPkYw4qQ2qNk0Xs3tEnbCx5ajSVEf3DZrJjoo8+A6MxqxSBrcU
K83lho8YgDBWhvQiMJ76OiBKujzoFMy1JBq80qWiZCzXVzGA9hniMbfobjHrhQr8GxTvLyGKva+r
bHuMr1ETNF95RuSIG4xmQf3h8x10wloIvngGjzeHD6tDnHoez7TVPJmfxRpnF7LY4tIJFNfRL/lx
oC63AEnuYtdBXeDRNCKChYVV1BdKmc9FgItjMgi1/tQMI6D+CTGNJM6Y34W7itYPSjXx4SQOtjbh
rdAe8s1PLQqAmq0tKZNyN+anOslRi009m4uEWhOoEyCft6daksYsCcZFgkgFyD5rGKgH/LFxTfOd
xyi2SwZPCPnpze3Vg9XA7QFl3Y6nUpOWWXXLeU9mdFTeZCylsxieS+hyHUnmTt+2SLSZVmrf7xV0
DMr8c7B8FHwDK8RxX0iw6IVkt+Ek+DEDMDhD/yOvYA/IbS7jJXKzLy+wu7M6V+4fqrZZ2n6sJ9A+
A8/4NOixWtKE3izAzxySYQ7+DKvRkvmYrck4TmtvkAHOCFFYSqMoNXTA2Kjr8TamZnD6bNW+8P6L
vtRP9SqZejkyqEjw2UFXPLV/OXS+ju4scAhFqRx4iKtUgSZD+Dd8QXIfSt4bufpvphvJw/k41+sc
Lu7lLwUBH6TOFGDFhpOr+nPxZc66y8W+RM87C6RtDeX0sEPvZnEsEGRv41tBL32SaW15cJFx73XF
XeroOW/l06lEMaybm7eM4DOEhHmEyNOQh/qY3Y2DiVI4IYcMFV2/Up89OFMquhrmMbcPiWEThgJc
7ZlfBer8lYiMObZZYYMXdEW+BSPbZX+6QDVHAaIhF0ZgO6Svt9gaJvI07KxIPHtTyjxc1tevBdQd
uWC8PRIKPePMFzVbjLjZVnXnApr+FdftzldEUADfo27K4BsGbqbKz7/f/3os9AX8YnZXNnBpcygq
KzEZnDmWiw0pMqIMrfnVM2lVWo2G3NkAyGciDRwB9AcmlsoAkJT9dBkwMJfa3MPHGtYr/rBHdsBo
Y0BUC5HZCVy6/c+wUXjypWq2PJVLB1AKvKEIaqWw0zWlVBS56quYDoHq6jV6ZIw7mMq1j3eJOfwM
+qDjd+2mPHWa7UJKlNDwUWIn68W8ysWojdeQAGRDFvOz33ca4TXA7d2rp4T+Kf1jPdGMu4GE3qZ3
Z93xQeyYMvdB72aaVE+dV7UceNm/AQn/V1znHCPONIL6TJYd/GLJlMWxoZWegTJSmIGab4zL6Gl/
+d1knsuY7giFeF/gguo/jIUOHU/9shDkZiHyyEuh1reVJURpRbAPivEg8h+LGVfUB4/G/RHIm7kQ
vLd7OmxlclvuBsQQA/NNB6t2Ai47chq/wU4NirG9B2tOzEd/Z6hd7JqR8W2J3EX+X8lInvpa5hh6
FAD92xbu/BQWKWL4aW714C4tOu6vK1c6CIVE0pCnFPuOkKPDZl4sDz0/tutZzW7nyaKFYGTT/UIM
9C4t/1dnhs85KPOqwC9Mm8Vw3fp/zpmv/Jpne4fGDw5kz6y7OkhLrZUfOwKTFcJTfAi4MMEmll0d
5j53+bq+y8BhHAgbTEm5J2hT/R3ingaExo8V0vWATEgzOnE6JzqqNnRykrcPmNpw3G9+ZP7rjPng
1/Bhzei8sJZh9tL0dCinX42/iR+A5kz6kxbeBae5Tavqw2pL2w57gd4ZDx9/pcgW57fl+IuVP+BY
3x5E0gev+FPQ8CCvJZrMVKtgCgj+w9h+R5Vspy/PwO+9cb5C47xKI4D5+bG3R7K91ybnxpiVhVKK
KDEWXPdoqSAeYvl1+J7wpUTNppnKClf17LhyCNFPIr7uFvgJ9i1oedGeMwJEm2+jC9NH1QbR7yDd
5qy4zjlyRL88jsiJBHonrNq6nrJh0FVBnWucWBxskR1ca5+uLH6PzedAbePzc0QPBHwWIuyoqulF
qcsd7smhi47YFWEGm7M107Q5xF6zyMr6gsvB3n5JZW3nVtl3T4vqQK5ayc6lLHr4TL1y+jHpk16s
RXr0oBBpjy+LsauKAvQav9kO6TDul4up++tPfze4dOOsSqXKVxCvxq4W71aXV7XvtPUrPk6JjeUc
YmnJsgyKa7I9RHJ/q3+iOzztg0gp1O7T5nEt20o/N5O8VVFmCttpXxl3K4XWLSKEzj9wHMJsAvD6
tgUOtae83k6M/P8tG16TWFnyaWCPOx0Zm/rXHeG7+oa7wJhDAOIUR8zL61erF2gwrg8Whnls0NX9
dvnm2uH6wQq6jlBB0gdhw1qfg+zL1yLYf4Uo5qm2RUi5xRciAB2x+2GjvjyBLkUxkCavy0EHO7oG
W0Fg0fDX61RXAulNx/rwJ0Z1n1lNN8qQyzl9bTbwsLfn+f7IbvhUphhy73WAzjCrQ0SqbJzuh70f
8ehJjS6bEZFDTAphZbf4hpCyIfSoSRmyQ4/J8711UKL3n9xY0W3CC09SK1jutMKqK7GaqlH6zEg4
wQhTumjTmY1SoKwvRmma8ZYgfhAs6QddbwGFPOT/AX84XpOMdT8jGHVNqEHCHmA2WQVj4yxWwZnj
+HlpyWFshIQdufpu+B1hXvaZ2AOXLaDZmdhrxvyoD8eyn9BhOY7QZUE5/Cif4lQfzLJbnvCKqIur
PC8CPal/NL2MOibvRBmeTQZK1K4W8j+ypNAbZOsBUgMixWVNq/hX8/LBlCB/5gBc54FiJOzrDX8r
bqoLzapCKL+TMHrg6mgHYOwLJwpYr3wB4C7rafPHO1y1/pYgH5h/JnzeVFxfL7aMYmYGUH2HagZ7
h3PEeUTW2m//vJcZMAIKQ2uez2q2EKQm03zoe9uJKvPDKfJtlhydmwK0B5UCNP/d7IR3DO1cKgEc
1GB+xkNtGBlbKnka0tsU84OrMlBR059eBl2ys3RXkTMPD6h1uXXDrUQ9KvTaBIy4kRDeLKgSdc6H
61OFkd3W0BS8aLNHd2aFQ8bq2UdOpE2CB5PXGFqf5E8KPPUqwmpL7A9LGGSGAlUc+IWNP7dzU8cT
RutTgjGUl75StaAiLt18WelcnQOWNAHH0BLjpUqJ0vGZQw/fGm8CmECEsbSaaSbM93/mI2w78Lgo
oimgdVLe6uCt/hoExvkn9zKhMB87c/aw1cqFnwpn4IG9H7fgvDYBNf1lnfPdc8IeBmy87FTQXO8k
72n4GeANy/fN3WkcX01oCyJWDO0WhQrG4GVHzGvTcB6PVMJIN3sryRgnGjFIYMK6JUwHlUQC/wVk
l+UaMJxXTHT09qlzPjZl35A9GaoYK7vuw6zCpJUqJZvPppUynF1djCZIHiMjPf1JzuTNKimPE2ta
YWs7vHsMrnmMie/YxhyJu+1rcfTmJACrS0H+pXZzxbbDH8+SdAOtEuSF0AxJlASTs6KkGM8WpDMX
yftMtPRY71GA45+d/TpX3qJPXebI7+VO9CH1GAQemlbJRPo+uY2+F1NffhdXqIWQeMc8/SnCFl9P
T643aQ0sYQAcw+jmj8LRjV2rIYB0TrNOaq3LNJsrsVkclEUGJk5LBswkSI9q8J4SmeIeLGpo9v63
CHQ++VjMVCGyg20z7WU8y81goAgdhDEUGh0fDLh8C2WoTBeJwLeTK2qWRM5wvXbwpBQI2+BEtqfN
y84u7Sn28O+iqIlyfirN8LrHMdm2esw7mcHCf7QpmIx+CkFRB2X6pSl6FDJR/PCc2CUdVTs5F94H
YjWUvKBuUky6d15FvjQoErgsasYhinj72jwfF/NNmZmBRnRyFhncJS0PUHbEDxbTAYDEsWT2G6S1
T5ZBpU+kjzlYEivZI7C27UkAl6dLPVXUrKqiOP3KHHLxp60SZOYH0UZWTChyIeJrbzJPncuAaLZ0
BAEUWpT1RPnhcvCtV9m0N8nOyNVvmAnmi4w1b+T+4zrVI4gpxlkw+w2HmdpxZkkNwbdE/6OkAf6p
RpPeFxdDW8xQbJnv+GBCnCEDex6PD+2BCsLvqz2H3K+RHuJNE+txPjVsm2nU2DvmXxzNP4RGcx9+
qJKHb7zj3npD/XweGnx8z2rS6p7il3GBf5baR1tI/iX2XngQmC9uDCtvHsVJmgMoaN0SInqQlvAm
FlMryeZtxLtu/1AaSVJTewuzBhudBkH/FXqSEWpV+XGQBk1FgtiK5VHKXsLYGGdx15SToHzUQrPf
sFPnTw2dldpRvrw7SGFBC6W4Pb3i0F9OL5UsRmvJxh8iE+tJMze2fLCjielsc5LHfcY6oWZ7w545
sBtWTB7nVmra2j/Kpomi7LRzBPGDZTNwiK7PKSoaxYzCnHsa1xP0KryMhJ+0Qxe8zseNvlXM71Jy
NFJVwy5LWhJfjTXmnFLe8jLCrRQqj3grdfX6M5JQlzx6cSTJednnZygDJDLsph4an7GfwF9suTtM
JnYSHuK7jZD0Ol3TZ/Ev4n7lK/DuPsxwD3D6oPr7LwzknY3tnFp0UdwOXj6Atixjz2fnyu7Td5AI
lI0aOtc6j8F99nrhxlKtTCpogDVVjOp+pNd2vHc/S8gU5BHHBE6jF02nmKXt0ZcIqNc0gatRqfXs
hf7/9a4/56JFqlTekomWCIDXS+qyg7iguBmRmXD1Sd6Az6gwCrdddSWnNrQbgIHCPgafCYwBr7tN
z3YF5wykTHAD7Ih0uO9KHH/51PfRQ2His9rfCuY1B/Stj5NrjccCLtToofM+3mgNzNXhOKZqzRit
Mh8nJwveftoScGNQAaloYfHHfg3TUJ1Epu6ghysZYQ4mKqGoE5kYAVbHnl7n7+x/LDDRjPEtzRxX
BbME90Y9sMJxF6CInfZivaC0YYQ/sp86Yruwo0MKzrVI+SxwYiuzSsANp6Yn9wrvkrHhL1UUGu+4
reLN2i55Gtxr7LQ8iZXPQm7FP6IAVkxqslLDAUx+OaGeHwgTRInEulgezT94FVNDS68VIT43Dmla
vMZ8E4CtIZ/wWJwJWaxDSemEVQMGOX/rMNMQcYRMZxHWlVZBPIp+6BLxOPBYNU8yElZKf/Jpb2C/
QFpSnWzupfc/YSrTSnyVzTduzu0NVV1rL0E80+nvLVHXVmSVtmHI3tqXkQlqipjHBQhZQyRnvXu+
PuxbSH1fB7jk/8TF1BAoTrREfsLUC+KMLGB+2Yemi3QheBj8m8rE7yGAZjcTzxAzrPeRJTcvRCBs
Jyk1+1Xd1sw5mmPu9ZfifMvpIgM0798LilqU0n6+ge39kr5dSK7qNgY+gknMMze4tUIjvSVnMnmF
t/q4+/WFAG4YJ0D2dmr6B/5WxWSfqye5Dn8l2+S1iWW1UIZzXp5dtXzbeUn8bWjGyfwbiJfJzEwD
4sw0tc/eO3VNyYfwIoJZR8Y4w/nwYVdIG/0/fhcOFzRUYDG0TvgrnN48GeO3TM4ecnMlOMgjNSI8
BVmsrhuxe9eeC6FmE+kNQnZqf6YnhbejiHk4JC344v/H16zC0q9las7o3HATeGRN2/Ze0kVjMSkx
2OLeJ2p2Ajz3kpYLPAz+B2hAtY10dwGpo79ik/z7xxEkW7kaWD/nO4AlhUdjNe/l1PYHTWI7ak2J
pgMvvns6szuM6eV7lWh+NakbCFrlh06NRqisD2mR3d2GtHn67Y4bXrFlJ144f/6/koyaoi3X90K+
6mcPyTRCSiKd21TraB0JkEpu13BlUZrrkal09xkrZeOM5l3z4f62x9enZGJjYy22rRNwOqlc7nrs
cVipnD4r9DcuEsFOBAooaNJS0ThHSqklxpWKPegjEjjoAcAcT2CycOetkjTYfPKH08tcuR45zskh
kS0wpEcFflwGwwYiPXHcPeYR3vMX6jlvDr0lBHzEVd32MTp2HFlIUvbPX43YnvTIXpQL34yy8Mq1
iiDK4ix8zF9QURcHOeSufxqOU3tXnw8FigjCq5Q4JGqM1ElfI+Mr6bkzp5iqzcfpVNDjVqUDXFui
POXmLLfsc5VNhnWpsoT66xt8k2uK9/lXL8UyR9RZkp1pEF1qIpMF2VBFztgIqyd10nmVG5cqKDZd
wCI9VLeE9XJ1T0dB+x8lfeWPq371HEJNEPUws0acB/k0vyPTAQ3hZqLuFYFxbSoKjED53q/Tw86V
rcs86nTBH14UZ+wey8CurXsbuHfEGh7aH/+F9Q3Me7leoRFMU+e7247VUy49vah48NLNkQIcxtIq
iS5ZpM54Czr4q4CbQOAWPUawM66JDSJ4z6szuner/a6TmWE6wffSrlo9g4gg/9rkT5C25NVgrZZP
4t6i0NcfIJ1YwunP0dV6cioWSG4Y3jcixd+KFgZFaRAF0XwZ3+L7sNoqNVKbjAWkQGDFHS8QvpnT
SaQlHIXHBQwbZ/24GawgpozbMtYNqP5fbyMFIygb7rqzhYklNTwt0HVwxYnDlYR9/HKpi7VsJQ5V
2J7REr2lwg6CZ9OeeKeITzXwXLqT2M0txMY2U3TMS37k2ciNt6mBFTam8PaGFXTEFs+YZWQnIWsv
0VHruFNkTNEtbaWYqlZBl9jOIlQUK+N+/PGxLyK71rWQvJoc3LaC5BkSOuhwxFXCWAXorRMYkYE1
z16wElu/TuZrmE94k0wvmnFQEBYzhPte787E6p6U1fw8U+eKaJhiFMQXJI6Lo8xMxiEkTvCphUBA
WGJX9/4QR8waXuQhgqNMO0qFwcxnat2AyyGOAKWWSW7/9IUHfwkwZlfIp/H70RIulNMU6NzNge38
qrn2zEuUIJk1pgDaCmBl5vY7xofbGbUnPXK1TSutmGzVS/ucqWXCaNNkWMCC2dE2cpK+HxXhIwET
lHsPLqiFWA9f5al1712g3Tt3IKQUMHd3SpFlgHkwD6BdGDC9Ri1Dhq20G0puQYzTtNgsk67OOVGk
fN1mHh70ffKbcAJkJUKNGIhLO0ev0NENjeCO+Ek2xLSSnz89osB6A+yQJtoPWxZeSsQU3VRnodBa
QRqQP7UbOoIS+0upSzvlzx/Y8s1Y6wSqlsVSeCFKHTH9hGqyjMBe+4n2rB+KBlvp3WHz78leyBm8
Pm1xU3jHo+yo1Be4ilUVa5I7GFnUAncKg1Kc06x3+1T8etS3KirsyVg1qZ4pfYzuFweRy3o44ZbW
1ebQerUe1evUY8cRJyj2zY3/yzHqdkE6x3lbzpe5X0OkBwcje0Qj387qI1FVz3h2si3JNYZvtEuy
wY0Jck5ITy/IExeJWDmHDyiXKBtYvb2S1xAaUGIOm5ujSUcB75soUbApDOIfUqrrxJ5HRFyLcEjY
ouMPX/kMrjvdpykIXHHccmb6sB1LSQ9VOQs5QiixVMKLXiLPA9XS1+sT5EUOQSlRSPklgbR1XNrn
jji+SlpYI9pFnBFyYDkBDmNzB7Dx/FvlPVu/oXlGjuvYpkO22f55S3zHyiOwGL6WdxPGnvGuHXGn
nlEDf1RVXC6rqXz3EtRLfZ2BENlQubRquSkfB8wNfYGp98LRxhNPQ23BDz0a8f/2jeWzhR2btJ16
ps/o5HGHePxD4h98AtqN8NBZudTltt1k2NzvRw6c5ann57YUZrzJOlFzXZOtc+5PPTqqcVaWZDI/
+KQYHMYTAl1Uns0fzQYI1Aonju1R1v6EM3N6nPPljG3EGwKO7RyMl7+tAMTjlusx+sXJbFnfRn3Q
OhbsWt1U4rtERol6rXFlrvA87dOaaTLWUSCiaBKI1sy+aLojYpBt+KYxRMv5dvFm7GcERf5h+yM3
UcNuZ8hS+ccOTH6W0Hy7Y0oA0Wq3wUxbFWa3j9aBa6FYeVOSIDRNj12Un9EuaYAyMLnZAmorW5n/
SlEknvzbKAnz0o33muezXtn7vNC2Tw7lFDe7LUVg8MMT5aeeWXw3vH7Rl/i1IZWNiHLoiKkNWWob
WGkSVInn/Tl4ScRdCrHcqfib3e3U+7HfMbJltBctkYwARqJPjoDmAYZ2iDK0h3UjftCzK3XNGlXp
T3JOBmgymptux8ZhQhyY4ytBDwOQATNAyo0wmIJc2Ga/Eip7tc27TujFgkBCoHTyB2wKlgtrUtLw
JON4aiR5pCh4Y0RvgcSgOAHeUMKAjswlMAYD6HYiXBptf6FWvPXW2q/d0ZsCwl8whZ8G0YdKqM31
YUuuLcNLyRsqch4LEMwn48e1IEtLS9rSCb3sC2vLQuEx41vjkzcLrtxKBkBW2lp1pSoyeyn7d8p5
EhI2KcywZrevR71Un7S8wTBn2g4eln0dexMgcMDVFkQLjNUku5H2XCbuFImIoMpfF10Hpq/dDGYm
ntugA8wHNlZYab9itzGDbfdwZRnJ0gzoprZXa17TWcTx3Al7Dpk654ZhpBwwvVSFxuwLTcFqHvv0
w+hMrWzS24IaQT3py9H7qTMskucMEcvdeppT+7ImfH0FUJ74EvYwi0f3DiTQHapGVJwYUTizfdH8
yerrZpU/cBIAWnhFPmNZjm0a8FGIAYI42wiVkeNFQsgNfw1T8cUS+Qvq9dKm4Xeh07riO13lDcXP
pv20ksTX8gjO2xAFFZGzZHIch6o14KuS+TPk0E/eLV1nzJn1uX+GrYALIXwhWArKp3tChAX9jRSf
F3gq5CTwvNcl+frsTPfBjVvKmzT99FcEi0rcNGrRHkl8IziEOCVVgJi2XrZS3mMAfmbAFv2fBCFq
KEBbiP4NLHPxgs30+lrGzxLcgZpukadIGaMCsX7avbxrnY/beSZ05rx52akTW7ZtKLZXma0bfBt0
IDz66fk5m5aTlWvu5kot0xI3QwE3rht/K4t1mNoSaHXo4eRGMiN2Z8VpkuQQzMrr/F2LAItKxWeP
K3ZoYa6AnZFeCpKh//7nvXdJ0mq4qNRQcbwMaxB79jtbFdZ+V9uhxvEo6yNxrnGyswD6zvXbkChC
gy8xCiz43quuLrfEf/y1CgLMMyX7rSWOWwOmD3PelV+dxZmfor62orYzeFhP8IDlwAZl0wyG5T99
1ScE/g/7ChPH9/9rCzpFlq3d8EceWu2SGK+Txh5DWbe6x9nl9SEyrYBqRi+vTNfrTzjaSEOFyBL/
MjPA1k8FGgipJz5FGA6j6Ptv9Ycv74jGnTCyQhIQuFahnmbBO8aZlsLYlkEo0pA8z5yhUN24lVvE
8ZSwn7YEL4VvfYKHxQUDja9rQ4wBV9vSKllw2v86pYNJWARw6vTCQuUps0/DD0W/GJffn2pjke5R
/WQ4v9kd/PMcVl32ZKNYhG/y9FoeYRbZI7618tN4sU34mAn9LOThz8Aw/4qaTojuuVxl1HTnkDFg
chtJ40W40NjItp4+F/Rvi4yV+V+s2F4dZl/4IWQpBj5eM0ucnov3/x6uv2Cbd7rWtVl1w5Siq2pW
fzOyyDbcItDqyt2fmJslOJJVnniZeMii6beWck4Rbm5PPvq6/tOdkATpqvBW3ZRoICj/2nFFtD+l
fX73yLF1haFP9LzQWTtGxL9YEuz8gL/9j6XcX8MmIPyudF4HVXYqdSmD/HcOVU9OLGLCyk2eKzf3
42HlfbgLdUXhLtHPXYMAmZC3C4hoovmq0deWlXYKpgJ1QcwTlJ9Sj4PQxX1L0I0BC9ksQlZqjHFY
5JAsOVJf8+911sw/4ZrHNcpcHmG3tLfgPAKFu2zLPf8yFGSoT/Zpl9Fke0dpnSNib/aTkcl4DFL9
Fn/Hu53MQMLF/sJAeZfXWFm4oxGgUSANOuh0ptUASRmLl+V/OJTFQJxE9pISqZEcGN4PQkqBiJNV
6SeA1TB8sd9tFyhH6j0mWP2fAOf8Xvd4Uw58Ntx/mRfws5dbfyjRUw3nPwZ9w8O8WKIebCwFSnH/
IuclEA9saVAb7FMxxTl1+KFSyB30RqwoMwAbaqKTw16iR1emgCNwAmCF3nudF+rZPnKLWUkzIvWh
gVkWdJzTOTqsIl8fY0TRJmDApj03YWsEbRmR1ruiKycWoJjgooAbglQj6tfBWXdCqy2NszdTnPjg
kJnjJU4dXh6j//bIOzN9SArm+RPGP0u4eekMZy9fCOnmHdSAaW36de1BMw7RUijmb4ZZAyUb8v2g
rZNZPzlIg4m7yYDUjLfnul+tZnmyT/ZDBDPdv81QhFCaow5ajXa4anOvHJBw5Q20JtOZeAj4cpkw
9Pad2iWte1LjyL4AUOFXDIWDJrNIu6kA/M4SPtIB2u6pDbHCalUMyMpTGjs4SlRydiobDyIaLOuO
M281ok7kGvweOxVfg3hMeGfcagsDa99OdvF0ku+nXXb+Ii0BuyhdAVL3lkZmrYGQVO2qEPxsjptQ
Vno5KBWcwF08kJg708i9Ghpf6iAdY6clE3zmGvuDLuw766KzCn33m4Cu2WiANNBwbpTkZtt2d943
g9asT+caIoAgCs5tnW4NN42uh8mBaC46vFSyiXqmHA4ITjy3sEbFPc4+DicPqqxHPO3GBIe9LdWq
6DdvxjzMpHWbNTfpmLAO5BlRwvnfkqBCS25WZhvqQw7Kxf0MsV5syoi3Vwxd/P8rXocuBtqxPAH4
9NlAPnGCYXFW6oOvD0ffYZFt3pHXYjEY20sHZUOPsytyG45KGGQdrXhhlr9prM3Y8hhXLDCwyWHJ
FUBiIA1tVfqboSMELn1Z2cgvao1Z5iN5x66dJe2/YLy2QaotE0/9dxG7bzlb1Xsq3uoHdus5TTRU
3/ftzaiezwokEXkuAGDzeVh2PoGkYLtzVO4dwOh+DO5yIaXFAKjz0QGZE36vfIxAuGewGBgpKUCm
eKu9M45OBGRkcu9LIp0QkIMe8SZdH/1rd7m8ScWq+DeRLU1aKkgQLMGDbGrroZ1OidxlCmXrQ8OH
TNrjGifR0jS98zwb3W9qZ8FviMvC2V+Bnoip6OCrDyJiIA3LxUYTEZGvJ0ruiF0+j1gILY2QFq/V
lR6ks601GRZgEG5OkZ5K7Mu5QcG/7y4Td8BdSPJTLMwMn5W0qG8ty/oxYosovPme2tiSZsqRYg0h
AW8VBsHaFn4J0uhBvME1K0Aa/0Vf8DbfVu/PwwtL1dAwNIUOP+m11cZLxMlB43ewhbAfZiBGTTpz
9U+xY6ejvux3GvsGJIwuxya36tm1BZpOHdU7FO0lzAkOOHwcRZpMHDlyqS3xj4ISET9/4zGe8yRh
GJ6LsO0+R4IxcuCYZz8OQw6wAQEM/cUN4DeatAgDJZBFoJbrr1N1YS3fgg+N2i7PnWjt+mJtgtGH
uczRDBNuR0U98R9avvtpVUGHekyiXzLND/a6zg/Ha3IqN64MDZIsykGOX1jVY+apnhSiCEz4zCcu
9UPtuep4AESyjGn5aDMB53X3KprsPYwNeI6N/EhOn08muUa00UD7Qc9nSn8BN/lTKoZYSzUXA94+
f3jALlfMueF9WXnNggBxfwTznS+jkA5vXCG6uKxTdlHyCmq2Pd8m7EA5ZOf205IcgMi3mL65kiYJ
QUoEnLN7GoVGtomPKg25AQEFYczcDZRcjXnwUswfvXaYLdgD4leg0ewuCIGYez3OG7KxY3P/zEKi
BAsbBTO/YMSlg/5feS1V8OhBAW+Bbm3seY23pcOkK9cooWfHQMuqB6Jn6PEFzKzoc19OBdNBZifO
mfMJysOHF/TrziQXGywc2Ja1HRoDn5922TkucJ9HALf/qPCeViP5zw9kQ2MvdS+6MRdXQgWtLe0F
hKVMEO9o42oEAYNaUtGsF8Cyx+qLq+lNY1UBwwldoJieHU2jJBrxc+g/3De6+gSc3sPFalBH1Pne
l2zPAkLc242eKUhoXEjMiYTmf6BlP59dAClnGA8h6VbSKX4pxt6iKb1jsDDjPcxkyxiE3Kd5sJNi
c09+IauX5JQa4J9frLGO9x45t2xC9i7wRNLB/rrX5bVi0FBe/jQUNpQjW4KDBnkSObzgTWnEbSa4
2h8IlIwTat98hf58ngpEYrn4clo4g9YNi1v0Da39mm7lL1vY9YQlx8ILW1m5L4HnCTaxJoHBuYs8
+fIj/7RA0zV9lP52ECFv8ABRWZQalZFpIujUc+2QwIeEEy/G+US7VPbMGOlPtykfGJxbT6XU5u8r
8nXUq1DnipUinpXcKSZZ9gustWiYl2ulIu9l7HFDf+I4Rkyd3/A/0uo/odjmcpjoyul2KI1WSB4e
0D6cmvH+ZKdbXN3mprEJedllVgckMvmY/yxQkYzBmf3EAMYyaQwFHVfi5PGjvYBnQpbXbKFRWsFi
GxFXxfjEDVSgt5C3fnp2Zva70oqSXlrtLaVxufm3rZpOOvP9o5D1Wqw6p+21Gec12J/SAx+4IiRF
ps5Q7SSJ/oeTTpx4hQOWlGI1fy2u1eqnFQ9WWChFDj1OFKEeo2fYywPYyP92ZpMFJtd0YxIIJLq9
trwqRsE0n7hFA+3zBEUHzd0lKZoT/y43nCM/DaQfAZiDbQfpZq15upx6D1fVCMoqwnB79xIk5Oma
6chHCXaDTRrvgVHQxpNAhB9IUicJmDZJjGvR8uFNHNkWA/WyStdM2/adUt5JmGjBry7eC/3kKaYr
NPrn2gAuj9/EY6a/AR5nioUqszUuCKvGxny5ZqRtXqDG8ucpFNpGZpFjOiqlfuhRLPv6p8TD/QcL
m/g97H0fAn52XtZOAjJSYygQY6z29mop+EYbWa442fa8tSSdMP3wi7DFlmqjKJsnaYxjjHREhq0b
daF4xMggvyKRe0WzYWw+CUaKKzQsiLYM0JyE5Tp8mq91KAhahLKU9adBWxt932z43KG4CBqSHayw
W+k6p4IodjLks72S51ICEwETCjP2IcBUYWCwJ9L2ThWMGpa6Sy+O8Eocj8iYpUXlmCkcZOB3SV/A
X0mpyj955zWgCwVQIUKzlPXZYtJkXIv0EBTD+mW9JkGBR+eqhhF1SgqkvGmedHOoXPoPwhHYnWll
hVAk+MRfUxx0wJmNGIayzRrFtqV79aGEfkFteBjRKM9wJol50yRg7H3wNaPfaTvCqpoXqO2i3vgZ
EvoZu4mS61uTMI8nUJU5w0YBAt08tzcG1yWQS+awMTfGbQ+oPX4CBBdHLzFsGsh/NE8W/7e3AE5v
idDyXveO5RE6q4Q5OF3v9hlp/kIA2Qw7r+VNp7Jcz8BQQ+H0BqW+BUDhg1J42ZEhxNpLszIzgI6U
GnPcaEfHjWgOb66Gwsvx02dd/zD4w5R2h+8TLzL1vQZVkRO4DAElPL7kPdszYKVxCnV4YKAUA5OP
Fz/TuiVySbE9Ww3XXR7GidDEAjMG/mChc5JEq54s7I7HuV9qMQonsXup3IOSxOrm1/K9GXeCVoen
pLOoqYhTionl+gZUpemT8ggpZXMzTiJblg9p0uNWMUlnQrXHzIipZxh5wrdw+azax0MBX33sYvTx
XztX7JZwylx0pD+4Wg2FcRhqL04hH1AqQACw5a6KhmONoSLLTXYHRyr8JLixxe41ECVT1wBPe2Zk
CL4Nc8Eb0Z7vtPXFNPa/7U1beoPY3orWOu+E+ngF+i0GW9m95VgDOMXjQvee8XEyg+BsgtRk98RH
LPWh+0QkeXWY0W+og360+3sbmDBtxA+2ROdjF1PosXrW5cIzhjT0zlW5E4DGlioeRAHjsLGIpMKj
Lf4NJzr3tco+VtQa6Fkdy+6WpkKGDi0Cg1T4tYTZhCNBRwxSSJe0RVNKW8jZm3X3zlmKaDVrxZDt
Pfwmp7xVdUwOQ5+3HcU4jIGmGE+HS9yzyAnRQCuCgOLsQ80dF96cOZyKfcvuDuyZcQsX2mT3hxRM
fw3JgGrjke5ysu1c3M+XEmj8jjRbAg+PYFhLustrsHy8fuEgWAWcXko3dvNP//LPyPVtaMq/QTG4
CjQ1WT4SaBq1feKhMD6eYxdYZpYDXyc+rVJy8GLOwTsz1vAszcjxY7fd6EhuU8aIb96tufJl7Tj6
2OPNMPBXn+puGOOshTc0m6BXDNJmR7Acs7O3u9zmuePcCaZF/V7Fhdgaik4QT8KY0GnL/qdYnr0h
29WCKJANcV2g6iB/NWWcRScD/fGwYP0Egjcvb/06vIvEuPBvbpGRs0YPZ0RoslPNebXG0jcymYeI
LvbKAvh7Alxi5TtifckcgdL6uA5+G4ISDN0DmtgDC9GOSYi/cC4mPAtWezlHWau0S12UDoqdq1AB
bPp6wsCf6sHYFfm45F5XVOv6G80AhluZWTk/9GQIlQoP0XsrJqZZwGxDml69xNXJtXi3ZS8Pd81P
2erUHngmSNHKR+p1Hjx21qlM5jiIe0irnONozMEq9GsFiAzal0+j5vc85v+P+sHrwEOpYBabJec5
APXThiO+gPIWPqMGqSTH9a0Y89t9swEmks1orskxlIxceKjy0cZUPGgZgUsoBEVHSzYqos69+15Y
rtThlQZAZmPPahhPm2ecv3u5+K1KX9bZIec7ceUbuS/GwJuqQVga1BnOVlPVweIzR+6AdtCP7aMk
Chdw/x7asaX8GPoOLrL8AZ+gFH96QTRnyEqrgFzkZ8yTxjLnr2I1axjP3P5kwdTzAlp57Ld4UP/N
U9W+emuFbs9rI6G9HgWtNPy9hWN4LKKDfENlv0+25h2woymmvXgG+HxkyPk2HRGpuqDbsco2DYAy
bRvjVG/XK7IAswqYR2xYUA8mUzgssJBg6KPuPByyUxtz2FMtkfWP6DtqgwjmTIUsR+TsW9gnMfn+
CmoITsb/q7FtSucPNNhsONZBXWUzr9QaQXV/1o/n+QNGyosqbOczJnygUmVUIUPQEaxHUXI3I2xe
4MK0h8Y2puBcqbq/AH9xEqjcMqSKbHerlPQXkhzFSJY99xJGRw0U3HnRZdxXtXAM7SjtUpevwgMv
rQI1BkMkzUQ1YxRZgkTznyk5pC4hoxzxIa2bjReTB0t+0/kvMtX3szcjpM5i653cVCoGIP3ipVqt
FPVhTaeeHa55W33oRZ6tGFo+4HwTc4TK3RhfPJrGx60ZkfMK65CBZpttJ9RW3WmPQr5zrOqryytW
4LDgSdJxAcVnfFcBgT7skIRqco6gKsQAe1cZsL0+hWXI74xdL0bpoSIS3NAVrE650E5fgH/gjd3Y
HetySio4QRZq45dwgdf0YGcurr6W2buJZEI1MXydlLZrzjom+O41kQSHU9E+k+3MbqycaykzCIGh
ju5K/pBtg8jp7ELFrIahwNnIZz1PV05pXnBfXHBUUneEBpbkO0Nn1FIndkuxpMCV3fSD7f4stXbs
J6apJSiVAU9yFsQ3+VHXbAdFKOjgLu2cEKS6PA6N+ks48p4g9d3B75H4kfaGcAZdn2kFDFZTDKac
m/+3w8Mo0t+7GNOF4PGUuu9eIz9/QoooTtNfb8R1H3quFjSpJH21fNqdxRHqvjbnpyI32Rec24NI
a6n5njPFbmDdYT4zvVh2HDv/uNMwKpW0HJrPkO1lwwwGsE6ymEGsc8Kpk6Fg0IHuDCoervCMIwA5
ifxUm406VFujHzP+FFWOWLC16yU6onyab60bCBx3Igmh4T9ccgd7GL5KNgqxvh5R/0OucwK6a1Z7
ow3GAuaBQrhWS61V2noWdnOE+/7awr93Rw7+NkpgRSPGzdFyE6FCjYtuz/QoXyJ9Ge7s+kDkllEJ
yBMkqktKFUxVbJdsvHDi3TgIGNciH7iz++5SJK1f5OaeHnT1ksdRgFaUph6k0jiMJJCkXF4HQCFd
9+5hm/bFRlpfKZ8Jnu2GVdUDUr0t6NweaaENm/knd3rgJWbl77cfkjzAXXcFDryvqnEfJSqcLuz7
yBMq22lzJMgRHWZpSnGH72NJk7uKQ5Bf8UK/KMaFky/m10cXpX+Vz72x2I4svgkvW/UB0XTSDa6M
Fdo8jz76zO/fJ5rwnJP4o1sw41K0WbnFf//w5kISueaxRYmwX4+9pggySwZlA53ZMVfsyWMhfkJE
qMaeBBqOtzRbkDcii34ELHABBBgCtxNzjPXU55RoUHhSWfr7/dIzYSOcYDdHPljkYhUrpuhr7W3m
+DXkL289Rsv6TX33N9alQlpgpSFwHhabp9LfKoM0+YV7bqKCuyf/OHHz6m8kFlNWTRMOHKxX2UGh
k4k3LgF5djTzvH/ZNxl36MdboC9dalafdCGezerfKdG8NGSBWxd/KR7gCgyryxIw1s2d0zkbhBYS
Ixn/b00S5CqKEJQ3vzRILqVG9QE/Fq7oWOhKP3UMSj2RfjAqtitHIauchBk+RsUePRIi+nT2lELA
wAoRbPa/CQfTHBSFfYIwvJ1QweNeh1Xpuww49a/0Wfl/Tr7Ndc3KOSramPBP8URI5sBsmgttTC7O
aYSOcBurdLJcLnqtqISr8Jsy8YPK4eAVN77GwMAB65N3B3DCIobBe+HUkFYmdztevT85bWGKNCsN
G9Sr/inTIIhxyLEjeLUPYbzKBo9czWPHNoYEKna5zofuI7LRZzyQt/KoIJWhF5E0h2JhQ53F2L0B
RHaC4ccNBN72PZQZtVKT9vlVsQZ0/MvAedL6i3e2tvSPMfkLqbcwRJP4QTB9dKeUjYwfbVaVB6ZJ
ot6+TY3SDsKWPXcoPUL3lfTEqu0YKUza/8ZUxbQOnpDyTkrZApMi0O4McC/XGpd1b8ZPTFuE0etN
zXgjFzjQhRGEj3D/tQYeB7v/pByj1w61223RHBMAPB2NBYmdSZOjRSsZ1Z/Um6bmVL6XgbPeLBFD
Wn8iJwiQc0u3ORg5SIMnOySt2RWFoubU3n2sbu7pE2Uv3x4YeGN3ucKytp/4F9pv9g1zRBEYXvU1
8Pq2bwCQouyABWxGPcOhbwmHRBHvifyGSVzDFtf+hpAovVb/d8Gw/PpiCKcFLRO551b+v1BWop2D
GbUiN2j0bwAjaLII5f2IFLvPm9Ly3hsog9NP/6mvTwPQgsyKyJ9T/zLQdiWPoxx/fTk7y9lE5p5s
InvX1PpbAH0pzWs8mdi/o+91pCAyUAyKbHnOXpEiPvq8TeduvXsUInxNKhkDMG/32ai2QzgWBbjZ
XiZVuYUGEInn4RxqNFTShX9DzLUfcSTEx4Ivbrbr8rC4RhQX9pSxY7S7wi9fiLXVJeBlsjsDb/uG
tq41HDxZQcspDdujpctO7awGuFmCyvVs/X6mI8BWE6QxgZf7pc3fE9jR/+JXUL2EpMEbdlAquFCZ
tfZmR+1pci4yF5N/JJ3e3Yj30pT5F4D4oDBBrFvmk5NhSSFgQSgzTJkUraPXZIQ+bljxEzBzSgvD
K8N5aHQhJoK8x8IccTwkwH0x3su5H71vt5f198C/jOjJm9dA+TZVuUWntwz0c3+CXV05rJRAQ9Qk
IUyz1CshTP8PcuhFGYYVjGSdxJjvtb6Knia1ARIsoCC+ogpUko2scL55Lpv4NcPbIA5qxU2sqJNd
CnS40TvnN755B9L4eRJYfWIlo7zrTOJPIQVQdCieKHXxcq6F69nen8ea124+dZ/cn5viE2k7x91J
LDyJOTrIoOHUWR0A3UXhUKngBqgmIPpJBVGDYGZAZIrIN2Qw/gsThnFgrgbTs36uHrcalV+2XJOa
+4aEc29hjEliNXvIVymG/XJFMwuD86UFO++M/DfXYx0KsWWVPnbOOhuLUE0g0wpAYO4vfBfSqWRk
Ou/dL2VyqsITU48Xv3Lq8lCJeOoXqGSLhvL803Zq+vfscFw8MoaR42poPrbD0ciKOSwXJYP/VvLo
+z5shphn3q49G1cr8b97Q4ZVscVZVm5PPOtMhdxObt3i+1sGbUeWNux26Psb1fwKeD95Iko976rk
Gj0ph+SzCAFusBg/YdoxMslkBGFIqXLnC/u6jshizNBo9cA4WbzSlVum+vSrTEQnKB9fnkEmlxfP
S1szlMDSd5jRbvALZgFa0FT+euPZa8A3Bon8lZE7vzaeg9ehVaLOZDd0X6//b7Wbdhp+v22RdBdE
whoON6fF/T41AAun0L5SPFoFyJX6g+whN3XFgJ0efneiWRMFj7WXaNYgD45S30ZX2OMf7FkyqyjG
qJWg3HSjErbnDN9z5ICnftVnMknVEIgUGHEYW4yty2dkQwPwaUgntgBKrv5v2PK+x+9eco65Sf+W
97DnJ9rRPU3n//0iHxLrLDhJ196OoAvcttu3iz3NQKEjMMxfOfx+cz8hVQuavxE5ecstrbD99z12
cTNfpOUumE2MzfZZZq53gO1BN1MIfstQL/XRGNOFAQHFJ3x9PMT7Sv+I129pOmh38Cat/mfdFGJn
QgWkBH8SXoiv2iGW9pB+wtD93Y43QwkDydQ9uS/JQB6pRIbe1SLnznZI4ljMh39HWNkrnlAMsHGx
hIXvLQdwFYWah78ZaDHim2rEZ7Bmkt4q8GE/eEue6QqgMBLRC5rbWdPK0hpu6kA74aPtFUh+wja9
Xq2/2rHSISjl9U/eXwFZykFLgWq30UdAEJk+2BeGeSqSqebJF+LIwsl8L/QKOIXmIPHrGFeklKGG
wricYINnh7uzmEtbOue5XPx4wRhfHRCwaev7G88a0Vy899MAWoGSDTb6h32cdlC6KERVmALCIjCu
925dcOEpkwL9Ffh660JCdk0yjlAEdmbMfQCRKVzCAXq5iyST8WgJx05ynhSIpIUsZgPO9ferZQUn
ECVpew+hb2A43cXJvhnCvP8L5u8v4vGDMdlF2VXogINlcJUra3SqY7pPIepEv7Zk7C62EFo4L3TQ
DNfVeP4lQX6R6nKO7w3BBMpsJD3+hNdRvo0nu4JTGq1KYGDWTGtlORzXDEKHpf/g8vy+HP38B28u
ds+pMalzFDML1ap5vq/hZLa2Vnngsr+fcUGGTJouzKz2fpbe0Mp1wdBy9Xe6vnDeJb/TcUYGWjSQ
7vHKfPEgJLz0SnOOyXaiPm289OWEY0YdGtke/31lnNMm8jph2px2E0qNrCXDW8xwPvzCcfL6mM/b
VW3qI8mZF3CPJAJrioz39HSNDG5YSquUXDoK4R8v3/TJS/afXYCUYP+kNuPsmHiiikpUzMXdsBLT
jGdDouq8ojQ41WlgTeEHBx2q1fFQsyyYkicTFLC/wCtFF9b13jffySfQmR1RItWknOQ502iJkVs/
rCGQ2cfzgSRxj7aVlhKEzsNb7SY53SlZV0GVwJWLQOUF7pnmZxYN+9UPXto5CVPfixBLEZa5INAI
CklkD+VtYXQFXKf1Fz+VYBtf8ScRQ6fdaPshP/zdCjnsvhvLXMFgjiSMQGohEW1XnxdvDOcm15Rs
8ZZ60Kz1sO13aHG86TRab6ZsV/TMjTxcAiAuN57oauUYx3hmrgebIyKMh8N+Tbh3aOKlImzDQsxe
jS/2AUB3cT7gBnMt6UWm4gM3igBM38Ybj1o/c16sRwvErRKlweY/ongzVM3epes3ko+eZ1GShp08
pzo9jZW8KweHB8TiBUUYoH3LhidM8mumEJpKzH4mOfXE5ji0fII0xYrZ0SrMej13/8V5P65UyB7K
oKQqX6ov4jmf7ykaKf/fdzrhl+cQzCCPnZbgk4Opv126kgjEy6mSzwQnGOEFybUDFsrO/J6f6JEf
38mCOxu1/dMyxjFTZwdDr9SBuapdZ1RABTVD9Rn23Q9usVQSCju5vVEmq5FipZaOERDo2GKBHFEY
EX+6dmEvkaljfvrY88VAnJJZGbPhDXn+VpGwYpk6EpcHm/XZfJN0FUd1GGyAAqmBC55bxAc1UwsU
hlOauTmzIjxfIcXf+uO3hFhcOlxTF1AmqlfhCBHI4bTOk/rBkKGWLXjLzXLyULZG5MakmtMSrl2J
XJF5zZp+Z4bd1BqHwkLTzKYfLc8jwe+aPs906ALbCUVv/qxRl5lFAJs52U/KhSeEPIjusm1XaHLc
7AAaKN5RMRA3yYtiqZ3gBs0Er0yW7ya6eLxE55nOwpBM6mS1Yz8KkF1LK5KpPM2lj1ZpYwJJGux+
mJIdxvggya2qtu8XJwLDsq30UkZz0tK3V5ueA9RZqrzG8asc9ubjhP2/XzfKEaoVvgMo3W5YGRrT
bnkeTCu3+vdIWko8+8IGfAzVusJzoByH4xAB5lccl702wqDJw9R3JyQGdlarHN9e84zofRKmFHlq
id+Q7hfTYPVjUhBfmOy8mzZbPVjxhZA52ApXr3mt7RkW3MrOHhbRfsr6d2MzcsbtVJ9bO4nqywQb
mgW68zL76btmb6scsWOVycG09KkEFiGC5Jxhq6fEM3yqd00rDNhHKTitm0iNLv3xKwTecbeXOWkv
mD096AAEg2UvmyiNsz3SPp5gRARUdcWg015Bk1HmPM+hSvHPr2xWwFdujCwJb0z8PP5kpNdMfRHf
uxVsGGUDpJgxuB3GObkHNVr9T2ZIgn9dobaRVhebln11831lSWZtK9jSfXdnSeDaP6QAqU0rpOGl
U3fBYacuo4zDVezLe3apoXE/55U0oyHb5QAW73n4hFHdRyZ04GVjPOdzo+fETjNaJtqa3FUWae2b
D+5xTzMshTCvi8hKuXJSy9l88FbCCnQQxw23H4Im9tOPQaBMB7FKC3NeFa6xbpQIkSo1X1fKPdwI
inwqarqlp8PGWKaBofb8PbcWDMHbAxYvm80u5UF01W3v+r1uTUtKBpEc3QnABZCVLfM8C0/ji7eX
5l5rF0dxiT7j57QFc7bn/aWQoLmrJlqu5Yp8MqoBhxEY4S32w8xeYxCA1cjGmYA3WOiyR8lxUjr9
VfPuR1YWdCaGgdZE+UFKCk8CkR2V5x6hPx/kFPn2fGMydt5Yk2GewS2CiCXtXKhsABDOViCPiz69
dEFDs4YoyVKpgo0G9VgA7HK9bUMMXtQ47xKM28SoFKCE6aHnBf7Uyx+2DRFUK5pM5ruAvb0YiJ9e
n9PQLIjjuX32mG0/HS23SmvW7yc0VTgd2wP6afUC/Rkij8/BZWjumODrWbZTtNWZg//xYSpWkmqe
7S7pxOlDlW3Ds5UwNnJTjBhROU0wINmmtfKWqj/QqEltj0GA+EUvny6cc7JbmFsW6zdoO353pXP3
D6fxT0tsQrQSaZIGos7qFwjFjzCLwTzXoh8XljzLkiBdcCZy3jvoUBZRmhjJpc/8YNiSnSUgslQx
KfSIj3tWmXMWWdbQKFGwrYzfNWYsbTITJB+odDx8PuULWzEzo42yGe5sSuy/8pCTYlPxV3WvglLG
IscZuBRWH35nhQQX4YhD6KwBUZ2KfZEzqYg80vR3Eyt8MhnqrqLKXFalsM7LTWudDpv/BwBFbCER
d0jVRa/9e/L9jHNJXYQaHSAyVu8aWEvRkqZDIXXrhZKAxkThJpNsiwnIM0ySrIXcoKm9OzOPP6ll
x/d/wVXPY3S+Qo3owv8L5o9VwvaZNnDWqbLZXJ8Jj11mmcR3ZKJuuZN/a+B+3pEGfodqVApe1JaP
vMLhqIHbu5yUtHE0FdCYBLqjwIq06iS5FASLvqjQ8qlkK70+oU7x3K8/qeq4TZhjITjcGvLhRAx3
12F0J5M1DycHcoH04Zo5DfxX/mGVCJtgqtVSd4CvM/5kF1OBMSyr5s2WRa9icnhxrko8SHFknWec
kdN0zYQ9BTtr+wRNWzN4ux0FHS3JS9K/SrrI2woE6ox7XnvHjIjFu6P/4rr8Dv3cfjqhE/7E6edc
1YAtHU4qQ5C8JwAZJRvVCCLGmDtPB6W3WBK6Q3gKtYDSkLURmcMmFBDUbaT7wflY9maJASoaI229
8+z99B/tBcc9J3m2TCxvPpeJ423M57Ys78aKOFeSxPslqfl352wvlHLhc7Kbj5+aVV7qK53A3u74
U8SKhlaLe3v6G2TpjNhH5b7n8VtHK+3N4Rkh/Sj6s6wUAZfYfO32aZoxcTwJLeQa/ba5XsgLLR3d
OSqv3W3JEInuhcJ9qgUdSzf9EYBp9nCZhMTUgYojzce36em4JuS3+hpX96q6W9E2LsNvO/gRuH3H
OxYUDtSZ8lgxLu1qFTDci5VIDhyFw+ccBQJKfllM6sjYVKWFXXdeuJQne1JyDcoZIh+r4ePs8Iz9
xVDdHTZCy4PPRnWXp6DS79gHEIl/imlyN6JP4hDKBVVDCi6PpI4h3aERHiWRGhcRNXi7C7AmR60Z
YImOFeWoD5na0XXSyMzp5esGHTz8haJPl4QF5885FBO6Q2URoZ21ZbzJPlxgqh/e5cA74ROsoaYG
zHQ3RICANQLooN34zMLUuo9gjytnyCvjnmLZQs6zPpxfT0Hae7n0SovGG8NidfBvyFQiHNirlmDv
oJ6NeiKlNQ2/nT8viZMMkdSHOZRXKenLMOR79NUvwgt7l5W2kYvckikyl3JDUE/KR0otQJib6EAz
/OGfhql4RT+yAKlePTiFcWO1J4kPyPbwfd/UPuzdG221Q4I9f1zMjGBxmc2sQJ7JFXsR+ZI314vc
TUL+/IIPgWAlXx8wh4dR74+H0PW+GGNl8jsSsCHNL4BMi0yjD9oLTkfdyem6o1stX0jRKdpr065M
U/8z+vrpPYQ1TR3Z0ymnd93AMXBPeT6NaQPnXbPExLU0F2RLpqv6eHMoFrYgFTFaWsMb1Qy6OlK9
g3eXxzGNZ+GcctQS6VgO4bf+mqFRqL6JJbtbYomw/Wv+Y2FPvZPeI6pWtzWDU+93m+D0EGkRpMJp
J0nlr9jRozRhs09coCcTrlvyp5/8gVh7un98rmQxy8t2YTAcLd7sk1+ulYN/JLjguAq/MqCeb0UN
awjfFDohg80+tpQj3yaH+gQVzOEuQKEy7TfD0gR6ON4nQD1c6gGi/VNMQC1JGBnqHsAHmkndEYnO
DJ1cd+FHp+MZ+cONPPGdr+avahd4jf9Ws8V2wW0LVZ81/bBPFZie2RSI33SIVH9p6CCLKan99B/s
83Z7uknlbR4GgJKjVy5s3SqiPAjN+DToS80F+/IiJ9eNwe7M9Yj6lrX7X+OBOhet0Sm8ewJYU1yt
Fgo4fX5/ZGPtG73m1P/dol8GKZEzRm7nni/yy6g+IctBfY9EYjFXmnbpDKni1STmOrzW51Z+NCcq
Tt5TXZO2Mp6mTuGomRXGCxf6mznBhxt6ZxEAZ10twX6h0wO8FjxyVyJRRby5MZWoYQMafmuF9DwW
M/f86KVaqs/FDWrrV6FX72Xohf39V81T7rZFZjQnEpIBaKvojxNdMJmTUBooScsGlGCsqvz0bZga
U7opO8SukxBjDrAkGJjcdDl6HgLcam2DshqwyD7E+NhQ7b8tPaHkw4Ap621MGx6VB+KrRMnPJyBN
GB5TtiN+I1GZHPoP51L/1/fTs4zAMjYnm1hJo4XJlfhp4M6CQGWig060ZcDnRDEYXfsqOmkmImms
ACbrkfsZ6n4O/ijT297vLqfRomQScDoVQqOVK9PZjBvXUje2y7x+2k2uknjKrgF4nnnEU3+N079b
Q8suvnLgBFGqHWwsaa1uWqBaDQs5EL8KgpmV7I3gNQn4ixxHt6eHNh4JRbgn1I13FpDoxx3KKw6y
zlqMMdmepWl/bVnphT71XTKuBb30B8UAeyBS3H8j4HsXTyF+myhxGMzCYFDV3LVojTFgAJhMw0Qf
N/OowVjltTVr/3LyNFWCrA8lNG3aV6YDonJwOHHllDWe
`protect end_protected
