`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DKaw2YF5X/sI0l9aLdTgbK/M5GUdtEMTnIFmxvSMohXCNpaRunL9ipaA59Dc71YrenIGtec5QT4M
zCoGKmFbyA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QRHRuF+/6jbJdc98CuDuU1RSPkw4Mrd2rWInSv90clZq9I1OTAA5/xdv3Hk99Vg2prXDV3YjNqoB
pcpnTJxql+YZ6VAzN0qCk+oUeO1cCu3qiinofcBjVXCdgYxomUKUeE7FJeYz3Js2G/kJGoeHFW9U
+zAl6jadwyF9Jbvv+i4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lb7wQIOJLuT7MorOQ8eHbXO7nLYJ4w6DRb/CRc0KXgD29tV/pKu8nH2e+iVICJbGwJJtQ3k8P1j/
LscOU8Hk23tTbvsi/KP4jYIAhUNpSlUfm6H0KJ2yht05tm7/nGOSq+YwUD5ni46LH6TZmw9wRjLo
RAHSpBohLboc3y/hVTXta9kQmKPnqAmdZWZqkVyyS5o93+63/fdqbFaxxtwx1mXeZDQ2+2zbTCKf
tbrO065IQsNhLqpQ6GmWS0y4Yk762FiY/PW8xLoCZ1V1Fh8ocFk7LKyATUlQjo3T4vsNks0JLfh6
k4wW0gpjLf86zBHim396ye0D0jCoECOhPpGtaQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZXacKhqAwgw8zLrWO0Oej9oQ1uNqsfSW24Ju9AdSqiO9hJgeX3QSs/Auka01BXmxZF02hREfAK/G
6uXtwOuytUDW3C0vu69znjuzfKa65iqAvitXfuV2wV2SBDUohxstI576S9cHfGPfoJ7tVzjIg2t8
+fXxMYGWVW/hL5Dt3LeBc+ul5BEG9/vwugVmMP2uMG9nGEtDEQeLb7bWAsdsP6jyz5L4K49swiWc
6TrDCW/53r7o1y18s7qcumMrH+8e09lZWlV7gV/qSGCmNFjNoXkvbq7X5+RT29nF6kaEY/1Y1wcM
sqDv/0rI3Yh5PZatD+o2YnHnz7Es16C87EBZrw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pkb010SLYsAhKXcWm+QlAA9Be33Kx3pWG3KQ8c4OXZxiNI+ziOzdNGDZkUALVJhYeeODAczIsICK
xPobg5BZJdmnFjXMkYzJiVNc7H8OtQ+xwCOlZfGQy0nG30bs3aCt+0ciZZz0ed8EJ3QfOUNUrA8S
ACDctQvzk535zqal7JGqVOcbax0rksASegZXl9TYHMAWSFXsQNDtHG7HCq8QaEGySiiJnEz1Zygi
CXmAaOXrSZ/75eRU/jV0Zmfl2uX9M3RD4WyT2L0mtTPVI1Jo5riNKDciMqi09G5yCgGBizlVK0Le
ynsKW0Fvo5j+TrmGuES2+DcsvwzxQUmrQ9n9YA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
saU9xQVocYCNVhmm+/jaIKt7f7lGDiBCwD7GUeN8jk+fV3dDx7VH8BXnwqh3bO2UtgQTq4TYazR5
PsEJU9lk5Y+2uIztywixaUOcY0t6PGvi6DZ5S1UapcNaqz1GzVDJNMdFrGWeodfXgyVpIeng6Jtk
EKceFNW0p1SgbLjlCjU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbTosJ4LwLIDFDsIbDQWyryoCwFpua23V6z9HaJa95eQ/VgCaYwQRc0pJmp/UgRFI8GxRIcCfLjR
nDQiDTQUzYsgXuFi39wSqyum1ybk+zJc/c0tfa3zo7fAh7WEKBR6EfegxJoOfQ6umn8yMUOq35ku
5cQGVgAH0mV2j7kgcszzSTcMNu1shLKlPJejpCdXAsAct77F4/JiYgr35R62Nw5TiOPHxLGWKlD0
S4rOzGqDzYI4jb5eYbnrBMtpHWXse9ybFZPj47SvpsioKcFIHeUE7GrNOvNDQPdNPahScNll6gSb
fa6tuXH+3Q3DQNGg7RW23POGEp2w+WE6Kef4qQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
VpynYjFs3lHshMpL59S7SvDJd8vc7dTEu8GdHtlN0PlCZoXU2+LM0NAqk5r94gmgb+U9bJHYqo4J
anpfqNNXMGFUSYS1DemQJtS3jIr83H/ssGaHxgCPPM6q0E6mvPTNII6Y8T55Eis+l/fyWtseLZ0t
CsctF4/oqDFgjLiK1zzo2fMZIW4dLWuzGk07XBKPT6Z+THX79GPb/mzGPx/rUjBl+SVhd/VFXWMe
3ZakdzORzyS1Y+9wxtF5QLyq3Q1oBu96GbC8AcLVhB3+ZZHak+fGU1snn56MBbC317tuB3TS9LCJ
dxWlnLcmDrGOXQCm+f6+YroP8jq3a5/kwHTx6iiO1MMsyUOR8GIEfrmPLO5tHh+SffLIXxLGi8D9
zkNTHvy3TumHZiIUt4I9pfnY67w9uzcwFPNcdII/dbZyt4FNsHVp3i0CIQ2q3maegpMA2khwkzyw
fSnZl2hPf6V7ABVjQRpLuso4qIIuxpxgrwR58lIn1IoikUPOjm+pVT4zo38aLs8pILLIU9ObLG9G
NJlCbIHt1W1y3Tf8V2OgO8ShQDeiEeAZqv28iE3gaMfrhRGRVHH2l/WOQ1lISV7RKMKrkCuzmLRV
RIEuFcqxuo8BOxbhsbYirPP4snl78Nn4WTGj9hZNb5xaYm0URvwP3gsnfMBzbd905xuW2NkEkWpU
p9w5BUZdwRbZeJRrJOhVUcq3SsHH7U3XwApsu7IRTYpiyHtW8YjqnHnT1LI8wRqu0bwRrKRXLytr
5GxqfaYZDV4c8SsbdANq3eDKZZ0QTNHai0nb+aLdBttEBtbUDpO/1ewhicLJ52W0R+qy7TRO79ir
0AYqKsfuTROMU+IyF81+3y5wfRpFZSkfLyCqOeN1me4mRyKXDBRv4IGtpXRzAxQK0RljLafw2jc4
jLIdY9gUKcF9TWg7/lTgJSwwxpIAzhTXTQzOHj2AEDf4LCEDZos1uDMENCRZ6DwNb09UVgoOc1q5
YLQE7twHuL3NE3dlmuuWCLpn83IGJx0GWLGo4LUMWwyb0PTN/qfaG/pSCp6DZZBdycD2tLcZyM58
jiS766isaqwcXRB/8UU+PUwB8zWVjlqMm2tL5YTytNp7sbj75BpA+j4lHf1fkryFRfABEXoEJ2G/
M4Lde/48ZVn20wYjhyUFapGSAsqZ+BAyZo3lXMAw9WP2FSJmH6jz2o7/sK+sk7e9Am0pPzOpKXtH
Xf7wJq7wFwSwZSGROT1NBHN2onmTyQeE8npuOEx16gP79YuWpBs5Jovmq7CIxQUQwNC7toasPt9l
qzwM7DKMDALNJTu06mJFF+sJUz12YRsLba/bDsn81lh3Jc/C7AdFaXl4sfvaA9HBTSv6IMk9bHb+
nJFFwVz04FdBDw19bif3G2LXA+yXPqdPHisUiGAt8vChGxv2iWHmmY6pBU2ace1LBPZe3gAaJ40a
Ns3q1hMsvnPZZvZECC2I6XmkwLRH1ZqfrxM0ulA63tRckUiDweNWunX0Q3TNfp4MYmNt49T4sJlK
kKHp2diZAoJFVcmWzekVsO/26YYJEr8LMCSecSFx0v44cCve6t3xXmCLzAgAGTYe2xtIrZTexF4U
hFV8aM8dSV3BCrdTXd8uORBnAxB8leJYBnLpp4qWF8NalHrnTQjsBUafzJ9jcH1506qNBux2MlXx
dQeq9BxGmOnN7X7dvHrHTN39o8PgCzUD0xnM91gIRxfCx6kFo5j96ETdaVmUeOeub6DREKe0idx9
5rAfKRenrqdw/Sx3zrep2xD4GmjCq2pjl6DLadwC6r+7qK68HWHqODQFovjfyyoFa4e0t1ZfllFW
ZMhtsOjyqHlb+wt9Gl9uYFjNxVkAl0U1LbtyBtR0AWsInQzZoj1Y5t9Us8zHdOUBOParNkBqa79m
UlNPjMqL2iDgLfM8cBlbVyUCv3Erc8E2uEs9N59SZ9iGP9vdqpxRUSDhZnydtjulIwSZ7PlKCFZu
Id83EPhZhQX/gVbZW/lsiVMo9X5P06TdEWB25/s43qCleu080IDHRFTGmuf3lsRe550yABPeYnKB
9D5OPFZJbGk6wRDV/HHuOLKcI/rrYqqaOk60hU0X/VSuqjXjp8aqdC0zXsrIQNGSPa+z1b9o9jhV
CBJMd1AnCawCBUloRWVBsdenG3/9S8hdLSq0fqOe4sr71iUqVIGjXtsOPKxtzu2zhnvWpdIRQ/dG
gLtkene2w03sA4DwvzxNVZ+7UW2ws255GgWNFzVvKdkLEQAWyuyO5wB7bZsqdg/vt4UKCDayLWFq
14ydcUb50TLEO1tlor4t0J/0izXUgDbug1h3XXxliSEqaTeaAqbJNTtojeGvqrZ7DpM851WtDlls
p9X5MnkjJXrdX+NNA07LIkHBcn2NHrWznSRB8GI/s5wrLGHXKP/bB0qM1sAkMw+bkgAP258zIz8F
i6rC3IqyA07z18NInYIuJmneLtPfE1/N8rDgKhNgmfX08EsO+rcUEfZLcAXKulzNXxcT2mTZjYNG
2P1EnrKH2BWmPg/lWRc4Fz3YTJmlYfEQEUumcytvsPZpgnwgedD+g9tcXibZ9NPOZXg96RgowyRq
c4gIDGWpcoorJjkIsyMGKkdXl7u8Qa/6kTzug9lgCmKVagL8NuNnk6OJwQVh2PYtAgJIUQwnDRAl
NJZyY48L04WqmdlgSBIrWR2G73Kzgvemru8l2K6fWNMII199IR7siJJx6y9PYzIDmCV9ECZUUZ/A
gtP8kGORULZG1fH5Rmc1iyAo3v+raDY2nU03gnngMQ0rH6YFxKTVCtSWRdgTPObYSxfJ29xMRwFy
vKnZJJUGfxLCs5vce1rnLqoohmZd7nIaR+4FJ6daWHhh6r+N82Tah1qJ38C0j4RJ5jjfszyQTjVX
GElNV662yjJL3yNmTrUkjp5LtRXSP4XuCT/00vRF4X1XMmTzugkNajp8pcyQb/9R2M2RCfvV3sXd
7farH3PkKovchByeoRTgcFU8j+83eue46ZBnTnQ2zqCFwVc6JkkGNRM1XI9fgFkfQ/8nJELjVe2U
+jTHY4O7Yrer3VsOoRS+kCNaWWMHn4XdAtm+l7peZqPo/tD6r558w1TXhCp1xlpr4Z3JhnDLLoYw
PezN4uQo7/Q+ieTBRO3HSZ+Lz9r/OEQU1n5dTatS8/RzQ3RYF5siER4g2G47q2PK98RMjG3mjI0n
7ZHbJJBitKoSU7y6NqB4Fw7QIaUidlMmHvrCI+A6PlC8B/ZwTokdrjQ3KdR+WS/9QvwBps4/Njrx
FVle7BVNEtgzYYbU4I3vhT1O/NKmnIOGhHNetUhKkfdXpzqFZJGHvupxVeklHl66y3ovtSlIsUk6
8NxT3/5VKHqtifan0+/p81E3QOgsx9YIo/hSZeAvjyC7vyLmUIKi7eeHCNSLM/6L7qiinrLEtLOw
nKzw69EsqOC/ack098VwKUNhTeKwqFDxfASR/h67RKKbw8ITac194InsH0xmMBIpbq9tFCoc+2IJ
f0Dt0I06+kakxf1/CFFJ9P0wSfhks/ws0l/C2MvIKCBeS/NrDmANOrOOsvmEwUzs5CWbjfGS2Leb
NU0jQSmQYPnb1jNkB8aV+iRm5KcL9eD5zjKlWlwNJgiglE1pWdfe+921AmEJldHJOc46SfUG9wDA
qKOPt3rKcQwiP7QrRG1kFT/ea1XS3BwJEVm20wqxQuahmzjYYNlEEmHzAVMAAAIjL5GW7Lc6UOm7
Cd7fYLLjWeMM5dSrVfKHN16IoSMjDRBPOiyajjPRMGXW12CEeS1S2Ss6AaY6l2SLa10vqETM1F9d
WvbXdnVuZAdO4TXvMRqy9UALzdr6YjuUF73v2MYCirkRje//UBfewiETbxomURb0xBknlIq//vEg
KeyUpuPB2OITyhhXLCfvAj/jxvcYkKApZK7U4fLwXL5J7m4CIoDM800PSa8x01SmOMcaMFzJxBAa
JhgeQckFt+vC0UrHHSrPGxZuzoEQoQhGIx/ZBVHs1SW+o+/7F9WvPlwxmd0PJHgP1W13Hi6GQyMm
zdHJtJl/qhm9NfTEGoaBfwFDvhFIEuUELISC+K7U2Vn/Ywkdzt0HHeIMZ+32B39NY0F4yF5tcaO8
I1JFZsNcQEvU3wd/OhdT7J83pj14Q3CWC1RimQDn5uiOIVq2Pfb9T2x1SJxR8M5H2hIdEE0YmFWG
nnYzzrXGtfxcpe61xYnzIoZE78cLKIVgo+O3tkCJKRSdkSaELBxGOSdWLbQmFtYglRuvFomCAL6K
TXN2REOB/mVaRD8RHxbFo4XkCkrjPTqxNL1mmKCdEonrB60OvtlIVgRxRlkbZ0N8BKHAVMQv6lN0
mHcE6ARNCFGuPwm15kcyQenNt2W2ZiAPrfqVHlWOf6XTFcyyrzWDJAUsnDK4FyI3d098Y+8Jb+FI
kwJRPCH26hFGKU0N0nQJR+WaJJec0HD8/yjb0TGVAq42S6v8MHG9UylXqwUw81NILJn1LpKlfuDB
E1+l8g2ygdtXiPk4riZErefcFKCn7vUviMxImVu92Wp2e6XPBH3lCIHERVvOkt7K+5UqSsGfqwFq
zXxElJO9wwTIkH0GNbEZLkdvcq7hUGWy1v38nbfRNYdJUXS1pNBgEHdOtfcqhpRV8pmq6vyeOC2T
OD3mRm9HSGul1h57k/gWFHn56ciE1ZVDTamKgvtmCU8iHokdlU5CUE16FWh60dKW9O8fgV3Risgh
XPSjtFbxJGHRdiKH3cJtuYBrRM11KTRwFi9DVVFd6Qm2UWSwTaWQlAk1kpcXK8Jw9WnScQDUCDdZ
6l56CcwiHHptz8NY9f+hw4gUSUkLBFU0IXtIzmTZBGUwtGlwb67FLPLxGkpj7spKDLurXkTxpfjr
lBAmRwmkI4nG2SCcDzbLqLYy7nT00rvrpVXJ3en20YcukyF1ZUzUbaih/jlPryX1EgLjelDzYEHL
s3+1Jli29m47DurkpZKnm0T7sKOlqvURAnewigfEsgaOvG4mxDZXgpE8edcuRpQvUe4MUKU0SpD8
IOG54cDXu1VqebpJTNJWUvGoEGoEb1RdKARZSMBoU1lRsVTmfO69IWjSH7bAV7AgiMqEsUROoPzo
+VWfq+nxrNmkEF4EtBHEUWC0+wSzyr/kpoN6ddEtdTYIFJxrees0MDKPn5lN4V8GMHIysrAN7N9g
CaP0/pxqBkC3GntwWskBQmyQJ7c2yMCp93tAl+BAT77PW/p70LomFZN15sfNWH+LBYq4Q5YOQTFK
tnZNEgYeRnDRyEThF9MbsDAwoNkK1KFdYlqsdA7zIZGwp7L24obOCG85efLYgRe9nu/fmlXUpS3n
HF2H6gx77sW+tr/TS52HGX3604a6ag9xLvkn4TcMKGFRIsFzD15h49qJ6tCMWrPstFHqpT4oA6rW
ew1xDv3NG5jIj1BLYAj/nZegw9xGUuZH1cDEirATPMq5oPlDlojYG26Ez9Qz7SvbcpYoqyKHR29U
KazGGWKV00o+i1ZQs8Bl982nlLOc2V+4zh4mr0gOLqNrrIJnFHkPirfPAGreit387md1Ojqf4dCq
JsKmFsPWPprkY1B2HywRCx8RN/lkfcFFyR7B1GL8LxnODvB7Z4FGuy2J0QleTnb0oKna+B/GUORH
EVwJdUCyEeikhHgNgllpDQN7UvopoNK/KeD/8H0dB4dLsnzbqoNLcltk/sOSGB6wfp+pPiPlCq8p
I+7mqXPeLqxG4+7k7zx8sN/xM4JccpNIJPc6xCrvs12jMoySi91MXgYkgCLgMk8HAk4R6Z6ERM7c
74cjmDtzBOrSVbgGbyhYXxpS1p55y4sPKbG1gCiLH2zwlJqojviyCoz89WD0YAmYR+O2fJp/tRlh
oVWzL0lIKMWEP4zQw387Rzrw6NDL7V8jMv/B8PaPXA1tqVdjlk/ZuiVPcT7+akFjB74SY7USgdBC
Sq/MVPHtWktGuTJ+/dNABiYrWmqYZQB7nOWT5xue9dCpUZjprgH68xYd5+HAeQkrJm7VQVSDp+5h
aBBV0NkOZ8gXk7dXpYBQuLpcCIMivWlEREJBr4eFQg71rgX49TDGHmYoCOaIll9tO5MNKnda+S+H
hsEI8kWiXD0QItL3Y+sinqAdry1KFOVGQArjHsb3JtcDGHqiUPtItJ5WMO2cPQfHxjyPRiSG95C3
hI7G2YpYeVnZT0B1dMbu5ODg6xsRAzhYDrsLkfe1DnvXgxAHQD4FxvlnXLncq4o2BA4nLQdP7z4s
4Utr6RtwbeZvfbX+WkSRfvVY3mGiJpE/JHXjk7bUWpRzyI90ZOWZC+YUdxkDqH8WFWut5FBTWLS4
7jt1na8wsHdVubCxXIK12XejM6jI+giN38twhw5JDL/ei4YjMXBFsRn/IXUWQ92IGgYeP34ALGtL
bdJGisDbpPoIEjC/ybtuCKtslU67fFJNEyuLVAiasasOENaFNOZSiBdbE+au3YqiRumt8Mc1oBON
ZRqDwZr7QbSEDE/DS+PH6zmYK4SQyZunuBK4hG5NR2/UGPn9BK7LeH/OQB4YfO7w7q2qxXcheG0L
omZVDqlGwoVOrhZxDZ3O52eHVmCthTSzfwt1BzU731DUxuhPQT0y2LuUmpw733DxGIFbkx8hKDaw
fEWI8GLgErE3jrvalEW1fMgvvsaFjQ1/+Tlnnt7Jdw9IqDeSh3J/7JHFI6AvXp+kwOyub+0RJWZQ
D3jUWEZ3ZdIDwr1PB14nk2O9p9nXRAgw3iZe6Xlnllt2m+iamGvOeFMzoA15mTJd6cWhnOVVoFTK
x7WGgGltnGMhwWI3OWFAixE9hoJv0ld6CY6m9/RtPrMz9JKyioLEygDyKZa5/pqKXV7hiY0keqhX
6pTzTsgOOBtLDkgHjOz7TXx8B0dbTbAGyNblY0SLaodoxV1MqzVH7zM/Ffa3/qkzcu6cHIKrcaOF
KFEiiIIhqRmpwcsWlUqkBMAI6bViES/9KPhwMGRAUKEZNjm9Kog73j4AvsJsWiWZsXUHMm5FODX6
oHmnMp0gMKwpXt65OBuTvByt7ZQE1qeJ7CmpSAKiGBL5vIEr/SZgBbmjdUmPO5ae+h4hjHJaxRpa
lTpMKGz5V6A5ZxeqHIkmDDT+hV/U5WUqb2hUfea0wYOmS5f4FYTmvRIODCM87guu4QmDn/+yXcZD
Aa/0VvJFlbirLNvp7Mg7svv84Zda/1GBWaImK+J7saU8E8cLVwKuJJ+8QjnwXCxtVnevAfDP3GQt
k/0vSReZd07FVWm96BZh4leexZmctihsHyEORtFfADjxxpMaoXJxrJhhkC9DmE/w6HSp+mbRqFlc
hMhUHqQd69a1aSJ8SuEe1ppUA/YidHyu/kEB8G6Eg9bWeLdfp/q8t59vAgEFE6TgjwmUV8x+jgdP
6UEv4wENpzW8IIi/NrDy3omvEOBjhbHJo4w2FKIZzrQxoDS74nLOI5+de4pxRD9pN3TlzSAHK/TC
i4FXI3FJ/UDZVx4wsw6gIFuxBEl8BOA/6HnNPYqKLCNr98aUf3g12NeOtocijCIIrX9Ni8PMcUvs
T5Q3zaRx3rshDEHuklrDfb8kQ0Z62A3eunJ+PNGmfnnBT79ti2FEOqFXiafICM33mSv9Kav6qt6A
MXJDNobxADflmATic5Qamp4ufJyD0xcoVHGfafxoHU7ImWdyM/H/tFTGQYYHdZMdFxbLViZzBark
VLPXlu9R1R/BD999bPg6uugxIuNYwV7BrXost+EGiIrdLk5RjjKfkNGpE59zvCyXlJFfQ9yl0gdu
1I6IDqlRHYwq7Yx6PJOAuMG9t6M5/YELWb0BaHOqttcaVadqGnPHK3S1fV0xYXinlvyxOgN2t1GA
8vZjFxw0f/MbLQuN8k4GADOix43EXaa33JWIltc+jUYBJgsaZplByhAyxHIyZMfM8lTcXn+HQcJI
M6Sga/zPA1R1+qlGwWNNm+XDg1umdgpbEL6bHAs6vBtzc/g5r6aP7jtutZkVn6m4VLfHK85F6jYZ
pgsV668YoQ/uc0Cbo55Cl01vXc8BtcSH/s0SZ6NbdylxfoXDQ8fG2KEYmf1++giseTKWdpdqyeUr
ZVOBiW53nzgWOf0MWnGA/pMoE4fwZqMWgxDzaUKgJ/DTY4zG/NVbsldUa3g3a8MQKVlsf/wg8ORO
bTLZp2ZqH8+CZkPuRElWFv4p+AGDkky7exd/MYytpQsjJ/TGGi91rHn64PEVyZtm7qVptF7Eegvd
XtDHCBR/GxJDyt01DYnlwXbtuicd1EQkJSxPNyomnLTHd170wD4/S4wrp6YEnqdiEPSwKMK0zvxK
i8I0lfUN5kFHrQAkhCYglD+M03+ln5QCOm8QmprmLu00ypcuasjMv8hJXZfs2Xd46dnG/Fnu8sy7
grGAaKhGeJzv/H7F52hBgem37i/Dw4X+jgvEhpzk9HCsIm7CjuXiOUjNHxEHwQC5LGJZdp6WqtiN
40Z+lN440kPTlAs+1EGPdH1estDI7vIjGRNlTsoxOoKHqO4kp0U6ec01ksW8QRfiUVn38PyNN+Sd
Kf6SFvQIB38aw/D6X72ThOBKsjJr/9uQ3k8DX80+MNCDdHVkd3UYl15LcyJcwH7XskIDNyH+UP6h
kfqkxIluQxnrBtp5Ugpo0YT8qyMiBJ1U1UTo+QJ7er+G+vUj/bGu4aYs+N1s6FHHZ13yiUJICUgX
itAtQAAfD6IuTxJwKo7RwQ051jX6SiN8ZaB/mO7W8ElaR8t70kzP6WJXKUXQmxkRm2JBRdO5P0JW
RaxNJ4rVcSOCbVRetly1Fax6LQFuq25PiuiF0bVgN07Ziue+hSAZUgHJhLgoVrP2v/LKPyVKz9OK
uHyH/PTuxG84EVG4PyYBRP3rH+KVXp/zwUmbOHHhztYfVTVAf5OuzGVYrqifelOwofcUTDkfgioJ
/NddT8bitboP6+ZH1+g2krdlopNabh50lpd1eVNJDemJk5GqIa3gy/P8SIdF/JFI5B15qCUtiMbq
Uh3RbwOgJxznG6/BgbfIjXBuZGReTQ8T6hU8a0nmoHjtLMm4IR5dFFwbH8F+Din41gIAWY9g+MNX
0sMgJwnhAKsXtMVQV0EziKgYcROuPkxl6tNwqV2msfiZuHCmyXOJ4clquPwA3gLYIBCfs43FP171
2bbZ9j9sP8RQyVZQ17DliS8j5eDbjJG9Y2gOZ8xkYCXOovwsZzhPTZzMckfmSv/j8lmMNzNpRpBA
mtfLYFXMri+x76QXUTYXuQVrQvGsfIOIhLuHk0yu1yv1c0IzLc/Ehp4iFf+8b60UW5un7vTFddKY
tdDIagIliq35pdPIsb4zO3oOJyc5HkPO24kThFLsv72ZW+/SQ6Ni/3ExmRk/6F4513vfmZgm9K0J
+dQNmzPb0V9tMId9FsV6cUFzNWEW8ygb4Xek7USx46ByiBCl8OKkDcsx8XZ/fFMTS/X8togyXL4m
ygc7S8rDPoN1GNgG9hXKc/A3yFehxR5X6EplQ9s5NEMgL9hUnYjSSJzFbyqCMRMpeM7kkrskUiDl
K8lGUSKgaPDKcqRg5jmYzYRqFqkW9rQu0C+qpx68z5VayNsDpRym5eG5BdoHR3mGpRtjs1NuS4Mc
vQ4The0R+zCZwGeVp2nzr9MinZFedRqoAtJ7qHcMCS4/rVrgr23mTIA5ezjh5Dq5gZ8AuwydfS9P
KhNdiO0obM89SqPOT+n5U9b9CPez1UYNsrOBeZqSyjFXnUTw/bTROyrW0AYrdIcx94fLZAzjahVb
FqyoUdMVZYRq0JqvuHveHLph2WaLhnS5TgyRUIYkqYTRiIB9AQleHXcRI7nVUHDWtoF6PH4+4sm0
gccYwpn0BB935L468DHxkhvR8jVzz0PFxXsPUZukxmFB5Ua75StkBqNsk59wNuH5i+UzLMOv83kK
JXzGeHHawRjmqNOoCx+YHlMfcaC9VCORslmpHl0c9s9qk7rDFacpYsl8BrqSvGTvCd+37AsyWDld
OoFymJLlvlad3/LUqJGIdtfCnQn5tnT00C6OuPdvcydZmsd0wqGkLi6LvUZCoEbNwEjJ+x7q8yG1
qHTAia6RCuIq5o4zm0xvYipj7woCByl2oU5fvl4gzxt4kgmzX8qKRn7CwXOytc2fLBq3vhP/w/81
Hr/7OUY06mu9nJW89giOz0mPoW8HLVDyoz7ZivR4u+Bkne18z52Q60HwZzodkC1Q2oUXAA4H3o7T
xDeMmE6uw23Nq9LRvjf2YQBuWgeO7/x5aGjl7tXjCQJEoeved5gRsAPPpeJCJkzpNi5ygR9ikvTI
on1Qt5Alv07vFbfcWCbO9qTjyOYow+2s0fcQJ1YpySbwy9kmsMhtNfJDQ+HkYkfQ7yMJq3QvcCGN
EwE8+L9jlLWp4fGmW0faBd9hNbfPnztiaZ29AG5auTeZmdNbnWvI6n+vJzSr/ebXFGamjYwv8we5
RVzpKO//v+RmDfbBgB7qjW7BFNGi1pPjv+HjcNBi/eKC2NMkWCyOP2uLsuYjRvKhFJ+Si2D9xNnV
hbBG1CNOrkSnL6IdkhdSfbdxi20zgohBA4dN2gDtfVUWZG6SBs3f4RxARXjAToTxmscnDFqFtbZa
Hge3OppI5/y0meAcDboHzXD7uNBjBvHd/LputJ9fWoV+S9IhpdWypycnnmKlIvIX0qUgwUGXVJd7
cVm/FRmGf8yY2ExUN77Jc+PUFIt6aJYA91d3KL0FCRPASTLlyYJNuAozlOpPsXih1NS1qteFXhKo
cD9DBa7o7XCUc1+h5sAr0jo0t7KGsDkscD4ZPPc2orBYXw/Z/ZVXFPYWqA4cWemBsM18eWagQI4S
1K6kZ0YAczy1ufeyOre7tR1IpnPSJmSat7zeKGc4wVEt2bi4x8LSxjRmaj8cNY8NA4BHiEXjKP6K
z7D2SKMvwTKRZoMaDglIRTQwTANusfb1qQvvfhBEBAB1xscKUqhO+LjWpLwiSa1mj8XfHZYi9Lnd
5PIS4f3SK6D6433b/KZoWfpcE4Yi4XPmVy2Buf+2QyKEWClmGPCwiq889p/hgZ0fJV0HbBZQHwIq
asD4L5+S04LvkKJfXLouEzFfUha/uhJ0E3d2k2G99p7cveeXPkUO4b5aAOGIFJEC2LyFyy7Zptge
Dsmql2MUy840Ff051FGASridRvRZ/lMRNMYteIBi/6l76Mk/1i5WnXf0mB7RS5GCwNV5XU9ugd8Y
9xZxSHjYvQDRmwn67/QpYwqxz3wnVTh/Azm5AMNW+1oUT8OxVAASw+rG/orHKu17NYI04DSPT9rn
7OxcxBidntUsthSEFeK2aUUrEwoQCNa/9659SxDLfc45wb5g05byv2gpfHzVoH10fFXi/9WxMigW
Hk7yWfV27d8vRPjdf80svB480z8yWh2R/jvxyxWyXlr/gCMvbrLUKDmmOhGhcgxahtkN2gU1AQdh
ZGwY1Jo5UUzngkUxwqyA54n86aL59l5qpNyhXNUD5ZCXU76s8IMi5KpVhgv74kxZbxUVNWZgeuzy
X3MSypGwcfEYB0C4MC3HOav5j1FxPzztD6BhyVi/yuaUGCDHU3xPL2jKc6eK+uJNCUF39DL12hdV
iBMHI2w1tzuKk3njTg/Dm0QGBhZc/pp/ODlMOYLz3FdZpWVVzA9tjGQsYNTm4o01pKCHsZARceqH
RvhyUu0U642AGAD3pVQz8E9R+BfnmIGhrrMBkCbPJuqpDBVZWa6tVpcTgR1xycKVw2XHJ1Vzd7yk
nhmvN0gQYMJa7dFKU0b1a41J5YoP9CotTnc0PLH6mRpGI1D3ljxqJOJAk6fT18dFrld2YAJAxIif
j4cIH+cLjv9hXGE0ldtwLKgZXbraIlFMGpykS8SOyuQFf+nPUpmON4MXQuNVFE7mZV2yJlD0QFId
DWft0i4Q+xYTdFrp+K+27Le6375IGBzrAI4cTRddxpDCiTTIMYlQP1f25KtG62vXw9I5G3xuIcDw
9sKZR5NaXDE5ERDGMoUHz1kJsUKCX8pCIp8E0xPjgr709POXCeEyYaPEEDiKaTJYstb67l8fQ3Mg
VWy7gReB+zAqxvAj0As4k2gCRLcNBFL6q28eidZy+1WuGImo+cPyya7kpYZa6pZrvVngvsn0AuBV
0z0/m0utTi1pXsHVWkOe0FdtjvLg/k95IdDh4jO5NAZRMFGMAz7Ea6kTtAXZe5LbFUZQY42ZKiWj
betai/GfR/j8zXtzjfIHD9unGwhEItnY4Nm5MQXMkkgzQ9w6GlgQXjw1oNpLqlaJ/Q1wfVZgFr2V
7mxAESEY9IG+go/u7k9ThJ3m7HXbuPvJyQxLQRgLFfCfW2Hd2e8rUlVMRjKE3J/0F46gXP2e2xnb
fg4GDG3xrVzZ/5XfIpIYNEp9aJzVaLJVF3uZN/vpUNg+OxKsOATHFgGyd1SaqGqN1jWkliiquDZP
0za5D1RG3t6ET9L8lBVIQotdFESMdqCnjJqzEpXFyHR9rL7xwWjgi2gk8Bx4I3n0I0oZIxyIEqX/
vjHD7L5cBriNEgHh7wbqa6NW3uz9eq4zzPt6eUI5Pufniw8v+KiqeVrYn63eFaGXUyCOsTsM0zJL
T96p5FfShGBjaW6TZGaTET6VcUAKlkjPzlxJx17Rt2sbOeWqi7Z1bDKec75LSmx8N+fOrDYtQKsC
kCM7lAL4J3+HTTL7lHY2+U9npF4iW1q3cBGlibN89kYrGYyjXA4D6wDPB2fyODjEcANq3x0ICWQh
CmV14MZA0AArIprKjF+GaEBoESOEA+S5X2V+cEaCxcDl0/OATB98QgEQ8eBWsO6gzhUhDfmeMRBs
XIVEhRSnCJPg4b0e0JGh1cb8/BOU0mpLc0CfqypE+1FkkSHdHc/1e4CUGv60ccGlciRqOgCNAQZ9
bsYI6TOidzkqdTHqcSX+k+3ODv4GOExtWSkMMUatP1zFBbP5ZRGvrXprEVZu/J3UQ0nsCemuLNlU
saY9+yjvmxm9FzyzNG7MvOBppnYXZRNmwh7sYYaSMBCbLuKDSs4AxYfLIB+CUJMzv7cL+u0fsjB1
tW2rT9ux78fXaKA6yqhhcNBDEnYEOn+rB9bIlLnE870Qp0WlkMbVQhcvheumgvJF0/0Am4ZIWOcV
iA55oP85GsPxf0PMrkGxo+bGlwxhQrjczR07WNgHiEoOCoXwVKChlm0/iIxaJ+eZakXOntgrhEH3
2lj+bANveLstoFGIRICF3pvIJCpEXyxghrdtFz5LstK8Ala4WVE3ZjzW/cF+vLtpEh+a6F5gWsXz
tdzPOVqXfWVwldHSM+d2TnV4t06JZqwrzFYI5dnG+ATFoZzcGpCMgd55GZUlR83lXb2WNex5d1Ry
PJygbDXNxB3s97QO/81UivnL9J9ljZ9EHg3SNqBtq2wOf6xK7Gja+mKtKaD5xva8LjUI8kxa3jqY
2uA7Q3Cjfz23iJYPdiLn1D+zMc/5VkguHrBAchw4gCMpu64WQAyltYjcgSC242FdThtbnXtu2g4d
kMGNlLmK2sBZLyoziOm69/qjg7ZbVtHQi1cwaqx74dTvRhL8KnROCMCq9ziB8PypyFmKu/iRVyZo
yEaTxhgTxtewVwkvAD9xebQxL3uGlw8CcPY9JIqD66O26KWDl2YNToj7SzOvgSjCTG0HdbGM39/B
z3Hh7FbseNBgaMMqvifCLHt+YH8NaKHi741kylVKyl6vklZCTgR5DpG7dkv+QjeY0HjrvRApFKw2
sZarMyGXW2/A1Erc9LewAy1IPT5jhpw41oQ7+5g5fgibX02pr3vGVAqAkfNTb9HOaBfhH2u3v379
HVhja9MbTAIxFBWqRMGD5Twhip6EnzwwrMospFMVA5vHvIhSEdhlXI5eMibUBiS1usyeOgHZ8jqQ
bD1q3JmZDf1WRb9lSIcot9+he6u6oFRtVpS+eqYPvvhslBCvfmRQ9bU8xvAXL7nrr8puFgmOOzRt
Gt+we16og4sS9ILFjMv2nl3CWTie+tAKXsrvzUQgFgEAJKWXsK1+hTFJuur151EwJxwxtWGJdygo
25jA/zqLpQp3lMeZ1bua109/kYDNmZW/44xJBid4D/pKTkhMrZ7BaNqmrZ5OQ3dXRABd0NbEN7Nm
itNrErjK+L55TF0wMzrV80FuJqUymTtIeU74XBlpz231/YaLw07NsEPqgx/R8Flb3aLq4JYn9jQa
i3cZpSfWtTvfF0VD9JmFVDOIh7KN5QkHCOEdEgQBWbFQjt2WlknzXVZvBg/P/nFC8YfZjhGMakf0
FkSAdwpJpLyY4zYxatZsyFV5qUtMUTRU7kYEAAO5Im6qdYRaF4QcyhGI5LLEUn3E7hLJGpPcx/wu
i+HgManeZtpmO3KjoQ3cE5LIjREWa6NAj7u6WOBKI7DH4EM1+YSg4LNZey8csq48QlOuQ+AJ9KRu
AZt18Wc91Su/jH9yFgLdU0cunyLNg+Ozzvc1cCe/M/1WdPaSm1CSDZFnIsul0XJk9I8cMXeBgvlc
Nl6pRTuCX9dA3IrYA7D54z0zqEMQFaV1HZYWkve9XeE9HpvIXhH24dZx2ssRoBJShmSui3xmmPYP
EtduTJ/KNfsGVTldzRIDK4ZSQoShRWDOIPwQsPbRKKFvcbZoe2Sa1BYZpfuUCebcaf7XTTKXdaWP
pP6/f+hmi84rTlUXOfSQvOzwmnSiyrf0s81mEK0q30LFChveeDfexTo0gqm3AeYGhMiFfcUbqnAV
eyBIfv00oB6sI8Bbd/6B2mjMV0xONvPDyL9jt3+0NtVR7k3zGlD33p0w16OYPEH6T662q4fQwB3Z
mO859vocPbA0q3RpEUTCrx5yF0Ck6OimhJeodK3ijM/SvrY/jBP5KshZ7NizpiXA26/cTzW+cBTd
qKA0nrftVRNhNk96b5NYz5ht0CpYE68r7JP8t/hn+l/Dk+UGUNwPgMHJrT7bS55nvIDloLKsKpP1
/VAHgEcPbyS9x0dY95xPIUQCOTgWKRUrkCAlkRSxu49RfXo/fn6WhlBjA/UYbfYRZdiQU/rVAvZV
PDSVLD/g/SfBZkQOwmA82k9WGavCXcz8/M/j+KSxxHIUUiXrqbhOHBGWm9yAaqNQw0fNg/Y/e8jV
I6K7INGEVXhZMIeR/e3KtsRNce6aFbAa1g/HNDakJNDB5g1S7qGwVHWRSrAOlnY1kKyzBRQJ570y
rQAn5LxgRnZe42JNJGD4r9Edx3iTZmAHWQxj9yTaOv04Bk6httydIRLsmuL1mD0qlfvoz+Hp2yVP
UM2h5S/C++0UjXxZ/+6gEJWMxz/tej6eK0lcJiat/1ZkBOaqp3gIwSfe7c5aU79lTY5bLqHlQuUL
fz4lsHGUh8L8XL0OCArkcqyoj6004g3gNll2c/XFUYlTliDSzBemh24tFQ2x41GaZJSaRiA6M3DE
Xiakgsnd6vWsMdXVJb9S6hgeW1swfSBlS1neIQORwr4HvXIxYx3td5Xixa0gIivcFhSxl2jiSnBB
w3RggeRfb27d99X9HEEGtLTGE0JCida10pVnho3iSuHzUdHjj+OY3GzKKzZSreyyJ4VUaG3g1gWz
+tTIbiYwVbNzM8/mW31Swkat6OJEoMp2sqFUPA6ZpgZQqyeJYBJmmLpUJ08ojCIbMQJYffZt7upJ
nSqRT9gkkpCpv3wlvsMCFcaXYl9MRXsWhpg/YkaQiGCEtX4pG+03hkbOwdgGGI2IhqR4dEEmPGNL
KxN9rBftGty6rjyA3/jGTSpYJJpuN0ixR3tra0v2Xk42g/NLbB/LE0aR/kAfFb60WAF+EoCEyltz
TMLtIjPEQam59N1OVkb4rTx6dSf/sCsv6tdVZNnATydX5I448st25a7T5BtOfyAlhDZSrfD6bhl1
AXgtWS03cQW256LbCKWZ3jidxfGr2Kdpa5hA08OCWCwfJyhM1hSiXH0PAg1euhLXvMImz+JNumtF
pD+u8yXZpYwQyrsx+8i62eOMenYNf/onhIlMZxlcXN5KrmIQGU6sT2xxAyZSXQEF3ExbzPiFHWbs
CAVAktI3Y3RUNmzZXZwSTw7qgcIm937Vha8/KdrEf631fiVh0TBShVCA7V/t92yPrrpYbrPMO08V
nIKIzGqtxQJD1vRnzBztD0iyZVEmIEw9TWWYRcCZeEtey7LHUTGKP6KMG6x8NJ3wM5jvy9VssL+9
Ik7wTvYUsvx0+8TSjosG34Mwsrn98Vz309QCarFFBpqgsOk1AKoYeaBdQcee3x/BDeSmUBp6zEKF
RyTASm9egiJtEEOUuerOooPnChF4sQWqhOc4hirLh/PcBbY+sQ6cU1hGYLLqFpruNWGScjUyX6FQ
KJfi+MnlBt5xBRzwoZ1PADGpAHTcZQH6vEvG9hxRYWhFDIawY5UYrppOV+W7vRRLQngNegQhxRDr
PK8Z+74LpKTcss/AUUku1F/vnxV3yQVSV1Lmige4WYfc6nImEPGXKqABieFsxEYXtYpDY2K01D+3
U0y+EBOoXaLaF+mdLpoHXTDhk2km/bwK4cyCRJFkyQw7pIQshpYmVsYAj4Vlxsg8UJTSM0FCKheD
sIAthsCque24cNSZidVYQf1lsIKWWZP6fVE5uSoh4HW9E2OZovRAY+Z0v27FiHZLLeXN47jdqPuV
iipJLtr/2D2hzMSR1zQhJ2X8obDGAENtfWsXYur9/ozlprab6G52+BfXLKOpnVA2jdT/ASYphq7u
bk0xFgsTh9xwSG2R3I9Upsc5d71txHO+VzXOG0ZnA5rBPzOpSJBTSFnSzq74dBhpV7D6bCRbrWAE
RQPPbrtUoJR3NMPvbGOs3UC2r6PML3fm3/a/QE1WpbPQGcvR/j1Gdk5eHt6iF2qMM4PBhzwIGxFD
91q3eLIBeJIQcB/wX3w1k9/8CML+3ov3UZO4mhPYPzNEYqjcaf0eST/Z2juL9Hg3DCjkB6tjUR0c
Tur38QHPl+K6Tj+DemM1W9pB8msEhiD3ytkcDf0rOtAutjlKLFJF+Cg8Ijjluonirc6KntztE6A3
56Q9r8iViQVvwDuFOZKeCuX0S29XpgtJwfDGuDaSR3iFGvTI9tLxa8guWLtGoVsryS+W/JPWAkdy
ond3Sd5lCid5d39oV3C4HxJMLvDyXVrSh5MstnR9k3hUWaw/tW3/+uOIXWYsjgfqDMzgo5eG3mAt
eWJnbKvaV098Hjznhsxns/OA0A7zagljg94IfMFfc6zNT6otXaqXBanASJrMb8td6E3ZPYnpLmxY
1/GXzdz0J2D6NR5h5QDL7ashxCi3zUZrG7YDRMqcbm+6L98fOCrNfV1IYRqv3+CSnUVJJYCh9v+Q
HK3F9AMN2ZM2obddNoiu0potUIb/4K8cDbYZFMR7r6mNIllSyQrX3UkFl4DqgA64XWdK80+Jmvlv
zQ/nDbNoL8ShRSNArJUF+HXqAYBtTEjTyFLWeD0mXcaDsA8U9FDT9execYfMz5C/xwuJPXtapVKQ
R3rlGq2435eibeSb4dEaNYDxuN3M2NaTuaTuNIy9wUElAnIAXSQ1KLiQ/dVjoiwePr0azgPGMd+F
Wx9fqNftlIxw3J1BUt4rpBjP7Qv4by10r2cnqlgaWa30ZMTWRkNTqYe5/3gRfJVr7gVYgzGoPQ2d
HuAua7yfBFpkGkg7qXbIhUVnvkTM/O60C1WX2T3uiNcXGCN1YRFLzZA6h7u0Gk6S9xTHBkZpalBV
NyFqSRWfLm03EuwN/nr3XN/IotxPzGc+7HmeugHs5za3fXTfBoGdcx0hjf4CVNwbo44xcwAymXpM
SCV5UENNvJDxNWUzdQBkvYX4gTIz/rhF+CBI5Dz6vsF2kKP0kJUuVyVo4ueN6HplP6YHXVqQ2gu1
Rd5d8tsApXZI4Fya3Yy4N72byWGBqpA+D4nGm6Gl0a6qOpfspy0uyegieL0RduKaFx2/TBz/LFMa
ub21NwK7lLDy/PIsE0aRGacsz88Ejogxp+SZsexmQMgCM0AW67ggJP098HuSNgL/MIxdR4PKhTf1
6ZK9qaXy2C1S3kXZS/VsWQwgTppyRJr3XJG9xetRx+A+6AzirQWGHTDOyPm2TxUkAi6PYVLl0J40
N49gc3ReF2+R/GqR91jkyCQojhx4dU4sK/DWNfDhCX4hLqfgpp8EGh6IVdmgSvVTt0x+1UESV66r
3BOQBka0yRnZ4hWHbI42K4YIX5xrWl7FjonY/qkTPdfDK2F1FVF7aP+6hayjq7cxyAW9NDJ7C1Hs
q1ZgqOTFbgekGGvqMvgniVh1knoAoi5/rO5BUPUVQ6KxYfJZx/xw1fCBWCMV0ZuSeRFYU0bteKKe
bzZMYiRq3NvSWlsfoClO7HSDrZMF8WaM9wLGIdoYn1jydaqkE+fUwd8eVvmBHfADxfi5GJPC/i9W
nYbWKN9PyvxypPLd74ScTcAWRsB8ypX9MS4ANO5BPAk9iMJ2ccKpzzn+BeaBNz/u+NFPTixDt1vP
C1c+40SFhNjd1CVZdt5pv6kkj2SxYMtxhesrFCyUcJXtXr9zQ7zHjASH18RIMLMgyjMVHyrc4aR5
ufGJjGV/c/LVEFq5WtFehY2GdJNgDF2HeG4uQ07AGTxoHLROaR3nDlQgawN8q4iCGR01axKmUE+C
GEzETP2ykRvlamm/AEcEJanuo5eNdrTA2m96auqGjXlIrls4djgeXRc8t7AmTy5oCT40C/K3M1bZ
044Bx65h3BvUyq/oRSkOrT4uSjziTGZwT0keox3W8y0e65Odpu1rNH7kXKpJbGX5sF9aXY5EYV6k
UPUkevB6PAC2mNh7khqEGtZwjS0/Afh5IUg4BnzEihJBxzi5U6ysAkXCsfdbN9ypi/e5ZDnhZ3Vb
Dku/ez06igDGv/xWQsN+SRIJ5ERWRf1//2NrI6qeFGZXO3jzoa91ALgzUYiA9YO9nfcirpiHjU/v
aLOVFi7yiDNMk03dh//DuHWFqvgTDRSqSrTa1wjzOdstSxFMT9IzORZrEZLsluYxjNJvjdJPp9Np
R/u0+lDS2/ityUx93tDqdbLyq7UbVSH91HACNimuHI4kmUVWHgPaiE9W3/mfnkxkKTTQSshr2jCQ
m7k2Xutoqt4yvbfeaWPuM97mHd0FIlKCLbKR6R/dzUbROUDydJoRi3Ay5UOy8uDrYyBIBG6uHYkT
U7wUBHt2764fRXD1lwfgZMlPt4f4/IfeqvNEgyXl38Ec+ZiDSXiUNTAUorz0GB4lo33UtM+cEYp7
NewQk3w1krpyY5ZrBeSejCECE+2hwez0WghYJCJMY7frmTTbDnk4c1djEuxlDQFCOSlLXQMKZoPN
X5PnPwnRsha/N7a6nHkhkrI78Y8Wld5fnLIX+bTGIc729dSt+1v3D7gtpo04/zk9VhgemBnAvSM6
xVFLCbIaDil5S6wy03H1T13BCj13Ev6UHlynyFZQBcZbp1QMiMOtN85NDqEvZc4yrYpLLRUVGTaf
srLnzJitGQFADCJYWIFg+mvCigNAUgNJigHA7ZR3NnSOUxITM4xv8c4cn2GceKxUo//+30sEn22e
2vKgIawlABkdkKQusGY53nrTNHUAu8tJP6vh67dRlE5AtlByA4IFIzCSI5zqk30HWuoLPlPDL4SK
yL/p5cQFMbQK+54gh9Ca8NomO6re564QgZ3tT/A81arKaku7VO7xQzsYfPHjBe/0IsxqzZWpA1bd
WUuNDCv1Uxb4Hu/1MSAt77TU63GmEkAKCiMiyrK2uahVHlXWM8eyPmDyHYmIzPN5Mgyfts5v08yD
vrvUk0EocvBf8z8OnYf1T2RsOYNTfl17LrKdQJ+2lJyX3+cWXrt13FDLnNIJTqU4DWq9Exvlfb2k
+DKUyEIrDPYOm4YDxJxwpHpJTfNjixU4OEUm6BzZALXB5J6AZM8sQLlP+kpITililRyGQyNGJRN5
Tkg5sLc+yIWg3/LBMl+kx//dQFGWT903W5IAK3w+yhAcBjkjM7Z//70z3JoSNvtq0XoLu/3chCTN
4z42ibfkNml43greBvf3ALOXtZuhT09iRDt9Se7jeAyFVi7UBEef2Imt09WC2fJkkW3+st/pCLUb
TRpCdJkDgfA7qgtvAIVZrFQO6oEqr+NIOJdhfTBYjG1qFGDApa7doCpgMEmRM27R/k6F7CMXqv1P
ILSaddjGtGovf/BoHl2I9WZuxSsHpbSo2vHxBot2qhoCjpli6+7pMFxgHbFAWU5RXpUN2gDxhKXB
TOUFX7VTdcUt9dYDAmLKWJupKbs9GFzukGNlnYvVLeQBZa2K8idCou5Pvf5wL0xm9lI/rvIdORMZ
IuzM6FFtFwRPzLyxYyuRrI7RgK9domf4m5oDGn4269SqAoIryY5MC6nNBFwu7ibYPl7urr7FxbHe
hnZDuuYuVmBRiUf/A/Ma2bXgMa6ZHYrEnjWSmv9Ebo/aO5425A8JWwMEFFMB+70ne/lkF/+ZQJRQ
pnGF8ZCBwlPe59bZ/sQaI9lmEYJ53OGpJl7fnl/UkZPe9xN11hSyVJ1mGghdb/lo6NK2TUyERHQf
6YK+dYLC1/KhUCdThwNcWUBILKXAnVA4D4VJYGAOshU1BAMfNOvMJooJjWtZ8hy/fHjYXD4l92Uv
/wPzPjTNMpoMZ0NNGORb4BXfngefIDg59goNzq7Vy8P9SrY8roC0rjAAl84RgO3HvgHOz5X3Xhz8
vV3srKmWF2QyBUuikqtaka+atWf/kVsASjSw0Lumjx/zi3QzqaTePCDysIzF+Osa9gXdIMrGfmA5
hn4ya7jBiInVWnASBO2naKC9lUxL+gXlCzXL8lYTJ7QvwoOL1/rlrct5QjJSI1L8FTQ90qYJIqUa
bQmsDv4ApWckM3cQYdQDnGcG52V8kXtMoFRdxZs9azrpnSvhd6ImY1BBm6RXFz62ZfMqHaZFHSOZ
fTLJap/Q9Rx26MMAOILhcv7gdFzNxFRVmrFJxlxX+6noqQTYJY9+a18ZmEwmcuqnf1lyDQz5G/FP
TGiLTLHkVEyPY/lpplir76cP0qWfJbwp1/YPNAe+Jl+pdqRQVwSeDTul/2TiyoooAaCmzkhtUX0b
DiNkg/XRotSWpKi/F774tO2PLzRIm4dPVmucFSTna65znrdMd+sloy9iulJnPbLnO/6kPiBFxNgy
GUmerIxZsoEyJgE61QkBMac5ItcD/C3ypn4dcTKbQI0mG+CthAEE+YCzmgaGn3eHit37Mq7v65/A
53AGxrKrI1ScVRCHJ+krz2QaxwRtdMzCX9RFFxNRjGX90QcTbiB2x4kUbelJj8/eJ0nNGsOGXPlM
CCCdYmVmETTM/jzPOut0kuI2S2O2cwIDCbkUmSpXpsA0wGp53+kU3YQUlWswWxZUorbqnbXJfEOV
hvife+AEQQlPnrNm/AK6BewCWJOutwoaFXVgwcVH0h5DcaRl947RxHSNkDVdb65LdgvyjBzb16SE
K7G065kDpZoCs7j2cEuLrSUJPnMHRnl1CaCRjHE+n0YXyHJhka9Z7X52l87U89J1vckFnlypgtW4
ApY6OHPzW840JvRvE7f1f8LRna5KaJ2s8QBRPb7bd5ICOLaQEMv+QcMCNg5CYlX8mOzdl9vFYTC6
cPOgiXht2LyXJ/qO5Tpccy+5EPgUU61H/egkpTOR8rVH42CAY8A9P51SonedijsK//Upw7w0xbAO
MnNgIgKvBDjx4CeBGfYKyPIx50a644oBLQZTKtQaDt8dtJUjFIQLsm2jKefo67p1GyIl0JjawKCr
/MI4LLhdkiOjTeQHz40dqt9J07ZepZZs4dntiDoTWCvm15/7EG/run4aYVnUxRqofJU94rVIo759
mQTNMWW+T+A19PfUJGz3m/GfcYA2OXYG7JsTQtx1fck/klmPb9MJX07EinlgzscCjtzU5vggjF02
21pm49+4n7xXyfNes9l9JZw3XKI6yccA2QKJqBmEh70Z+7hvQwjZsmgU4FskRLjsiEfvORZcc+bQ
P99g1qfU9Re1266z/5jFOEbemTscJQByaP1h6W8jAdtctrlxo/j70nDihkGPH3Kn6bcs0CF6G3Us
by/3YtqDT3npnduAPY8wgM+eRUQ5dECtQc80NliM177O4T6XFMy+jsVYMgzPjA/l442jgcdpW3Yo
n9ss9RoylF74pwJnaS9GvM7R9l8H0EWCaV3fmeSpb+KaOjE+vnkhdXhc12z5phcxtCSksSTDkDLA
SqL1pt+kQi/Hc0Ca1g1lfv655dvR4VmsZ7qPimke7ZWkJXlPw6aAL+JVJV/N6vmV8tmI67IqeF7V
3PZpva8I7H7rLZcGdBGx0pYHiULRZF/KtT+ns6oV0DAwfo2k7D/41rdg8s0WpC3vVE7EPPrFmvsH
axXmO6s+Oem7bcrU2TpxTep0WeTrDVv5HFAXjIvm36Vm/3I2hMTHEI4frw2pDFqonnpWUV6f2gey
OLacku/6ieiwy7GA4tuP/qfxEN+M17ZF11RU7I9qL2H3Ze2av2LRLuO0vm+5aD1qe7hdJakrLhyx
yNmOnxi0nsw//77Lg7/8Vrc9MqlYdn/irThmEwt85fFc514HlxAiipuoEDpz6+42ml4+u4K8nwMu
qFi0u2V3hIKM3jgODbe5IqM3rzg30p+++B5VGm89/nJaqKbIwPGztnFP0UTROr9LeNF5Bs9+6+Nq
UqTNzE+JcVGWfCXCoY0WKd3o+9q/EgFT1m+PCgAakjODAz7HJDnckW/6bh3LWpo4gisyS73NP1jX
h7oE/phiy3rtJmewD8HAbvpbsOsOT2YEtvj5tKjClYqG0OJoK206xF3P469UjUXyfqzuoNkTWB/l
webZxCbUNjk7gw/LBOauwsNZjc7QRwf2u1QRJCVC8p7r/5TJsPhxppC+LvdZ3HTL7gJOXuy30TbO
JpUXDHQ7xzWDNg24gSb1AGKCsubvE1MjsPlffrWyqiLQlqNEeKqS2DjGt2rA3B2fxxACJc/7t60m
eES2et6yPFs6rlrinuqC2dK63vy/PuEfjv/PvCooy1lKCOcIvvXClPK4WjR8MLeZGiICrReYbpUz
yJZkAKxttnbI3hIg/wJmr9oOBym5GYWlc6Cox+ZVm+wNsLLV3gZjJS8NgC0pZY7wRBMQX/hrLLWH
8fkHcmgp3bYUThV9wLMl6gth1/DUKcLNNgEkv0eqEzNcCjOCsQL2LFj9sGVoq7GP6Ai00sBE+LFv
fywbhFU3OWq3Hww9zc9D0FDkLkeh8Yvpk9wiriY4wwXr5A79BmLrMvMk7AP9h23lNj8IStfw3a2u
IlR/9/OkFIgPJuc8VEhnvy+8RuzbNvDxFauKfoxdTN91YFFHS1QydeIZTc14oQhM76KKXePuuiyn
Nyx8MMlMm4BJCZZtnVXQ0+3F6YtZCdctlP5ZR6R4nO8FUKt+QH85rAv+ZSNDNhY3nfCkM4u1E9jl
86KKpaYrxdFe+y1/a7YSCmWFtOMLfetgDoO3FYm4PQbDKXMeo38I0EbM9CNu+A4o1807Ah0GbBt9
JzceHvJqoCmXf/JZgFWMv5il5rb78ZH4ForjfeB76vXhd4cxXNep8/d6HKq1UOHjcust1EFvfi1E
qgaBhAREEYAGm/4YUzehkEy8pNtfUiDNxJaSUk+J0oRe14WVnV57ML6eMvnflv6tjKJpIAoJMqcR
XZAKa3cP2eKKdou2xutnuirtaVD3bWY9i11qQiAfCzGXlDP7OpHCXcihZco/jsu2dzVtV2BZSt9v
GR43Z6aaHoG/NWltLMsT2Dup2JJdhrarVlpYtS7895aV///Lq/nMRflE7U31fgLXYBM8EcYErTcc
WdlxLQrfyAvW/zk4iGxLCruLh+k/bhjnJ1ofcd/EYnf8TY8MsO0x0jnhZbGEIZ0ETrg880SG9Va3
h1dqn0yBGWhOD5U9cee8kzP/zdlcRoM6lj+qvUS3Z7K3gBQd92ZTo0f34JkUj5SpOKc/ouB/nVDu
kKuHDkUHGE29oNJSo7OsDYnPoSa2nLQTfF7weS3BGfXt4cW9+6OujHZk8YZps91QN5knTaVISLo4
oCyCDKhbkvpdnn4WLgOJb8/Vx/3XGc5etBmqtChK6lSuKFsdgKZ1/DtkzmSUThVMjgq0U/wOGZIY
iBCs9zJ/O1rQ12SgjoJFYDgcTHyXYHjgibaW+CJVgIgCftN74yygGffHSv2FRV02JFBHJANvz+dl
y2cpaMLjmsIlhVK4tzuu1H1LGyO3QeqxUcP4eVNYj4cIFx8YCJyzzW2WmgdQNBp3KPFKAWk9S7xe
HA4k1guv7vA/mnwwAGa9w2O5vN/+gO9z4iFDD6en2RB56XKy7h0ZmODo5+ws452SpcMGZneqydgF
8H1vvc7hInv6RRWlnRIEF0B+LxmwrekfRbReZwx20KYTJbzqKVoCqfuyvE3afdBZ3bG6nY+8Kljr
3d1KHDqKfWGJFeM0GBjmau/h6a9+x/VBODLo+WlW7/DOghxYKA77JJRRGzBT4liWZvVmwzSQKeNd
VFlJ2Al8HyRE+jse3qX2+fMkPj9jE6ZLzRqmAHpmjwF/xUS8hlIEnZhGhdVbE85oAQ85NUB0Myos
7jWMoAKtgfxZdXw0Kan96OcIu/0lvPFtxw/qlI0BomIyhPYdWi4gvvn/dVwsw4CdCqZpJRQqvo6t
JpIj9XmonVj4PdSX2aqbw96JI0OHUX9UAJkASGTunWNMJBrci84fc1aW2TNcTIO9YW4ihJPAZlWe
VetqCAGrdzx/zgVyBFspVRglNM5GwMP57QUqKxcNcX2mSLuIv/Ol53rB8vjJ3vBAczn6fsU3VyY0
tLN68DyQCMBmuXTD0pBSbi4sldmfeKfGqhTbYcYoo+gdvX39pFRSKq49Q7HG2hxZzzl6siCQMk5C
s01zhnymVKW2dTiDL95y55Uz7yAilFxP4lLgoJoAsmwtdtiUkZVOuj1LF1ST81JOf58BZucfGjPt
KYie+qEZPLPa7YJixBK7tX4Yh3LJyfYIEtXuoK8R+mSEAWLcMlCvr1sejTQWIAANgJobq28l2h73
pj2hu5R+8SrrKhcwQ2sWrJmPYQpXloXlxKmbBDjFHMHoDastjfLPr2yCdjyKigJB6HzKdl9PRViZ
fzQk88j6thNAwKveO1er+VjrpXGaHNw7Ydb0/tUI0zWT/HunBR78WTdh8A2ww92n4T7NP3ejYnrs
ILA0vPy4at1+WXLd4KljyNenCM6TX14+mqFHkKMBuJ/IdmaK0v/dLB+r18M9hSBw+uoIBOktTmWj
PrGozkemwUwLsVgc8AKI+kqVV/HGEdm3sEv2Qk8Amxr5XtcOyFkbc/jK4/zyOqr4/T38yJgcgw8a
qBNYnS/tjABQa6DBT2lVH0Xf9b2bV3A4NtO3uAwXGmqrj9ZCbCoBizeX0pBTui4hEqaY8SyLx0/O
ZiJDJDa5vZfS7Yfbeishw988wSivk1rJkwOf2iwPLuCxJWOsQrUcfCMsgklO19Ky16Tfj0aHFfi3
SZVDsyOKLgNUu9oSC/2mk9RcDmUpLuM3fl6+D5mwNUxo3CJpf6v7yM5vzAuLVIbGgcUYlctP8Lg+
VJHXXwfYm6yOdNB2ltVbVm3LAdAzEcCCqhIXT//ppAu0yjxvnpvFEh4yh17kWXxWKAKXl++nUEMG
Ea+aRhtGN8ZeYLb42Wj8pwRbnRqfuAbdqjZRLwmZK9qd16KRdDM2zd4nLfHf1mysvmMy4RWz6Dmg
yI5JDzHSSRbk46rXhOZMHeF50GazHdDAcjcPPD6Gs5ff2i2CO5NR9C1jyqSsuMkfdbUuWP4xg9VU
a6iBLocusTB9kRDqQ6S9LM/Z565xIm+ZnfdDxxUITUOr4HqIXd7Pme6LqjniqbjYZmFzJtPzh8p6
VpsUDw8yLi491kMZsu120anRkjT0RvWDQnWJM20sJseBeCE9lzj5X3dBHzex6A0Be3Tm7KfKoYsl
W05WeoqcKZun6dPrZcPAk5KB7OnGbvhOGAF5C3bwTHl8du3OmsV8RbAQ2j/mHfWxHyOyw7W1uYbG
1w5hQ2IElmWK344IgFTxNht5dcEC39vKF6BdFGrYKMb8mYJzHQS5PNqnqJnZHyIP6+zGEHU4Gk+a
hhJ0W9Spg95+/6RFWKQIyPvaK14VVZKe077gFWESYQ/vopLO0Zf7e5W+58VXU6vladILKAL/EpBU
Vs/PnxVBW+MPgEjlNqd8eLsPzUXzAeHo/cG0//xV14dyA8sDuv0pSa2JXcscDkx6YK9BVklAtQe/
N/W1ISCX57o5tGCDOMCG7uRtqTIDHe0NWuUsTsn4uQ0rs5oFF008/toCDAfIdcvxmIOWnNp1h9qE
hX9WGd+u6AOydH1yUzg1zL5gnSTyGB2QQXmP6BYjfiHCRLYMQZSB/fpDhDLh/Qa008JMqyVETn8q
fL1xvFRRCey0ZwR5SSzKCdsEDkXGssOGto7mostJ4NZVbkWDRZxmMGmft6OWoHHWN24Q12FLEpK8
ZsPS4HpMWHoqtWlVaZNigV2gJ5dAacnMR5DFeArdzeDnKw5+and1e/LA25HQ1Mn4CzuJPR4kAWsQ
rgNTY4RXtE/jDz3kyD6sNOtx29TgO71s6K0ZwHCdtsFHCo3el6usaAUJ7f0ETGwHJvJaJTD4F53/
gj9QTv5zYTqmLEjAFHvokW//3odVXyNq0OkSwbTw33hnzYmeBb7HgzTvGFxi58RrbEiijTocaKbF
4bR+3Y/4zC0Na1ElLzD5m6IX9slcNVOnKEACyK1metb0C7SXTHXHloFY5btR+YzoGZ7UzI9dOsH5
HKsTEQyPV/2Ao4my6XnOZiR+1C8e2o2JAl5giCA8ESi4Hxp3Xs6e+uH5Rs5ayf0nuFd2RUzWpyZE
m8uFkhyJGoPwLDKfz/d0/yI+b1SW+kEPu1flrgE3RemtxkeLHXdcxfBzJYJJ7hte6fUbe5eTnGjn
R+539N8lOLy/zugPdSRw1cjizRrsGIyovhxTvjbKZD8gaIyCsOS+E99FSXkdAJPWrRzAvl1qyG2V
pBDbGJJpWLO38SBNumHWVUVhZenm2zar4aB62JoA/SvRJJv6sMLNni3I92Pong8YRH7glY5Obc6j
A9dYilbr8vPzcoGMebQUYx/O5eRcZ6T1v/6V6GVpYPj/r8X75NjsVhFoUYZcfC9DGvhbVKVKN5Mv
nTQrJ5qyPWfCl21AaqQ/xYES7LOVsActl+pK7gIyweY6oQiyM0/zchjngdSANNip7KOSXsVJeY5O
B4wdb1nuKc55Lh/nww4vC8wXQBYl4f/RsW7VH/YduDMmDKtl411Ca2OMG69Cyn9oHGKsaLB8AmZu
TZV+yyNpR4lVy8e3MuFcVgxZ+MxVIBPQUmhxmSn323246u+MrIRW9EYro9tM2IMy9oDW1N+y5y9I
HuvfGbnp5CWdhT+sWHpAxBcMIkGPOlkEV5HGS137ztxFWY9HhIYNwgEsePCAD1dQyNm04O1yzjBY
rxLFXgdeFbeNbpsEKocI5gqfUpLAKMDcMAqnnT4kJVgT/POFBWhDJUeCa2cD2mJgBhy7BrjMfFoX
iErNf8IN1m94YpJvPeomc9HsLOEBSyQONfwcajnWo7jnaqw3XwVU357bnY3Xzup3Ue8wJy6c93aV
fLOk0z9YiVVukaOTdTykVkj9BU5U5Ue2DTRl89OdM5H/+5XzU+gCj+wrA/EOk963R/YLNbEdqyZV
Lh2bJdaOI0R5GDB+2oIH9o1MEUVTrxCJKVRZKRb0jMdZgzFyY0Prl/KckRjOHil9H9xGgJxGYN0c
aXi3wmwpUqTUAyPPpqQE6nmclgQ0yJmk9ve6DDRXlFBaWV7KtvZS+qwcaASoctY5SJspFLJjWLKM
uT4zv13gMMQuo2sNAw43tsQuUqrq1FyUroLs37oI8WZEh5tOE3pWfF0oaj7hXA8O6IGCVm36oVHr
5c9g1qp4+NNW/Kz7/bhsAeT4J2Phq3WfGrmnTaERipJP7DNsY2TGjmdvv0nZCMxljxB3wezgmODJ
4wSdIMZr5vh+c1POV52oqj6g58Mf9BlmhlXqEepEV7K77+yQ2yJIwYqUnkt8O6Ot/NiNbL2PVkAW
1iokPF7MgdFPNbMtmpM7aR91Eq71dt8YzMBMVEk8VCleHm9TFHFGEfNn7gHvrbGaEpkfVB9cK8cC
ARcErea08+6Zil7Z4F4nkzdR0V+Ku83grm1aw7R8WMf80ZLt3cP7vod8F72ZizrLgF1Hgwh8+FYz
AR7dZWO4A4+/bb14AJgKPnb0/qLlQEEwzxbgWUGp89fikTImTSyNm6N0q/CRlVD46so1G4/WTRji
StMhL1yoj5DZMzG55cLmwKUv9r4hh1ZCCEBGE93gOJyRAEUG4YtfnaeNw0OWJa8ctYR7Y1K9ieY5
ApVaWWDAB4a9qsHWNoifJGZOFNLp3Jko7yUT93c2sNq4nvHOzcCBSQRX4lKaJ1gY3oV41j/YP8M1
/zkH8Yw/Ygml11yuGYimAWrFxMtFxDr46e5AZ7aOm0PwabK+gNZsKuJ9J5HgR5kBtbrGAm1VblAa
K+RYP5jBR1Rkp//20vPtVra69lCDVC+1WJ0jILr8cy4V9D0VZQPDwvUl/wuuhDt7CC7shTttnFMW
GTTXQ+GLlicxPJjBxm5Jzj6H800hZnOE2Fu4OJ2cHkybDEVU8ecpyFs8w3kTMjWsy9jjNSQzNRWk
DYqWlFERe65Geyzh6y7fLMOdL5kXhPWUgHbGnGlpeTGFpE6Z8U2eZY0hBF0EuIxAhOAY7jTukx51
gnxIYEQeewOITCxV5MEhdn+WSPX9ECTWeH1//36cNEm1EjVNq35wXPEnA5Wv9yIRJKq2MsMu7KgZ
XsiQP6NOEOKhMnCwyzj/HSUmToyQep7+5TKL9xwfTF/u7H/NJ1P9srrZ2KM5lgGXB3P9Ayy7Bo7z
NjILoTmMS2lTgfQNY5ozdo4TAWB4y6T3FBcgd1TEOjqu2ntaih0lgORQKMg3PxVJwCzwq7vEOjIm
8dHI/aFlqlqzShE5V2YqHXu0xjFOaEpwQ2mQn2/gXkPgvfQ3WnS1HulR1sMaFtFtv5VHob+Y1NpW
T47QMCZXFm327NqIknsLiQOyzPcTyDvMJ3BMnvw0nFsmCfq1c6IUUUjIjDwdIaTO9bqoADLroOA2
lXiT0dEBw7VrHi4Js0bqCl82bPZ/KwQ2BxxGESjzEi6mHQRnf0id/MdKTCGIp48pHM3S9PYFqBJu
IPWMWQfKjy7HDLiX9WvVmKe3StUG4vJgL8xyS+/GUACFz+mNow/hqLe1lZruRP/NZ0UVt9IXafG2
aixKDDHhVCLEk1HxXcQ9f6CGVIfePcDQL7Og4+hrrUqbpolSLQLAT1ZHT305B0n+oE0Coe22/alh
/DpTHAwyOCXwPdQRYw6Ms0Hl63VvE2Y/B6Ec6X9H8PmHB1smvjGBLpeqmWpw92nDX5Pq5IFSPv45
+sb35AJb2Kksw+VMC14hRMmoAoaFudMdwf2zHyFhhjqAnTzSIee9UhMkNI90TbXlPYdDpBFrLD5o
o1YkeoxHT7oWD1uVNdDrqS9G3nGqBbCIVmS7Pkd0OLjdEnngrWT0iuxgCtpmicYKQrDd3QFdZgi9
KiRvlNK6A7roSjrT38qhSmIAgIu64AjhsPTVP5jLegSYUeLbYBw0ZSNqTOBUI/Obxj1GlPiUNVGm
+wxL/+yYuEUrLRFnv+FepyvfIWvn7X7YhdpetuU+7cYo5K8eTHrqZXwioZxl1gpJC0J+IWvDxuI2
i/wZziD6jK13Yo2j75fWswQb8hswVVgIjtpxK/sX+sG6js2t4huSsV/b6XD9Fdk8YJahIRjn58Va
fyCORudnGuezUTOaBX2/w8jD1p0y7rOZkXUxxsS4KygUI1i8vUZugRtXnTR+L3WOcz2MGUS3G4nh
fr53c8/r5Jqmeh0Pkyeyx6KitvALZXdjeIDztLDOj7kLywOdFhBkIV3rhARpHMO6y+firEUNyUnb
pa6LulY03dV9KvWB9TUhjLhGqrsk9vV4hI0LrAW2GrcHshICSQNpHGU1eakJheeAobgBi4aT2l7a
IpGO0mIeVR9vnY0wYCpzO+UVf9H1En5NhJa4ylynCAolsLl5gOmVrAv63aOxO3qVzEBWj+lh1BE0
KzB0jtVyOYgg5615g0ae+eGFcMkzj9DXlO3LkDItFv1FHr8iQKc1INCHcV40damctCx05T/te7CX
TlyZi2oRG0N+jwftNwFTweE+kdudGgdhIgV84zjXXIGuxkB15uqInv4ImKqDy8LX0nmjWegYE27Q
PNAwBaFm2UpZGJuLkk68U28dNkJgWvjK7h0kqH6+SsVeEq50srASpYvd75htqvEyLXzvlLwOQ2hh
AvXIVod+krOKCALzzMhIW04iYDwljAKxnMfFkYGEApSi2gpVAdgdGIbLUDmTAN1WywqXXaNCMYRA
2AMOddytsZH34sxYiIq5cJpF/dpTQx/COXoltd0F9m6kUIphB+0uJQfFIWIrpw36BdPPfKHqvK0W
dmcIvAWoE3rm7y0EfF1LDwgb/Zis03NG/wxDoXasKj/7dBi3SFJTMPpQ6Nb9dWRZqjL3i8oHCLFR
qG880vuzTY3Ka1uBqBBY06vYCT+lOANfQPzl3dhXPLnDGM8d7mR9EL9ZTfTXOOlSDbJetwPt7Cu7
vtJfvzseNk3Bk09b4Q5SU5KEt3YGjQ4cX3lPlP9xiMlhKoc1y+GHQb5fbGq2sgAEYEZJrBjO1L+B
Itc0noNT090C2JoCIM77Zvf+0m5li1Nv1fOyDjP5cRH37oDa/eP0drvmRpOvUFWiJfYq44ibHHfc
jy+T1roOeWCMus5Gghk2fsLJ0fZ39IMse+qDqOsmUFh/121WyFNcU8nNbNFkq6aiGSRO/OtfdnGG
pgGVJr+EfyXuIXbrVuPhT3M4Oyaq6aqkc8TALXSCFoKBLOeDdx2DtNvPlVuweIFx9HIlFYppg4My
JcDv6nVlDWqdQFJAQo4S9zQ/d/5SaO3w/yP8JgRfT83a42xFrkwYaPNpDztcW/CtNjeukHKRTszd
PSmVmIiBlpUMyDlvdD2AGEqP95hYGzguI7hQo4tiJ5kA8SVriDx6/6erTMwhZDGSDLaKD4aoC6TB
W7p+577UwyCID2jWHqrbLKYMm1KOyELgkIlk3UjlZboABFckpy5YVFeAjZAgsCXHywXtK6TDUWPs
dDApushpM43lqpi0l5a68IBKaMY6ffVMBdikhGAg1EKtCaDkkDGk0EA3aHOnqkhBqgHxp87Pu16P
a8z7iNPWERZz9BNMkeLXXU/SrrakUuOvFLmmuic+F9h61whQPFm3NXnHKNzxgPl1ikYwXChbnzNg
TEorLJ3GJBs+Oyhp6NLIs+KbZqODLRqk6BkjUEGQnf7OoMMSuNUhQExCyzKQnEgjpG/LRuMbMA5Q
EStaoiv/GnmJv8xer+PCbh3PBF7V4djhV1gQZYa6wKQqG3UcMyYx0YmFQ3MdoqKXU9pOAQoq1gV1
JcT+qjVqTmpcvwBjZw2QP126SUR9MFpk6iioY+MtfWL40XHtZJWwe+3LYzyjbmd0RQiI8AzGmqMD
3wDAaZi6hSzEQEaM8gpd1IVfJlx8x+wWcazh40bstn6j85s6ALLsaI3oxorLmYbzJOuv8QAQ9Mtb
Fl1K1A6EZ8xdCjmUVhSoJNpw7UM65FE1vD620dWOYA4AMc6dTVyFZnhpceRfAaSkVo1e0ruqcVKQ
8ckPiU7JcKz5ZvhWxm42Zquz7a2yxKEYm9Tcz216TpUGXnOJ5s7LmGr3w2AZIrsI0kqMtbI0kuR8
d++qhAeTkO7EbiP6s+0uKsnPw8k3fjO0H9e1nVCg5pGdt3xg7B8fdwte0mDzupWVaHh+zUU5boHV
NLYUEebSwsMJV5UpXV29E9mAz7Ny3MRItgi7oxYfQwe2c8VzbV3QHVVh1GojYMJs39pTmu5l221L
j903lxWyI/e5mElvEVS0PCHUZLxff377T6o9WlGmJAaqsAA4hiYl35vOPjziTypGvnuLl2Jv8OVW
VoVCPT2deN3N0WOeDOvpFtrsMSvbTEDN+/wuJx8ju88qEPsUZOCoVi2I5dyJNBAiWZDfbOeJN8uv
boI9XiEIp5SkCil8GnEvuO6bKF0WijokZ/PuK3PmsQKmEgUlwOyl6pk2pIHq3bp1LXMhbm6IhmXG
Y3QsNo8lb6IlEbsXohN9eRekxeU7tODc/x+hyk3/CN+neR/9FPpqAfxrF+zlcvEHRsDp8RoLrA7v
FkE3QVBT9sgcHGo5v0VmRGpKLSJNNk8AWsf9jDdVS8i4gQ5iPSStjETm3PnmGa2HNXJV5D2cljKZ
YwGF7MAWsUSX+g3MtMhOWNRZWOG3bixBw0Im2hkNKSChdPF8Fi+PbHs6QivATnPh0WvtkiwMIW10
2tN7dBI+N9rp+9/1VXut2SBX1lJwoAPwFPuFATh3zNcZzc4rX3qszm7x+9zkjNK7OGMEIpn/sQUc
iL02XAOQ8Wv7OuRpthgLpZW1LLZ4hB/6AimJOwVPtf09TaECRguWa9uM40ztMZ9VzmouK3H9oake
Gmjf3W/c6Qd+agEZiSFedWZXcC4LqVHtizh5Sf/iHHW6OdqX0azBOq/jKS/VOvhv4Ye0Eu2vaX0l
c6xKmbEwfrlJIFnVMDYiW81GMg89JjWMqXoJlRXLtgomkH/lPKRMkuRBtLU/F5WKwdzltin/aCxR
2wC2ccrZTMr/k1uXtVnAAyqIo0UwNy/ZqEop9FeQlD1jEtM/40JjV0M9F59QKdBcEWKzWz/QXbSO
tBlQezQCSz8C82TNSePInaV+MDgra9jRKesRVB544x6e5cInwHcPL7HQcQxBYzBZWP5RT7vDRCB+
wVRI04ljvau43uW7dcJe89Vpp7UUjfWeYnl+356HpiKsMvA6YI+I8WhRyTXTJQJXtsGhjoX5hmwX
jBGjFQnc0co2Pz+9m8rNnuG7jNXHfZE9wC0lSpgM5Hj7ebN8SaZkclKZj7grke40bBZiFyrzH4KH
s8DW20+7oQR+Ocycr6vNw404ECDLwub33j0Ts9SwnoSVm3dl5ozVYkGuIT5AUxeWWjToweg/BONh
XdCoIQX03WQzwwvc/5OXpEM3kHwYzHIG/CyGUKmNVw7idGtGT2y/MRZzv5btzEE0WIoUgmoe5sP5
UyuVDiOMeS3i2Wbnp0PYwfTzCTZJohd+zrkEucYjP5eOaSoFwA3f9uf7nP4xAn4dJSgZjfP60Gvj
iMz+Q15UMDJadbYBni07YTAhE4J517B44n1OBHAsPds71kxGQCSTNSCLW/7R16DIMm6Q0WwyyELw
mppyU9Uts79eOwJcXcdG7Zi7p+Z4RuIGV+sbM3jm8Wul1QHpprqAW6lqDfLsCfHM29riVvgVvX2Y
7dasKFpV/LzAXSPKM1bCwy8BOqMzh/K+mFz72dI297zPjMFl7qn0B83Y1Z1tmaPWQECTLlG+BeQa
LvgLMerkl6mBItMs56C2BwmfhRJc0tUlDgV9OuvUcYHdrF9MGAGrXMNdwAkG8vh/bsGUPKmUElP0
lgw8tQjQAf0DBa29O00Zt2Qspm6BlXT5WR43Jq/qYhadK7ovb3uN61SgnSgNqlEFnqOsoR2dTdT6
381APteNuBQkvkrrXiECXXN7OY2kGP3/g9SHiG2WGDgVLLqFDlzhKtjx9qVN5qXsdZgbA6lcD/TE
lrhJgMTA+RD6wWU5tD4f8lyskTS9gxxKbus7ICCweksCLxIX7G24BQ0081hObkzVrHZSd8fTnkkp
p1osC16O/KhxxUiMDS2p4O1Y/9vCcTsAHNijbp8an7WbO0oyE4G4UR/sBv58dN3yybWCBJsqFw52
DIJKip97E2V7u6JhZYHjdYWSGRIlYqCfIy6c87Qry8HbLdV+gNoFZD/g8wZgznKkRxNMF5QfooHi
qM/DBqwGcnyo95NOes14QOaxQaHrUZv/Bmb8YdWlbwPYKBk/mGBUspsGu3hoIZnwzA4U/umnVo4A
w2TsgEL+p+L56PEiamaz81oYKqFrV8ddz1DnvZTB/bhSch0KEla3tDkcBsv8yCfNrCX6hCJ8n1le
vsapwQ2hD1OwQA9R7YdL6ckdmS+zmHtPM5GRuTUkw3Er7Z2qAkP/bkqzpmYrHRfgWZlmIZKE9Ni7
RCNSiH2nvk2wx67d0sjFUpYPV4bRa7AZZkrtp7y1VaRrOiG3VWaap54AYPZbjVbNgiKi+wUN4v6T
LwM8tYMXltrvCSDJd6zfP4kY3dUbkGwRPgd97+CugaIUilq8Zi2+Bw1sFU7I7XAxQFE6Bxv5OD2x
ryHshdGhozkt6jef5ne2CyksIWNKaCsgPU9y7+sfUXxQ3oBj3poVrOT0VDH/43ARfeyMW5ctSxR6
9Yi3DTfMpxFp8x0CPar1Cz5mO5WmVOQeu3qJ7DKcnYhZNXC0mhQdjDTUdaMfM0cmaMNZfBoEnfHV
TN07AbY32UEIo0Bu/q2lerq01ju0+L2CScVfmmeBEY/qIh8bScXR/PH4VkL6hOXvDMNBsGPibjsl
+O1Q6e4j9kkdOfe28hzPd9RxIB9HbCVZG8sMrnKOuNXgWU5ovqot5ylwkbCxVROs2xYOLvmAKQJ2
Bc7iRAvuvlt2dOmJIeKoj12UqE5YJseWmBe4lQ1wg1ynEQHQZ0pe/Qe/A2PrxfjvhtZOyVflyYqo
1/BrBrUgunHwPKArx6GqVd3x5u+C9VI5QJrNfFLK1oJYy9ktIYBJoSlSvD23uU9eoUE8PdwlrL5X
LeIeLDwsQT12o3LIVHs0wy6S5IWEArqFpBtyVfErZj071UTcyVdDBQFbr3v5i9665CS3xL78V9se
qLFPqB+UjdoRrynjgxjAUrIsLU0xAsLom+3/mBgNfhj82IMynOBEaS8MmuprtxwLSuuG8itKDUsu
1yckHRn3pK38iSybIKk0/Wo1O8Sp60o0pZGKFYqYdcx7N10NYf1UJjwE8lKXYexwKyDpZJ8HnA3l
Mlis1Kax4PISr7dgJthrxLUTsb7OTgFwjp1A8/9shzitxnLllwQT2viMbaUGgfYz1N9bLbbVWZMw
FYHqia30yUEI01wgwO6cCGScZAfnmxKKWJZ1rd6rieV+2YwwyVSwCX/Qu1WObBrB6Ia+KxI7z08b
fLCUEtwsF+pnMqux/4QDChdVav2+8poBg+t8nT6Zn9H85YCCwOv+lE0hPotdyQ6lJ5fTf1yWStBX
Jd28kSJAShP2h4KHmMoyM929FGxQsg5Gd4imXaHnclDol+x9VRkqPIgC6H50xyHaw0F5q66aIe5D
02vV2iKWPocM/yuuE9/OgWwtyw3kn5ghzkOpLD7RKMGb8C5ODLsZ3mUBSCLm2JPyn8zjK3yDzoN8
Y7No5gsPK4tVdyOe8hVyBvjLCUS//x2x9F4UXve6+aeKiBNT2/m1V1/xGG6UFtFB/HY5DSyBo2e7
op7816Shj+fQg8qiA9lpJwvJq3/MWv30Hu5uTwCn0K8yTKpaEadUDJKG47rjA2k2kiU3ZKlGRbZA
x+5bxmPssYclxBL1VaQuHMK+SPYf9+LjNWpb8Oa5OlkBHujzbOhCv6xsn8z5zMQYNOmE5pk5InvY
3OwduDObCf3yfZdVK8xsO/R2TcIPKLFC921469H/FXC93UozKkTptVgNvMhfi7pUqzzWnvz4Gwkw
kxYw99ttLUxQpcPVIHOBqssbDsMWXl/vgOXm4MA4juu/ahY1gH4sRv74ySpMMoaAyjwVv1qRUJSX
vlTgoH6MNQzR3wwvxRGMtONIEoOvrqWPVSRR4xES4eKjdPY61BnvUBcvIV7DEHvutMWjB3P9Yeme
wL6ZZlR073X30nigQqptRZIrWTNH3ECJjHSWXrYLeUXmBDIikYy5kF5S20YPJ02oJ/XLeaLYEteV
QIBhL/mjTQ9QDlyA8SUH6z+1rMgxnC8ZoNWoUQdDxQVKItc6WvakPQiS8l/ui8AZG2xQKvgx0LFD
DhNTyDsz1WXKfr87kIJ0DeNnmJUgas+Bi0JxxApaLoJHLeO3KPaS4COpv/lee/hpz8zSDfMq5EDX
wj5hz+nJrko+X13y+ggx6XZFnvjG0rDR2qOtHZRfC5BfmSyKXMg4/kvvK6aE+vxtTT46+w/oGXmu
ubm4E7/ZsCjJzMspD3sTf9KPBtAH/fkAVqjVLvu1FxTKoWMvy3gK2kOKll+K9XES1Qy5OXPmFzcT
OtR3MOBivWWell1N69MMyzO/WLBb3X0Ar1IqMrIyVEZb1EFaYDFcOSorAIuAZY/MQc6gMXr15Z8Q
eZXNCFIlrSC5PxN+VbSZuB1YxCckwn/hytOC1wFjFgTgVDWxvaG4lNslxFuhkGf5BtBhvBfO7Rth
nEvm9RrXTvwjgWgT2gngBX8muPKa6Ijw5US1WPg2Un8SAkb4EBEH/y5r4joFKpmuN8/cz1tR6Hdd
j1JB3eq1IkgN7PIu9Rfq8osgor7gdXOLbw8sagYbbYrAcSR8D/rNxFjIAOC53YkmbeKCvVGCJF3y
hQab+Xa2HyZvnlQmIaeie3SdNCw+MtyobS0MsvlvGrL1qMcmEXIvewFQN+MOtIjvj9CUDsy6hWPR
16Li+91tpLM6KvSEB0rro2MH3/KL33PQAgfHTS1EipiujmCQmgCQWM3Qc5nxcYWKQiEyHu5vOEaH
XYkEBvzvI503StGDp+citDtXhUN8TghqQErjcU62DGxJCOASpB0qkU3j7VsvtDi4XNwj5SIWmytW
8w+yDilS9cpNEqKWSvp3W/eodpz7yWlA+GbC8FyMSC0LDTxO5suPvGkzyexJgmEjEkAssH8qECI2
DwpcPP4yEVrNUUqGDMfV20y1S7VoGhBOKjtITcdbiBn/VEmIb30oie/ewrfzHICAsoWtVMQUvsnP
3aFgwd8l2nqJwzJkV2ic4iqQ1fZ1ENaeKm4mkfVDmZFLzb3iu46wCZXiLkMbsiqs/yFRE5IsL6u+
Xc7DwgbPw0CT4COmp+QUctd6srGH9u5XTop6nv17IkPs4FDhceo7cq8l2CxRReJpZgPulcV6M6Kc
sFrti4jABvBIaHpNVu6eyd4t3y5OLl6G4HCmNHvc/YjHzLR+lJBn+OAp0rP1ChLYNzf8lwEAh1t9
KGx6VzwEYx/uCY2Zd2QShBrfTxraEXLo2vrFZiwTeh00LSgS1wCkmdqXoEfT/TlBten8uWCc4keL
dZ+tnicl8DEzdI96O+z9uqSX8BIBUpMqP948MNsiYZjCBj47QGfH0Rpbz2PiFJbNylcS5QTXiCqH
9ZXcyMcQzd4B5yWIzvcgvy27FbUW/QWZKrlSDq2w+IF9Bs7d5GoNhp4s3WioUZHD1e53obCNvR6R
7V3GkeMEoYLQac+vjyg+z/dfU6h2Q3ZP0VsDLhXEuN1SpVrwnhRPdbJUcxwq3ehIGDS5QRXhiqG8
oDi+b1D75UTXumlh7lLTFVS8Wh0aQ4/ERzqUwg/XrT9ABkZ8B7Xe1t6gzD581f+mjcJdlcWM7i0T
69ZIkZzPOKuymsRZRiyRJt49pmucs3rhYkptv2LpxPgMRpx6gLoB7Uk2bv/szn5fVlYhGdrtBGAz
5KJaKI3A6MaLls+CsDXW1Za05YHl5k/b2FaAU1Jezv6p27NrNeGk6K4Wesfp+AOaBTZgqM0V3VrY
DXDDZcmM2sCArNFgWN1JaWyACogtYD2Jgg04Nkj2zUq0Jvzo6aQ9DipcSJZcdDOBBkpeCM95X+0u
VIyVo6OexOn8alg92q0tTPxitBZbkcL/f8I9KzrFBZLXVE+Y6rnjWOfTVy1P3sKxlNUEi0LWI9L8
5uDDHM4TjbxYMIs4jkb1TGQ5jgFQk+qrRfGY4BCGtVajLFQn1JaPyZr8i95M8Kjf71ewD8iCwksL
186QsvkKwPtLvcuGONwY94P5lzYeUbMUkYPsqY5BfEqQo0Rk5VY71vUIYEPVYfHZytGmI47a7vo1
3X5W1tdnSAxFoPJdaia7oz6YIvkkZ58O0/TOqFZAizInwz5NjF0+d0oPDioVX5yc7EkYSgUZLUlz
IjZheHslc2KSNmUe6OSN02F4tVGyZ2qedkynu1dTRruVCcoeYmfCrx+stwdWJpyST7RnNNNOYCIy
3qJFPQSpb8cYGvvjgLbcpuc13aGR3JoTu8ZKX9vzKWOyxS9+m3hu4fQ9FEctEyfio0tlCwoFjgZX
Cof0XGOgMCy4q9/isgXT5i9qK6UElqo0o1eZGAl+VqoOXTOzaq2wxYL9/xv88yCZd9l1hljbCYmh
Qww0az6BuE9l9pjjo6NtcHgT1deuSdUhLAaUtQZOF9ANsDXevcMAlvV/5tqxi/BL8cXVKrmgd8Sd
PX9vi0XcxZYZEWSvx2rjrDG6yPygLtR4G0kjL39dhZjZvn3M571Cq+XClb0ytklma53ry1zLekWT
Or0KIeJVOTo2l2hP4/0dgy7DEeWQ95xvVDK5gaTkq8EvCBZAVSvLP2zW+/OfEIXY8cM42nK5Ez23
APxOrf5FUB1jaILes7Rivy4T6PdYrx+PfGn+FCrc3MFNCV9xuSXfQxxSxshqQeBYktILBCsav8U0
FZKZhW3RpFXdE89o0M0dBdIHB9Q7hbtlCOC5f9sICi/GBKCfb1PD8os21+lgS4IfE+WlWA8FLUaf
0eTJQj1/g/+lIQmzOW00jGus6ghqzPPWyYtXDsxaPPTL240gurf+LC+UJb60zqMss+TYulMoDlGS
Vl6TQNo2IyopN7/yRZL41+CdNN50sbZqoivMUP2bSslvxOuo06ZTZfH9JXtVe1P7yPPVkRY1YQEw
Ev9f6fuYXeEOjgrJQOciugtnAgo1cy/S0jm3aO08hf24lwcKXZlvdGc7S08VHtNQFHOjZvB1T7P/
pI6vuoKqFXB2/WibFkKCwnOraoh7W0JBpIe1fO0/KDfnBVqNMxYHoMAIwJ1jiJPsXjhewEIa2OGT
yH2omFsPRePLUFNtn9u1qX7h+YGDRuYrvMmBfRtKUvGoBCOwRjjzkbfDCl/BV9NlWZcchQBzjFKA
VS6lZKFwzsCa02PuTjOms0KYuTe/ANJ9xWxlTyJObIIP8gR+6J/LT1mYN/2jOhNP0gIU62s9jMia
6MIOQ+exaEywFhuYE7q97qNHo/wXF5caeuef4Wtv8MSZaGyAIZ3M/Uq5JM/DRRSLo0znI5VnSO8P
0RBH3MEcWhj4LTvpUaW+abJtiUrXN6RCuahMYzDwvSJoLeENnb3Y60OhITe193j2Y66fB6Ndlqj8
3tC2oI9XrsYvQzDziUIvUxOYgGmV4QpNeAXwumSOPzH1cCRziaJ9RMcMYA+78LDQmvBhuV0nsIRG
KAM/MGknYXIufof+cesDgj8Y/aaa6tW71lbusV63BHLNxrN5mBYAhzlC3DMJ/1vilV9cEhwhhyuk
8eXhr0FPLYGZoFmSjV4J4DStKb2bLBwat1e6sa9vsPgBFgqOPe9LjwXZMAMhysVjiNv7jo4oBB41
XaiOCBbmsQfSQmrRvd8s/cuz8pUvpB7ltrq+VWuwp/G9pZcp8riYklQDYWKS8JZXXeliRlRB1GGI
+EVI7gmMklVQGcSH7IunD3sbkFEt0gELA+/5H1vwZFrLUfzT9s7HuuNXnRvlFoaTBLZ8qoTxxbWH
dRhYRrIMwmR8jsbptnWM3uae5PXmcc6rhZCY5bAhrGSpvbyJKo8YKFFLG+qZreoelC2rUEkVhf+y
uoeJfS+cdLnwBvwkef3ImWs8m7KU1QmFe8V7oKOGdYcj0+4v3ZRDlp7U2Jy1AAKAJy+lIFowbTZv
XkSbAMUrieOFvo967lWJDJGwA8RBz7hl3T8hJEnHMwOspp4IfH7qiRM+nJam1ovtKcDQlHUqD/Zh
C2sgJe0HPbeyqW1wvF6XKBHLK+VIrQOP/epZz68oPCngrVDRthcexAMMWkLfFnMAYI/sdFwr0Ra2
ab5pCxCxe7KdWs8ee/jxzd+x3FI5twK5WJT2Y3ZJWSB90jsa6KCk1cuhdulBoAswiODhnb2/pc5Z
i61Dgb4M0Gv/N/hzzkrmn9ziujmm+25HgjneSS+nkGCFn1eLFV7D9vXoDGDi8plBxIojQjd6zhtT
KkJK+DhStfuEFzv9f4/e5V6hugdIGWtYeWnyLw8C6+7P78ry+uTo8O7W2O6xwi/mgTk5lpAGPtea
zd77ajU2VWKU+cXn1beM9L2kbwHp8n+rm5XhnHRST+sCLadWYzNE+uKX2TjyeXG3duBd/muBuXa/
ULHKsxepOg6A0r8AS3kEGnsJ3PhFt7XvbZqtdvzOqKjX+4QJ6ha2RY2/K/1jKTmAwbQr0FHIHzoX
LmUXwdcYbw5pHddYcHFIHQ/PL3+KtHtIOCcIjjuoVukskv9ViMJhVekXL2e29pvsSJ5i1thEq0qZ
6nhn8pxIeJ1Ul0eo+DORhYj/X2y+U18krvmtLl/u30q7sjt5H9qT0Dn6wS+2PFEIVcvTLy9AGreG
DpzulgJ8kAXSctO4kLEeAz+MXhzWmSrU6Uubuvs/v0GTd4Tu4/J/zF6QpjaLYu/I5pjYC1ylNAQz
rWUvRBxTXhWNzpinpInHdZNBT7mouRuiGn1loSQp16RpILt4kHW/OIOKd7lCmun3qZWejgQ/yQy6
keRfl8P3vJHXwLGvnDHcteMGRkUQx2PTTBF5NBbk3V5RD7wQ4UKF+ejzmAhwx7Yh2xMLSb3Rn6gs
mqHOEt/1IeGegks4BdSyKcVhWzDv7X6IeT5OiK8yPbBMA3kZEzU7CA3k5qFnOII3M0KU4uGqLm5D
iMWwTGU3jhS4IT6uz52X4DkF3zTtakwlI63jC8cIFNu9i2A3mgKEPM5FyZcQ3i1lV+VE7zTR3VAK
+EBFXpP6clCB+b3xFBfeJ7/vsJFU4blMd1xOcnC78TyTqfeosb+pttDBn8GaWLprPjqiX2OODSUs
UlykqMR2DYnnbRyBpJmm4yTsq0BXB6ZLWO/PSH8M6DKc+y1s68e4nq6YQXvCHn3vUxF0KaS2QqSw
kDoAwCSujCOR2c4gSgHSZ6G8dTzYBpCddj8Lumj9+orLEpIw05sTVjWBeYq10o73IzrlVWgNYnUw
cnrrUKYihQFDRDK9CfBGFEffAn2lkNNET7JLq/WALZ5OPKMsT7y89yXZ+iL10xo/ZyfG1dMSAuCC
EGI2hNOPAOKeJ1/Yf9axxm3BI4dI+PN1aqtOKTdUeQlwajB9APO8MRtavMysBkehhRxKyBfJlbGn
p2suwXiQsS/8QJ0tHjcjxEoTIjzcszb3Io21w5CquDQ5es24PQoffdHIvQERQLuqIEAUDFA5Yv7C
KHlzHw4lzEKEnQbCtR2IvG6V7BTIbhcVl0Eyykcq+nGorHJz/mWo83ShP9VUNS6fjNe7CQBoT2Cg
x7l3B8P+p9jaPRHZstSVMDz9cItMkL1P75w6llWcigwj8JUG7I88e4k0gFY1w8ZHNkQiFg3VID9u
qpF7nJ4GVvkM+ELDmP0xxSv/Ytikt3/xAqpjQN2wZ+/agV7LfNAr3XhQYsHvtRtmqSQBFhPgEUBA
VVWttsARDt4R3WyQnoI/KfNKKU01tpzrGcO0Gx+K5QWA7EJdynA/80VSaQXNSR6HQL2EBDjRnDXX
6KQ6qEHYEDp2KHmLviJ7VQ1YieZSgiiNVjgc5bwwJl6zgXp1AlRKa/LhPeRobg1mayeIG39KweNL
CaGJ9fYRe2tV6syX4m0kJPevXj/3dRUk5MfL1q4mUAdZSWbr3cxW40oN6+Lx27Fdx02/g8w3Xun/
rTLAQeE67XreZN8OH6tpsjur2nqhrZL5TkMS61F/xXplJjl1WqQf0eY7q2b1aAFxLZM1pJWfeEqx
6Nr8RQPDmkB6totzMI8e3BD7yc1AOwrAiU3yjtE8ecDVT17cCEDEtl19wycKOs1LitsPPB1sqkZy
fH/yCDrd80Uvmd8tCsSnh/vU9dsqpAljFdxM+M8UhGy1xpFSMFIyptP8zIWjiX2iW/aToD7EWZI3
xwkhNPiHtaTujhTP+QHAdaQ9Uxq4fd3p7VdgBJHFFtpgKGeZK2uhTrUqon1KFqVXODSxXVCOtrsx
xn6T/hB8eF+lNB05Z54vBH4kzfISF/u5IpZvlzie7jV4OAdiT6owxtKz9HVlKTRs/zt3D48jSBCu
bM9ynjXRWUEn/pLuLXqX6gAQ9WBCES6SCpWfIe5/B3cseqEZiJxnPot9p5SddYfaI6zZI3nozmZL
GFEWcx6q6MEJ+LpSo81D60s9HFz+eJmPafvusxwcBj5y9/D6lN16fIkF5SL+lLA9Yp1jtjJtSH9L
t5v2083n1ZA2kns8ywp/TvfvJ5fwTmX7QW3dw+bGHUOTNeGZBCqt+MRbUYy0L4638TKfo7K8tYyg
c5RYwPblPYKOKwZvjXGW9oGTmhJ6NE26WO+vx5jpQvG4VzSWRb0TXXUIjlYxWIIfKg7/PFvUa9ZX
xQriXYZmZatjfeIHtDaNyJj597nUkFQ5/Jl7v/IUabF3UwXFtXpgxmA4fVo7LCZB7lq1vyJlhClk
FnxaZ86JYTsO2dHcTMwakJpxnH52jwyPQLwxwvuAABzPJDvwc5m+xBxnEDLZlBXxaN5uYyj80uCV
RxwzWaCzHqiSAeFiYzPPewNnJGbxnkfjfxReEdkq1dDWh0XjWqqts6/U7OS9cE9m48NubeQyvTRM
wMGW2kRQWU5RQZAUocHoxwOR/SMTPgBcXinFt9YYZ+SOvA6rugtgD9rx5iJQOnIT+tFUtFIFrrZu
7/GmEhWVPdfZm2IgReUz9Pc4703un1nilJ++ucMQ6wCwWUQ2/xwXXOlRsbqai3IXLMa+gjRu7FtD
Ts//UFsyg9FxHSTR+RAIWNTAnJ+l/ghv613BiQ05DzI6aQ2jAYdq3KU+lrmFM8TRxnpRMqhdj2uE
bqcz0Kn2YMZrMauoMSAMX/CCIyvtXcD6hWh8tYxrw6Xi3nX3tDByUUUCyhK5Ed5A8Pi8B3knnUy5
ghHK3wUpG1bMq5OsKXa9Ig4ZM9QSfcr+Kvf8BUlLYOJcdnKdmEThvh16xHS6yWTYnHhGf2pI1el4
OGt242w98UYCFtUTEaAbyV7Ih0YYCGqGDEZadsZU3gd5bFeATRkB/HqyEc1Iy+ZkIEMFs/hxYwyT
F4EUrMhpU69tjUxvqjs3YBuGJPKsRmidcT1gDXsfcoEm2rMy/dPDLdREgar6aQfXAMZ92NkWKoO9
F90pK79lf0iuqqd6BRU2dhedaRrjp+Tf/4OLbVoNZ4aMACynZi4Pz3A5VxPFySDSRn9WTeScq3UN
K81MFW0ggdX/PtspOh6R+l8hS2njULzltClJNA4aflvT2NhJZ4ksa3T3h94zIKTusI7g82TAaOGI
M3HBxs8i7JseJVirWb+lYfzmOZ6AZG1EvdiHkXs3Aqxo+8mOAw7+zLIwuK6RqziYbIku3owYyu7F
7e5rlpz7fTo6eMAusGkelRb2x7w983uVKFJY4+2ir95+LW4YXiTvwryw2kD0UE7UW6AA233q5the
/cEGc7c5+dXuB4ezOBBQCK9bH1ww8X8SWIGS5JXA1dMYdXHnG/smW+JQDAUIxoJON09NMN2z2uua
Z6jWHFJzxHB5rpEfs/Dg4bmnUDrfbeLzJjzJQfATfebnmYAM48lYvrRiQxuomEgd+L3kAN6sNNgy
Z1GVrqVJNN2nxlQZnACwdUeTclwqlV2wx0ZlQI1o9Myx9BceYQfHugAog9D/2JWEiB7HiksD/6xd
/3JSwi1hSMixQY+W1Wv/ZzwZTJrQO3coSG+LPOEd4B5b5cmvwOLHPK2J5CsecqzA+sng71jw5DUh
sp1fxqEIHoR66vzN4lTq2sXPQ+P03pmXSyrX3EmKFfEMX0ynywv96CREchMFkoO2sRpius6EzYJ+
sfTrk/sm2yqWYpjSQfIbV8fMKFJ1IaoTzLZ/Io2BVW2RbMkzriNXlviFJ1u3e/OW98nQxUxou596
g5MEmzsQwb5c0DYVhqXEixTA0ImPP5/9nOejA9xfvb5obVSYtavNJb5RIJH6J1hHsMKsMhYVlLU8
0o1PNmSAtjudMYnkXaVEdLhT8S13G9aU8EzEX3xOC877fb2REzoPS8Qul2mO99sftoe8mjnA4OAv
BLl4DeUVRrCqkGYFM5hizZaFlZ68u3n722u9btHjvQy1bLDx6SYBgDsm3yz7eJYI4rhtrYXEcJuQ
69FAk/xvcY/hyNLyHqggKOm6qcUKHBluh/f0EyyJa0nOKmE8VvpVpKvraqXJzAuCXf+lxJYL5jzz
ySZ49qfuzLH69Y5WDMoIWyHW6wbNKFGwMqxqy05EQZN1LcEMSOrQ7TnE+VfLQlZspla6K4up9Xv0
lv2W7+8iZzyBiAspD7EQxGTosBUp4Gj/SFvxdo0+NpBGNC6i7CEbPbI0yOVybB2KaIMGxXtW+/t+
yBRDrns9AtBggHevEwxAEFFQGfNiErmUIwu7Ay2jF5rPbWgYzFlMIRxPW0J+VLZUa48ie70kcXrQ
iGm19KIsGNsqbkcVy6e81jO0LnVAkpuQKuLbk8wLDhc03/ba5UNn+j7gp6K3QksFtyk1HamUf7lG
BF2iFeCmhBWnpPcplyPkzX1zK1xdkrz8hGzJvwABJIwJ71NvSp2ThkIlmBA2MEfLnHsFRjvrkkqk
ACAptIjU/0pOZ7aAR9oa8J77Jus+0ucaIlo5PMdBItFHiQ8lDYCp9gBOE95J1PogynN8llme4W6f
UQzjSu7z5Ij1YsZxHLqSbG6v7b+4QEt71Cc7C4Ec7Tk9bJCKQBbBv+UyvB2aI9JeXMcJhi0jebRe
Xp66CY2tymMUYFgfrumSzn/H8r25SqVmwMiy7SydUWBRbBEVrmnn8AXpZzdni7j+5QIo/T8jMOla
O4IPg1HEV4ZGQdfw2gcRvFTXgYpOAXuoRLSNClp7drOu9t/EOdl5OODo4hQVFm6597fjmxCdZPGz
FcYYMObew3P42RR/ZwfZnovcL2KoYTwvV2qKlxTgCoV71zsm4Zgm9C0Ik2CYHGTiFZJpJsxEQ8vp
kIoB4OM/Hhle3e9N9Blxqyl1fnsD/sPtlnVu0AE1K1yUXXB+J8dc1PMDmspBzL7G3k3X7+R1Zzre
MDI4frQ3tYXW2GbcbQ5JmKuU05zY0mKBaAuS7At7Gj3Y24KNrASikffhHjjqB9TrTln+L4Uh4DcM
m8hAKm47DqMM0ihiCZbFOZA/hf0xWREd7pJSBfxsP+kRqdeUStUW+jDhQ0RANX2odfDaxXFHmV5t
eCtg/azdR3OIGCby1/z4fB2fzEuqMpM7E3jRXB1KPi2cJBHnUa+EGm47sYTMJBb6uX+wIPNBAlci
NGF89uBCZapUqu+JjJ6Lvcz2rQimTJmreFYvDu9MfqRGFxmM055RAAz5QA9NPSGjrwqZ8rsGj7HA
CZt05RLsMJ+utn7GFlUZIi1QQChqZDk+Pgo/cQDUcgEWv1xMwgC7JknlYQ2KCqWHmRuuVCNR79Ag
Gz7lKv/2QaX+U64N31YC8qh6PxhwZLftQ5NNnRDOJ/lZOFCXU9UZdWXv3govCMaXsu6pgxYOrtrX
k6eadO3+WiQwlyDZnq85+DMAo90OAv5R0zRYW52N2TubTKR8S+Qcv5Eu+6S+yPtbndh8dGTQL730
mZtsEt9p9ilIob6UL/Qu4uXWf+eZxyyWzEOUAqEGFVGMWhdukPFHIOc98c/25FnNeRW9kqVBHCA5
veqIbvxZPElMDhI2s61U6Y3eAv+0tw3YOQRBO5b/hlv/rK7xiIRrQpc7trcQtnKC2fKydSFyriIf
vJQl94dQdI86v7jon3jPrQp0EAoH0pjopTM6F0atilb08Zf5lsaaC5Vuv+F8uPVmBEBDWTrxdpaI
ogVr4yZ4H686DqgBOuMFsvzgfM4yOdWcCy1gXW1+IMyESfpJ/jIUrnKu6+FUu4kd+tGtbBnqZKEK
Cl53uGIYff4egEcFI0Et2XR3jPUnuLjQ/Nj6o6j4HSFQ6WqjAZCMMNp3LedfiCrsj4lPK1gxgFri
OkWKQCfrttDbujE4NA5f4W9kmBtPJZ6n56u75LxBBGUN8opz7uZxF01zKzpUuETPUFsmKFqpbWF9
I66LC8/Dl8Yc2QpfEDe/Fwyw/PS8n3oYfdEE2hDCOP4junHaImmq0CW0N9GbSxhqgIDiqbMHXzrN
eTl1szbk4ZPXaazE3EObZrRramlmUAcPsDWmPDIXFOeopPRhpD5Lu5ZmAmCi5Y1LzFEETQgL86wZ
l+BetoT5MlJlnd0+ciHxFlf3GUXktGLaq9TJ5+zxDeYSMAVyDVUkCXrHR6zQZPY5uCMuoCo35hMd
dFyfyNAft2ryo6KBCgTERHAGMs+JU5aaU7PCwHQtPPuTmvZ3Q5hMQpdVk+Uksavns9mTlBB391I0
8mzPIga4CG1nQWcxzjhueFjUPAWmIFuY6QNygLQFiu6PWqeCb+shP3hriSM0bnBjmFPcVlw2KEA/
YGoHah1JLDZOjL+WMs0pQxU/yFHe8N08W55MFhY00Kda3E51xCpor3+c6gpxcnBj2l5LyZmzP43t
R2oNFHskvGQyjB0/kHHwJMR0Pk07DogemKjIHeMDbgDPLQFAeucixAal8XenVxAUf4iN0dB1FhXh
/If0UKsdcjbe0yYFxA1TMV0kOCPoOitlgeFyPe5O9W41xINr3bzS6q3F5GtDVnWRMvdyFFnSxRho
by6jHUEg9479cfIN+qf5P/spde9C18apumfrvQ5juZX36FtAL3hIVyThD0/LPtF6U9HSJNR2F3Uc
hvVlOH1F/efyPjlOIvPeZkxMoPtaxKa3D8Z8QxkAWL2ruRPoGFZ+T1rSb/YuOAIk43TTXRlfQOFe
wOh0qX4W7wtt8hTgvD8mkvv+Z6hGkvxIUPl6aIdTfLLMrZvYsnKpt4wUKPizcG3zpxHG4sLdGUu3
lQvBh0qxvHXRGWzyVxE1KZGvPrznZLVFnMmMpbujmqbnWv/cAgIrHKgUGn7rC6bd7A045Nf80FQH
26/dKTWLPl744XH8UUxYFWAREElo1j+wuGaBbehioMRocpj8+xpAEyXf+UwO/pMXd24y9UelenEf
l+nFW6u7PLcuzl2KgNS+75G3it90e35A2W+HB3xhRCvU5RaeG3gxgx4RHvUdI1AItlGbA731M+qS
cMkYua7PbWdC5LkU3YW6+U6THgxKIo6BppyaRCmqENWht94ySoeyd60aNNBDIi63MN1sozWRAO4B
sO02STZaTzbP/rzsGE4Lu38Wgw6ATbvi/nWUcwpzW8dTu3pHlKt7W5PonFd0iuo27IKGDgTiELea
YilWlFqZxc3hJlmRxo1BxTaEWiEF4vBpW5C6TTWMpC8voH7uQDkb3sS4Jh5KNXx55U9gykjDD7Vp
2xj3ARovzmwyo/51bxFn10l0fxAgyGFFn4SVCcl0TXZ+GzT9filvQODaYqpVnDCU0kjB6sJ2TjC+
tEA5ZLEoxCUX7yejA8gpedC7MuN7Ohp4f3OE5jCzyr8hwPQ6H6cbnwS+IkhK4joubkeTchxQd/uv
X7xTjamHeTVpJIvOLBF7eLWP6uftsd2WJIhbHNtWSct5IX+73mFfy5XSaU9cu5Ig1tO6hWhARavY
06dQbo7WWSQxH4o1k9M9X4UrrloUbEsbCJpLB9HYZkz28Gprr/RG8x3XEUYUi+bZD90lksXX9Pi0
wET0lxbPDnYEYRzGvEhN1Vxw4BcZuZUzIOXS4WQqLtWK3nqu74hT/OcLcnpCKzmFS4W1O0BtPKTA
u1TS+ITLhU7XqsQ9P+BXBNpgGLTc86ObutjtGOMere8RuLF9o+4W9+qGWv+n+oYcG++KPxj/KQj7
NuyfRu7Pjp2HHUOvuekC2Sz+GNE51FDLd+AgkVziBTbFp1LQLkGuzn0RBb5KWFZVjYuKop2EZCDq
7jEL8o3V9Nfmw3j/Agtc5h/YAOri3rPLocr/ote2vfkrM4jLi1lfo8AeGHN6/6fxDRs5gOGgmeXS
rf/sg6ZltdoIgCgqwtaBj8hoxm0rzxgK2LyU0QU8hBOaIXgVnhcOlqyfjKRdKdk7sdtiFaeL4eld
Ir+adpXog24ob04W8kkAwlXQGDHi+gwt0DcEEJV5WRNaoPPKcISsLnCi1Ih6oHXJ6N0DSMIo81+J
PK3O5sNlUp8u2KFbBTA4oOtSKZNWOdXSmyy03b4DsZwg3mNm029uTUExHAX9HHRh4VX9e6/703Hg
wD3QzSvC+nlZ08hzrULbHDaYZrdlwzcavy1/c3QokH6jBu9ysTx+YpXL0xE/3fNmW7SzNYbADsts
NZotRssvjLQMiSn0xkwqt1jL/oPoXt3ixixgj8I2qp9+JW40vz8BkZ56xTiVL7sF664hn9sOC9kN
1iNcHGzfLwnDklaAEN6PIuBPwCseXLqXC5bexQ7ZBRPZN6u+utUgMmIoOgfPoKgq0TGrKuu36ntR
DuTGuf0c32FfeqsaVS7RSbYRpDIpO6Gr7uphXMNBdSCtxAPyPAN17LYPGDXjoX2XojXpp7Fk3Sqt
9jTrT8xDFojlwWGCeP9rH1+cqtF9d0pJxYcvBwAkKNc48K0ht/pX96l6/dMbUD5Ik4ECfzgcXU0K
ire082S9RjTBs8x4A17hK7Xuv5PzpUvZvUO2bLOQWDw2c0FtqlJKUgL9xmEqhNspVmEImMiUEGS5
zS9WIjzlTMa9opjue+YC0LgBC+3yagNbHasWG5mpVYiffJH3ZTB25TKFBNl4gXXo5F3KN652K2y6
5Sk9YMNw5SFlYbnDbrI45HUexrMhRzBLA1CeACk1yEI+YIYUOt70tAJn09fVMUCOlNRBhrlNfCc4
1A5xaZ5evn7zvsiWyJpAiodo4E/8j1r21DtfCE9f7UBk9GuBCb+sVOOIKSa1qo84C6yoL93S2rMS
c053b/pq0QJqpS49BMvU+F+Z3FZhkTTqvcihEgStddsRj8l7e4Y7K9QZxTpO+I1XYxgcfGGiCwmq
h8h4V+IuvOuo2et50QJoYtDmI4nkMuHM3efqqiXDtcrvWc1Ff9T65n5lbZR6733E5g4GgpK0xWhm
nJ24B4NmGFjVGV4/WCezq8V0J8h3Ff+25710DT+leZAFZJCBqxwK5iIG+3f2r1uY0nj0apWZqXr1
uV4iUvl2OzUGMCaX+YNoCggXEo1q0inLFh3peywomEwjr56DYpQQiPOOIQKeHe0LUuVy9Ee+zGdY
2bXq4Q0C/GXEEmo1IbXvebTgLksHKTBIrWn+9fikel8Xku7yfvxMGNn0H12sKp2biI3wL+51fKdp
oPCzjnQZSo2vhobZzjpmDUBcoRSvDOlUdxYagj/YZhjqxuJkcai73ndNNgZBut/d/wA2gxVsds1p
7gorTn5KVplC0oaRSugef4zJxSQoIN3k4FWRHgtQV3kxFqWy9h0lGcMRcHn6rCUToJrym+M3TMqA
jMl5DCk4oto4IeLVS8iPYirI5/Y9QH9lqLrjj1Cxk5nO0mUYCe3yPCfYMdgE7E0smX67DPCsQPpz
DEw0aFyYNBoQRLX4SDjvpvGi6CdHuKfIvPBk/C9U/kaNCBG9E9z5jK2/wf4xjCw7PX0YryBZh2SG
acoYA6I2NqkTUw/i/kzEaveUzQuYfHa+FyFKJ7Z1d0pgtps50VuhQKR5aqleGh8kkuVImlvQhWRa
5JIFnqe5n2dQjFh1gp+wXA3/d3evvG4Xn/spyfLiqGJq0t6fV0btaYX1jb8JfmohzzrUFvVy+qLx
Pi+iaqZeW/qQIC2eE2HElvaVqMxZOAM2nTzL5QXT0VfQHSuNTKt6hMIlzaS0iLrE0gQao4MXyV0u
76WpLpBj1d9h3H2UIwOKLh5cJk/gdFl+Z13gjKW1GMqozgL0z3TS4CmC975aGc+9x1/IEV1Nz/BV
AM3ch4gpwucpj5bYdlZQqoRuViFE/TmlwL+BbdXA2MWMWAtaWZCpBHU30+uL9HK3t5cbrLbVD+1Z
rJWLTg9SEO0Sa/LnQc/ppoD0s+7RRiZQtPPBgek9CXldKtxA4+Wg53niX6BYV0oWx9FxiAF02HRu
Fw/BPw2hUmfRyxGuiQv9AK4TY4CeT1LQ6YH08f8nyAvHdaWKG6Ukfv6KNDljUlczG+lvYCK9r6zP
O025nPf86s1vsRxHpcthxjcON027HnenPnnKawAvHCakKRQbnkOgXyy+N1+ep91yewSrhsloI1Vq
shu1EZviSt4N0g6d2U1FJ0Tiw6fsquZ8kWTPOJ+WdlWH1s+1P1gtVFhxsvySdNepyqLv8br/M63R
itHjshkwQD6kmkloLnx8DKYEKMX7ymVdkw9t8+58VEG6qZ0ZFnIMpbvCYjSjqOxCtco8+C3NPLiw
YaCM/mZi5JyahyP2k1E6bOeeoERItw7xD8O77WoWLdjUdlJMMg/rL6NLZdxzWxS1rDidHsVmorRL
LxL+KtUmTU+caJexn3dScUJJtIcB7b3doQYJeh++XP5eu9lAoA5XquCCR4urg+oLp8vNDwXbvH09
MyhbSl+0kefgocFdIqXe0oghJNp57MeEuer03qN0wDebF5F/Os+EUjr+lp3ksxEhQ1zMOv3SayUm
lkPsfPmxJECMlkdVADF3N2fpmIqqFTcg6rFZz/nYsM+vVZn6oTltFmrVcJs7PUngvUttb5dHNgjR
em4J53wnBUvTTWJISLN0CGvwI2tqkTDvotG/+2B4hn6pTnhGvomyCq/z6y7gtG3a4Q/wqjeNkRpJ
4EXcmqnJAh4ta3dk/ssxxHiFyIw2tte9Zvl/nLW++go0Y2VqA3YLFdD0x27xmO9HundPv1nJ3IBb
YOWQ8tK8gBPDYEE/YKM17ScSHSW+LUamNcQwNEv3txPhVm9FDaU1qQ/qBi+XbH6i1gSOdPtpJbU1
M7nWaHu3uxrIp9zuW5mq92KeLNhdDx7zYbyYSEvTD/xHf9ZJKwkGaEVKEK2DP6XEr+nwgB8vKaPS
T7h8iPIkI3V0dund64Pa2+oeQudWHNnt3XW2mBS0TtWNzXpfrtxjXNHJLCgvD+acWMHC5nm8flaU
/p0sv+0aeoMj3ImvoUo3MSxvLEp5qRHm86WDUvw25VA+AgXy0h7vkNEr4NhdOsiRynXWwhcEYwVH
NH8P8zy69njPr+fh2fgNicbpywPJXduecRgYQj0eKpboyRqHZ1DKmVMn8ak6NZFVL0Mpj12d7J2b
eL9yPcJUHTHIjZiFoY3LwwaESPYn834Dh0MFSVQo7gQ9lO5MnIWskbMS2mEB0sPouVxJk9dcdJFV
5cTSXhD8otCQ/sRK6dpc3JTCIgeO0+WAtmtrb/yCgSXgnOoysXaceLqatEsTix6p1/wx7GwCcKMP
WjBWUDiVKFG6YUw/88wPoUxv3NP4iKxFchgJO6AJk+cg62wfIlqL2uvOWNl+mxCp6NJrU4MuI+Aj
EghwCcx4tH1G33/uOh01OEj8okTquQWZ1rW/MQ9nC0r/Fj4CcLB5JdBhRKhSyDh8ID8C5dgwz5DV
/CvtBIY5bOXKpsNHvcwSzfv1wtmKCn31wZDJFVzdyAmq+ga4Fm81feey5YPR7yTfSx/BO/NyF4be
JE9asSZEd+I0kyI8dhOdvBr8j6OaPOTbyC/rsiy31/F9ghmQO82ulzPi6xu/j7sqRDmFDc3vm4HC
Yn1emleOC24mpIgzKBJRJh/5XhCwsNmDBtWeWlCI0XjD3nOW7U/9Ek5Vox9kH6c+oSo8Qr9WfG1Q
qhMIvYoP6aXQ3AF4Su5/wpnjn3jyIX0/rnquOe7xsC0eU9poqgyNarP/B7R3Ynq6WRH1mDeV0c//
eNSkl4+tr/rEmzK1DplV9i5Jf78WFpoU61hbkO50E1eEKHhppNoJO8m2g+CGS741pR8OHK/d2vcL
Yogqa+T3dzq1aC9trw+7KJQOyS8VsPZPFMajfJx9iTwi2XEK1aVsWoLonyRV6N7ylWd1jb9DdDhQ
y1eLQ4/QnFlf4X0Slpigt9tlNuNXMcqHqxJuuu2/B21mnNpCvPXG79UfMBM/KW4EHWfxng9QUDE5
Ha2nBckIfXPL+UQzg3PojgRk6pdcHpj2fn5G8iNOZLn0ZlLrECOjfvF7cNyKX59MkbCitgnF6+CG
5NWd5zDW6EKxR++bKW6eW1Gzp8qNs0U0DnAPWSvVhUAOuv1sFWUz9t5GP3ceh7hEsQK08lUnqv4T
wdrDnp7+lBvRruxW3ZAzOupnO9o1UhRj2Fm9bx/C5PXDMk02r5CgnXgpREuq9MKNpY9Lp2gGzOON
zswJNUTbifU1UD1tNFNni9SfWoHem3A5VZn5Tlk3osK2sW8SVHwWgtI3i7Ii5l+/qWAK7gRWOHCM
xhtp5OY0YK8hb2qY7awECTwhi9Vkm/pIsl2giBLNHWdMsTMhTeOyye+bDWndGKmhcOUyDISy0yBn
SVAapFHGj0yWLSkwX5b7ZMfae3LRcCEd6w3lbALguYJqVBWVUxPhA24omSRb0T1OFvaEGbrPjwCT
ZRKikeBiSUhfmgrN2gb6t5XxLceX90cWPTa3qRJ4gVqihRRszFAM8TGOAv1yg8k09lXJ9xATX5A/
5bfGsvP2Lp6pmapHpCkVpeTorZYyEQ2XRX9zY1deTwLQsQPocuHDbJH5ivyfRgctzU7kAxwGNkmU
JrcVh0cGsiekghZFCKymiw28qPeIwaZB8NkujU8p8s9u7mThBLkcejjLMDXgavuR2reYOWNMpU9y
Q4sgkr1EQ6ND4/WbqMb8B5n3gLWoMhYj/ScYs+KbxoyarrGNaSjEJBvtlU00b7zf6yczvUrAW4GH
dhh0b8tvOQZUWtWQ/BBoWsw5FNVUpNo4SxY8gmvLymwdV4sXP2MreAb0gisG0VhHqmu52NqMruL/
y6vNptxHm1PN1tRLJ7zKzthuiP80mFKK+FnRLCn6XCcvFJ9qXe0Xp3aIgZDCF4xo7swYFcrpRsvi
MMrEqQapRxJyNqstAqMV04w8IXMUDt0JfpIK/EsCP4RoyjM/Y9aQqnJU1zxt2rnbYKPdAzs+wgb9
jUogH7rTm/i9aJfZXlaV9kC4Cx5lmmv4IfQfQ2JPAASVsjqnuf2Wyt1QDlPcTsIgq1/4Uhjp8PDh
0z4vHssOESLvT378yzyEEafB9hS22uOC7G87f1SUhyERcUIaCqSUUTOvPCuZhgXyVx+2I95dQnFe
1Bo267pqMWuHevOsT/sBbHl1BHTYzhp52Hx3GXzDDzhVbfkhEhr/aD6Qno0kqdlboyxXoEBVPKMw
BMpUY1KE/CaBPJZ7i+EJ1eeKJ5nceQgMZaVLC3l3s5f8zLFxFJIZ3RobyXXqkU/PH65AKCZkSBQJ
GzEztxoJL0t1Vcp3J+AVav+p0yrnFBtMmLq2GTZkr9AQtGjPXR24c65uDqeQ8BhDoYHDQ5IotQCs
dXU9/LoTywLwUsjma0fMH6O0oQpxjMOQS6Xx/sNJ8C9gfRa5E3jLZAMxJLtBnlKq6awzkQ/LQgxT
wg81ALspzWRk+LqIS31ZJzHE5NLQlt/qyVCoJrZ6QfetAJ5Hiyh7qae4H97kSsm41cURypwFM+UV
vPc+PxWXgT1YPAOcPFSJGpQzpTkdUQJ+ViDNZOUjtIgRwmJ6VY+D+hAiL4fyaBnu3ezbN+zusGcT
osDoohBotFH9vqlkKgOp5jfWuJXpSyKeTH8q0somZlrb/H80RPhBqGEWuyFrlA4zEp7C+/kZ2tcQ
4d7iUDZ2oquDIu3j+zGgf0u3ihL+3YvaL8vs4nfk0u/d/u0BQZzobTpLGwIcELnUtt29fTch2v2l
yNoWqgiMR/m/4y4j2Ci4nZPM2jfZx+P9OGDaJKNSyQNAeLXVzNNLA4/nOVdrfJbcJXtiMIft5Ko8
DpkW6KKxc7VX01nqSP2HSK2iS/TiCKN91Efem6b9/abCpPqAeBbc8/RvUooH2cZ5X7flfQisXXpq
b/1JVzxtNBN+PvZtWr1/ARc4CjEfLApGwwgEbHDJxkOFFbVJRo0O/LKyOqSIpCmhzPUOzx4jmSkQ
8AigZk74BwYonJC/2hQSTcx52ybkF5Z3WfA7RQMqvoXfXcG5g2kmj5EJMkuzYyzYZJoT0Rc3QTfM
1ExmXJ7/+RB8zJOe8k66ODxbs44Mx9isHI1Ovm3iiEiG+nclFw8skKKN1SpSYnsHQAtOq1EBxBAG
qia4D+oZOv+H5vT77aIDpOBv9m+YAGETpRxyK1kZHqiIyr5vUE/GzV0nZ++ltQbP8P7X3PvAxCif
uKKk74KGJK7P8J6EhMu96E6S7YlXSQKQjNHbtoeTAkCvbxmmtUzr3+BlVXxEKkEL0kkW1US+q70M
VkFF76vS5GtIKh8jARw1UMnFIEugUAVXIZD8drrMg7RsbktIGU9+I93xl2M4Lmy9lrNCPMLGZ5Uc
WxlBzp/6Z445diVKuxBnbOuUkM2XJ/p81suITulsSo5y5J9+/y56T8ldzNG4wyFZfEnvsSiNR6qB
ug6tEegu7nsVa71Y+3iiuzsCisa5Rq1rOnE/Dh/UeBfT/JK8l+YaWv5hHTaRlHZVK72vHaCD+JcB
jrcpDIXp+h2NNCKZ5fXYSYxGemWblXfwk6auIKjvyXguEjAqDrAiw2C/gvLb0vXAr+GnKWZydGdV
gTp0/75TLjH2D0vwQLdMahL6eeuN5nQD/JwYirFV+nANK0Zqa3RweeSeXg9pdO8bl1ly61zJk/LO
bDwE7I8NBWsNDMM+dtPwgMlCsVYh7zB2hCngdhum4duFlaZsXh5QKtwCB4I8+wEbQRrH7j1oEQzZ
dlx0Lm/1t+opnjSXBIfRrfALxe93IV9Lre9HmjynWdstR6o/o9k668cBl2H8lahYFnqtG213SsXO
grEgIKnptw11XATK5jZILF1ODVmY/DXKzvYZqhhQgNvahkeJG0NxNnRifCwbRCjwGZ/kdQArFtR8
NkwSur8wMdmnFnPY6ZfBdFbCQa76/0W6rbypweCZSaro/ZypRtP92T6Q8EqEm6XOmWkfO7hQnxaw
xIiCnA7h9vv5VfRZoXDzEjReX9uYSh8cBaTW3Mu8G/bkqITLUphV+b6jO8qPl/XnPuhroIYZiqPw
uD3ly6EhMaREauKFh5UP7XRYnqOC2O5QB31lxZh4JhnVFwygPKs/JT8XU6g4DfDgLy4uIM0lxE5H
KlCPW+4sKLNXamXODhPT/+9ffvGUGFM4IhKyNJV2icM21oAM0jHHolqM85L0EHIM2P8cD6VFOCkI
U5GOVBavTKDvpJT9jOvs72j14U5sWYYinNlEznfZ5TDTO1rTpz2yQ2M4OFmyepwQaSSHVeRBUCRL
gaoMKcQXGFWojjH1TxUqdtD4HdUvMQ6dkfujLgFuxrlXA2FybzX0mNYLqR4An2v7YtklMK4rEQ4j
OFHeNsmqZo+OG49WCXGs62KEVGboAHKZE8Uk3BIkNJSzZT2+Bl3bn9eqme6oEGcRFneMiCgL2LG9
Xx6OuQzVSdW2VE6GhpUBA6mYruq6EYyzxnqJr3PfX0zNNk7+zLrd4lzlYL54i8oetTbysS0k9CQW
kOvQtHSr0149/ghZTfHE54uTiMGHXzyJ+a3kWuIAqJQYNvbqXkgYphF1FZlhw5kV0lM4Q2QZREFB
sJ5dKJeK3Sn1tQuksuwu1R8X38hDQ/JRm9UpORuCITbOrz2pYnTgCHEB6TsWB0d5jS0hgv/IL+7m
QDKq2iuzn9Ifn1KfrNyelGj3DHgAStdeoYrCQgga9pjFEjoHvtyl0DHaFDUUWFoileKrnD43tFIa
yK1Mtbs9RzNeMOpeaJ5afl5Mnkh7t0XRpO8CLjfGDnkPaRIaDYnrc11mKIvPSEbWKrtvr3JDqegK
ZQZ8+4Jswn0ShL0MZH6gzBGkrRwrj8iBA0ki3PvMErSoTFv0Xr+80FHhcF91LrLbapOS/YM0doNU
6AHlFIb43Z0MlxT5slf6Z680T7J5wfvi3JDHW/5BDpaxe3hUrVyEomHtRTNJKPXNA+t03/PwOijg
kC0436AfxeLWd3Xcx10LeEYCzvciwd9PMq++4yKtpv+JhG/19IdVm/J6GqTCzYNjUOUbdV359EQR
f0KKQWaqP4SSfqw2wV+Pyxl7vYCouxYK/5E8tytfUpc/NqLWNt8Z2E6UjqdpyGayK4N1YirkTm/c
RHuMWr9k7vRBuTIHU+fvQ+aE8+DiRnOBRbFW87Bp8MM4HECgQ/OuUfe5Adcz7b5tmPt0BceeRvLn
6Epv98h1EPRZDtRkUdH6Uge3MtYRAd4FjXEC4OBqqSU+P4zbdPVdBoYdnQ8pixeqAc9hEzQjzjPJ
PxbjT/cFB4yjcr8IppvYvZsSBNOXH/6RRE+B/i2ryghWi1FGXh9O4ezCOjOIf+I87vbLVLB9xxi/
9ZMekMVrXzEIwcxhf5CyEqV5av951mnZw6U4mW0/nad2EE/1SCaQEdLNuA7MBiaSlLHWTJsl5ltG
w3GM7VAWCP2/i20JqzUR2uXTqMqOMDnylb2Kp4fhLP/46lLju8YlpNROdZr2lwsyMYO03Ydxwhl4
+0ArTaHyZU1YMWUxegxKpZMuyC6fvpdWZhy8Fs/HzEWYHPRTfT6Jp8z6haZA3B0RG2MVljLKHaep
dSDOC3e2bZoP8p+0DA+PNfiLA4SboE8ZC3Dy1iUuZAEApLV7sSAj1v0u+DF8FQT9o2JeDzmd1HUv
dh2XyAOPo9jH3OBccnERUCwGeCImV5VI/DsWebOiO2GFMoWLtJkLQUjaAUXPuyuyHcXI1POmlGGW
xIQyYTbBK2VlnMz3SGCjY9zCuLyNNYe9zMIsXOyjYJ0pkzrx1lfzLbQGKs1VQu+C5n7ScWi5mSO6
uYmZbYqHIO5QGmnW/h3uNWXD7CcJnkVBmuNeVe5Bael7lqH4AqPpykuEx9rT8yl6xHlxHKSzJqpZ
uwGnf1cLTMuIXJrPA1O0sKcIlQX6JxAEBtW7shnyQT3MPcmz4Oz5XxuMKyyZm2MziaKZpuub6pHn
MdFujQwFUBwLv2PJpuCSmOLtoVBcqC73rAXi2wBGY+00hsU/J14ONLCDrM6UBR2xkM/biXo9dzfx
qZsqmU4IdKHHNMm50WWDuFCXIZvKc9UFdpiSQOVnsiCzrc1oSFzDq+7L4kYyQuYTmwyXwYYexn2w
YY7iXEFYp9GwfiDhX/SYbIm+G9OAmwJYLrM+kYG8C860gjlZ6SzaNuNvlxFUdOIJQ+og21mHxRUa
qIsUeY5Qe5kZ884h39imzHJCAAa1SoiCBGEJR7dOHJxwTHTjvt7MLfOez85s4JQ/8r5LISKkWMRT
IsJD04TfTaiXTtKA/j2t3BOXTJc3rZgujl+pyILpLC+4TeWXLM0HoBMtIrniO/PMSXTXqQ+vT1I0
T3OunbtzOuWGpbTUv7ZYgjp13TMENmT9PmJ2Y7eK/lr2RAMRAjOYcQeEgG/LTimSDiyF8hL4LTw8
uoRuaHAP/Y0Di5jLX9uujrD9Z5Eqv7/WuL7yOhgCrTDIYkoSoopCfMmIuFohDdFeURswyVs854g2
i37JQkr1YLhujpsoHD28dXNMhMrUe6+Rkb/QIiAX30CNshW91G8G5Xj0/hd3936zg6MDXqO6bm5Q
G8CjqAwj6Pq7FXddBHjraqoaHxr+7LKX2alqQCfal/5CpQQvcHEy7Jcvd6QhJWmzKtNpm9RwZEAD
yA39oPWx8TMBbtj3EHD7w+v/9p/+x5l3N6kNMM2koukw1O+vwzfT3MrYE+7MPuGFWB5TJwMkjMoi
q0Azdy5VY1vlvozWviBS/qhVKVJgLKDX+wiHolkqKwd6TTFzzEuFM5kCdVnsPoB4XYf1vdVmosnj
hDWJEnuwBgg5518GxpELXEp/A/jAjf4nUyxHgaOaTpIlCelbfgfcKMC/2DdQ9HpwuR0B7dr6dFbT
Hpu0Q4mlhYYGe2g1PxeR5Cxjr7hnPBgEi+ZmmF5a1g0aqYPqjnw5a6BrTfIq2hxpG2Q8UbQB7awL
nuICjfKHaEQlbaP1473hvisMd2BrFWfmz+rscDSpcPf1+l2c5V59oWq6iaYWCp3/QUcdPKWzkGdo
MvjBLgubGuH3ajYIrqoK+jGu0ztiY2JFqe8hfuPQ7xH6SNrIa1mfypGZw4lv63MtD6gGdHzFgdQm
wNlcQQFJD6B5EHBs0fFf4uQfsV5/98jPi0pxH8jz0ViFw02g4+nAxNXY5Rhvt5Cx2VhMWXnLYTU6
QtyhOQQRcuEgwofEqeZaouAbM9xKhPy0dlIzDlefsVYOUizYJMXFmNUqevC8t4YYt29jWS3Ht+3C
jk0o32lrkqwvaGAgwBwTaByY5e43seDu+77/slFZiGPvKnL3UCz1USTTH53qbKJ0o3KCn2pR6Lqb
+df4shC/t0tCUb2QgbDyflZm1s/ZmtgsbgCk3zjQJADvq01EivV1I3dHYS55kJjTAKd7NeARXDN8
MP0paFJhp9+vipo8g7n+B21OjlaVLtpPg7dUdHeOAP17dmPkj8jx14cAYl9iTfOJLAFPQEQSlp9A
e5XPTstSgMn7Pxn3lw8979s7WEz6v7esoQjv1xZ1IcCVg6n2CdWaXsSH8I2JmOljOjoICHhnviOK
30KJZ0D65fACJKTi6D6ZShdFK8g+5u99uYzgvhLiTv947lhQOtkPQ5pFJRjaURJgBFUKrkji2lBo
Ouk4eo+BlAfi0GWJf4qT0r/ex+ZkLCmzkQ+C43lN01SgHCriY9OCcAGHWaqKfqH/X53hLpBXnEI5
3siVcM21p1aNKQx3DYrBkdQmWPSX/JL7c9D0aAWyfVlpr5fJOB0KaMWmvJ2CoKqSqRDCuLcr24pn
wANf6lPXdhGKs2lFqVJJglwVbUo1lEgv+VoobHCNwf9WXORG1aySZzig05vyGNksTOpZBJGsQs7X
C5Rv6KUaYvPe1HbE/QmdB/kkmeok2wR05kE6YldnN9z+2ZAgq1fDAJj5aOS3uPYEt8b0bj++LjaX
Wa2zv+7kO0OUt9egB2J+Z4N7MejiJPriRqg4hXAEwZ02GjR2cjnX3jneEeW/iEabx8c9Vx4rCr0k
85uHxJsdpciAQ/ujXJRVmNe4rFlGcgOdVewvvZOFDEB0QVUtFTZ2p2ygHeyGiehQ0SILVXyFVJO3
rqV4tOye3t/7bJYOmaecmfxEW9eSzh/hYgUUV5em+XmpHAZDYrDsljslC3Jsm+izcoS9atJcAuVn
35V8UfDGKlc3zxe7viLMwQglY9BGBHoVn9KeIBlS4g4OD4WPftDQjDBpwP8cUE78A98Ast0i2Cl+
EzyXN/Aj/0x9gohW06hdMHo9wUt0tuc7bHIHAic5cQFGyGwbM5yDHZpaG/pxkaeh8mtZ99lDvDUw
2ywF1xq0UkSonxZMGsfPi6nRom/QEWY+zjx0+w8BxiAWsCUbG5JSRBWfGQxOERN4XZtAMI325z2g
IisG8YcJHYfdgJw5L+cTP8BD0xOUnDVQOUfF37r92BFKkyApzJCOlicBao1cFFsO7Utx2efWZB0Q
ZtrHeeYZCb+zqwK+2mCl0+Ke1mAmprogzSPe71XDgCSyEHw8tBvEeou6xq12nBT68JuvM/C0YoKC
mOSVfwMx+zM2wHow+vPU3y4H7Bi5nQMZDvGvoIjccmeQMjTFQhiR7AG8+/9HurWCnqcsNxJGL8rg
pgQgrLqSekH1oKJX50Tki4zHelLQLjcCyrz/+2kuYyd3bsq9+U6lY/AM/LCLg51TgzDKPkVVvkUH
mZCa2LmZu9ezFvbAVFRsuXs3/TQW7H5sHXcUj+oRRcAbV9N4hLmhKlgAoSH2BXyYeCALJ/GcZ8Sz
S0EacSk+RCOxOeAU8fhMAQd80Wn8nIz3ccF3IKrPhCiSFNAVSGWiFagvh3KVFSlvyl3k0MTspgQP
GBque04JZVd4ZlefnDHVrTQcA7Od+WGvnDavnUcc4JpbHFvLvEPZAbJvVjVg84+4NXLl/MA6SDiO
ihh12ulHtqEdHR29GJSCB9wShc2BdgidHZiTjnQhS6w/KJjz0TYVe9T+EvkWsBEwldq3KviASHe/
DEy/8GVLhaYhOf4zAlJ3SBLfXm7u0J4/qHpQCBaO9w8APTwtPTjIIf2GTSh7U1iO7DucTXx2AhLl
pjOF9Vcv49xR43XISOQP62TDOYuaxJTEQz688clkLT0880/YgcgTc23hM2cG1SmsavlnlwHnZEGO
T/WZSELi0V/QooyQAwGj+iEzpQOgssoqDRGv/87G32Ovod8jKwTaiW6hNWPitLt0DlH8C4H7JhNn
3jiBAfguLxScsvqmbbLQpwJHrat+KGrBn8T1o9GPgDY3wGjGyWlfiKcwDLfqFWYUig7+0UCN/HwY
FjZRi3bc6vw5ClTPNyTBxX6nWcfL+0dYvQQ7YhyZEs0Wl/oUaaWuSMIypjCP5gsDHvbHB89+y1mX
BtUBD72cfF02Y8F5G80dMBPrwxoa7RYLECLJmJLtowVm2PHfpFANrwRy4mt8JCjVjq+uQ/xbDzYJ
bQvq2NuU3UtrpUDTDm8BOwAfWMt5st9xOn9v7DIii0LIZbe+QImLKJFITAtXnTQMiuDojC+tQdYB
4903VMMC9qyyZoHJ0UisJDiuc6ehOt+ToULL7e0IngsjaA+7vRXvKnsBj+k0pp55jHmeWyX1AvHE
tMiSXeoIvNYUU43j3/mBihkKt6WA9r80mWucaNx1Km2cq/2+ambWT/nZGsoN3M+BnSCatucIoWKh
8+u+DAHAaIveSV4g2S8/Hgj8ve45QdGtDi2h4ONKtxZvpdBKhUyt4k36Us4o0izxtslwRUrxTzVl
ECPuNmz9vb/4uCTTdt4NObvpeUyyCb2ICGh3F2aC0y8DEa/aMEhjtGJauq2KEV6z6hLnbKV4bBCJ
pLq/0e5/EAAguvhkjyqGPuGMvbGP/zz5ON74LeDs0d5tpew/J/h7Zb++ZEtpFQ+8g19qreTu9VUt
VhvSq19KKMh5shhuuKSIJdWPuh27y2BAKgV/gZYhjxu8rKkxdktzoukzuzzX1n+aIsZroc5J8wQS
gXPhsZgidE/osuywtSXGzbMeXSWt2YkKDzij4rYiMlcb/PGSacg2xOg/XdmBfPEBGDn3DkLn0kJ/
+3ZS5L93ypKBR46HaaFyjcoh+HyxEBrfab+yl8wpmwkTHtpzaa9Vfbq+jIR2PiO/MztdP1zJnJpF
Ds0+6GqRg3SbzurTD6GkfUXdjYqjV3WvVE62bCtygSCVbzh1zV13cyv3gZg3QsfT4UKsfjh5q3qQ
PMpRzv4wkyMMLPIPDtFxcpyUPR05jzsihZcbIAuBfVgo7ZqoNFtpKqvhVy9CwKSrB8a0CM5CWuI6
bU5mdAVBcdKb6g61bIPmiMCJ7Btw20aoCLVttLJPcmKnnNuhNb0NBJXdEPmSAoPEBl/HPmBPRmxD
tvlgFjN9Yo272yy7IScv4MiILIw67jg183axekXJAj/B7pI9Vwl6Cw3tD3cniCn4XAV2GxkiGmON
hieVKmwB7WH5ayhpWl0S8UI0F4/Tq+CywnvTYrXgSw6Btzo5ilXF+oCcs9Dvy8Q22jQMLZMJAoRt
QYP41Lt+YUwDeQ84mCn6+tmlQFnKRUflEedGuHtO0+2uT0XIOY5RVD7VnjXlJ2I8reuqHzXSpHB1
VxxC+NeoHm1ppvsWH+7F05jTG/YM5cgtpvT/282PdhKzzHW47twauxFK15Z3DEkF/2/i1po3bukY
4YcTvfwTf5yaOTZQM+qwxU2d0oe6AUc+nSdLTt/ptzTc3bsGRrAuhKXvDrUI7O/fIKt8y/ci1ovk
Og4zY4c3a7jjSkBEElE6iP0dc1DnIRWbdkaFp0kURCKkZzcAbGfQnyPfKh0Uy32q28O60ahw/aO+
s+jGGBYdBqacfyUrG/e9Xr3/AfLr27lAHAZMCEZ9xbt724FOgVReuejZTR3qY/0z1NPuNuf/93Mk
m3dOzOY6dVSanqEukRPK3LbeYM5YcGB2AI74lHN/BhsYN0qsdGM/LXEJaYZMle+Kt9/PO0bY7M8l
2tB/ACH8ZszPXL91EdWSkkLAF8f0KFp+xLsSneaVK/LZFZt4OiOPREEKEIaq887bwotQu4p5+FPm
WGPzmG7hPn/7Fc0kQHLcg7jGL2m9Wzsrfn2eCc7yKlZNDOFzBLzg2Nut992VkkUqDJ58l/yBvTMI
y2aGXb2i1rr4414MRPuUsjbMqHqCk50jkhv34zeS1VMFLrarS1L+siUxMAmvGYy5/H5g8hnJ7f97
Z5wBWX+qbdzSIfRyj5pnisk1gXnxFauDrjc7G1anuDxcgh61zJFRpFSB4kDets51sKYDtKxLX2Tu
pICXM1ka1r1Bjotv4Cy7rH7y+dm55175DKq81RJ1+G/K1NisKO7+dgMw2L4W+kjxp1w710ZCGihh
9QceREFGD/e/pgZvSAu6Uxt7xXPODdrKXrWUdR+sL8yoZfjoCzU5b0laBmHUvBdhw4h19PYJ8mh5
HzaKBycnKNg/zD0JzpIUMsPEs3/Mqu/Jm3QnsbiFql38xzotmQAq2vDuyDdyRG5lz6RGqAwRFwQt
n8yjhD1sqPE74yBfJjqevU2hhpZxOjKqFGkWCgPgSr/xJQnyBsMpdGlwrga7ZgaaYm4pELEgmW9R
u95KQsepXfkx7j1w0WFcaBl2aAsPcQsPXTKR68oaVG+YKeIdecDdJzJXHwxC7b8IGpQzOtW6wbsj
C2DoBXRDVvtgwNJINz4b4j4IsmXuRYMG/bS4k/M/NWaKF58KhO4A9UDFjZDjbXjpi/ZV95Cb0W9v
wUhw91EvZIbWbYHft/0ep4awwRzWCLbPtGM3FmFc9P9AyXZIqiPlnR3yYu5mIdw2/r/pxxOXAo42
OWCvdToXCz+UUW4XWM9Gk7QMKX+iHbkDFfwtYTxGK4R/gq612feJJRbo+dnpJihS8gY9ttScRozB
ZV5U8s3QtQFN+w78Xe6rqrhewpW3bEvyvjUcuJI6ylbSxK7FKEyMCBN5kjNziI6OwDXq7cSPSD3m
EcKDfrhsKm163aXlJY6sdbxMTL7eAk5iO3YqmGdyZqNxAR1/MRpEJxJcCwgBK38VsTQ86GVxNF5i
IDfoAqgprgYIIosrgqaR1IbFwmY0rsIRGIO3h4aYsHFu8DXIW4iMwdjMf2U0pRBVdAOMkKsG0oGf
TtooVuKgSAkofN3FuVtfICgb5JGjUw933K4GEmE+EzMoY5wm3AynYYKdUMiJzyQF2BADmUe68Qtc
KBTNIEgMV9U6ovHpTkWaoKUc5v3CJaofX21KtUk54K6SyZ1sKCpbpvUpZYgaGUn2NezZqF1/5PUV
FAtC+JYEupa1iNVqSfGRXoJ4SG45PaSedBKz2yObY5YrCMsm6MLgRJXbv5q5epxYon4X5yC3NQk/
GtT2OaMPjIg6IVeV0dz0/bpOUdTyOKYvvMo4mgrfR+xSaE0ByKSM34a8ENCjmm6PUhNhKPHp8GZR
BTK5QhwqZJFS5Gl+brehIDhjdqVGPFvEjQE68rUKw0iu4O4ek4wlWmgYzZkZiZgzt++6MjcVeHmS
iq62HPeGq8OBnAs8cXWmOIa3DVjw1mQ0L8bQQVrC1Nas9iQ0/XOlnkEJWJUeu3V5iUI/sBTJQ4n5
kNDflobSUJ7mvP7m35I/CrhxGgUtYs62PemPovl7wf75n2doQjyUq+W/u3FhCgTge/oNXHUtvSQy
mWP0ZygmiKIUXIYrlhp5+b3f+d9BI/pHBnCzFrjPsMsCo7GPkJN/nBiORh19tDUPQXuHjstbPVdg
dx45HU7+LG08ulRD9PTGm+sqANY5zuhl/2N1jovafl7zO+4pUrRmq0tY8MslxiaNUVJRuQGflD17
60GYi5273vaDV03ADYZF4pi7VBR5Mpe2FBOZGkoBlSiPXpEYRlS71urxGyFYqOSRcjRxWeDh9Axr
Ws6FRQKAwzWpXOneN5ax/51bK6fM7Uv5iYDSH9tRDa3M3AXL5io3jIe/f9ncSk2/CTl/W0WnVkZf
rSId5J0fCEUDlnE+baLTph26wl6JtanbZeZFjii4ZPQ+LWdFUh0rW2BO4D65nXhYMHSyYiZEP4kV
MSts6nQ7KSzauy0jm+ATcILthpvBCxTcIMFawsit+5dAUhnoWCmu2QGtZz5Z40jVdcl84QApai87
0KT0CpUubq+rMZnOF6qaV8t++c2oQ1PDb5rBXcnMWyoPWp4w0en4HlbrBF/z0qM6qvxEdZ0XVBRY
yAqyxkc7WieJ4eNk8TQEJkYl5R8UpzgUYPXNHj17juc2JrOAK2Fhap1IdRo864slZcSvf9nZqu9L
bNIiiwh1dokqzma24vwm18NKojoFfLnldUO7fRQBmOva89+w8MIvpsqqDT/05e97Y9/NCFwPP86L
onTb44xbQezubJCpQWXKzLNe43IU7Oxgaa6Hbvk7ayWzBwNolLhlYsNJAuWsO2BNz1VSqp+1yYs5
i1wgSFavlCJ4oMMuGl2HK7dO0pAkF4bOFuHAxKl03n9pHw7B0audEsjQgcLA7vJlOplrTMjdxSPA
OoolgXjjeSVRyGkuPMCjn3vnLPyYMTRgqiQv8MOUJC1Evr257j7sb7GgkzZyu370G1DLH3yxww0C
L40wGXNrm/7h6mh/Tz6LvoJt8s8Qwa+EQJTNe4qOM6MQBvIf+QmbnbMHwDKEJV2NNTV02E6VJ7Ax
KenAtrczMFF3UCRV1idth6KFn8LFLj7lnyCkai9cOPMo/jT8N29lQvadj+kUZjIAOM2MGgxYKhhM
S9Ad4w9TXKQFK+l7OvukhxJ5CKFzkVB8OrbGzdPZTn7rjxmNcV5yUymuzGlypyG08cxVvbz9THdY
vmMcHbjHRZ7Vkwnnn1AREevesLAgWAqwMM1G2eRD//Z8NHenfw/kcvlBcX+QRXsCXm5gme6bVVZb
UbgcYaT4mE16EVjN3OQ0JmtHaDFEyEQPTZVSxdcd6H/qR9N5YpU3PyAFVsrr5Opb5gx5r5phroP1
EUlkCy6rzAZWLdwwo1jcajwixHBUXwy2xmUBBNhIte4qxe84vV+p/p0o/N0N4MUc4Ndm0AgzVEIi
83nnvYjB/vB9nqDkPfcSLJiuci3ZTgm70QSrvTNpxOWFbuzsf/YqB5YVD7xHNHciWEtpMDwusHM+
ZwdsT395+36Qlq+6W7POZ3UPmdeu8SbeOiSntzHSYrLOud4AIZq+NvPkEKNrKK7rLlnEZAUDdY9O
8OTIQFZw0I/CglofZdHEkK4GiFsDNH3A/CKVWrCpzcGEcKdA20VZGP7YW9W2zR3IIapjJXbRe3QK
mXohWFBP7aI6mI1+ICVY3uN6/3oBn36xiLBONNNPV/bpOHbGOgX/vT0MhleP7o8JLOyRzsOq4hOx
QrQTibSpQ/m1Crd93RRjtXHWr4VUclMLjEIDIghEKpkVzkLj23L3/+GZXYWoD3jB42dzxsxzjk3E
VumpdqI6g2lrzpE2I7rDV5pUA0cDrX0CNyc2ojJJ6N0Hmn4M6eE8qPvdYPrTPaWsF/wwADjrqgWL
ssYda8yWYxFbOFUKVxqugx6CqaD9D7bWqM49Idtxb+03VdwVlqiGL3v0z7sqt04ByxVqL3J2JeeM
8/65Fz3gs00mnyAvCrznuGPbGVYZEFuk2HXHGEfU44arjaeRafhzOt5YZfVxnVbn2XsJ6+WTZqUo
eqNu5EguU3L7G8pRPPydHw1OTO3H2UahT/5noBNgoXTOqrf0LRN6rn0Gkl2jula2Ls+nIZxTD1Kq
q9/VX6B3zl+juYIOQYZJZD/ZQWjNZIL4o3EVyCLurJ+wMLJuThwgR6N+PXWw867KzHeneaoKw1fK
DCw8fwI9GSRc2gfc6nFaWysdLKLDaZHbncykL91cgDgK/jSjjkzqj7+CwWZVopK4p8CySIUhkVLf
XsR4LOP63KPLeE/MDXYp/0fvYy6dsvNNKuggyPPnb4yM2At5k72MiZUurFPW7+wtxJ9IXse62WNy
T1SYfDD9u9hJ6fwj2ID/K8fWptSfQIIrt6MVqQ6dOBmvki0rUhY2q+27ikifjAMJkHjP2lIF66Bm
m7HNl/YE6QKhojx2N9iQ+TFZRS6qopXWqsyySOmtaswdsuCf7vY9O1BTj1QTGoN0ZNLxJRYcdMsU
lu9NGKa9DkFSUXmc9HPHFbipJUODR9sVYavvD0mJJ2rKC19mxhhV30Qou/NGbdIYekmmq3mlu38+
CTICI4vfojGVpjClf3QVKYPuqEiTuFCdXDoXADYtjgZPWYXkxiod2XDHX2Bl8PvEyxdDihkfEC4x
tvlUOcLAbYTD1vLbM3/Avf1GZbMVAcXHqqlcxqop/NDRuTkLNoEFjXCPuNCEN2HePna0y9ZMrC+E
PTTfrFqwSBGOE83L6U74rlRehwj3OjqeBIO9hGuwC/K17JfudqE9HdmnGMpnRXPkzh8QadS+nJ76
Wyw/gZwlmICSEP79UWQDASwE60Tcmvmd2ZnWDmuvOBX3kqfpQN4MWkg9aWPegToTsbCGGST6vkiZ
QkOwpDNBm2WcLr350KUqcGBn3M5MIhLm0kuDfvhRQbPh2yGv3s819RVZn0zQubq9OrAKMU9CdmDj
hfgQM5iYJpBeU259LDZ+bTramFT7PjTIcK//YgxyHpvmYppTGgExow6js0jROsaG4XBFGZfPgyro
XgZxfrV9V30d9IRAcB+CN409RgYH/87WS4w6VlSRG3/ZHmVvEly6ZoIXsI3rIiuRFF7vQHJl6yVu
xHsOHWcgmwn3ze+7p98gAIb3ujjE4Uoarp0hzmvS69kDAiHNjyWzwQstwLvouQo44AQNIbrXfrrL
NqMdz9BsgLDCaFcVvTJGl97/zefUa8MeCewSF0bcR9QNpjSESEGLEtwDcabpdMJ90kdyR0c5NCJW
ht/dJeFi7P9fpHcqaAFSEeeKSeTEAwjrfDTM9sTY3RZVsx/d9gPcx6RH4ATp8Se6Bc0IePvOBn1y
0y9BeQozug+RMZxNyVVmlvd0wPfpivQL8ph93GUnLu4nSaPbpxBZ1tOIJ8fShDRfw0RiQGeKSt5I
QQSP449YPkW7iaqlaBq3Uyxgw5P1mAs/E/nD4UksFuZeKXWeMrNTmXZ+c+F6Xlra23doCGYfCaYn
xxolebbTY1+DGfq+dn3zgE3fVpMZ75hjPs8vUJg+ZjrFw36HWyrZbK02+7zajjcA5G8BEo6HVdRp
OA8LNArrv6bAmS+yGBLJsmKfyhLZn9FvIFZobIAxY/6u9Fg/mglUDDsSH7uMfLEoisnZaah2bnvd
lHhU6xAdsw68dAugVOWTgOM3SrqzzaPpL91nHHLJcvyaUQ3Sq0JnCcO401EaLxaOEcehUK1y4eEF
1czbI/hWXyOg+H5F8wxTQAZMd7JKkzdGLYucDtPu+CutWCyIgw/lfAfaCjMuTe680TZp0nIR9DPb
how14vDyFXiDHl5zVL2nQVAap9xUb+08E52vUvQl2/+LrY1E5RtrrSgUmQS5tuBWuQ3DV0sHOj8B
06la2GPFnvbwHR1xvg0mrCJCSz+Qr09O49QEADD7GEBd2PSl7v3i9bzB10LSGj1XSdZaDvo2msA2
xzrNObugxWk9gcEVeIN2yKpcyo6xYSXBxK7vM+UnaUE1WVIb9how0HP59nSjciVAqi8PQ8suyd4q
Gl+eLLuoaAZ+Fzv7wzjndyzbSACwLTFsLeR/yxwnphzxMdbzf45RSR3lTFRttVH3yY4ICmgDkkcC
kT5NuujfeJkJA88m48elh4r7jK6ARYPDbEWvTokajwxS3uzXmvEkqGXE+bofRy04af3VONFk7pli
3Gqtrcvo9EFgBXcEoBdkSrN+rfd9zA+ZGYnHImJPhN1UDUQaxEtz+SOKSvUOs+0+sfzJpqZwR8mf
TNv5eeJSKDNNJmUaXcbsK3OkARFZtfeVhiJNbOGTSXbvzY3no8pkf3GYQifjsfu5C51LxEsDGr1S
j0uBLMpH0SDhoLrtfMiUiOUfQcjujJOcxpsv2WDmXscTuCpg4FSuwsJkGfZHjVAM4VVGsoZMRgcr
hRdosgcHSj01FLpG+Ow/T/qXNBBXw2UVoIcd8IVa6AfoqdN7YAaWWcs4Y5NEAzxMAwkFNJ5AFUu7
KcJDYnkLe/dNFaqJ1sYZSE2a2BN2V8zrxCLileiYc82ssN0UIm18UHANWE+ma5fOwVbZ2ttmjIXf
yhAVN8ga3iDsWhZRuUhSQpptzXNrNfvvaBVJt6xwiMD/VuROOCVOJR1bXvfQynyfQMjXzaOVmdfP
p1LocILiGURomsqJfMuWxjYUAckph68GJGSygTYuioJDyGikyr7QG0qF+1ZutvPvRICViNIyGQp/
PH4ef+h36uLOg+rb3Dq8DRMU6csZ6i3inH3cYJfVvq0lf0upSL+2qSA56RMUcHGK9Q9r8OIvVScg
JlqK7RcSqk2OLVi4n57jYhGawJBPyQE79YtOI3AVLF7w7GMHgHm1zAHuTzelWadPr3A2VzdIPYoD
USWX8J6W84hyPfr1rKG+8U3f5XoowZ33iN4K3GyPXMdM0571qv/dMah5OkWZOIUwiI7Q7gwvW4ze
VRa3OkUjll5GmgfEjJuT2crWIrU9/XMKivDv3aIBWFi3a2g0RgcUZLpl2lWEfRKlE806zNYQ3i41
amGJTGHQpMR9pzRK6XcITFxBAgO7fz/QOA3ujpVbzxDwkmhj259KGdWO7Z35qqyqmJbhoNRn0N2X
CPakqgeEqHzo3Id3JRxNutYE6tRD9N/zttYCfMO/T5j95BnTHGsSvyRJ7J2fsaDbOZEXQE5k66cH
zRiNiCm1Mj2/HkNogxdw4Ct14c18QZLCK0WhovjlNpJ1kC/3v9wwdAZpHsRtr/aNMWp3xaU1++/m
5CksfTL8mdVMtYV5/2/eJ8WBm9xIQM9m5XexjgfNEdgm899pP9cU6p/YxDuoMDrkCrt8y+Uwrt1w
8jn4XAs63oxCCqhPLAOTsqRMzEOtCsAAlnfQeY9+gl06D3UIitwqqPKZE5NwfuIcpIRjEU52QC37
EQObQiiKPiyvvYizKceY6MiZI+xT8eUnqOAYM3E+JohjehGbm2qWokireWZFIFrYz6WP62//wbc1
HvXPAhvejc+JjVyUs6B3oEA1XLeO0DcR5JxYab7J76gWeqw5hm1aJ1AF9C7ctgvtnKbedMViVru1
NRoXkf28qEwS9CTTNP2K4K3f7M8AW6GxKpwBVOueG6ykwQuozuHQhhKQO0Vp4rRbIztdXfGTbEmy
RGXaYN8/v8n5I6OjvFUdxTWChlyBuOU/YfT9USyX9rS2ImiuU+yTid6x1iykx4f0XUZBnkhkBYji
2Nh58yK52B5ww+upGJmTmZiGz029ElPCLSapcYS3ef7Wk5asBGPyI99X9gCVJGzDcVwxANrhTGkE
AoA+4a3HImcf/7oN1wt5hkczohNavyueAlIVdqxjxBJig5LTRLeLa9tXqMkyG0uhXKtoBqnvT8un
s+arGWWX19q1ymGG7Dc3T3lMDQ/3KtBTHMcL6gHc8UlZVfgMIHYFzNT+Fwx/qWssqPNW5ZwQFHo/
98bWidSTOGwHP07tuo8g/K3OC7ITIjwrHXHyMcZLAOlB1XoeIoFJIIL2mo9Di+wFOLHrtvjpKvsT
8LqdhnXnuuTCz6wGITLdy0GDz7LrZbEzjANi/PpnELAgfcmNVKTVMpIFp8BIO+adCiEgyCucNIc3
sRUuGt89crb5Wpi9MdhuTdaCyI+SY1Ix2PzINd8SFQIsmgZiAhc4xcY6beR31RHZ3KlcYUnMPjgn
ooeeVgQkKgWxpUQFAVygKekdO06kDj6JmPIpRSLFc1CAMIdKLIKzd042MQkJrp5QxlBIZJUyH6FN
/mPG85uIAmGXWtvrl0HSVq7WJ00b12hgiiwmnHUIZBffMcOl+tOfl4OkaaVvfD80KsdazVdxjha3
XT+w8Mazs7FNDs7e8DvNLWwotQSMpgIdduA5H2LjAvPESzidzZoc1xzebZjU3JlgftGrfz8/f9Io
gU5zY3y72yGp8Sz8MSGR6NPUqIjz1bcjhQk6CJOWphf1HQPN+YiLCyQSjKXyWQkaW2V9WN3sJkVE
2+n1G4MG/6BKXDPg4dRudVUOMGAQvw86yikvLSflPHcI06lDFmOaWdtENaQuXK7qkDf66tlPkxfm
v7kSHyhx6ebIteV7VIGhckRryGo9eEtETY3DzCq272IZZiHaEwsl/qxbOFTDrCCL/7j1XvwCd96l
M8JsjI4SBqTbM6D/HpoiNXG7PMqnPv4g0EmcvKxO8UtN7g3m3a3rlSLIlmEp8UkuvSlqNOpTMrl/
0uK6wg+A+QckkwDtJ0uVXpt+tLWyilyKjReBG1vYB5HCuPsrIbl8ZNWbtJvraXA3hF/KmGQihSzD
6yVLgtB0DrDurf3X3+dkxCKwBKOIbzW3Rhn7apj4Vrx4aSNA9o6Ei3V61vLMxC40plPcd2kGZaim
XXg4gUYRvtXZc6zniXA6bOnXOGWv/A3i+K9MF2E9rqHWe2wZ/xdmRjO4QCOSbQ3cAFWdt80b/4T0
vTlP9kGv95CGUnOAk0yEgUAU6NQeyhOihfw+mAl4Y0FBmG4duVj76EbBGSktRp0srkp2699Dut//
beucYSsfoEGlPTkiRLq/3ZqeRz2HN0SAIdhARktjNQXHNThgANSqcZXd4EsL3+2TxD7Or7t9q18y
QbQhf2UFarYRHFH+GQVNQ1KTfCfGBktU6WLyVfiDQaH1R2K+ZSXYr8KSNthJcAaQfskaPWGMH+mY
lcDeV3vPl1RJkEdGS1XZw9er2l9WUQAgtAPlJqzYgzDXF/f6cwBnyZyL0UhkzF5oS9gT5TvKPa0S
jTl0AGYpVMu7nrYDLD51NTJ9b2+Bg6UQ3IQk9l4QAUKjuNwq0zI96VpoC4btYUbnIHgINpqcsXLt
8JEyYMj+FrOheQ9jJGsW4OEAVSfh+5XNRA91tVeWLcyOFWMJSv6dQIhJXcaepIWX9XlgZfWrgiH5
IqALt4h/GwYjnRi0A6M7joRb5BGHqSjknWi69wabzH1cig+Dza66HLVQ7i3mfmlEJKutT9Cgxpbu
z3EBpRXTm9QAl/dhb4ZayYB3GCYCcSG3ObjGjjnyJjmZdifMg7ZPLxvlsarwuDXQYAUhd8ZQ2XDD
PmyJsOKY/ETb1I4IZy/NDzWxlnKO8w0URq/XHmCQoEMMl2kdtKc1I8QRK6tHWNN/DuoSKcH1G7xH
C+v/SG4zSInJEXYdS81sJf7a5MzyAGjOgmeYANLu0rdBQQPPrcVvYsFfXrCF3lslx365DPHNfZ8r
Iw9TXHYm9A5/cz9cT9/HdzfYtLahEqZBHJsID1bUiH0rM4t4AzFc/VL/V910doxtGP2j4TiEAZ6X
0ijfSy9djd1UxlmtP6pi36wtBbq8alzZ9JTI+5kt5YdWGowoJ73tQISrYHVgaUFUMS9t7B9KN5AQ
TFpsf1AIwvNPV4Mon8A1Jt/91GfHGYDg3pMr+SNap1wFFq9Cfp9WvCVzMYso/Fbx9Gxsl5A3tVGb
G0sYYLO6eYyEei8wrIR1yvwhEo2MbCW/SEaYfPNfnC9vkXKEtqMgw4pHWPCk7/FC5k6Oe2yJo0qT
Atkfv9brtF0FVOlkvWBxbAci2EEHuzvLfYVdJxyrK9bzVu9wZ66FAUQ5xP5M9zbfFbecxflUijd6
6ETGj3PZhTfZR5xgr6bzrTTMt63azAjqKFnPEaNTiJLr07t8K+yqYiP5kmp/FPEw+s+VMNt4SoQF
hJsKY4wecjWHOu6ajroJI5/s11rc+ymvwMWPWkzeg3nCC866tuE4ieevgul5Hta5oyrXKcOW5VC9
wWL+PRnPjNNAP9pAiZx1GvSmAjW31toTA+hME1FYc/Jg7ZB0GtehT5vcggVkrRgJ4I5voJHaaS6Q
nvzwlHDCJFiYtrsUMjdYKOl0cPYX9MMc6QGSejlLmkKjfo8EreoyveeYfOBCbXCzdf3l/UpTUPUf
V/zWPt2MtetMOzwEasPuFC0MopSmZqRLY3jJqVRW59LWBFnhRUJHRUDQnboqy5srwBtBsWN1IPcp
y9I6YhYQV2o8J8hcKQmUWs0eHKSfDv9TcoY5GhSFKfUbYKbnYujs+643ju6NxqR12jVuv0j6jQqe
0HLi04Hv8GQsHetkrGuQaSr5fR04S0s/oSjdi89BaehlXS3ut+03DPX0LArs3ivF2sd16JKgRIDS
kABiXwmUEcRPW4qMO/sor2KziNxHWj2X2cNd2nl1DseGq6EzG4VXZQ5js6O1dk+H8BFd4JfpHSCD
4Do2+5MEr7v8Z38+W9adIE1YimxMUpF18srlLUC1JJf6GW2CruQQ6hnyNgRXdHHJt6E7gTWusSdD
UNv6cB3iM+DAsqK90j+u9iVSU/BloyCTVZj9U1/wFdfSXkwJEMcyq/p5JWU5OVyl+IFIbLtHgGRo
McWjxF3OaZczxHvr/bE+L+xhqyNOXld8bZS1K19qbVfOQxcRLviot7GSwmPD2K4TwpnvbBwErWhh
4or5u5VU7Tgnog0Y+AlqGyk7tfCbqLXlvnjh/qvlciaG63jWJlMA+I6VXHGjl5vikpjeGH1wdVl4
u09BFxpK23WQCDZ9w8WyxYL1VJexC5BpKSbTIXWC9+NiB9dD4A3OpT2378jBUvms9f8pFF96po8C
DVLaz5AUiH0dE/iNlkXpdF1/DA12fcLhsnBeZmHVZ3zwAP9n8AeGD34tTI2x1L6afkkqemvlxQnM
2nfWtNuolk8mUgcgZNl00tmQyneU7z9zf5aQfmfL5E+1ebMPgCfFcp0kBttOdV2dHKu8drSgYgBI
jgka+hbLp5wAkHJ4LnrRJnEKmLYBS86HAE/PpDOLgtRqB4vowq7c7ia24fdv5BtcR4/hxUMpKcka
pCkuoicp84VzVcdEfP1oI6su5fHyI0TeV5wPC4Ol3OlZnt/qvW76hF1lVDaomvRDhoVpXK+7JCOd
ylnFpfPWH10UVcF+LGn2WfNQjhF0ydLyXA0fInN31UO8NHHvA0qfhEAENh40aSIJ0cbUzCMHXDFZ
PyZqF/KNT5gvYLWW+TKmSWga4L6aj0XblsZ8ijWA5Fv7wfc78cAPTOG33kpss448ikQ+FKp0GmaN
AXlwVhOSTwyUJYL1suP3fyHqPz40jtZV3IO2oEl/iV3/MQd2Vc3fFwt+o/r6LxZRRxxYirPDzXkv
aCuUNmMciytWihyY7emZwiG3MILBYpH9t+ceg5NHslbY7Za19MYyQkygo2i8hsFksgKf/K9wJaBK
4Mw4pGo8h54iZ273W7gEAk7VrYHtdQ/ZczyX+BJBhQSopFbwi00pL9ra4s2MVH5LZn3ceVBjNbSy
LihA7jY3a9/q3VEqb9i4i/PitfNcQAMBwxQddwPBTIWdEZm+g3e6UiXZe1wFySL58BtouysVU6CH
AqLRzEqn83qvKkNjhKbydQJouY248V+QgNfLHIGTH/qcljj66fh9EXuBlKX0CmA6p63H7Gyfivm9
oVscGaZsdqtItQNwTg6uYa2bL12kiae1d1Yd/7TjKCkb1LhGNUuxDEQ8mch6VIByv2ox7iWZWqH7
OgkR0wn95EGGD9W87T6VAFyMDUp98jDFAgNXusL7mKGklPwZuNjDyugeXLwx3jJsgDUQO9zShKSG
A6vk50WAz6PGaSaS6ni6ECtaOxxMrhwGDVbZs+4GdnqkDFGHRHj6Wi/Nxt9cxAqVlEwiViUE0QVL
NCgg/CT03ZV75Hr/Ru+2MjO+E4bOxs2H8sfmAKid40hPNm15EQZmZ6JGB4AbJWph1aVovL7E9it5
UgqAQdkkK42/iT/37qTayo8i8e1SyUTcDIWQruSb9VcYMkBIXi+t//r2e1hZM0e7D4LzofYNdPv9
+kkThjp3mLHySJeoLcbpf8ZXPzr1hqSp8awHfkeMStRQL5qswsRkx7IyogtFXB5eW4C64yAqxAlS
539QDuQokmWQ7XR6gxLqFJiVyJZ6XJAQQlsjEbRLgEUC8YONtg9K8tEsSLd05OWEuq69FHkOPGbb
7ksUqAc0UVGgQjf+mAhPcdhSOwIeS6JpgLku79NDbLPfjTY6Qoxf6P0xxQ0h2FzFiUPHirJMzySk
jQyFE3dY5Lra3ZxmH4T6rnZYqBn8fpepkGlJVbQBHncq14lZdDsx2/Q1MoEaeNUaP4NnCFA0sUQh
OlaYGCQB/ms08hhkPNDCGyKjj5p+nrzyKU1V5nho8Zfaw5uwsJMFQNzEOFVCnyQIMDlHdKkwm/qu
l08Th/xEW7ySCW+8TyXB+LPrWFlHZhUHmNPXMrl4/x/mXRRsoQIIVP7OosHAcsrZjeZrgw3LHxVO
iDVgVIjR2rcD14zeMrPWQ5l7eLWm3KbwrMEfdcheeVXIG88WDP9B4SOOE2F59DU1ufoMI+6Uyx0i
dJLPg7VlHv8aBSoilzg0r/cXvvAfZBxIQjhTK/KmBLTEp9/Vp4gdtVl0ejAZB5lE9dMkoE01gWvR
d9ofH7WvennX7NsiMLlI/mLy8pG2ItP5JFVQwosa5bGcc3g9KAkAWICBdkz1XmuTCed4Qq+Cv1LH
c8tAumboRRBwApa3Pg7he/37EK/uQcaOAlhKPSaVpF6NbDn7Tr4NhlHE4VNUzsdvbvqIUs4UfXLm
d8V3DJXT/oCwTVlOt8D2TiprIX7NsyK35G81t6shZMBr/zjhnCO60GFJgY1rDST+69I/TJ0qP204
pQXo2ontZutQfosSp3J7uFuHV7VYNoFw9FN3W9yiHKuWpjkdcl0jV1vWC8AAEk+9naGzz/UV/0M1
vpwpeeFOXhNgbZFqxXujmxHUMHBMs1Q0c6BRAlzw7Kv3tXh03nqC/vN3SRgJQqzIeUhFsG5ghkAk
JxSznxdnCP45kKi8OXAS1Y1T36w0C5udvpHKXDi88oC8b5UstHW1Bi+Xq7C9wl7vL5Y/Z9f4Ffvu
Pfp0BeSQuxeiIcRSQFy9ZtbScpPrP8Xgpi5/7zmBq9YZYLJEXPb40so2bS2R9gtIRjF/tTI31azj
Yo9bAxTe/d2ypb/GwAJz3s/33iC39xzMH3esVumqYPxNoWd3otTXWPpEB4rqll9seBRJa7DALOCw
k+gmoUu2AKjimck2IUoTMi/61K89zzPYWLsHcZ+uo33uEN/ILenbdJLopYSRWUzudyw0hrX8E1ZL
WhPbsSIsg45GwLolm16JWVMozDxc00aCIhD1OpMVGVuNFgSn9ZpQ6iB0vWvpJ+jEeQzuyJgY7TxT
H2wbkU1aLrWmgvDrGVE0X9/3/QEX0es15x4f+c9uW6I8bn2TTVY5dYnZj909A974FVb9Cntz7Xg0
TIJNSQNczEVB8gIr12SDJe1hsrmNAxuhyPc5oZFRjF3xBv2Ji+XTMyIjv+kB0Xc/HwThWGkj5tLJ
F6AmS2KimJMohg44lsrLY1wyrhsWnyIIH3cLdj7yMgXx5XcTAQdq5A0AVbg/ln0PdGZsjztX/p5c
eeNRUKWvgSZwpMqzymaSow1feaVGU4jITH5ME4RbQEqashc0399+vutJRcoWxyYjjfUolaxhNofO
3qZ0NuG+JC+LydQQBmeZgSgH6mX5uP+mYgUStTxna6uhhCoIGUx7Wrj9BA8a9/XKvFDiUczne12G
Hke/Yibs1gDvAWX7PhpqxGUgquc/VfbCGvANCUXc2WwFAxg94iuSrGkZ0wVuJYQ2BcLayTi7XoaI
AWA6GnHjbJhkYFNxtTQel1vUA6xu2+rSJv4shqe2pC/gKWFHlR/+/yKIMPCZeDsIH5D1lhbPuTKj
MKmewLVBg+7sirZcVtGWa65cIFkesLcKrZPNo/NapXN75b45ODV1JIojG1T5L+O3YtB8d7wkY3Lw
eWOrlNwc67UwJ1cGLMu/MnNDQjabYjfsaZGPHJK3Ges2d8gDsxl4V7I2YfiuNKqyGtzKKWHaMubs
6RBdNoIYzU+5E964+2ukHiKeoujEN07GCaX/mq79ADwNtM1imSoewnnqRBBCX9GPygh84zHUlKLU
S/1YBT8we8+hXc6y059/MNNfvWqewq9SRJyTcGqrVvpgo8D/RzOG/nilyVCme+cL1dBGVuFXLIQK
qRGoKxVaDyZEA9A5KdF/r+ZOh1P1stbFdIN8FMXia9MMErH9o94qCV3Fnshs5s6aeDn9Yx0prUfX
Z/mP/3bV7QTS8hgCm74/GCHXv9N+wORkscyo01NGFSJO6eLuGx1Pu+cwmQxOZsytqT396N74aYTi
qJXdW7UWrgggytc0xdtP+LKTzgMFlsxVocdi1Goy757eWintTx0jgPu2E18RvfehjCiOWUJFqpBg
65B+znivZsGvxKiEisagaimzsoV3STcevjGVwPc5OoM5y5+8OwJ7izOjjClCM4CNIaWTat8upeyj
dF2kGJkWEOR6FwmYaccBIvs1rWgyG6uhJCFROO06ptAgzaCLxsIGWSm34Qo4Et0gPlvN+VSILZT3
iFPnFv4W0062GwQCrJBqFHYXQZe1BSdTIOQ464bGRK5mA/ZAG6Pz4G/ix/aCFJHNuZR+XeCDsPIr
wlqNAsgnOcVI4L3GW2z0vpmVu0aWTcafA0yFjj+rDGdxBive03LVn3uoG6iGuqC43cHWtUkV5mZE
oGoGqO8rbY6o5gJC5oh0543ZGXYh0U/Sc0yJyWBXLm8zFArfu+s6OiRWDHkecxk6xjQ5f05TUeEP
DOuPotlQMhagSOcAuxJlnGeEutD/cbj+i3NYE+EhWEzCmoQYen8KVFYGCnpM/ceA6pzyBlZVC1QK
lfTALzPft7szFpfkv2zyHxUjMElp3PTS+yeaGghgMDjBc7ICXMbKo8rRb0KZc7osdLOeGD4Ju7jV
LFbR+Afu8OBtJ5OBJ0HuRwmJTDdvFSCPr7+hMt/mU2IOpjWHyzqPHyrFj3oEBczmPfGditPK5TQW
M9TbaLVhQcSDy7RK0oyTzQcsGAOW/SbCUyp47uuFrsF/aTDIzJWqbD0V9Jjuh05BqXzOqqJFDMhO
hTmgpuB8EDJY9zFWscTZsJxJO6Qrla82sIrGjVLrGNEuqw5XY+fyPZ+hETs0Rg47WwASAxVtfKF4
sTq0uF/yn3cbqlq2M6/BxkDL5DvW2na0Dn4Q0UxD/uBXbuKSAgAscL2M8tH/aOuTkEN0ZXlwtpCN
toIUMlKtPF22kR9DGEpXlljJvQF361GePp3rYe3QfbmF+W9QvAyOFl2rRfmRjVhybPdBjs5P/l7I
gzXxrkHESuzgXhO/dgW95VLvMr4s4N5JBsbDyJYuSfuRgnxra4f6DSxRMZwfwLdARd9nVnS72AtE
ytVeD77cYVoZxVnrz20v0lv8P5339wv0MsH7dR8v1Vqlbs1MjZCrJor2QpxdHjc1pOh/tKW70tzA
B4swDQszT4kmexp82OI0MPMXEP2OlMz+3qt5cYdY18TJkoYKdzSveZpnsKU5E1cDHZUuSqeFfcId
ZwPfp2e3nJ3qCsylr6JqQLZvYsOjQxu9BTkaEjcm1HN4qTHrRMi7dvof3pksxZ3LsI/eMI1LeDNL
wOiwChiTFBmk7uZgJL8YwwFTaqJQyKxjLKKaNfQnXmX9NxRgQY/7Dj/VlPBdlO5WQjMHrQwLtpWL
S+D+AjMx91Stx8TfiQWrGWCRrpPEB0RK/M3YVKulVdcGiJGHpkP65ldHYKkjJP2YUl4qyT4lCDdg
e+5f30zla3vxT95azA49FVdldqBpj3Nd2qOf8Pst8ljg2D+pCi9mZ8MK0WPSPysLFhmuhL6ZWAq2
QuBArCQ6giMooTpm1lgJxmoe/Zi6KhXVYpYdR1SFeD6z5K58n2RGW6t9X6X8Z4IqFtA6ZL2rnqG5
9JNa45kraB/1sC0nx1NO84JCw/TfZkfVFBjasBT0i3OfxbyKRRml9hBEbgwtSn9Lj2/EVKWDtB2l
+C0lVQqyKrVPCIRtTlGgo3XfkmNDnN3W/8/3CsDNBEt6F73fQbLW+xM92ZPp+geuAXex44/taRbO
KLDeXH9bhRz/aaZwc5O25OTmIsfVMikOWmqbLusqNkz5q2p1I9xG6LTHc+QTXBRB2jbsDB89m1Xy
OsO8iA5M7/Za9+qfvRF1bSCJGdoALBXmwZtKDp9SrEWyWAIuU+MxaPsUh4owae+9vTjzKPtcLpgR
StMRVaQ1cI6q2Z94ixmim4RMjeoFHoQPq8Gw2i+4y1BMIJzWjUvERV/VzNZt+k+RfhlHGZXTlc1g
dEfixXXOEgT4/GT+v2NAoIVVHL3MZZuUNYTgiSzp6jepXLImoyPrQrGfCJXIfRckmKSquCsnm8Rl
QSLuhrvGd9omai6UljomK1YQsoI2Y4yjAmyomT8gstAwSclZ3HViUqi3tRWA4dE6Sni+BhymoqKw
wHMC30KwY0ryLZLMgx7xC7gLmDnPXSOXYBVTzYjxzWFnEC9+Td6UtuNbImAuXWRTmpPsAcSqBJJY
J01DrWkmmbZKjZnuD4+SfZ3XSlAwFXcDObpNdyvWcUdP3NT/pGmYz0lnSUE3nLnCr2tbShM4Xgb1
leG9Gu/a1QyUi5tEBVMBqkBKvqygAaYAWiNAN0+U8d2P04ySEPWF01gFBASxxgrBf1BixCaZUl+k
/58g9kpt0yoGLe4Kqyv3uuUXyKR5M98z6O57UJETr7E/hvRxx11cyY71MmMb9F5jzfFS0M+fDn15
SRNTfGKJBZ6LnMmFP8B3w4dTktEQwOiri5CEFuqgEDYMqs4+GiVwxykGjtoZy3V0+A4iFUoZh7Si
Jdqni00dv5jq2gjJ3MTotHyym2h9fM+IyjFiaX4zMsAOUDXKmjbIgaMNN/jlitTBq9K06dIadAes
tR/JAWq2SfnxT6enDEcJNUFosmRWqmLTmXJH6YLy0njN7VzIcKjysmNeMvFBG79YoMgWBabkU9x8
bkJ1JScZqGvAftLb7GYzkjedOzi4Q5PETbDTZlA1gR8cNVDePsCbJIkQNA/PqbHqmoiMoKbM7GEB
fZb0zUdHCr74ZuWEgr6EP5GYyyeSCPUfJG5k2/ifQKxdVC/kvW9657Os5jWxQLwqqZMtgwqocy/g
wpuATz7jIJFzHZvFfi6mEyfUSb/dr8Gjixn4kjZgvYD85jUEQdFeBXr3RNGNH7xC/+mEIvY3ld1u
zhPVVzDtYqkMJzLNKYpqKHYPXea/4gF602MWqqN8ldQzxQSmK6gK0mUujrtFzzrnk2D8nAbdrUWs
BFeha7YpKZSCEzF0H4CsrOkSv+gGrkOBjrg22PwUsZzfi+SyZjce0cpg+KVnlgGuHwntWteiftXE
vsshbZ86LHFrHLkqB+S0cN7ItXViyJJ0AcnGE6doIrEowYQdsORoBKLVRR9BxcC0P7fLdUE+Dhsy
eq0en4aB07FW2esD3YTQcZlUYoceCiguY1HAr5AI9Gz3irEefrBXzaVnXr2/iClzeKCD0yDMGI1Z
vl+hZCtmRDiwzVh4ESnw7w2JfnR1xaR1FEytl2sb3OlaVF+v0R7lLToXiYo5lHQZEHDtQl4RRCDo
IklV2ehftNMsREcvpnYddpka33ZurE2w4vjIi6fGlnjYAqkCaln9OTxXIfVdTYcPLuPxIeQdEUpi
upazC1gsXbXSMfSS3A1kT8iGieu62nsC4+d4NT2QUTRBwRkA+JdBxdz2hhIg2FYvqP8sDdRgkpoJ
ojOgilDwbHeH5H5DJcvqCIAWo2pjjE//+rj7Z6Us2RVK0JfG+cinFFUgzN3IHEvrWv5I00e59hmp
n1Uckdq+vJ5AHXr5boRZ019GP4Y8pmOmKseK0jgPBNgpFcNySGa/mFDz649Bl2bPCbGX9jzb5QIQ
cRkR+eId2Q1UML1vOjkqgvDNhI0z584kXgwH7cvI4tx/7pjSBVTlBEUU9UYmnQ6tyw3ZR//Cwl8Z
gdADsGNp2n7P6QQM5IoNX5ru4a6Axxc5toiayvGgdoGTGU49iN4XMMAJHecY52scsfHnJ7cxH0Y5
nKXmsmr6fYIdt8ZTQarB32T4xwiLzvC6uyLSo2xaxTz1/gPnURc72CHVkFPn3qgnJBe9c9hFH/Le
KjheZjDgmLKhvaP+6YcxbVOa9NhSt3vOcEGbjOi8AiFQTWfAt4/YefNjZJ3CIno6b936CqX2Lk/K
snGee83HE5pdVjbHv4yXV2/2JETA2D8hp3BbnbtkxV6ksv3TtazqE8N0p2o2Ssm48pDeeujc6N0t
0n0tfNSH5uQ/JGexnmfMf6WRGKUI6aNKL+zpUL3Idfu5jnKZcyoXkCiMO1+8q+ZbyUSjtr52EhX1
GyV+oRp0LQNn3hEs5YKaZ/Qih6/o4IP2WZDyFAS4k6Zt8ttvEsv0BkZKZP06muQxJh0jyinL6TsB
O2KUMZ4tammd1N4Jzja859GnxuTUNZMNcpgs2EY4Gf88YZkhDMtqPvgCmolVOfsQMYVSS8Un5N+Z
ndZO+pb5bsiXFMNDsjsPFGRh/xP0DAUIumbQ3+CT8OyVygTtQGmyUhMeCBTYsIUcES6YwJnvz+Ih
gMW3AxpL8QyojE8g8aQ16gAWHUZsxVgaHOBfslLa+EjD5gHJxKMW1xTPgS5mJYGdaoNCGh1RsJGw
FhWhDf45cVabcX0hKmltz8mDf2FMl4fVBUZVo/CaEBUlVnfstdddByZIQMCAKiK8sjUeQkyDP0yC
W/VNskrBAKVzUEwl9uJHsf9MnBQDtM4coFCAdKYmoZhgn3KlamzB+ekV3Cdkc8vsBG/j0pkuEqfF
QU1l9RuDKq8qwFnE3/V+9HHOIbY5+2BxgTRVBzaKcjAU+hkJZIVu0Y1vZOQahoWShDePEtolFLWn
UxlK6LAg3UlRKBGhXuPri3MtNb+7pAN8ntfeLXpZFGX7GvTk4BQrdq0UVC38Xho8AWFQlHxjob8R
jOWKPAifs3YXZJ4QqwmHPRBTrJk0k275hPhrtOfdGn0s2uSyyNKufjfpfckKpp5VV3+knulkpoir
6yl38kr6dRhzyvUrLVKcKMd7OytqoX2Wux6JDcxRXQ/ZhOGFeFV418p0pQBUvFwjE5OleN5q/dfI
ge/TGO8FW0m+uQAaPWv531G8FzHfijR5QDWX3WcbbI6CPF0oUkBHjRHdwhwSE64zjQE7TnPIXCR1
21SGjmZB9Qjho4drTyW1enHySYQoTDREEbE8OoJQO3aiJRIlzX4fUSZP4b3VCHjtIrMQiL+Wz6Hf
IZAAU+eZpQH2cZttC7Tf4BDlmdyS6kLePXBZ2NfUoQgjliHZHSmqCxYkudvX+H0L3xwCY/9zWi8U
+Wn88z2S9gXeH4QCRh033KXOjojtK97M8nV3kZ8o/8ryzVv0TQOrP1PXWE1HSWEULbGivSUIWXpX
GkxufMkkrKp5k/I4ODUHX9dijG5egDMLZUPrQaGyPSJQwHBNKGBsUypJ1+IfVJaAextLvOpVC4Cd
MnAz+WoDtq8HBIJiVxUwi68TVv/sNuocOkWNQhpi0u5WKhS3brRY0ycnFxSSHbA5upVwm+clEwZL
YX5e+Txo+mULw6Vw1FUAVY70VOVB6LdseFNtFDd3mtv5+e3r2/HY4fpqYKeaBXwUbJ2kuhSZGKOQ
KzTfh4K9COc3i/fnpuqD04inksS9C4LQmfb3QOGJrHwcZ9aOkK/ZGLQwzduXJWkKbSmXV0MEYAW/
U4+2olFDRFnTLMRPvG9tD8y7NRHNVK/aWGlrsY2nzVnSHxfLrLF+f8IbgMF51TFa6nrBwrRz9DAz
hQF4q2yqHoS28/WW04460QuinjUd6Ko9SDOGMZ4qzP/SmfAvq4bySq2lc6lhaQdfDWpu841R8r8W
wiOLT6/7CVM1fq/GWIgGkxD7NASoVkeoYNBaRKfXJaJCm7og4BoUf0m01UbD2o3AYoSgPjn2afMo
6yZGeJV1sqkpjb8Hl2z7NUbAF44uDWuEnu+6EDxxYJ23PsWkU/fHq1oP4H5uYZ96ExRMQ8xs+Ivh
0z5KITl+bLdDFE+Q4m/KmlDqcl0cG+Z0iExLG0jHspwodxhfOY/xpaQI6QL3oaARDf8MVV8H0xBg
zWCZ72CIlmLZ9qV8LzfDkP4Q+2pv5dgI60Ac9aki6zwCM3Hdn8pqbKuHJ4SsNzJORARG0HTdqJkD
H+PgVR+vUAEDkWeIfb2FJWbazlx9yql6H2Rpav5zD2HH943n6HYLL2GFw2ZsgTQ0GKh6iyw1K7AB
SXeUm5ir9F0AjXdR/HSOmNxiSBV4xy5d4vQ1jAzj5NdF1rQZvyAuXYCJogntDGEA50GPAn7dtCeJ
GLhNF3PSmCnLIF+gxcmV71krshWUooQtYoISWjxF+29s5L5+qBTfi1unH4m9qAdTaCUqQgWe5mvY
LyOZ+Ym/YLugNSTIkLD9SPQFjpRR7UMk4gS734LxHo0TqBcbyGbM7SpICp36n5BhzyF0FwWuWSyP
AM35B1C4ohkTu4H/BT6H+K3SfChtuEXBCBs6yrRD4GCif5vHawOVAXsrdsd9RejfB8yyMdgz7O28
66M6nKDIkopvsY3iIOdnoHwUXa5gXGzn7lNs4znYynYLrDCj5TN3Lh4vo56C8Rj/lg3Ud/QmzpUT
ijZ/aZaigBrPihZoeaJcJyZvUSZcG/1oZEWmFsk2X4e8FpXVqr8xCE3cAs5Hd30eMdlDN8+3+tks
K8uS+mzvfORE1dtj/iGYSnQwE4+Vh+fpx6ZaSxXNFYZzl2jwGBbtV6WxFFT4RfWODOgPsmBmfMqD
kRLeIzZ+huR5VGIdfxo095/fzMgN/+FbGGhflMKjr3q8idPNoTpCH+v71LRfrCPCfpaPHDAr+3Qh
SwPv2aFim6elRPJ5+xKnDdNm2+nq4mxcBG0t0JZQV234p2JSbwO3CXfaGQKqm8yt9Wc83x6g/vqh
QKcYrxRlw/cCRath2oIvhzdF0QrBmao0AY8AyxttsV5VlmsWHno4TYSw6fGItnwe8hJsQcXPQbxf
7KDWYehKv7JeArLY04K6kWbSdcKZcRRTLl+AnR2XB0RO5Ig4tQFYtHGauh5CpTaearO0pOxnjNQr
MDD0dtxsJ7xSKZPhZ8lLbcOAFaIwroi3wPh5M941xERc2Enuv9NWt+RGA/jxFLHM0VcokJfEthKG
Z7E9ddXRWA8mEtE+17iTKreoqhkig69R9iOxoQHz5NNndca8LnM1FDCyuZXGcoyliTIZhdxUfUD1
oY0tU92Zb/NYuw5Y0d+G8br9cN4y8FKWfJWC+KnwZdc9VHRcgLqn8gsjx7egiK/zjudUIa9q5R6H
JcRaY5TXLj3kcJhqhxiYbuD/hCIMZ5z9Wo6snMNq7utGdh272OfYr8471LYdzJH7pGYGMGSMMmtI
i5/TiCABgV6675GL8lyfYHFUQARozC/+3rDIrE6aUwdh9Q8jRjNFuqDh38WPJKkRirsNjPilgdg2
VQZMzrbr85mVQOdWFMnAaxKpLYldbsqoV7ItRbiTh3oPXwP58k6ky+GULFL5I57cd9SjglE8oTVX
J7XiYJPDbXgG2/pNqDdv6CuMAmgZbFgPR5B/7XjWZwRomzmx2yNkF0ROoScqhgKEqeoXzKYG1X4B
VEiYc9ou+LPdzWbNrHW03RaPscyD4I2dB4sEEk06WvY6LIhlEiCH0U4ToQBYQKqYNj9e6NL25zRF
4Mixylhn0XQiBqKlSDhnLxrynrT5B+k+h++o/TLT8/tqAf/W0jOK751+6caQJjkKxduBiRtDONFd
khIGBH3ICTS/nifF6JrTajtJn03vIeA06fsA3ddrx72eq1ZLvyvhdn5QIg18yA6nRe/5y2lP5Fe4
G0ESL5SwQ96NYQ90HDeoTE6RylP333cOEfeW9DEXR1nq8FX6imRXBjybQcNlNx9/A3vYrjG1pfCD
5ccdwYSL3Nr5BzHo04Dh1V9C2P74NGh9J9tX50lJdEXlpjCkF9hXZojMUCQS1IfM50cou4Mnuad2
3TmHlDKikEQC+TPBVy1Cq5rwWVRbQ0tjbe6RfBnGVOZFW7kjYkEI+ALydCMLgMMbkzvW3wvion+P
B4v6r4VdhF+9vfEgvvCofFQGB9s6Shu/tSM8+HVgbJaWnKwevL6+OEHnQTeK9lRruvFP947J4PvL
ZWQLDq8/9gKvOcDV9k5cqU+ElGamPlb71S/CLMDASb8PXwq2Rwl0AnIrYKuchHKqTtSjXwdY47Tr
5rcZY5UGp8+UFOn2ktpr6hgyRanoOHETNZq2z0BLA3hYLq0RmSdKUaVQu2NgKRWCTiLLcKRHjlq2
hFw9D+1F/w07A5TXdZWIho5boGRkZvMXSncspiHXXnvZ+2ei+rZplGVqBJE01a1pec1L8hLcTVgy
hT01w8eALIixP4eYXyZvNF50XBF2QU71CTls8CUPHIRGamya+sBLL99ZdspCOxS4lRoi/u019Er2
DUMnKL1npD3N8tlw5xs/VSGtTzHXlgjhFoaVzPlAtGJTrF0cinhiGzV6SJByxZz48UT02O1A2V/F
mhYXAmY1n0NOwU0qgGFh5ozAC6u3ECTb/IP6ABPpBbWcHEhSzW/NLBZe9MdsrL8TI3tyGITH7jqv
PWRTayaRkBl34twcF55NtD2M1s2cZDUnDu48I1/bItMet5md/tg/nsYTEdHDE8z62AaOMCmMUpE6
yqwR+JhpF8XJxRMyX0tnLbqv00z26vyXWF9BNH9hxdSpZhHpwGqu3b7erq/Wik5Q5stdSZAlQ7fV
2rrXEMabbOhIhixVZy09XYhrNPwlmp2oTuaahNF8Q3BbMM7AKmq/uYEjRmZY2Vnz5gGuqbl+NUgu
C+V/eSFE9gBdkBjlcGHt9cmUd6wouePY8+y7Mh1zWykg9uBJGsR5tw8i+HlPzE5O8vsNKPYOqP+Q
8NJ8Spz/R1UbwUJctHNIjie2abxnLWmEyO80rndswPLuM+Otok2Us7voRqIv1PN3oMrczcRP7c2Z
M6CvQuI31+6h72TiadX2svkPybp8NiBHnOYw8sgleYnsP52QeK+UZtnF+tNbIJ+gyk9mef/+NcyY
dvad8M7kRb94kq0GLiBeqPZulHUyTEdKODUGKG1nBG7U+F0Q6rR3YFuP2NxAY0OpTp4L1rnpxjqm
ppxi3HFH862kFbYEWytv+hVcwJFSxQzxH4qSznetwP185D8fDUCW2miWwdlNAPzRcq99dttHdTGy
zK3Ni1uYUd/z+sBmNgrH1kTC9sLJFEjddtJg2IodHk5qY7OtOKG72MiSksUuFv9f6MXE5G62KrQu
AD6OlU4UG6tY8R3R46r3sSHtbjySlmJ6DE9/EeYP4PBsXi1bc1kAdbCUWDFN5EVweViXzvBGP26D
KvI2Hz+YwjpNYU8N2/l86GGpH5vW+tBVh5ESb7Ynb4pSmHmXa/UBEcOww1DHbbDB3NyaU5nLe7ey
fVHAyHx3M5cI2JuyFkO+67QVfDcUTRC0SCl26LYkE9lIWk8R9oQDCoxJWkctEVzoL9cH5KIpi3sN
UvSAzE29phRrUAzCzsqqrvmYFU1TjZ23otFS4Q74Bj8+rb67IZkFNpziPJoOLkJuMIcrVHzxtHS6
9B+HtLD6ZTEk0Q13jn1TKWtJ/9WAWsEdNpUWc/EvCLsS40EbnkIJZbbtqL8ex2yTSb2GL+afpP6H
b8X0Ei+ft0mwKl2rhN+nhTil5wxMKf5z7Xy4bh4I2ABlDC/kbY1Q0W59ADtcemFI/TNod4tHm71g
e0/kbZUqsfEHHYS6Tt/d77WCqvQxgHBnIPvEAkO3p9VavckfMFX05ctuCnP8ILla0yCgcPrYGFNb
3/Hch4+ImCoTl6pS6VVT1BTVjqmNrTKy+fzBQZ01bcN069eiW23NguNLrZlTo8BS3r7QzraCejGX
eM732f8wjgNGd9/Z4TVlxqGNHL4uSIP3qFp6FZfZrHeY2ELUGhTh858PVgi+0jBDB9rBBQMzxurh
KL8PyBbpQrfwmbEw5AuQWvIxbymdZJB3j6/rJ3h+uNnwVIzfhrwJirFAVnHbbk5WTLQhnSKFi80f
T1eVXQUHCRF+7NM3czeOLpSoUCgfIPnSJoont2M7J7gjkkoTfsbnHfyBNAhdkrSCV/PEjuEMqOlI
rx8/gkBudlmOdvrsW90kGbGAC6LaHeddQihsCZA+5lqt57ziI82JT4qpB8UtUK1SSZPWl3FPt9dm
Ybdt1OYVyS9jb8l7bFWhz5qC1kepij9ZWSj5M4DWgYsShoNsMPJUxpuEXinEo3IsOmZG0/IUdOOZ
R/5z0GyZS30RVgrLY1vzvLMCaA+CjGCjNzln8V2hDR6ULoaQJXmrhnI3djfEuizwMDBOa80pYHiD
UH9tvHSGOC10JG40CeOW0thqLuIwck81Y/O+W21jr/tiV5lO1g3U3P9dfu84z7O9e1Y0w2W0G/Y7
33VtG44lBaLWwXK4yxSGRC425+0YJj4fA66lXEQJ8FdFooSx0X/jUmG2sX+6iYnxL9EcDwyr5m8U
UckQC6hRQFpmAw1BExxe66z3HXX/O76mf7eaWU7krrWj59eJIMulLCUXv8UHr7kHC+L7op7vSjzc
tzySzQgk6zCe/frmi1D2b4B6N6HgxTwUFrEmnjIT9bB+WaJ33eP5+Irw/W2lEfyr1yOYXOeZCsOF
9uULcg1kLCCHAqLZzRpgRA1g6UhAkC1wHj8j1hSg+QOGJHU1XTDpbFRLaD9SeXmcrgMdYKWFMIyo
O0nf7y9onZ3Y5ML2bc0vLgeeomVnzheitbE1WP76s9gM3ePZTSc2HixHBTvEkZm3mkE+uoHdwNna
vZ9p5fQ8kS38C5g7ZLC6/h5I+M+l96ksM96EZa8xkMOWtXCqdRCRRk6KvN8rHSJ7osdEV4lgzMhR
6rT8znOeZxyA81zLqicwEnl9p0DccT56o1P2k3qlVpEijhTSbDJHsDc77ZXz0dWhd/2FcayCKR6Z
VRyYD5juwmRrR7PFf2DvpgQK8ua1qHS4/O1WmVAEah2I3OE+VyDJW5Dnv8JJqHPDFA23JV7h7hG7
13MOa1B0z3IXgbnsOVgecM3yrSMV8ade71sVj6z5xo/SLyJRTAkE7cyPGyqnmIFHOCF2leTJ/G1m
m+iZZrXrEgy6r0o+RwBG+IsxzqO4sHEmJ1Az3uoQq00WyGOev1DBfAI5AsGc3U1cYxVOV8R/Bthm
yOhHAl8NF5r/zjy2KTU/dlnvfPkB40QzLNMnTebrh15c3l7VThyPFBbLAFDJUQOeBcFYMe/ktKsM
SRsbXz8FFPc4q9kCbRG+6cz8NXflavSnhC/q/JP9o0sLaGdZjy8JRQnAHZYjA1ihYsmUqnFJqlTP
FsZJMhJzwQfmgtUUdwTQ4o6d+aoe7ONP3aoSC6fEvYgZzkYpoAsKHY1W6E90y8qRRkNBkvqcSbYv
auMM4q5juFKIEuRnO7k52xfiPqETFMVxML+Esp2svozyeNJ1l5dw2gM+/WqzKuRmlooKiRA/8tPn
yrqW4F6Wtkcfkdh8nzs25B99Y+5H+Q3+HuyHyLWcIVdHp8h/nIGGWAbZaW7IUE+AP3BYcESLK0CA
MtGcJD2pFy+zr4fykifEffTiEhYMy7QPQhuJlqjoRSmTLpiQXxb2IkM4uQo18zgmiRb04NX2UwVo
jQ1Dor2bxJ0HqIeCerV9pn/bob6HZjCc3QKaIyMHZUPw454PQxk1mrJxVKPAyVNhLTBDNPcezcsq
pXyVJTGdSxuUhf4gZgiQS9llzolanLG+ThkjKqE45Lk0BQHG6u1OsHgdVZuznLxP91VgZdY7ww/8
Hex5RNmAvSNxg+unw3fD5/5G5c40LZ0MODf6cjVf7VR0MJxL7DOC2vBSRNXzkp04V5Jin5KTyWJL
r2l67nnuE7ov9cqLfSVKNKE0wPuFxRppxvY3+dhB6qF/ssT2uzk9MARBGVJQk6c4zf+tLK20oNuC
NIx05Ie9KTRSDJyA8PQNyyEaDBzOkO9Jek0HaaXD0sC26Ol7Aq3NaRufPV+MM0a1IOpXU6vJmzju
kraLjzlQsJ+T2SoXjHowhf0aFNQNVmd3ILTkmC1EkmDHAO6BxgMqUATuINtTviBn4YhnN/Nro+zv
OpX1WZBoxf/zkA+g2qW1WSPB6eggTBiFdrJL+eRFPE3B0kwnCO/LJP437m6VuGrVjGaTMHvFYyHz
C3/mQQEyUCbtSJXGzYg0Xff0jddiWEcU3y1HRJ5P0S46yPToU6ha0qfYrpApxP8o15Re+NbOT/on
A9Tq9q/OJMzX/j1xJhRBqIXI3QNR8M/dzqaGiJZbqUR74iBKtCN5/1jMg9GRSMGDOOhTguwcDO+L
qTBoJvkoiR/qjcCDOHz2Ex5jh3If8eOSIFzFZf3z6P8XzNR9mviVEeuKfFgVZwc2bjwLi+r9Phrt
SClOnJx22VNWHA3HbjhJXLY+yLXgDA8zYS6zKgr+99xXoIk/xrbrsPQvi1vNpQiOCCnCAwxrOLHi
Lzo90+BuJmvlJXDM1k9rudfX8Yp0+rqoBcbTEQ8NrvAUJxnPyEUp8fUHZ0qI2+s5Gre3nzHDHL/S
nU8++cOI7cZSgp4WItarN/5C9W5f4b5LdojB9JYu2aXEv3a8T4lQ/ZoFRgdDEbyRFl976bTCWbCg
dBspVdPfVi3TPdXxYJLugVbU327eoEQ1fTxDSwlQMuGIc5oy+3LiHCxXT1C7tDqdULxQAQ8dW8cf
HOIvN4m+jwxrH0Iq9su5X57kqV842SOTM7lQwWps+Y0mw6EB0Dhe8r8VwIuLP7naOtWO7vuECEk+
+mVjq5w+DG2vVOjuRS03KB7osjVzCA7W4E38a4W3t2Kp9GgEpAvJbFDcPjS4g1V51yv3AHLtuCcR
2KvIRSRacPo6KYI7T+MkvPyrIYz6fAo/ivfxjMQm7m29d8Au47h3sRM8pGm7UtbJFo1cZ422jZ1f
ZN4NsCs336H76bauztMSZ4zfESj1+KWChfB+e5cW9XTvobE4Iu0HnCGiHoCENLq+DqFqYegWNX7H
8qdh3dokXR2y4TI20ml5av44brA9YbXowSSEd/dXylEaJ/7VyqmZi8+vkD1v5TadYAcxp4S/nB+R
jrQUxFLD6qDH9XkYJ4INjrFuW8EZJEu22HLcsC10xQHUM7/GRrkVWf3RxJl0Z4x/0gWFjbf/6+Ha
m//ruTb8KTcknFNlgj81vIitgV3eH2X7M++KilJmxCfG0loRL9ZrFKqJmp7zVoTGuGmaG183bsn5
a/41GJT4oa2XXByAwxXmK8OW/5CUzmFGP70xOV9bnyuOS4pozOOxxYSQz1H4Dbnn9SHNwQObIhFY
pRxCiXy3OYr0in3x859ZQdkROluH2T2ieOKZcCsoZT+AGu9drSFtlI5g6RWO4Ygm9f+5KayvSE2a
Mo/iQhhOkjg4Ape/6+qP4i9OhNvMZzZ5HAvmp7enpVillBhLBYUae5qBrhJXmLTMSSKYxRkY12r1
xGulgunEIq3B5FpKnrIeVihAmkUZJoq3JAIbLZsuzonEwZc/KICMMOYhOZA58RYJGfNYCDNS1msh
+NN3/G88gTvdgDIY+0OSvk/VOYaQLtpcTvirsjnPOzDw2PT7VIW7jqzhf6k16yYk4/oDo/EBrxEU
Euj6yCw5rJjiwxsv7MGIuEo/42lbvVhrgJg3kmtoCoCtz9midR+hp2zPKtyamGhq8dc9+lK1KFQ2
STrahi936WIAymvgMok1YwBVJT2iyVfWUYiCjJt5T7Q74UgXT9QXG792yjNjQjlqfLlX/T4EvZZO
A1RR23+YXOqmh7NkQJqcT7u+DlqWNxrnU8Rr/TFa8UvPb7cJ5UdWXcBd86RA34fCE0D4TV8sWMY1
qAvUBHfJCcMuM38jDqLn4K00O3y+6UNG16P8JBKMlnqOnnHCloZHu0Ts+fuTOQjddF3CjHafftdv
GwzxekzBpTIJZ6fESNnndSwMEkjlFR5taxU2zve4NB9sb5inhC/1QvLQ0iaNX+Pv94BoJ3xSeevd
QWTQHmixWN4P1Zb2yqP4DoYO1MD6RILlZPBeN97TfIOBnhkBeiXmmoq8A1ao86B2Gs99ePtOCYVg
DoapgElmhl97HA6Tk6SqImlYx+8L9nfSDWupkiX27y8/3t6qhfmOy+j57PxoyNOjZzgZtDHWiNJW
gSPI35254YGxDb034h9rc0WMMQc72kP+lhx8mn1yGJWld3QUw3ZSrbV0Kh/mNrhidXmIfchUjVQL
+tDBBkFjuDJtCzChN+h3eXfNwAAA67BLTRhF61tAgZUil9wn8vLbjNv0E/+/7Rc+lpRz/gX9zaxY
/AOz1OhYHxKefLnvLiwRNazX0Hs47AgSMRLsl02Bxs34cnKeVqhOBpDwIl484fUWQpDNaBWCVM6W
M38MX8R8XudBa35RGjdaXAC+S8TzSc148yaPT/RK0sZztMcC4EwDeAm+4DTvl22+xPct633RzSXs
R7PMzQNlF6WqqmazHU0AQflVwwLUrp8U6NTyItiO95ciGi30pzp+6SDYMHf3oOPFgkRq38CBjFJ/
/wWmYeINEXbN2308/aDhzP+fUUA/IEWnfbqP9yTXdcyCmwZv5thggQoc1fCOd907NmR1AtCwginh
D0xelb2Nq7qsN9e/6MwC2BKaCdVybNykhSnSaCBhpob0hb86pChhiIudo+FlRym9glp195Yfh+82
yD9ND1ebcX+KYPDxPcXp2E6sciBpuc9f7Hmd79Rq+peHBAODWZRSSO4JIy5LvZmuVkG8l3z1s/AV
cpRQShSPIbSmd/bRS5wVQCwGZlaOXg9qa0A8kBofkzPlZN8MAg9GThzfHXng3mQqqLDzoMR7KrTi
kk9rsHEDst86rstQshBFEnlwUFpwCgnpcWBFzsimK0h6BDiHsDvYr+QbLGlxpCDtp3+flU8uLhKn
5QztMkXhVnHAxE7gUoTyimiHDifTXoixUuCG6gY2ozLcBUvMPCOpmKgLnUfG9gZWfYUCgKyGjEiT
rN8EtVC6qkFHRBhfJDP/yZSYHr0Vi2DNqhlbjB/kQ369x0x+hiPBCfOc/SFQ9+Yj0TDdOd3rVsnq
gX69hGps/JiiFyKDrhGIQt4nL4xuBSxs/q7wFqXHFzn64xYJydGVZk0QNzE2/zgVOrVWgg673pXw
V5FKScGsg1z6iKDYv2KYqpMI0iAnxj0+4b4+HaWEMzo3O6WqOBrS9uqC2tnU1tqu7MFdDlGEIPs+
fYGOYSwy2whYdHlsvAM1fFmcgbuYCNU0bvHA1z3M1UyoUolaeBZ4Qv1wAshmagnSMN7jpF/nfznm
e64E1LqaeK5zIXTEw9L7hYVkxXX1hG/c4HORSmS4jAgCJHsaM6ac8QTkz6+24juEHsj8rb4nAKRe
//U1+xOWk5lkGbYr0yHyyRnY5kDJkXvDScLmpT8PNgPfq/Th1YJrlFQkf6qxnmj7rzlmlyWbCjGF
q66UGHlOrThjG87NBY0E20U+dB8T0PFg7XSbBD9Oc2dfzyMK4R5kNvGdlwxdenZ+uJ8xYrloHTeV
KBjP/H+mENrGviNP49OGwqw9veBOW2Pjr48l7qhzzrC/9rW4Hiq+YzH1tr85Q8XUL21J/AiqtzYL
9SrU9WIX1m8GFKRJIp2zH7a/egMlwpksNGFr21ByF6RU//GfMgMDVVjNSBm1OmHSmmKNKUDc+bN7
RM2ZU5l92dd+yzx/c625mgdB0U7nsYMs1VxCYaIRCFqF/v6XjLsH/I88R++9nZhPy7yLEa18+2Hi
wc+ZAX0bPWjab2OzG8wWzTj5WNENBPeH1UQ6EkCI442+sgJArM3nSMmt1KXqBZX5xUsFWOeYKnQU
NyLAMI/mmg1mLdX+5rZu5kO+2Ak21bHkQugG9CHX7l7DpEZcdYWgLoR6A4LdBVEpWRy8OpLKaKHW
nVn/r29khFipeyT6uoW/fNcxP3TwZwD/AhNC0O4aVv7LOeE+j4ysxIwHALhulyARiEEmjkLHof1x
XTdsOzbvH7lIuu2nyHjcrM3NXJdNmaPVYLES8KZ9DphedFRCz+vcH5vcmB5kc12DklJPk/l3VVGT
4tBb0ltFyeq0NYV+FLZy8f+24pmoYPuOoW6LWShoYtjQXN7jhJn0MnKs5MpctrCTs9Dn5l/Xt+uD
DBvaHamZx/LShtzyUeoxDhI/536i4V0Ijs2HCBxg7lvY0qPl9cMOH5CRFQIWT43dHKonjTAdBhVG
1Hsd3aSxlrim5KfLAKcar4OQzF7rPlR7XNqt1qaQ2lJ1j4RGN6EpGX4WuUdVPwIYuxjKeLgd+eUR
S/aVJiBJ5B87GbcmzlanXgtcL8m3Y6OHD3kiXyXSGywnDKcRk0gWXBxgVr67WWh1MM6doIBanHeR
xwxvXkjorGrQyFVuKYwBWSC5MPYQunWm8hZK26ttThQhFNsyly3YFXMBuYclqEJAUbB1aVunE7aC
7mg2mkCkVi95Te6IIV/+aPhFdJor2WildTDE/D1XB1zP8iF/9attkGn+ztf39zA9KqxS7LquQv81
kq4gLC45dGFz773/9YZRl2rCqUCqjc7r4Rja/PsplceUZh//3w+JVsQI2kylv3ruSs3ZlUZn7NUH
73SASlEjAMeapC83bEb4PdEhETG1O3Uz6QCM5BXYQJ2VR+2T2c5uK4QshMlrEQH0kQn57EYGTbpP
yf35UkUx1S9ig/EY7uieJhEMMJymG+rAbkuXCHlN472Kc/xtDLwcV9ffUH90MlJtbskrkQE5RaqX
U0MWGaTvxOrVnFSDqXRqTsnq7pMWUEStbEGOLQkYqO8BGiws7MXGJn3aZsR6yYk4eSnWPNgEFm3+
CGvqz50RgIaQzdo6MLmZO8/uh/DWwwpFf12G1nJOFAFbKS/2szd6tB6kSQAAXS9eFQFK/zWUdHbo
HmMYUwLS9XWUpaZnFs3k3L6JUdzLOvr/mXJyfqN2X/B5nJRYlHHSg6qUsczekn+ZUsrU0DoAebBe
viYRXu1hnwpD7lmeFP9osUm4U17pN7X6RvlmmJIeSCrFqlevQ+6TO1ZeZ76shm0Jqz26p417q6sK
moogqkt4GK26xaAEA3Hn+csDSf/lQ6PUGi+fhcyqA5+PjZ2Ca6QijeN5WItPMEHLhS3nRVLxhLQo
EvbBUBs4lr1XTR3DLdcEIAlvh5Byg7p+ckEiO+pBuNpFzl/vBf8RFUkSJ7XWw1uEauu5uTJ7FdJc
wVWcBbB9esOvURBZn2LLjLBnKN1FmlpvjnRBfuPhu2G2myS4J2WXHw95tfqzc5JBwqTQF/98/7kh
AM5ufCHEvPdvjXFQf+P+pItDEtL4a5Lj5YXrb0oV7YRISnkvxVYd8PBzkSWwLvgPZ6dggcjlyD7m
uT2/+hBSVPc8iDpsz4jG64jO2AwcnHRYTYVyrXe6EM5anZhI5+wc0JboY+6+KSidyvYOxjkJlexc
6G4Ft8QXDdvVNeCOivfj8GWFgjaJh70Eb4y2rrwGZ2ct1LwulAhmkJ1btKwi3ObwjsWiUSxLtqvW
Caz0l/NmAug13wpRQ5tiIWEbpYhCicNNGNMknQ9fTSuVuKz5wBa1JmbsrE/80Ch2S8zQ+CFyZK8+
Z1OB7NIiVXeGAgmcRXPb1mspyv59dpdojj/dUktcQ1jwEYv/T0AKQ3l4bM1iFVTXN0lOZVl4vkDd
gC2Aeg5/S9/t0lEC0Rj9xX1GBvZM531jS1ev7FMEkLMPNOyYPmSzCpia7LG29Ms5WOMhA2yPXkQt
/0edT4G7MC+EAfAr3gtb15FjxYLj5Oi77BJeUrmf2JT/6rfQTq4zB0URLZWnWfV6VtyE8WE2MZej
fxi/868gxoH8xSMwopyuuiqKchGBOG2pWcDcz3TyTulvNX5lWuuAd91H5/vSsdOMHwK7YOsS04Uy
MIj+oNp9A4ENkCI0sY2dqou23gkFlGBINIOFFbkKBhh2OCNOWn/oXjn1xDiMKn48IzP3PYbSeAmb
Q1fUYVzQXlJFivDSbvucTVpHUfk4Q4h3pbKFs37MHJe0UZyFf+f9wHKUCgeg72v5gzgZ+TUsKlNd
Q3YBLMZt0Pse4fPrycZc7T0F+MUkKROAoGnlS1SGwdMH7sBo1FAp54aMiZtjkOBHvbJ3FHhjqSjR
XAEgmrwdJYpFGufyFehHfW1UZKgE5O+JhLSWG6vFNee2bPfpU/0cZ0+2Mw/oF1BmtSzHHZB1cl+G
QpbJY+dJxqSAEZZEgRyXD4VLj8upmuf8o2pamWtwAHPbInxqZFndqLzrlvpURXEGKXANEABCMWwJ
xSPjZHbmV6p9rCBvaanXEj/7RA963JdmEzm7z0iA0cGlynrYoIPf11Q/b4FA/B9GogHQp0IoDh03
zuotrvMbIxffL5GiBjt6oeupVOJ0dFaYO/knAwasbgV4BuGhuJRVKHnVSjKxOz5wZrD8cQspavJn
F5X168963/vDO9NPDIpRcanayKzDnPk7Ps0DiEd9dh+oA1SXZk0yfg31qeiwGySqID3M+r7uK6W5
QJJoPpcBJPXDrrfELPGHS3WIvihf4EcehiI1UgDWM6gJR9IX6FMgEe3lCF/tsMlRX7LPlVJcNRvp
ZeeOY6DPBlxJtAm3b1ouKDVVTzjtfL95qP50j7coFTqRWF9oQVi2qe6Eb9Bs2lw8bVlEXi8ehbTc
K2suqwcJ27EQsm3JXwmXiJWRzcNBU4Zwxpq3aCMVcJx8CfuII2B6YM8gcFlCf77lwWysQxSTBnjP
RWIOjPbhXXLV9qG4prD5M2hM02ffHcgOd+8HVGWE0E/k8FSqrCLMl6WTllOo0KTcJDkpIZyLhOGA
QylbralSrSkrdI0CSvya0G7rvlyEffvbaK5DSc2PVyLpXaO7AzNOLjWuTSQrk23I9xUik6yJR62f
l4KrOqds7UF7ofeQq2AQ6EE5+Vx64X3IblzhiKdUPDudevpuWjo/0otk6pNKlahmkPPpIne9W6nb
lG3pFVvszTWK0Spsj/2junYW2Bckb3RT1rmJp5COwsA1ugvYojkxzEYmHlCOF2a0A0nCQNxbF+Em
dhJeKkRIfKeNq3/JgySXldNnVSFsq6eLD+nvteI2DozZOELJDMUHiH3kUUfazwm+5cUd/PRho+sV
dYRTQqcV097F0Bu1yDRAo0N1Ws12i0FHIhgHEwvdxTxFozEh4mrMKgF8cO9KiQzzB2SqizF+XTUq
BtfLe+kg5FslnYWKQuG3tF6/J7HVQW0PzU56WnN4tUHkzeMMERGqEORzRElu21ZH3ZKqhGjfLx7b
8Ov/Rrz5vUzTWZwsf8zu6QCIbbY1mG/g4KUPued6D3508wEf+Ozb6rZWIcVRQlBjNBYMIVcpaQS4
BwfAKB+FNUswojB7pt/M6hkjuTiVn9eR6EWLi3bCHqrl80RgqQza9WeUYQFypEBRcGU8etqYLtvh
/PQbwndu7xUCYOoROkRY6qDium9rRJ2vdv0Vrar3jMo+csvmg6zNDmJCX84vt1TnDKFJem2s7oyE
/15Oer8wuXZTDrcpmdkUyfvn4fjci9afYmptPhqFtdatumAvuK/YIryy+uUfaRCEr2ivgK2+I9JP
jkLTXaH3F/f92jhrW4SpyQPKlmb5S9gMhLcGrSC6e6j0OJfeqokrXmun7QZ53ZMwxwIgC5m9dJqb
dUovO2K/YIXk5/mmT3z0LitYYb6DT28ciofvip6wl7IwzHZnjnQOjU3CYH6vlAynv013OpP9gPkY
zaCUWL4pmg9h0qVBnD8i9xywi5ifdFN1mTlExXLt7hY7Reirc4unJbAy09Rqi64TYMdjW9AQsCkP
nQfOFe1xlSSKz+HxUdMVLPKvn/x+wiRsLa8shmCuGLlx5WbM6pbnQpD/AcSh8sLbhTmEtaKjbxkt
61hjBbTFGfSZe5XhewXS8ReTp4CjGMCcx4X74/9MCMRhQ63XoFQBgLqFx4yO5YBS8DGaAxFPFYvU
qVhpaFPYQozU3as2bv7QV9m04Kz5+4DKVPSBOAeNM7crxIiI5gv4K0moUvwhXp3hxLwwKU4c24Q7
MbU4eWsPqXDVUqgI65EkgYDJSOJPLjPdMhYL5d5JGaJvh4f4Vj9Vx5jcrSFJeAHNAqE+PIUi60cy
V3OOBcMnCtVHAFYNJg0el4PuUyVWqDTjjhCPam37CGyIyPy9WCNxnADGe1Dag35HHHeKiAJfIWBm
bUh/OMoD4EVgiVGVbq3wVbYI/IzdC4O+6rzJJcV6pjcGNPH1tsudk/MmOTMipXLQGHRIA/xc/ZRy
qpc1JjlSJ+gXRn0VO0IidbRW0acEXNoy1i8Ox54CYxmYQZgq1gFgrPJDOWgrvhZ/2dFQeP7BbsnV
nwUoEu9l9xWOcqcUplAMehM0v+gvE5TXaojPGYokEG/MI5emnfvqzhtjq9tuPtvU4Kv1Ez19ZdyK
sqUtipQUDuGLrSyFM1nO/RLL4rRmvQ7Ih5bCibVi3YvXPE51ovZAeaCmOzuEQa640qIlRMcfJkQt
runYv9mQO8kJqLP78aGzFkQ3rkM9ZPOSN2hiDJWEtlqyDRDfdaBrN19xQ+bh0BSMUExCRmLDfEFk
pzhsW/8fExjP3WdyV7EfNeEcSxYy6URwEmSmYj3pumWhgXCloqt/cNkLEQxEaBqiMyhUyJhjqQjN
ocbVeIwAMKTk1xeSR9fNKp/hjLW6wXgIo7BPc6NkM4ZN+6ctndMX80tYY6EW1fC8YnQAsLiRZZ43
TwHUmPGRiF/yzmkd/ptsBuNk/7ekO6qGwOtovQ74pabLKKGktyj1c6sYQ4t7Ygse0ySieMZsfS34
FxbG5pJtN4ltydcTwkq9NE4x63rsNeb8325ZKFnlRd0uawykFiQaZWCZh4enmQh6zhKoPqJGepEY
1DmBvXOHAXZwZMC3xy3iJTerPkrzTh3waXqTp2z3o+LJqsc4F9Dym56hPfbnx/udJ0YG5b2SfQr6
KXVa/hrOFcQguajMK4W+5ib6e4At8lnWO713QrciHL9smyoHUJwpSOFzleIOFLzxcxWf+G6UQxOB
RRL/t3EBbXeCvaMOuqHiyddkBzsdSKF97SjuBE1B7N55w9uQNzVa9kulvvo+eb/EY29ieDbq4/dz
hpZ4FpU87ipHi4w/B9DVZuY6RjM8f+KE4b/5g+yYhIBMDkDf6Qrpp9awQWgpsXmn6FnZSNsbd7Bp
xfQbRlAQ+vedMaWbQK2r0HvzQjwkfBqUHYhBA6mvWaS30WYhhpxIKh90lmoXTrfkFD8BUV6Hy2XP
9c9KiLwglsKe7uSF1udu1JoznOsmkoKCn2iebwG81Hr5NThdzcgVG9ofrpG7WvDyNfdR1b/p0JQ9
mtIboG8PmZrl4TiSgy591DNAziq6/lfkr+9imc+K3Yldj73YELGIbVXldqxYXpm0bzyOLWeQKyaT
U4pECV4HGzCeZkLp4lWqXLI/ncjsshx9k8VnNar09tyhsrkuUoafbrPPXWG/PjOWOWHe4yb5zLaz
yfs7F66uCK++20egAVF9QScSTcW2tr73dyGbtFn5/dja6rqxJZUyaSVmZKfqY5wWEx/0Metd61AM
EKr/CHz+YZeVWOlnvFCQjaNjp48eshpBUprWHaAmvCcwhkUl1UQB54C6b++35qljWmbBwo8hJ13G
2dB0Yt6E1w6UocUz4BhvomECV9knKFIlJDDGpSOw68r3buP8aemNNgQXmVdwb0o0JvUqsUnlxu82
WInTU2OzZuxBcv+zArMiiGWnJ0d8N0NPwjU1QbAO+/Dzu/wpP4CEiRDHu/Ub+ecPCzUaTEyIUP8p
C6i64Yxl2H/3iTGaODBol3tKwXOhNVPPNGoQPglRiZ1Eg/hvZYiAmBU+ycM2qYCZDdKFPFpMZqTz
YSWg2k5yvITangc7tRkb4Vrm9mcKirJM2QRBtv/cKiJYsaqrZPPkO6kusuVXf5DZu+HZNlBW9/dZ
Q9DLhxRbUW9TE9/VhjbruLqhy0HNfkEE3jCnIR4zTuc/hSvcq50b2Uv9dSd77JqYNmC9jdBitv2V
DTO182xHFoSn6iK975cGeG0QAVrP5UzRgxJ3PtmBIGVWiEqcHvv7HMiQIfg2SRKAvlLEzBdViZC6
1nQo1vMF6rZGb1qefqvhNxQ9cgZXg6L64CQ0IczX1fwWzVR3lDAahxpP4sxEoLZLB2JPeIcP+Vbg
D5ekmrf5HunJ3dmAXzFrr/OSYUz6VHKEqa/MMgr8gTwc6KHGmVxHlaf4Mtu+/94gzHyp113m6qGj
nnFmsvr6Y/7EzDitZYYdxbbqlPV4noCfFIRS04vbIoSAJhZLb5mlhvilqQxSSm6wPbUU10xKrIVH
mPgBXasxOfCQMV1hm3fIxWk0M2fuBg4QRdAIpYfd2ck4Qny8rsEgiH5p4wQu1zhLJ786bCUxje+2
L4Es0WMk5FHcyFzwKue1Xutv+VSHa/4qy5V5tNIFkI+6KnvRqu46J40yZ/p/Sn4OxEh7qbg18fBC
ycbbk7IQ6YZbJ0l5O85ZB7vIVyGtsNENMVE6COpWPZbYK2BCMYpNq7jVQYOlwAbOZHtEHlQiVet5
Ap7mLpqtLgzqDHcSzJ50+siDNGO1fUStYWSR2x7DCXgW4BOKw29kzn0FDjdLM73AqlO3nspVd5xx
lk1l+Y63oI7rvFPcFPLzcPhUfb0IZjyaTknJLapyZBJLcaRSyo1LXGt0pBlP2Vj+T4rVXQWnn2+t
dL0ZWeCJnNWkozLs+Nr+1GxLJfrKJqlLvDVCV0/oSGB9aN7jljFSn5o+j4lU0Ym+0sO1YwISWCPH
YoSLTE3fzn7yGPyOQDicpvOVVBc9RASHXfUZ0d3xgQ3UuAf9lKadbibsiJ5YASGX5a974jAd5LWC
ghHRVQ6JLdmMhAmzHxXnmY6qLoWwZPfAdDICwr8Gtm6tCbuS0+YhvooCshwvZx5VBWexOI84ULJr
qGA7MVTHgvQVHGM77jwroljpwcjDoH3voyGTV/ozQ9CihpgxpIz3mTEmLporXUF0pNEke4R6pMsg
N12ch/cKu/9lxRIOkhVD0bNJtpzne0BSh4W3XhRO/5V7MUZ75s/Kkf/ZcBJnOIoCuJco4+WbuRpb
aPgo9hs/RnvCfcDya1BhIOwYfskvM+uHjVHq5NVsmuXp+KUFQ/ELoiliXVGLuLRxsR02xm4BQD3+
enedOAh1hWM581MJhzsVLEjD++URsHxHPIGjFci/ybmN8jHn8FFf4X1qrg8CHMcHku33k2vuDPRx
tXt5UXXCFMpmTw==
`protect end_protected
