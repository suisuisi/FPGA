`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AEKVEpuJ/c1+hRr53PizYwDoBvUy58TPDx++lq7a62K2FevIv5kMJIDZBatRLoqy9PCWzft7UfT1
1fTtvJDDfA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qAJxqfXhhM7M/8Y/a9dLg0bEcc1hCZzJ/f7iwWh6GX7ejtBeW/TVJe2lCoJ6nK0Uw4IPDtskMILl
k9jf8mC8SHSy5C6RXscD6b1NTvJ+ayNXanuVuvwVTzvkbwf9vFrICQ7V02Jk65fSD4AsMCfXd8qB
H7yCN+E+PgNRt8bdc50=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uqgf6uS5F2yMyJ7vS282rogvBKT5aAWL6rjc7Lp7rNeGHieRJy8Om+lc8TpVQtwh4VQ+uCTE1hg3
C8p89jaY+awmHViwBjUcMWIhWtYlCVSSYuVvUQs9MxgS1CmMSRa+2oR8CyNVaIOl0nmnlQAxAqfq
UWbsxJJThLpjKmvsug9pfX/zxaGRWcAYennBedlgUetAfiYjueZlEDtbNgx7rLciLiLU4dBAqzBq
ohaZjukX6teqYZ35vEXuQmK9KxeZ+cfxTuBqZWmYUtFy5AWjlw8y8S+oEWxJvvw7W3AJMtEwn+xp
OJNoWKmyiJ93VJDXw7K9ZW7jAVrl2Oe//4tm+w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hSGDkzMxoTAR80Xd+7Y+YAYXOIJDEyrLQjWXXQHSi6wdjrdxwj0s9nHzr4dzFo5lsSnvPipPqrq0
lc3RCPrk8A9VHhnU14lyNnSGrvhWf4EzFsWxqqjYxUBQ8GG5mhwyyF58+J5Q9HKXi2/XLzxwimqW
scUhjg4Wgmqer516sn/xWJHN8IyEgMTOcMGAcYljPh7cBXB5+Ts3ZvQaR2AGwitwm4HE0cQw1ELX
xo6zfFmD6HyBdb0AyGDrnCWHECWoGHTdNhnMozqOijGpQMZllpqNpq5CMl0uiHCDhRA36yoIkKiu
GN4dElvu553VWHEJN2oU2H8FqUg4UrBZEbXtcw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ih0F2aw8WNHRaBla5DZJIZrq4f8X+PePq/9TRrpHpQemeXd1MRlq8oiv2rmuTCuShVqEb/PtCdLn
RdLguGwwq4RVoLHETPLXdeKvthF/uboAF/yr9iIhnd/R0OkZ99ohOQhz1vKE9XhA1JfXzfU6pFF5
yKSSJ7dgNyTAnfZt1Z/Oqi9rMQs5XH/BnBjYaA1YB76q3DEZQwwR2RcNuuNOrbcrYyuBCJzD3vf/
9zvtSj3tDmpK58Kp8guVqfjsSJs/+sKrnO/ffETgMZi0CF/VEzhCP71f7hbA126QJ2WwD0ld09Bn
FWvbmV+pRNujnD7gyO+mHROkK9Y1b4Hw9K93vA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XAzZYq11tJZ0y8d1f99qokqtJm67MTEZ34t8cXcIHyZCjHNveB9CJj6bUwLBMIF0gIosSHNJVxhq
G1Fb2Mge8YEChnstYLQz3Ytih1UDb+9/YW1b0jcVh3oOWhTfDf1YtSWdnssj8kcdTVNVgVQRfeix
2P1NLM8j8PxAa/3T/UE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Uxgy3Jw6viJrQLUPubHImcyEnCcjMj6KctHy2rgYQyXaf40ZfCAf6F2juUdiJpGCNjJBWfOwKe7r
g/S+X8TMSSku6lxjHMOFP4PVGREdQHuzXDmxpgxxo66X8OPgUzqmVGBKFmB9THAPOw8h6WHZWQf3
Asa7Elo2gYrhcTXINAEMJ9z/JFOkfcBusiKbHhrLBa2MaUqp/plpXo8OePsHKhaHDp+lyKTjuji6
s3GUqF3LR/MmBC7sfhkLK5JyMAb237nnwOWDDvMT7LZ6EykWiqwGifLcxXRdPNgAC4Iinkz9pOxy
bTr4Iej2RTk5GyeQb6AJx1kqMnMsI0aFQ7JQ+Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
wQn58XydDnY9/upPaFq2OGr1AvkeQ5m0z8QRCEspJ/uLg8mY9EaQRg51AVeWZJOJwIWNH9hrGWVm
mz5kBO9rYjzFjCIsrro+wJAZvlPDdlnfivZjn57fd65Wrg4ufAyCg4l3bXA0MjQ6z3TtYFG2EpDO
Oh7E66bCEZCRwgleWw4sYqeQR8TVsmRCCQ5VVlASd/UPUVM+YvRiaGWc7cTAusuVvZeEhTRpkUVP
J5j3L+7mwCVsw8nZmQpp8jkdC84OtT/ja7mm3L0rZmlSOTNEdIK6L5EeXlwwwZVORQlSwMAf+xh/
CfZFFLDRpN8F7Ylb9MhtPF6bLrs6anfxuHjOrfJsSDEgOBbfNHGBAJ2tYLzpIyBVnsJSdxH5LaM+
qK8BJzKfK3hFOdeoawhloip3k9Ef7jnfGNYX5MOX26niuhvlDZVpUBC9iUhCaXrum2Fs17e8S2vy
TeJko6KwEFJAzkhDK1lxRTfeROyI34hmV5zZQS+h/F0P8FixdVluq/rCJxmSkaCNYKo6UopUoXee
Fm9xV6bGL0NOxjrFLCg6iAR4akncWabnNLMtLdtSa6aBRbo2PJJ09QTMKNMQH5qPUGMwiwLHbQmd
2FMP5JN0ciD8XylHGL3nZuhcSmFKjQ7YIchSHvve4LbgUzoW+DxCu7cfpoAEo2A6H3v1yM+KLfxJ
UUeS9nY6MRICQM6wryaMaTeDzboOW3P53aJ1fpeY5LvtajiCK5DHp5NY5X36Hcvi0bwf4Y1wKdOS
afnwNgHmrsVbYmubQDXXHuHWf/CYjt9n96+bH1JPCuutEKvVuewrrc5sfz7Vtb9FwCV3uZ2TOBym
2bjwvPMItJUsRr/viY++uh0hAc9mTT7K8aMD8EIaG+9WbJ3bm40Rd37ATyeTdLf9UMdUCwJ6fwIT
n5xTRtGg0UqmzTbs/v3yjwcRidhb1f73JvNQ+U4x1zjTyqHB0tvxSvpMmP3EbU25cnR4CwgQv8s0
NGqkpgt06hUStuPefHt5NlyCwgU9hDXUUjB2ITka0f9v7um/j84qYbSaKqkY8YuADdTYKx4xnu3M
XeKSHO5WgqknSrq35Ga86IcsaMkH2MSygrUZs+alNglvzqkNOCrJgCQ9jVrvqYsirpDNTvG/jWok
tsZBumWRaIlGx/zu3rhxhgtlNvsDXPsquYDadc1vgXaFP+bGZIUzg8cB5cwlT2SSHttXaFmeuYIA
XmFXoJ1kakKiJygpJ7K2NtPNYo50oxPQB6TwnokNTEnYzyZxl2Zt7kYqPU/6Dae1laqSOmzf6sux
0ztiefEIJAaUm/r700ryamjWT4qBdPVEqzJpxi72H+FCR/+ouxfwDTiGm7td+xGduS9wyY0xkthV
8jlZkqUJLsjaHOXppISTiUEddUkb4E8H4c5C5J/QsbWN+LcLJhVT4BVuXrh4loUEqRguMCUOSdXD
EGKpZWdNFzHd26O4X26DR877AgUGNXSLTM5f6tYHvOj71Hw/fKUTaxR1JyDyJRUIZkx6WlVUyaop
URZAa0TpFN43bTff65rYp5B3vuxQ9BdJlT6LD5esiNxab0tQRVvHXeiG53e2oUV7VVbFJXHmAZAd
O3Xs3v0S/bEUzKM8BWe1yh4O5KcnL26p6JESZVJFhL4EY/URKk2Dzmnc8bzEGI5gRhWq2unqnqYb
ZeLMgabdH/MSAWT+17GszxBqvnZFcV/ngtZMkvQrHFt/ucBd6bDRvh7Aojg0RcxbEIeWm2D92ASY
D7RbSOhJ7UN4BDT0gIZou1Iu9qA4fVuFGheRcNSELnJRqgTYdPo9EBfaatv9Z3JWHLhRtqP6oAWi
G1TygQYvod6XRiBAPFdOizmAPrSFYxuU6HdSfK4eYN2rPrQ9w8fTB7YGlrZN/V6ARkthV+/ZdOD5
CS522KchDmdKt3Xj8bU09uJpcxCLYTZU1KkcLlGhH+w2s6XAMMI45cBAh6Hk5QM15n6U39t7FBta
CL16SxmKTv/EZCS/Hy0WtxkSZ1sYbqZY5xMXZn9K3ICtP+DRP36z3nDl7CajX2o8K//sBpvsfTUy
Dj25r6LYprWZZ2wOUQFmR23GfTdDclrmPTlXnIUYnKhWI0Mz9K5tPSbY1wwLfuk4kgoxtW5toD1r
RClLGM5XJgpwXL1TIY88EuA/eG+EZeOKGSRMHFxpcqa0kjcDDwnH0/IFcg5J0Ze9iJ82tEJf4SGI
FUjaIZZN0a1FGr62CLgFg03XLro+5rpgVn0YN6S/MW+FW41wvBezm3oaNjQ+uo+g81enz3NnhBKB
Y7wCAZC4pVcAnvGXpfsakFhGhGenXjmyh8F7TtuvLuXCtScv/D1D+m/cCFBLDmCqGUogFbUmONIm
RRpL15QskkZc7zuFFLMUT/X1pylTQ68a2tSPkc+Voqh7Zai/dAs3Bkbg9VsM+FQqx+SOBbWRwVyF
YsRzvBGshdRSYaBT72K9FPgFjpAfkq9RNklmEVwTPRjlm67WrDGVI5b17KGo58/Q9Kp8XYeuaLCC
iRAHANXV4TmW73SU1l78aM1En13y2n9KeG23DPbcJiy0AWljgaO6W4AOBfoUgRf6zJa6iU/BjXwY
rquilCwU4iImp6H8n9lLiF/t4AeDNy/NtULtOQCC4j2SPrhxWqPzvihyhUEniaL4hG4MPdd18Am3
rkgHpAkfRcxixON6hrMcEwIuRXomJxGwd7+mkIlSReCjG6bzQsHjK7J2/MQb85tEF0ZDh3wAKvBG
xDhWDCJyNE1v/bm4Slq861pyMyZAKb/rHB3giXbVayHj1RQevTkEr4sxYKG+JR+GDx6pIuwjBfso
S4P5ccJONKxdc/MQCfytAWlmH568HCb0R93XkpRonA8bXGf+ez6n9+fAtwDAcbS8MTPraP6C7POm
fis9aBZ6bKJsJZ3CysD+EspaCPFtCUTrc78b3jHWCVFZqffbCwZ1YlWn0gQXb6wwQIeVo2EfP6F0
v478Z8xcMB1Rz1jbtvDgBu0AXDaIYBCLnUYJVY0LpJSYSdmGy6lOl2AcKsJsLuiQ+PZ7N9KKoI7a
qb4kbQHDPEUifR0pfd7M1QG3KCSvC7IFCu4MXO+R+C3IgHiRb6jFrtpFrtTCSp7Chdwd4oZW/VCl
UXRBOiKs90vYN9Ts0QHs9THhbDlzcTjwLosugdEgTEdam0DuEVPcPBIabzKxrwlVPs7keU01LGFf
mLD2e7+n0Glnw6SvvA0R0QOkh97qauSZQhKmarvWw3waNCZswA3Xkx6fqV/AZNqh9dTX85A+Ie3v
QajVjll7tOp3pxQaSbI0E2kr+C0qnWBtVTjwoRaQAzqxWZM8PyxXV9oYoBuXZQ4Sf4qK9CkRbjhc
0vxFPlueFTxa21BdUlVHanGil4JZPONHYIoQ/YVfVPf/wtuJba6e7K4fmm3MQq0r39dhvcdOWmCZ
sjRGItNdJ5clXmwzAWSzfV7glo/48cCG4vMb2W0l/q/2b4QEt+Ec5MYibpM/EJziODVQZM/qUKG/
Rqa8a/wvW14QBeAVJRBiLDb5ydSxsaIhachFSEIK9iPt1YJkqT9YBKVk568onthKnv1CZgoTUXho
gbZWkbsi5bkw5J6MpnRcp2G1WfMNtSz9u97jKuti4WYDZNms3HJ3DwueA8D0G46NJ7OdykRJ4iuf
n99lTAo3CnPDtrDo2AUbiVYtxhfjQ41DvR5QGMPLHTz8oGBwNm0Lzsy5D/w5yJ53uhhZewYPSYWl
lk26/sZpeJqvryePUxtuBspzmVhyZpdV0b/dKWbXbS5dmHM+cXa/xuHX8a5/aq2luQ5ASGdQGYyh
0ckl4SI38QySz9aXDxssjBNgAjzG2O9OaxfT4ytsLzjbKdkDQdXv2NL/un6mOftUkQZCUzNNhPkI
JQ01w38fw10uCg7swyBBaaLh5ruJc36l5CFavOfV8EmO8C0/fDPG47Cleth/7+jN0fOaDVGTY2JS
1LEB5ReyYTii1JDtWztbBnBFzLr76KiKZ3YHcA8sqpoqnz4sGOkOLaBwqqiWlJ+rkvMpMr/e/pFg
RtdYY4er96dOS0IbXvCuHlfa0us0hhh1elqO4nNGvrVGVK94Vbwn7AOXVFpIOpgTe67yQ/eAbbSM
xTVCdVBJEmzIjlifI6dGbDB3HmOoH4KnWbcmg5NNrbMImW7MnGiFDUCjiFe1JI0DzwIIUWuyUqDl
+qFoYGL9aHF8FLDAhv0BQQFrIIEUacxBwQ/DNV1RACtO1gAUrK833ichtbV42EB5tUv3uftsTY+e
AOEWkimopaBb5Cj7PflzjjJDdTIGGH0CaN9KWOtynmeDtU+wkDG2PQxjKkwgNUr9FdKhRdtz0vOV
5uRlIraBcm4IwK3Px6nqSRtBHsaqFFHnQfn++Wvvjg3GBgQr/euwP7pguz5HwOR1h3mE7m3Sx5Ty
QxelHr4fiQ+4AOq4arSGligMgv75pMlUhcE0OPIXc1iqWCBbdsQgcEL86QXxypl4vS/hxIClLLip
8HROdWsU8yIksM+LNip8cQJAoO+SQoDO3M/Znp+HDp238HqfSbEmGf3H0GBKvyHMy5UgOA/AIbNV
aDisUUisnCw/AZOjFbA2NuutbCWQnyUHxGShNzuS8L3OoJnp15tPu3RDfV0QfXvuszBDLHMok4Sn
7H1UbsmZkQnmNTOJZ0lrHzrppGNWyP76/VEWCJcYrkTuJz7SwhpLMl4opOXKaOCtc99119hdjaqn
eQQSegq7EUo/oRia9HFGMHgqx7jXp/BKyuAKqp0hxpEQ0zW9vZiIHqByN9K65xlfnju0NFoOooI4
NFZ+BrrEBcqPWKa2tllel/z4fEGwp/o2QijHXYo+57bbimnO6tH+nrGh8VZwBT+DDQAbXz0Axb2m
XJqgguhWgeTrl1z9QDY3pVujEjp2oMXZaIYENskhR52j7K26CT34Uba68723dAPD5r0899vv1zOZ
arCrNM7CPohuGT0sgULS02Ur3XYiHdeaSJ+2+P5JpQUQWkCv3aAw3Hj8YllLXYyyl/1qs/iT7QWY
dq7gnt/bqQUkqYoKSUrgR98mh2V+tSgSZGgq2SQ9FFwd7AjkXS/HTE/0Y7wFKWQqFqQ0XZq0bREV
oJt4VXU10bNuxacMjbOgF1LrynyY16z1RZ2cNVpI6uD7mvRPqJJYlKGSqg6AWVzsHd6PKTBcv3jH
ZMZ11AyasEhxux3zNCjc+PrOrVkIqWlTy/arv1UzNYMPGeeFhvJyk+dh1I1QVNoyK8rSFopNjfvR
OewRkeM/5GLNKJc7KAkCA7+LPSQ+4VZ6PLcOcMsaS8ix0FbtpgucY0DjJmHCnzYKJVTD8XFneWcw
rSNR1LBLuriMkXFmZExpa3lkxsThNSNc0vVp8sTuT6AO0S9+fYZmdf1NwQKvqBUPOKF7Ayv5I9r/
wM8W5CUkRLzDBpJQrJn88JsrlrU41k5boeghe7WxmU4Xfuq53IJXp/K7KkVXPVODqlEUwNP1v07O
+3ydEGlxiHtvynHidf+PAI23aqEx5DYu0hO/KorN9k0rY2ZfL0b4yRA3UPx8cxRC61xCLIUlFiPw
3E7f8phlRAuaBV3mJz0+ag5zzCIlG+k1pO3VaAZnuZhJgfhRdwXn/yvOB9qS7gqvp2XjLvj7xKYq
JEbyPfMzHimO5tI1RyMKgNXL3ynO1x1KfgvYP20IX38z+1L4Cj20E9FG1moc0pb00dGFCxWg1B3g
3ODc9XOD4qOw8Fs9gwj3n0USUXasnvG36xTP+YxogG7LrWGvGbUzWOz7M6qskHte+7aDDz72/ko/
GtdULlfnaiRGbgoUccrMO0IevDb+vjMJjyklbZfpWCU9l9DcZ1c40nmD2j69QmeCfi7RjOJLNqJL
fj/HC6DEJo36mTNkmpsOoioNBJL/Kly3vVGaPP6O6tF7O+AZOjcX4S654l8X0Eov+8Vq8Kj6DNzj
FXAe8uMUk8yYswHHsOFEKSARfb2z0ibyIlctfwaKyJNXUZXZuKeSALRFSDtIE8b8fI4pQ0CX9Qhj
V7R4s5BZMiPzblRT4Uc4skkTO2LUtxK3KD4RkZrzAfeqVdX57p+OHRdisMYThctBpeSr1DgpVnw5
M48VgiW2Qc5Q1/rOO1CCg0kWVVHjXKeCrwYv4tknyQtx0xNJn1bYm6V6idR5CyW0j+ZGj4NZpFND
YXhvEIDpEYN67zn2vNJyDwOIaOFIlv480LeCUQaAhEJilb7mwMqiBlZCHR6e3JBRQ70qHanslCbu
HIs/6OUukPxMPNLCiuAC07exM5b/UKFpuYLK2WeXTM+J4bCQQA6l8tGiwo7x1v8YWICv1I0SV2R6
bZRrcO0DrILIWTxi2pvhJooymiCSZwdabCyTFOiyYPWgIUukjt+vbvdMEA/s7IVTtZbU7t89JqHP
og5/pp9WCItOSDk9hD4ah1KKW/A8NP5FLoAwVFAn/olXB2Kl+7C1ZEtG0VTxmOS8d/hdZoVzyInn
CxBUZHpdFoqN3cMaLIan7FavDJP/Q9cxhgsrwdfMOmnxsWtAnsS9o/i7OT2mESujAyLNuvHZ1Tia
LdzxTZirM6cPCBjMxyJSndnqKMKlbyIFaHYkfS9XYuWMW6RqlzJ6x57XMpWq2q2AMv+HPA3LmKHG
Bvo+nFF7MinF2Akti8wJg2NwCnIR5JuQoFq5Y6bmOm3SbchSHZrXZSwtL4pOuUgzPdzhE9TDWINJ
oVsnDbTdZcMLI8KUXSLZpaqMO2PsGu7RRWEPO3iEV0stBWajrqUZuLJCpn9/gNUCTrnfC3l0axkW
M/c5T3KOxDuALEWU2Fn2CYEn+E9+/bWd2RvIoPXHqNUOolpnKsaKL6a3jyFgAIQOUE08956BBusy
5cBMhjtuX18V67i6GkCByzfKnKvgAhmVJZ5cmP+27YmjBfxwkCxhiwEXD7Y/1eLUX1M3/mkWBfVh
U5c7zj9MYnq7ocCgL/quhEUyQOht8siVsw+U/Y8/IbV1wHnzKCmeK6KEPtyKmQdDrNl9Ah1ELsus
GYGDhYGnojQWU4Gj9K5KkE98epJAEvQH4deSBPJei2jGTgiXHV4tB4PFoVkO8pu0D4NWkolLsJ2u
8qzqqSQy/A0Owfli9MauaaK5YYzhv6MNS8SeF7CKhMrrZE40CgbKluoC86rcSbyw1KNmkogSbflF
PpQUnRrxoLDPNcv6yoJIKkPxYMUFGnKAG5wSSzC0STOneu+h0xVXvC7raYSnBfZAzkMf3Ao13oY8
8JyvT9GJnbuPd2kvTRIMVpiP8nq3ZElluGwBe7/WSN1C59wNxB6xI6ij1ohZ8B5ExhKVl2y73VQf
biiKyVd6p37IC3W2Ai8sCouUoNsFUblQO8z1x+lTgiLX2CawvtbephdSdrsQrTqDtz3v0BbLuPly
BzmXRfx2nFJ50nE52tU9gj9yCogcRCWRaYZSSxG+lOYFIbp4Wb6nL/gov/R3RCh3YnNJXhOaJyV8
+gVt5T8WljiAOvK23k/D7SGMGL26TP6HDnx+qfh3HJeBTvA3TepzJkbLitph+kUCvoDkxzBmljvQ
XhcxIjmgfwsUENqLcabiOufpXtX1TsN39WwxMlIat+Kh0P7bXy1QCX7cP4hkxOlw6+lIU/oDbudI
ShOtpQc0FeYG7sknLTyHKfO32uUZKMuw3Hs7wD44lmz/Q3gDAdYH53/9GFxeUy9HSBns/SYooTSZ
MhsVZa0EFdq/+deijkKA7C1SmIsrzlQk9OywznTF1pvEYVHOrNSYTs7y6zC/xFRFO1nwpg9Uo6YQ
rWBgBpaSqbqDMndlLvdlOFIC2o1Y7AOr8B+hst+Ch3B4fetBsKPNZ0lwrLMC1zO9jSSREx+9pijh
XPZuBnCGGLa/wlT2Zuo9rUMuG/d565vvZoy794oEZBtzTtUVsCSuyZCZZ0ORS2DuLUVB4mc+8Rdq
LUdNosNZh+jaOfzITBQgX9WDkdZBRYXuw3hdEd6X5+HCMe0h41/SY3KOEQMwIDz2WMqOx/5kivPy
fqA5aS4CU6MzVoQzIcONJkGAkW6Pl1IMGeTj23CN/MSe3DkDeYy6BFi1YfPHGLmIeugo923JwIeg
k0VMyRJLfcv7G2vFYN72KYZX4SzbVH3QuP18gNbFpyj5GXDZEbM6EROMtJ1+zpcxJgr5+J7r9eBH
6yHeCZYGSdNeqEbByE0bWinE6bLAFIwukGHaJqOnNFjTqgg+7YHv8/Wrl1VKr3uQ6hCm8U3E8f8O
3sQf8Ayvw/Y9z8yPzxmnVN6qbyoFGHvFM2a+jBTSlgnW88BFGikicrvovl2EXCgLK44xiCEMTryJ
mxyXGkt5nwfqk3NRUHCEMfyaWRyj4tIyq9AjqKNX4HB0nCUR90y823CzHnLGcxuHGG7Zba5RJSTc
wHewPHQlPRY33AOwyCqy7D3vzj5yNjFdzsJZqYsAwBuMUaWODxUWPLg7/w8gopKlQvNZ9fJ5kJRP
0vPhzUDP35MxjiFyk/H85/R7XvYMX+9s4JgIwbElxiRp3ZO39KwM9hkeq7c5qUqhDyoVDkqajQAP
qLXh9nF02nWB8pZRYXBfgW+pB0m0M7Y81KWuJVOlMsgwUeJIvYgAhYtCIRpflPrQz/MYYtIUO/8S
P06UyA/NrYFmwWnir+XuenmGxwC/3VYabc7dbzhhtzdVgwpS1fGdTDmxbiK/Jn/B6jN6MhRwhn1Y
WqyX/TqVI1Di5FYU3n6vZJdwwzK0kA9De/osnDPdDw/8QNzel+U5YgghJfNdk0iBjuLsBVlHOQO7
R2OuHwSn2+cw5+9kgksom3CTGe3eJLbPwLfnfmuu9tbHA8uTWmNROGtUFLbYc6bpRm7othQwAUXB
WiDUV48mZvM4H5aUCEceySBUiDm9LFsSqC7bp34J6rwHPsnlOOBDw6duhtNPMIWzKJIxw6w7aKu1
/NSGnrCne+t+u60MGKMd/NOTBCpZuIQgioei0gw7F6inbSX8Nku/hPEFKo1fnGVFX4L6dgQMlxYH
mU7Cecf88Lh3Pa5tu9AL0i0vRZOQr8XMTkR60icVZ61/C0DLoG6N1piiIjwPArX74+wfNy3kTlGA
Wx36Fm+9X5TZfnpOW1sTAfjVNUHpUrejfPLQk5TbuTHiH/50XNlWrm0wpghDXONR2b65koOAwnkv
9b+4NrDyJOgxf5enuCsjr/OzRVQYTNjm0xlAxtAJ6ujeFq7xLXU/5iXHhysJ5Eat3xK2s30brs+Z
ZBiSGtqI+aFBBJmz5a/vtD0G4ess9nhdW8T8/MXBZgz5/dD2tYjxwA87f4Dh7rrW3Wbo/GFUp2lQ
V2j+tmZt1yEN7XTuHLQ1eaSFNF0Wb4hHJFPPJwSlsEuH6mP5hj7yvTByQjIeXNjcKmnenAW7L1/x
KL8CbZRQl8HFLOh2CNKyBARrA6NnJNmL/Q7ej7fV1q08KeVjAvCGea7UL3DVox/Lcji1JPPJKyPA
JHGUSEawb2oSBISrrcLFkWyZAH8pB6tkZVSQpE4+jb3UDVxm9WZklTUVRcq4AToJcAByHTuuwDEf
yo2ckQf+6oB7XESRLAyS7YJS3nPumWI4BLXtca1AQTTT/de8U87qV2p2bwfiDHNX1/E2C8jNJnzP
+F3uMiwC6yOl5DhczQC6vxbwVU9Eur8j4dV/EHZ/apedWEot+/aqdVWLyh3X3SsmpnTH+EVb52E4
E3xmM8k+7WH+e7YyBzg7qwcgzTeNwSsddOpfknOrBperbLLXYMtj5pGmrTpplXU0m99HmeVFKao6
wh/rRUBUDJKdw5vi8bORK94V9FY/3qrM11D3o/XszBNYAf34WqLtrGjqodk0h5v2RJ5R6iM4AYJ7
OOeI6PP3ZX8bAYhKjsCHGydYZJlfNnDa3yHjzIrw1ehZ5QlsFGkAmiR8nRfFSG90tqwsaiIcSSRh
vQmzZJmjcBkj6o70ao90QV+0+Zt4uAR19LHnChi8LRbS5WorPtX+L6Olbyl/39gha9Y00n7rm3Ou
wzicoKIrQicHw01T9N6fGevQCTGeIRIleWF1PlhGHiXqEJNPS2RcgMFEBJK2kgOFrX13hkX6XkKu
4f4lP/NmRAT4pxZoazS51pavG0D7ezlLlu9nLRCdg5t+mmzGp8VFd5F/XWqDjmGSw27x4VOvo8ts
WFyFNUvFtR3tVARdhNj/9qlNBcBVZQOFOO6ShQyozVuywao6bKICOw/Hf8//pasKdaKDO3xV6Jaa
xHAUpkjnHvG9RneTZOR4DgHdvn2gcE/EwDiwoCpzQADF2aruBF566LoOjixwimEu9QBb8k4pBJLh
wSv+PEJwlLwAjlwbqlYDg2YtDzl10eY0pOhOv4RPXTBnsVwBf+/dOtiZ/AHmyX0UlUACoADQpwgJ
TKGG5FAqugA/fnSQ9SfUkBfm9tsR43KNnXcnF35I9c0X0CfJ/CRV5Ice9r/fkQkwPAN1CxXy0BbD
3wo6Sy8WqJCFfJIp+kSSbkHRPKPBZrZumcqsQaZVcWoEp924/oMKAb39cjI720ZLKpJhvRn4UDfo
EyCnrhlBQylAfKX1R+Gb6yRAMDtZEF2mBB0kuz4hcvEbeLPwD6ynKjxxG2de+apQDdrvHkX74fJk
ce6w9uCN9A38g9B6lP9CybbbU4Nxy5ZwjxYSM5Oihca7UZ3heLMcXihTNV5rzsNtaBU7QAfIb/2Z
eDWPi7lTsoS4K7uaaXQl1nJmLq/Rkc6Zmrn1AB6CLn62uULY9VxRIiZ4yoPWZDSXH22pniGw3YAR
aaeEfxgXqlRvCHYznAz+Pgl4F20JeO7+5zWhZ5wUe8+Q0m/RB4HZx1+lkLKeJhM1SXjvW4rrPGLX
RPCMGAAPKDIb1vO5afSCG8FjSx9G/xLC5WmfF3KWuiQ9g8Dpis7fWvAnSV6exE6wwK02yNPUm6/x
rNyhmU7n+JbW3ASqZdHcR4MGqDg3mJeauR69DB1N2SzTu16hB0lmZvWbRbzUXKXFhLc3nPIUeDEZ
FhAYUyJbtf+Ncts3ENMFynJLCNXEQrLcxWAtVDDLcSYwxmtIOCnZ1FGy+COkBPnT8kHlc7KvLieH
Dq3Yw4dilapLqSsycpnUFsZa5Ai6Ab57Jp3Bc0uSk4zRK22e5bvPOC9aT11MGoq82opZc3S/d8Bs
Tg3ELw+OBhtqxrEZM7M+71D2ZIUvxn4RamgcpkV2p8z452usQQtJDY50dTkqIg9sfSMkXZe32glc
mJzxf7ZHYgL4HY5k1S1Gvtm872fUGmxHSuo4AK94BLieNuWeYakCyuKJkYaB5ZEqS8Tfx+H5vZFl
HiwL/ioIwpD/ZoA9Y5AHFR9iSwTlxwpV7J/u7Vbtmm9MeKglH8Z3itlFI1BSJW46esmDFBeU+3A9
HXj0JAkscSM+NDojVe4ktX3ifvjVyzWQT4YjkENLL3kdkjGhUmJuFusL4Xj8XBfZIpba3A6M3Uj1
7cIRLkg7ldegUouXPzKbuib+nGsYhO9QIufr7L1PZ/f67LkFcl3IR3ceKahEYuJbCghABjY0ZXgq
/oopoURZt5vNn0c2aAXG9IQuNd2PPjRMNpmUFMfwdDTHDZUOfSnddG95sq5Xg7NEgne4emNeNTO6
kaoJHs6aufEwJoPhppf+mDWjWT7I9THeJxJslIyUeyviwnt3Z8+lAD4TwiuJ5T3SKNyW3/rv290E
SyaH8IEy2rAnPZvqbWAjiO6NRzyrbLwIT1ofMZEHUgcJukE2zbKmEmUPFg8EGGDQQSCbPFEhiaDq
90vXaM7LZsEgvBj2vjYF75gC6MaA+vRzBsBWjyFM9iP6f4iI2MTxWY+KKMEn7FcPUpkWk8/pdLzf
x+RfI2eXU9GMQOc1geNb6ItGQJzdiLzFGfsKEaIBby1t42cy/B+S0srBEa+rLg1DN2kCyfjQ6zrU
5aHiJk8a+3fgBl/r9RkXFpqifginmzom+CoO/7qCzc0K0QChcBknptnStmn23mM3fc5Sh61z1BuU
LLPFNGTAcjX2qtvHE8o26SBaDW/FvR+/BVGrLNvObfEXlOEUEcx++iHWzNh2R0gAma3/mG1MdJgH
armSLLioLn2oguwUWGdi7oK9UBOssANQZcvWChXBllqXXFnRQKE2DGoaz4TF7S2x7qmt3nkN2XBA
yMJL4IbXZa5vps/3YqZAoikD0i6tlwJ0qDyVk6Epnk0HTwIW48iZr2VTZKwaBCqcrSCLEtVJbXHg
QHSeZplzaLXrsinhPSs7l53RaPAuARH135bRNCxM5IYoe2wgvOka2Mq9Hix6blw56ByBNJQp+d1T
mkJfx+bIR3wO5Ml+RugUPwsvw8ig1A0lAEvN9fGX1ZWDMMoaByrfAiVZLxFK0/i+Tp5iCygbZAFz
dYYejAhTtBO3gcLUCLG+y/78PmwX7LanKdAK3nEpBVp8tF5KJJ36Ll7TBLwgxq72wn+7Z+4xdjyC
OVwllIxatG2bnwtSZ5nHmsmQrP2CJr8noEnJ4BIlZYFyVsxV6+3CowN0eICFA4gLKeinnlnFUmXe
l+1/JXyMJIyIjaMfmwjSZRAObgcntXiD0Uc7F0NQyTVfbQNW2r9C0r3mO0Q53OaMPsdmiCY+2KHW
7HKosbkb2HguwePxRXib1TG/hIbhoTsQJ18hy2Bnv0HboactLmpUtaqZKMnIXtf9OD/xQl5TccUo
RG5Pqp2lNe0/i01FfhXsPvduHsQgDaCNEmdgkM5PvspS/3r2xSxWjDDlGKOVDfmBd+WKf/E2L1gc
6ftmRM8CsHji0FPVtWkkXIwTBwhE7WP2WO8b5fPiCyfy7ByJzYTzZVHNH7evt5PkFZWY5SjAG4we
nP1qkFgS8R8ZtHTTsVmZlBt24C2hJq7ChntFEqcH2Dhfyw+V/7UNr8ca5So15VBStmIkvEm8/W9y
A5R+pvFXQCkLG3idh/AFovf9bgwuxAOFVEquK8Pgj/D8iwgcghNQhI4/kPw5VGvLfrq3+/cth4VV
g2yk/Y4LAGhkgFY7ieZh2ylVGQUEVPXPe6K0vyCNlJmpp4gGIc0nM+21unwHfgu68kwzymw/ZxQy
AdCvkfJ8b0QrdKANU67TjL7NNJW4OtZQygsLlUL4DmiS+uaXGxJB43jdORwXSUjX7oZP/Y/+oxWj
95HL0Bj5hgTaanv3kwjFznt1cQJGSu555b08zh+jUF69qj4ZvwS/7PXSj4JOHYr/28XAHijxFAnA
nFZ8RXimLdfincZnKvV0Y4vEBlT6bcb9GP7ijd0JjxsSi9sG/bPGeDgF2fs7Q2I1WmQyU0cS2lDU
ktNC2FDZ+CH9Y42TJJd94/RhZ8D2NzgloLBc2gxfad+mU4hUd4BkC59SCnn1NqfKxPCBGILds9oK
CKy+8jfYHRTAvfywEINBs4A2DvNFCVndIgzpy0KLQmfRu/edtmeanmZUNgSocxJwrt6eRzjJrbC/
T9IHruv2/dqGFN3I2nmQKADTZlWI5ImhDeJnpaOp36ZXQIy6j0LGTbv3mefhPeRNgYlQq0Kk/rmD
VdV507LB9SvNRKWGOkuHkarEFaSFcuO3UzzWu2Wl9BMRqoAavwXlbDNdhMCOnaDOaBUa26qsusPi
Np157Ha0fU/IvAOxQIoMn2bdxlSbpJQolHkOJ7o6a0I3kmhGqUWzc+cnJs5ENVkXdFByRw7vVXWc
eB+QY6ww+hubqP6BpEX3N1y4bYP2f2gqmofGRppVZ3wa21z47lopzNNz1ed0/T8y851rUhiyY+JA
TQH1R9JQ/FxVK6v/y+HIUT3EVPnV47TEHK0tm55o/X4p+0pjal1J19j91PUAHlN+KfyC2a1tZ3A/
WArPCEkX0UbIuuePLnyQD3THXb7Ha8PoKOlvPeKNrPRnmjwH4xsddk2ny+3AMi9SbfjT6G4hRkqO
xfpoxE/CUqr4w+HpbQmFHfm9UIx+0ScdODCwb/jetkjq7WyE6WACBQtWIA0Anjkn2DmEYO4X+JJu
Wh6h7xGUmTV4QjtJ/uixDgvjPkegzLQFNUUGYsUrhsRDNPyvl1TDuhHWB3tPC21F8YbmtM6YwGqn
6tl2cEHhNe05/0EK/wO08oqvPEuNOosAydwuGgwzmQ2tBuHBCX6z70y43fL/9bN0VEynVS6i5W3R
kusT6onIuxdWMLtpc28FEfk1Qqv4N03hOamVHqojdMpFFQuQWbysFPSQ8KHEU3PQGBHruoDyCvEK
SMCKAPQgSGkrJI6nrKcmC4X+pajv+rRbk5WpSIEgjKYn0Zpvu+BL5J6agvz6KxyhEx1bVD3Rpykb
GGOQUhTtIBQ6O1bUNNfJpWWNECh/HsticfPEafuti0LT7e7PqB3lpBywFLKt0i6o+qe6aLFFZ1ah
ceyOfoVwYgIqgaJcknBgAJ1aeRlXJ7Vs5ha7uoHmpu7B4HmkcFLz1UnWgrBKvMM608iTmHXtCXyN
qwvgPSIFZqFLMaP1YzG+M6SR4CK3nJsSzLziIUd+2vcasE+WQNJ+rEixgDoaQPaEWZQC53LKyTb0
hfuW7Awxz/gaZDFHMDlqw8voeW6wcJk0H9grxz4mIc4Ll+zC65FfJoaYKaS55ulV6NvrzBcJ6wAp
zP47Qcl4/gJdUagN3OoodiaEdTMdBkI9qGIIW2fKOeawRNkOyuzFV6Z0zthesKrJj6Mw5BzaP3e4
xJTJ/bJ1ffrDLAT9xruN/3HygVDeSG9fxZZRBc1M352tYmlEwwkB3uXvvlGDg/fczePVOdNh49cz
1LodnXy2VFspPo8VMftBIs5lxaIHwxHijiDPGEOZfko+HxGZuJuhwXyfLDvrqH6KG0NrpEJWLcOD
jKgFxY3KjWVSMjOx33wPE8H+zOWFqQJT4x1nQ+DIRz7rOFXyO02JTl+F26aRliv8ZOXbgNW0/yx8
JB+h0o8aDbAbS1L0HVIvOx5H0xH3lQmFJehasqVf2XmhutbI3dQdjXJa05D2m5AbSohT883VqWiI
XIwxIrLQxsTa0wdsbYJ3yx2Dy0X21U2Bc/r/Fg/37TUaOXulqJVWprbBwNVBXhEhINCuWbJL4BwP
rKjfMI5Wwpzo3grTJaYAxERMc7YjCOgPU+ACFmgxsKoOj4zyQk3kdInmpkVRL5zGhPr8e9LfTE5Z
Hm9BLJu1zSl2NWt1Vqt8RTfKJMb+b5EsM47wm9GcoqgMsh3/QqAKWuOt56u5T084Oin2cWjsjPip
g9mDD733GqveNawSw4Y6Ki4kFSFiMHF/Kd94rVmA27zas4jvBRyHjW0BHqHSbvZWagzUb9xUOaiL
BCphOAQpuGjx2Oh8ZyniF6/g0/SvZCAWeSu78KUDO6usWlg56sYMH9F97F0t1bmLhK//LcjBGZCZ
V5gAT9Vfld6C49ctNRbpQBC6J6lWLk+0iQID1r3LI4oc60/8hJExAZktRiQPLEF1zubKM6feFS2g
gJL+CxzEuobiXIyKaR/WC+BBKUHzq8ubQzwbQB+oJshVq8YsLIPBExg7RuEZ7FOfNCzzj3KHzNPT
nAKycXtQSJuSotHuCtdjsi1ah3c02s9+EkAviko0m7k1cEJCDSU77Zknk2XfyWQgAQztv8fErsNi
z9ptO36varLZkOorC+sOcbMcqf97ZJG3Kt3XuXrL6jiTq7+ckFrtpUTQyDHz+35GUCNJbpAoxGqp
G3uLuL2tAjTrijsW5Unc7rPsOZaBtFSdazaZhf0rOg8HJPf/6dHF+y/ErpgbbsJFAELjSa6kVTPb
DUrJPQrJIUkqZA2SFrCQrtkUS9cYdErjPgZZ5i1jKlqgE+7yB3ddTOfBRPuXECLJsr2/S0Ds/c5S
zJTGk49OTAuzW/q6VAWUWlKVX4UrBo3BUii/NpUrPsg0DtTex60kb6bBRE/cV5D/v0mJDFB6VjKR
aY86jeDbQtsGlGC86Nngs9R2ZyRL60TQ/Z4RbxHcG4EJDtQWX4wGugZmPrQZGoQvuXNZZGbRsBpc
bmSm+dfsCLzPT9+b58qYmSM6D2HZtQ6slbXtCdvkcV0HDPGd8R8UECcgZ3OFPZUml0XqpcCFzA2x
xgfhu6FTlXiXHNHzP6oPnC8iZDqmVfLPLmmk3F7ufaxSQn/eBx7K6x6qdB5hVmP+FaMewdW0UDrc
QpCfbpAbelkpYDCpA/uGdHmCeWmhNv5md0NaYXb7i2sQPW3CsCafJ3uNcxXVVZte4zhfUz9A5Tfm
fz8gLFUbDJ1heOqT/l+oX+1MlU90ksJ+t4WDBC/UF42YVwq0ORJ6aACrGpqpaFessy1/DlQ1ZYMP
rj1BHkoMLouIleTM3F7bqrlOVFW0E+QmDiypz4HdP2uXEhj7MpIYB04N6muOjpweGLLwdNuWRmMU
x73rGDmsYFigE1DpCnmvQKktPSmIRIyxEvnb8MHAGxcKgbUn5Z5Y8TTpkz6rbKXxN5nX643KN3VA
nN+8lvvLLAZj5Xen3kAuzlEnqniz5Iwo5EPeT3kwI8CSsjQrymVwwpIacDcpD7ChqLM135peY9mY
040FN8RLrX4fTZTCE29xdO+5+XNsEtdn+doXcn0waxD5vpnxwkABi+gN9cQfIxGWBJgmxdl3jSNW
Gy7kISfb1oBkeI1J0I+03RQK4GI1Y6PAmr6WH5Jn63FX8sydQWES9oUoOUvE/J44XZzduiNEKuDf
1L07bHkoReNkqC1zV8LvYa3hqiLqxfEW9UX8bG3FSNFIYcx/tFYSXjOX8HriGxNzKM4Q4mxVWrct
dO15JGnyopK778SaN+pbBDKZ0xCHSgSNbQxrycPgACeeA6nn0opx0AOvH49Yd3vFlHF7NGqde6ul
rK6cxo00i5hyU02rLFluJMpiJFfhvxjsZFBJ7BGBrzpfLZSHhHrpswb3x98201K972vGQEmjmKL8
tUJ3o8LbsLVJNYNd3KJd+vxB9U/dRnPSZ0eDxEAE8atOywrFXy60ZBpivOjZAgZd0C+5saKWvuEM
MgxUo8Oe/UEOBGrRzHvN/FV8LIHxA26iq7NRJeysoek+bEoELzTzdXS9b/hVT/ELbkMrWRC0BBxc
qqxLxV8GDSpB7aEnvZB0qiTRvMel+Mnqq2no9vcj43XNwCy1t3o7+ALjSrtmuBz1eCFFxLONmyvS
yJcmILCEB2344hSgxbteY27lxP0ZT1WMUIiGDh85bUTj4zWFxINHm1xAaKsCR33Dmg7/jcUEDAy3
eBy56BulgJT9pY0CusvkqTQmxzdod/XwoS39J1SbSn9BDHIfE8Bx446mkCeC8Y0BnK7mdkHB5ucQ
9MtJnPzTQigKd/o4AsNhWeEu+zPH9wOCQvaVyTrabxNLPfD19VLy4z5A+UTIgagcg3KQ9hAji9Cb
BERIUmv3pLDNn1jtWsgrjKiDlETZzgseZLdfIuhgu8Hx0Oc+clxo40teXxSDfEGBbiR+ExAhwrdy
0Y7sAf5gYZbfKbtVOSps5h22jBvrv5BfUyjv5lyjbtzyJGnGWd+LTjrBcOjV9Om11pc3PTyJvKl3
5amsnMTyWE2JcvR57PdsbXph+S2Nng4PTH2JryHzIqAJfYRDM9hc9MoNWql+SiM5RgnR3TDTFJta
Be6Eg8UVCENXJZs3MDgLsmYZcU6kIZwzT9SmKanUpyatgciGS3t7k8mVK5H/qUIa9IVUx5XrchO1
6VuVOXUmnduFVR93owjNrg+n12giaHpULIRBm9vUVA50ClrLsv0GGf48q9yQPqaMuE4F/HKbSbzx
/1/xjL9SYqm0b0K/xK6YFUydrw5asQ7SXGq4S10U60iEjhQwtPCwT7K2nbFYXfGGkn/t7PqCgbGC
9orMTkm0r5YHiMKed9bEA5/RdBUEr7NUFSrsUMw+1H4ONMRD413LEt8N9tB0p4Jf6Z3qR5kD0zEv
QHQ9sH4PHo7WlQ58ZXcd6gqg3oeDy+VQVJRy/KSMhFFMdCznXLAWOfdGbqgc0iWEQgjskYPdA7ui
6fWPKvw1f4AkOEe5Dje/bgWwwnFO0MPLknLZfV8RcwWHwXoftP0W/9NtRv4yMKFTT+1EBTo5agOL
EEGlMUp1KOTHUvJm4IilucUvwSJgf5ftL+tm7odcO7PN0ZaaMmUQ6GjN1pX9JEbxuJn2wuCfXBYP
N+u2fzL/YWUtu307ZDsjOXo/WbJgppp/g9Q6Ce7aBto+A0GEsLqxuj04xGaFjX/rW1Bb7Dln79e2
3hlWMscny6/vciNRX5NuvLcpQI+21oKiqsN6VLyOmWQ5eupeyKilXSK07uVbcfCf4rj1jxOMZtko
24PC62hdPlz73MEOatUKW6WMMucMVanScg6jhjR7y9EJgvgT4SXjFKmoXhswlcB95lT8zkHOwUDE
fa847OSXUdJQqvDb//tLBL9c6Ocs7NOt6/Lzw+JSGOpYnKyeX0yTC0mhckhEioUzDhO+qcqZdD23
ISQOgAHl+6BvjDmYnG4xFl0sjwBI62joe5u/awDCd48pWxQIbOL5HvincfKfZNKPUn4oZTNh+lsu
RFyGFv8vWxpSuOAzUZ23AUBSIycvWxiYa9cpwyOUK4rPspM+yAbH7Boc+CTIx77q17LEtTNrNrw/
5y7TAR6Y7JkR2mrHdTPm/oeW9mpKj+7DgiYdWeQt/KNv3/X3b2s89BVYIFjvSIrYyV8913T2Puh5
kTr1wyVGfZJvOGdVKXpvGT0A4gn+M52RpTBkxaebk7c41ex1t31CSqKCrRBSQzTe73mhgQXqwS3e
5eA+f7/e3ILjDVuV9uVfPlPAs0lgofOpBRrnyqliBwJ7jjgia1NT2GyQJTjD2F3XO9kw4pQAsBq8
Jhp73P4oPN1GtWKdmphYr+Z5ealG/zODVgq7fRc6kcAXZcEvPYjSnhEf/IQf5EM0+/1k6OGHEEOo
/bswwuRhmY01bNMZihme3yaTTXnMEEk7D8UjMuW1n69aVa2OZaGVcclBGnBIs6Yh83qisCYNwcwE
MmiBLk1yEZJcUJgLuYblOCxJ6UecNqWAb5RAe/KEZ1rj1Cxa2nZoqvntoVSMBbwzw5QIWB3siYgD
DOCjnSbqZEuNCHzmRlqNpn5j3BTcEkGwS+Cickan6cSfSP4KkW/qVk0jPQcW7lPg3FizNIrsp5PP
6xrnnrvhB+tdtU1syO6h1DLfn3FDmDBheteSY7DuecGaLYBjZVtrVnsb/4ReJtjOOurHokO9oNf4
LrcQomGmHHRWSpHIRZRVBKiOsA3ALJR0GE8jTfpE+xNCP8TEEj1hgm7s5769pup+brJPQPCj3qjf
Q4wWLks8mawSeBJ5YcpYmQCWmPScXQDptp+l/Pg9p14pf+NRSZgVeZIx1HY8AwoEArCTWT8M5SxP
zAYEd6TTqXpG1YQgMbVtTtavjoGr5p42kxTIaPnu5udnpeufmxREc1KrJaopcxpc30/l0l3fILvw
zNoonlm0slUOFYtJoA0MHMGZiLuAiINoaLBLA3EeTqy5+CCEX8JJ6y53FYIMaCVPKdzNkmyVAtUm
AMONT/NqiwY1HHOcYx+TqpZ8Bhx/GMEXnkMT2p5h0iZgJKrwVPXN4nk4uOkG6xQEutUXnD3lV3TY
u2mwTstv8WjzbLpvblSjBKxefTdEkxTcGvVm8NF4Fj4j6U1htZai0xIg1MDPZAQkFKLU1U3/Ajgk
eJP1sWeOdfN8QGGIIqJ6Hi9Z6DHxR1ovmnqjva4+2q3KJ3idZmBS4VFdptxBBJIfsNws+umY82Gh
xxzUpA1nPeWPJxTg/OFghRzrcfSoj0uFjoCAcnKpVbvkmpKOCbboTddQMUIR+CRuiKgE0wqUSuCf
M+VqZcSXtu4Enxd2fq4xpi1qFV9BFG9OQF8GKE5Q+ywwFsjunMo9bVu6VISS8ZfET0QDDpYeqJ2j
GTTcy5EzP1qCDyD6IQ4M6nFgMbvZTrVmOOgua/CrTQeeXAmVKmUr4o5UNHXm8K/2alJzsjYGP62S
S1IEInAy53BwJD2FeFxiMjCLuGovo476n+8z764KSWm7W01lrMlPdIpOfp3zrT4iIb8ETp6hxwTf
TPbSbozVhBDg031RQHt6RJ0wOqkMvx+sq129C/5+Y5DxrR5TBAJhdTuStwgQUOHDoWUumwz2HaqY
WseiXJMP7JRLTHvSTeqPcevdVQharmoVJSKzVDrYaK4EHv8n64vfnbrBongNxhBXaGWMp444RZ3V
EVFnOc1z5JW/arqL1GNNLgG0jfHhkrx45m1IR2fvGBtoMkMIb50WRJnQmZ7zVqwvGFoQrE/cCQfY
oDPRUEa/uF/KJyQ5Qz9qOyZ3Z6zOuQZO5Zjckz8k4O+XLdKBixJf9vNCfG6aMcM9fXGO+T2tQDp+
h3oxmvF1Nt1cJqjkDZnhZOxrT/g8/4owfVzY5HdrkhYKC3CD6K/PtkacCZX/QDiwvLtjBWFpEguf
IZVUt0oEDP5YuA135PM/PUQxibm0RTJFLDK4chx9AlAE+I3Di0PiZvRBP5u9rwaJP9w+hRRerx46
/6nxeQKGyVYM5WJzIqgI4yJ+a+c8yzzGHER2y35oOVeszjt/49oS6Pt+CP9y6oxgnovG0JlyAd6K
GcpaEK+cnmWCECkZ1xBm5vnJuiSdZUAGhN4cxpX4H1Sg+CgEjQ6LI1jgHzP1hsCxFshkADGEsNkb
Qg8dW2h0kHCDiHEWOBWL0bbvt+LFXSxlCB3HRpf7Hz+2fLsmkhvFo2XdTsoLhf6IoSqfp8Y+4g+b
XuqCAvBuQ2uFxOM+FCY/LrltWgNiis5mTJu7PTvBgRG3wo6aqe+m4xLhhRyiq+eCWSLMqx6Gi9Bn
hkcD86FO34NdQY+yx1YMBN7FP02HFg1xddmgtt7ZVEO1KB2cSgGOJgxmTtbQj8tk8LUS7ZMs2NGk
5durVzs7i/G7X73+VSfTfSY9Zc5rVR+VLJinQ9SCmvELa2l2scRL4qgx/2xwOxhcf/THbzDtNF/V
tORy8ajmdCmUcXIoZd6DNV4BJgDb+4WpnrIq6kN9MV+GTaSQZk1W4FRyuv/UmTjYUjdcGJFjWv3U
mT7RhqhNTC6WcONIP6D6GQZmdvFK1zOFJAiHLSpjgtGO1khJWMTF+vf9RkBKLSlc30d7h4OcRTzZ
Fb0wdmiZMODMGLGt7uXuiF2SacMG47QuPX4DcjHuJYvHS1+4KpVI32DEEpLKMFDVS4PRzaY8soL7
AI915y+/h4TexmdVfV/bEuQuT6Kle9gCsF3j3GLv4eFOQvjFnIB4Xsj8v+sQ2q/yScVkhzMMlEH/
n0LamGNpA0En7GvgsDytRYnudm1FPdDmy4gF9KKl5uxhqEmL8Gk3OTGOkWmGlF8XJbt1Zd4u8HbB
d1fuSua7UZuJuHq7vgIqXX0nEF9nNNAP55ri/uFO6OXjABdFZbk/tCbQlnsPEFEAsRNjNvjmFQiB
E3lJWbTXJSFb6uv1su2jaQYAOBKaNQ8u/gIP8bwxw2oSCXblBMdUudXYiaPwwNonLjzyRaRc27p7
lkD3jmBS2kZwyx5xWeJ1KxJRaVFuyZLor0oBWklBg5FhreLMWKu0EWUkYAH+Sbxc4lmUizlZDrAh
2xPZsQ5NlDgm+LUWqcgr8SEmmaRot+3T1AyiujwbYJJhdpeyoDHmqT9NEG3xlMboYY+lluOypsag
C+6sXetMmffAH0B/wL1t3e4clH+E8uKYaNFxoPCsAh4+yR4fMS00/ihs/1+yeS/HK5PPpW3nodVL
6p24utS9N57pzpkfRBAfLVi3HEK80TfCkTiYonf/719m/J5BmILCykXa636ROS3WEOeM3UnvaeBC
e7el1Mk8VNhGFCyZqmbivjIgD5VqTkp4kjSyM4UzNBVuOt6NmGF3jLDLiqMTFyOEj3/KplQQ4S2K
yoRCtPgBJqhMTaN4m5YJsoDOw2kcXuaS73yuo5X72EM1j1d3pHIZwyjy6nqPUYE9+isAj5fMgLzl
G4KblIhM+UJ29403k5XiMDtlHG91hP1/GS4gI9DGJUgbOIzRW1NVprIA0LGYTTFQr7vd1ecXZIAB
7EEVCZsQ/acADMZFxlBgo/zT4b/7kpQDptayWnCeCtQKBGS+XC/1/3WcQKQfDeHnhoUaK/c91gNS
JcZ9LiRA1e7jRuvX/FQiHYzavwogMVgKOBGigqHQQCMoBtfyDRJMiwLo3qMCYMKj1Fp/GC2UYYcb
XSLQZGUxM60l1ePE2GDv2NIYtOjfw6xptJTDZVix8psdV/F8YJDcRproKlskutTMF1xEPkKaGnwo
0tAjAFa23cPxMjR7CAbMDG6VQyrFdPIYB6LfsUiZQ0PLuky9KSHUFA2hi8Q/OxP4CTvw6smK4hLG
41kJi8Nk0wGw9hEYP7mUSxX49uK7TSMS+ksJpW3IkNJe5NTw/5pMXHw/U8FgrZwok76Uluo4dBmC
01zJ/Kkq+0wsgmc7qc6MHD/E3js8w7T/PYxt5cgWhNcc/ROIBd0J7iojf4/tRFoKzHld5R9ievUn
k/I2I2QzSmQKdwaNo/n297UEMUuhFCFEsZyCkuCdja8p9LMJouLACrDT6G/6tmIbhWlZNzjqWvS6
QhCpCPjBXP/r4Vje6vY7k0rH9BtWXU+OOoB88Y9+UGZD2NwqYlbDcLyBT0hsjYdfG71NBVCcf3jf
XgwZT9GuQADHUx6eMcNWWrU4U9WaK3NV/ZQ5p1WbIzG2e+pKwnSGMde/twRSox+FZH3neZK4AOrX
BEnS004fsTaYCYtQSZIB5oRpQNoIIVy0UMi3z6rlizRwyCOAlqLNY6XEdISsZvtl920X66prNv16
GBtZnOYRmtkbVkt+uH+fQb2z7Zqdgjv/gNgI2tSQqwR3gB7N+Nw2CKb18RRoxqI5H5tPnnuFCFaT
R3YxVMGVjFtf3SjDCKfTSbYBHPPc8hOG3tMQuJwT8zf/QIDkzQeA3JBeS/0h435py7hv07G6ZbU9
wt52tQ8WjFrIvTJXL9PWueegydkuZrHJDbBnp832GS/1Yp6Oldd7wplxtlUoGY32Ifnbu164+eES
0hgZRdUc5QxzGQ6yLOU5z40/kpLJ/Ti4YMKIER566RwYO5jJEFq3vizHFJ9OV1Lc+SfNHB4lt3BM
Ozw10Dr3JUIZN7HEhtQlGpR1taWVqrxPvzhgIte9QGKWwjc9RQFPWyutoYqaNlcwobxUCXzEV3Y5
VUNVfdkETBYDExrQToclN1U2vXopzbfOkkPtW7As5nie08awhX/fIi2t2vLBhBYKAH/khAoH3tAb
ZhH25eSvvKpbVFd4Y8DeAC0zDiNm8VfOhFVArCTYYaUmFEOfIUA6pArvnImvrtBh2e0842vhRq39
nfFilmiEOIgI81jFcIkT0f7WY/2c3ItYaMfutp50k00hISFAZSBG+qn5nAVfAQht9oNxmjaRaNDp
AAQUX1B4TCtyrFJjmiyEzQeeT5wUL3fWotDO/566h+/8Yg4bB3aoDLS0rbhhVWRF+G4jhqn0RS0K
ukrUuu6cEa1arMC1dXG5xFHUOI+QnP8Tyndc6jQ2udKAO0s/zHEeflnVgNQmJEXzvhoMJt2c2FdP
tB5svshwP67EOsyb2KmXb/B36RwgSO9/h8sFJzjWRWImilgU+yHJ69OSnPCtU3cGeR3vHMzzV2c/
dzOCrQPpHSpqzA/kFk9Af3RZK/p0cOUXKUhz+m0o229lsFFy1IqvrPVpQ9e+WgWQ/kpcbXTUX+lu
vs3oTqwTHDFooalGfZMS+J46xVrHdyZgtWz5pL7E1BunN10HDYtHhjQy7GyXtoOvvxUHlbNJ8EHY
RNcBgDeQnFp6SjsIkX4jbVI0rj6nXEnk/JYscFZogDCHhfvcw2C/D3kTsFz07JZ2IXZY9QxsvrGR
+PISWtzZuciUeASy0iWtcXzW6xSShMk18u+S5KrnzjYgFPoV/fOUcntNuCJ6/egp5pzrW31AqAt4
vnzf+iAL7P/jgB6iJDa87t2SBijCq7zDGtogmIiuAC/GCvs0fRQRbpXvzeeZ/uV3vSj6wn+Z6mU+
LEmEKvC7F2n6K7oqVOQ/Et2EfRair9CCUgIEOlplelsztcWX/VGkGZ6kxi7Twdc4x+/JMFRJq+XT
vAxw4Tli0JhSZC/vESdQOnrbmOi7zaMsmvxiT/3ULh0P4KIvo31zwIuMe/L+Cey6g85WLzsBhHoN
kNncjNlnlGz2KCI/aHIRovqCIon7Rk0whpQWzgIwXv0Fr+9OigXkxW124oDdlvvQLUp0muG9VkZh
4NyLpBkSmR84P1IDF47Mk3z+ppcgAqpZAS0ukPRqvyh+NGl/UXqh4KZl0LLil01WLzJ+Nb9miFiN
vWucHalxaZFpg+5lDfegd61a/x6cNO6TNfOaQhAaLXxqlQSl2G+c5oAn+2XinOguN9+n3Sr+Uynf
WNbSwJNxRC2jzrQqxcSMIkzDQJF/KDVEGQQWZDXrmELenrsy79gVnrg7lzVEIUyrKKIeXRabXKXG
jMHHr2nGCPSfvlcvsNbyHo+GE/mMeQ3iYfJFQhdySp7Z5ifUMTcDDmzL1WPYSWWlxwIcNglR45B+
QER7uAWy0u+c3LkMt+c6id1QsXJklLLraDqB7rwV/W6VUQ4pbv2MWJCkkKXPjQbhsNFVmnXg+k6B
wTY2NYzTim1KPWKQAYicpfv2sXANC1Ff57yrE13rg/8AG1tw29dnkjZ5Lybuhj8Bw6EB5huo0Vx1
UjqnDQgYZZKS7S5es/ANbGYQ6BD0w0wck4eKrXsWcRRkbLqQvOuElTZKCt4CkO0x1zRP8onkNctl
DNQDVTu1638Utg2uf9A1/Sssdkih5wopbbz28Tit0CJnyXtzBjFRkyQnHf9EBaKJPDurK8aj3KYv
X0A4SFH7LBPdGO47+m4+MVHGG7elZJPfKicrBk9wFC8j47vNzO2c6sHDapnZuT0zlaR40OPi5PQK
4mfbwiPahdnYrjPXV/VRey8NlTfvgDM0l1+HbIhYCxotvokWcC4AN560kBohRgy0DhNgq+jEIbbl
cbs/6OEGqEFvFlE4vrJONSVPAHGWjKVXsKU701y22CHu29Jhe/Nph2tKXBjqkaHUdaSY6BpkoNsN
eUh9BKUahF5yxLSfffpt3mQlivbcE7aRSowa5MEAuGqmwa8/7mwtcrVQDIKyxVikNHlAtK1gKr5+
BeKjh5T7SBJaxCsPYhrMN0kkYbXgGQkbVRqG2uEYsjOj+rr3ebnTUyv3WpeDj9SS/e+6EJdGArNh
OKjYc5owBFCtLDnqMGNT+10uovjB3+QWx8+dTHONqXki6adqz9SB6peg7ii8ypO0UkE6QB+RICbQ
3Sc1wbBW81KqOdFJ/eGij82auivoWw8C5HLkEGqDSfLGEFFyRUc5LDyunQ6t8ozC5zZqPrUa8AW1
13obTMivKqIJAprRz5okLxmEdvhrLymQrkIEEZpwu7mk2QfB+1KCMZDV+NeZ7PqwKbsr/3R+0HED
opzBQxKX5s08WoQ/1dDzlfVSJ0WPA5YXlLicszxxR4pPnei1uo9PcwhV9/fXige5tp/l/wEyb4JW
tUcm/wce2FB//gmg1nJl7tFFUIfBBVaee3eybZE8yAGum4Fbdp+jJYv1Ryo8yEZ8hLzSPLAlWLSR
ZxIFR53hB/t7MaiRImABu4kFZbb8QAnpMBqcOcedcq61DGtnym2rsP1w6o6XYTkbUYHbh3Z6+SyE
MoRkmuJU0j3XkQoRNINo3VTn2OOny4uT/NR5UXGCDbNMmDs/LmSGh+QCH+6AkNEu2EQhiPVOIn9L
D8SYad3p1lDQuDQ35oKXywNu0b0NP07QjgdKekuqtJEe0MN4T6003XnRKb4cc7Dfd9A3sTXqXeUX
9nrIBsajOyzS64lrllkAR3+bfIxp7o0nSD4V/1LwU50ANId3Ybj0v3heTsP07eqE1avszolyNhbp
cBy9Hs3LgptExUog8si+MJ9Kqq9lLW6WSoP5RoFCAmS8wnTHYFJrFgCHxS7wPapGvfH//KBme6lW
Qu+7+Jj5htYjzFYYfznmxXM1qHzLhAlDXK2sGM6CWh8TX6s4CoBEGhdwn3v2ER8c6Olbdn17SeDO
ZImKCZBXRo4tImFdXUeN6coYTCP50fJCPkNSEvKJ3NKMGpUsyE1yrv1Ev1TpY5T2/P/BJvFBZpKr
XBSirzlkcN0Op82o/idtkXjUi53PUBbZFqekyT8MowbF5p0itkZ5DuFDTu03saM6Dv83p3TOWaq6
17xfyJW1izFyQ2CIRHeNDcIW6CTy5eiP1pDEwD5V/3EM03X7gtfVgZ83J9aXZGpf3TF+OfFVoxRB
XlwBED/AREXrrkiwsrtyI7uEJQNVD3RMoVKYl3DM02rseeQea2rBiiP7KONV1WP/sUSA6IfIF/2s
CumAZbPbdS7Qu/kGJBQH7LF1JHaZqkyfyVHkrxkpY5jeEobfOqIkgFJ3aIRHWK4qWH6sysgHv2zX
0EIq0l+OoLi/D7ERCgIddFW6uODRa5qk17JX3+duVtQHhVmpfKb3dfPzueQs+1PA036yJLvK1JuZ
ltuKLENjETNU4xyyfqyckHnlXs4qjsErlfI+oVEP3KhvvBogWMAle6TJ0vGr8An3gIHFMqp1hcI9
u137vlSoSgJpS2WxI5Xphu5bp+oQyBaAfrimxrULU7lOn05T2Qit32nnY7Ouyz4N84SCEicIOpIr
3QwJMzGh2EgbmJjUHrY1pLJLq/qVX7AZ/9mSU2iYhjOtarSc2y1gWbY+g9pArRwh6teAno4dXImN
eXDKyOTjY27Vgznw/KCzBXmvEc9NQGhwifk5Gl8040K+317G/fYp9PljTj81JVrbBOkCbOaO9O92
QopWdgTVl0zsSYys5lazzi6HIvf+HssK36O9kcVvIj7Hr9ByEvU4Q4bIxsxSSv8FjQLa3Qfl6nBG
5TR6djnnm4qT2UJ9jjIwnGgnDqzBmne1xN0vZ6Frqjxp6TDplSMdTqyvHFKp6Hw1lHA1K/NzugFu
Ts5B3+Gr85JTrfS6fZp9RlT0VoO6JnZLafClTcwaTd2YDgm6bNO6RmWRBNLdMDdaRGOmcAuLyLIo
k/VCWzdzOpXkTDFiqkFO19IMBdPcVjKUcpKmxUuM1ntHBi5R/SgbwHvRccp8ijIVoC5phNyghu3U
l3nbb6g/x1/kjZLcfrQeWnP1TDtJPoVs94/XxRwfzFtdSiboIn7kOBuRE/3Oz3U7PJGjCpleWAMY
bvSgvt16fIbsTMpX7soINOVZ2KjL4dbOaLp1fm6GWQMdzUVHzN9cUxsLJvHvNhfFUBG+qrO6sZNe
k9NVNX092zYnjZT0zIVmJh/CkGIgaIM0td7fCMyDxCW9ahSq1yjOPEUZq2eVUnw34JKa2v3o8lff
eGSAFCyhQB4pU/f8YE0gsyx4nFtZWxlu7gDEark9nH/vMdzGldwEQ5RHoa52mGHo2TBFxR+IpSc0
GleBufepjvCx7tsVMLLTQsNu3ReLrUIbtM7yANGaOJND05mjEod1PWQ6L+obK5pobb+p8+TGYfxo
kvA3WxVwpBv5AvNPNwHaM5n6DjQbxOjpgi0KoBmmFCXuQsVncKIolgsO4Witn/BzaoWZAKmhIzGM
ZF9qeTlKySAm1SMCxQtcLbqj0zKrEw8rI2JAsohjUo/DEP2gQqkZKS6PWkPK465IQsE8KoJ8aWv1
cf5zUT4NqJwo7LlnNvO8lk4aPKRbvBqyLoEM0fYp/dTmBK20vRaEqai/pUMVqM2YJcK2qDC98DJ8
6iWh+BHvSTYkqJSEkgyG5EtBPqiRVh2Uk46ZmLgkygZZHH87RJTVVJtPa+AObesv/AMdcsKCeTO0
XVV5+5mXPQ6VE1BUWTlf0LVfqvS/CSX6shELmuKSFBAZeczU2ZIU0CI7fNwkAq6vN5VcRrrkAofp
v64B5kmrUDPEbOnFIvma3ubM6+3mZydgQd5xTk8A2QeMrtrD0YeCZb3vcG7HDc0iWOxWoD9yc3+X
zC58tTlaG70/mf5yH65lfIq1uQ9zYw8Pijpqba9wvOPsrHF4Cqzs2KO438FBBl5/SzQDRxVm2947
mdaqdFiwNcfsjCCEsNlgl6f6jPtKZxkDsJjOR1mWM61A6BSMIh6o3mkghoYmErS6NKd3exaG3W7a
OyP8Y+3uFsDNH2prQdMUa1/BTT8H6sKjj2QDEYVgJJXlqKFPF5PmghqxtoqAEBCx47RaPPDHyB43
NPcFb85hSi1dLXtHKvhu0vfgnijgAyjKpDdM2PIuZR3+2xN19AzRACytrIFynjYvFi57EN8t9pkF
gXV/hRLvgFTJm3H0HV2gUWMxkYVP/nTZ6h976t18MqCPLLzaTz1yRLZurG8SiKnbDMICUmS5nzfw
oAkCi6QQriEsO6sM9ncYG9Rz31rImKTpNKTbIQucLu0oqnY9boQhzZq9BZMMdlAApCQwPtL1AxA0
PWfXPfTbqEINe473YBO3Vr5oHs8z9cTxMyd/ZIKMckJ5fGFpDpOBqSWZB0zUxsV+ecbtG+uUQGyf
J3KhS+eg+E9fFjlc241AA5Utr6QfrZtR0eQsNFsGTnVOKgaOLCL5+hC3pp9kmtcE09VUNlJIrBcE
Zvi5k0P7QEbRGWdlXoE9OZU+f9Ua2XOLiL3Fn+LuY6EzPTWzxLOT9EoPj9Oytp8i++UtZFMzOvjN
cQfrPD+KITTp6VxKaFMkJC9cSYZDGYdMsRgvDfG2zriHkzAM2J+ccjZBx0BovYqtq/KvLT6zDdc5
N5l3EUx6H/FE8LRcBHbICw+YlQQ9MKBS/nKUtySjWebUSJ7XYRBeaUfV79RmPfcw5U2RjfpPQpQj
EyPGLtHmdxy0C5cpG9ir1fvFAR6HPa3tonXR9SJfrQ8j4afJWQwmt0bR7jBDsWDq6TJldlYRhFap
62qA3ZkfRsuvLQHAG5NWdsjD6NFIePv3z2FaMp89SAog15eVaxEHyu16/z9msXf41rz0pHA2PDPA
r76U8gxMATRG7925u15aP/0y0zOAEhKjbnykEOW656ZBQRE/poL8zM6cWsWiT37GN2F0Sw+j36WI
IcBfuE6vPDTum1GTLEuUTKOHK8I2nFo3u1r6Pp0yvleW4/xTwCNUlnwxzIpDu/M7DUH19Czg/Uaj
g2KRcKopcfoyhGFy1v9jfQ3ZymNovGFON7YtaOBVJgFFckLINk9vR8+pMNVbNe6UqxjOrvReHCOg
gsXYQs2ksjCKSn/e0jiEREwleC6dMKLxwBGIS8mJfaXaRNNCk1b3Fo7dUNIAYo6ZpYe0DyE7McHs
YsOOaZEfMAiCUnxkU5/gOIlk/QtcfZrzB4oDrMLUgy2ieUtaLECARSk+1FwaPgfOJ0Rl0ORKA09D
i+rr5GRni73sdloEDUsaAR+SLQabX/71phCEkAiQkF2Qxfejig4K+NiajX5aklOiOXo4MVoF5hZf
VfAoodcUe3E3It5BCPRUzHaGksRoJ5RMQijoZ3mV2+65RSzqxpeW42YGwTYqwGlAFgCR+bZgnqnB
6O30taKpdj6TtZGrih9gvtE8lc5HC3n+pDG3BaEmtCSevi87lXe48QT20jI2okegR+Flg93du3CU
/n34SGCpYsOw/wzu5LsWyvk2SAut+LkSBCJADXQdlqKua2LLu78hId08GXDqKBEuahZBPEOzrAW0
syt4lQeuSdVJMn91XAdI4IAdPYu4jH/TrAlOY+4iuSyknsyZULs66O+pppQr+bj8my7BtEDEOCBu
Ir+YzEoFWvbSUhvsIoNZaSEHTq0vPBb3ByYPVzJ49wQCB1iOC24jmMSyeJ9zeKVpiQ18ZQyZHKhf
3fNifMZuerSFJIfdIF0hJf87mfWcbYHi7944uGZM+evooWsyE8UM9Lj7+hNtctr+zJD/tzwJjGIL
tS+fasY9C4H2sBTIAlu28rVx0IFNCxAwqdv22OEpBijXU6MC3Fgq+F+L3Z6FJhSnl7ww9sWHfBCY
orXazLT2zD4DUSotBm0eFjUFRk2o4Wa/DF+qF+n0z+fSCDic2BduWA8SOfahHz2NHD2vfvZVVgwx
mE/NP/nV4pd6vIa/rFk9j7dltxlko7lC/2cB/G8TLvOSlJqOmFMNYmHX9j9XYEy4308lbZdru5Fv
7+fYOmT3Jur82WcWYLQiAmPOeu+dlN46RIF13YlZaoc192OGDcqq8TC26UZTBuzuA7GsmjMy2idj
xZ+LEar6ItYURAzGjSP2Tbr7FX46HTPAyRHGrfR27gaQ2ssK4VlS9A6bkSRgrjRiEU/Mnw3ZTXfQ
Qs+PG0oIIY/SnqpdfHz9UrrBmFwc0HZfraPALRcMOtAT1I4oDHwkMKxpDN/WvmjsWEbZmI0W1YgA
Q3PI9iPlG3IBLP214aEZQGyNQgcBc9TF+KHYg2IHQ+6zkDJuUaGX/a/P9u/xqN88AFdK7w/55tn7
jZXWuZr+ZKnXkKkRK84dTaKL8/Ckr8XWneOdPh+V4Cii4wuByL9lcGjpisD61DhZmKfzIvRXTv8i
BwWQlQZPxQxtuzwQQc4ffypv2nBk82zyg8X+RnCWkJXxNyc8H9TE4cU7+W1Wc7Crj73cSO0pcrm9
O7cXn+AgAMwl6Rk/0fJJtnijh9CO1zol7ovhgrA3QryMJTNR2NWb9hU5Z10OoHuFmd2sxrcZRBb6
DnZo6uXi08hKzJQzsbzLcbm/kgp5r2MoHG9jWdPAu+NF+6JABlFVQB/D7ix9y+rJ3yOzzZp+rzTs
+/hjADPwa21cIO3BKUyN3jaxjqnOyrZVii75gQoqvlkzSmjLx/t6HVhDbKb/muuTObCEwBhlxaqU
QQ7Sdx/7IDHoBLJhJMkD9LB1OjfjqRS4O7AJHoNITqjLjkyNpeXqShXYLJVMFtlYWeqBr6K5GnI2
dvfV/zkQITbESPpfT5Vc/x/P/Ssdx7wrZw+EYMeUWamKr0ydXNC0NyHkVbmFYqNuT6mfa6+q07uf
weSNebn1BZ5id7Zt86p+BSzLBzjJef0S+a48uyhU2746s28P7lyn1f2deItjcQfAMZIg7HUfbNVl
5xMvIoGNBsgKsBFpTLuYQ0bmEHbxH+b/Fpiocz+Byb96obvhmAHynKibLnqTJkjQ3xFEobbbwmen
0bX2a/joKryNckNaKNqrq+IFsrYjZVI3L0Om5y8/9vFoJi+lkZWiR6xC8tq0wJPOGG87y+AOd9Sc
xvEBLraQwtpc855x1HxdmnB6OiU+Uk0zydli0KUsb88UHnVzkH44sELuhvuzTXkeu0HKAtRWdrSl
hKQ6kmen9o4fdnHZRQ8DuJxnRCNenNFg4eC/77h6Su+NxE8AfDeQNCsHaCxZdQR0Jh0qCSeowqH/
rLCrJVty+CBk/oaLj+vGAT0Kq0w/jBA7xuenwdw/MBdBQuaiVf5qM1KekBzlqJhvDlLtrC/KOPZD
okT/Tki/Nxl4NaC/99vp9UPK38t8K8aCt7cdILTyyLK3Mr8kgI3YCUy1RiSIRsstV4/HuzcQtnEI
WbxR+yC9OoUSl1vdukUxblOZa8QDgY28su9MKBZuW1djBkkmNIEjHyc94x5AJRU4vydLGaQWJds+
YpArIYSCU/vlHcAAHdVnOmVbplz2ZFTOXhOUjbHARC8AdpCixlRuWKAZAYmw4a+r9wShEek8zHEp
dWvQoC63gROJuEyZ1afAgQLC0Z0NLyimjMGviBf7If/UvBOKbTjjhzbSeKS0NGO1ATe/NCG2APFy
PGVr3fUoMaBvDov6wfr4sy20jvIYScz8Np31dOsXNAlklxm/TjCdfON3LREot9RDHzKFigfhwkiA
jTNhPe22q9Yf7pMuX8xt6Oi3Xt2WGLcJa/pgvYSOxEKUW54WO4fjua0Q9zzA9Zpm0zt3Eq83Dg7u
Pi2lgLcxnLxaXDEPfGyhunopxzPd2j1M9cf0lUyyXOV/I0P5/nllO9Eqy71NqLIyRHO44QmPpX48
y7T9lefZN4deAF1ocl6Vw3DOKWgzOuuwIKVdDEzwa0KnXeu3Cq5jVnGKc6HEUcF3TvCqtrQJcmgT
r0r308855H+D89iiHYl6ECC1fbblYaim/l9oZMSNWUs31Y5sQt/MnedEk6ZAH6zGp4sACSmvJNam
1p4QgyZ0E5fbfmj0STP3ymPxCj/S6ny2Ake9tYiouPt+mHubdXtjeZdqLZKweDIa2oZAE2bpWz2+
DSI/p1aYc03mi/X6mrKsEn+nKtmp05ko7wCXlcZ10SE3IPHHL3c6bSetoLOC9N/duYly2nsH1+cb
p+dcTLm7E6VWVB5jG+guU9O5krys/VAu2D8kvt/xC/sWQp06xFlu5jbpQ3MBHZmZgupMolESdYAn
IpSNErEaNpaZrceXmevMrMQuqMUYJldrmwGunEVJx4OusfCU6TWjHx+PzYRTGO/L6DehUn5eWH5X
nIEnBvdjlH6Tzd2awJHESWoXRLOecZ1wpoE0PsRI4ZZzAhblzzJHJmNMEZTAaTYSpFCPsPy+SUum
nNL90IVe5XGec1+ZljI/Ap3ORZEBY4PNc5Q8DOF8auvfg7lsy68iQHr3gfCQgRgZI+af8vkPp3HM
+Mrp4YYNwdhRIoZwQzaeRjLtna11edJI0pe/JoMjND3i1rybxIidp7G/L8k+QfsyPKYOfV50UyxB
AFjdtz5qRkrKoWnd6x63TMTTEn4pSHE7SC8bWuBriJK3aOjABbt3P0WUcbBotY1+iMz/KanTJBeR
VQFZoPsjyKCXq6fEsPdA0JNKuw43RjCgGWI/SrqZuzavv7qowLVAfsMPLh+gEnkgRfUVb6xebNdH
zUKtQPwirkazstyFDkIxd0SHImCe6z3Z3/u5EjpitALzWbA4pCDo3SjrqmrivIG2kkGPWSM6PUIA
Et+8pk7TR365M9EVcBa/cORmfA6HIof4JcR8w6M5P7b4Ubr+vHPyBnBSkQfkWDsku065/DcOAxXP
dpqYUZEhuIEjjHcQLyf/wAVt5wWN5sIHVVj7BwnohQqrS/r8k64YZ/6/Ypz/Cuv7NVsVHe3QpZQP
HNm3TVhYCEslw2hzNE3oJpEjql1IEAYfqGuB07yMbItCH7/qFMdR8BL2L0D43YW7/bjXS1/xbmAv
YD0rLDhOj2ZI4fQLDvPXYJ3zlddzp2rQlmVmWa3/yaaEUOht6bzWGQUi8GAn/za91ZhwKuHwyJVW
o591Wgw/Y+Ro5zrcpXnktmZwc5q82425CRAJjQVKHLU2J9CmB4s4duh9A78rtE3fYva5tyoQ35gW
WquOsit7Edn2cP1xDhPya2HkcFnn3etLCtLVT/PyAgsXjwehHtI7zeH1Ak5GVNRV2lDoO91maOlJ
dkZafFn2MGNNSkJpmRYeq/IvRNdHB5zS60sgueM5Ls0hm163pZOKGt2dbR9Qh1jgY4uY23TToLsF
ZcoJOj2Ux4yuEAQdJ7sn6jRdzBO6vfQ6EwxTmbXaq5bzcvjG9kmTjJaA5ZKIPvzO6yY4aWelkb/E
66c2OHopEitWpkxcgO64yj1hDXpv0slNBs+Ri9JQ6bS2IMFv8k2hyUKkOdmW4tH9aO1ehqLBDiz2
QBVSiWwiOL3aSVD6F4rVVP+GQaVUMN0SGXxlO7nwA/up716n1n6UbfHkJf29d1kK+IPm53b0oacV
1/Ei3mdFnTVwQKJB0uRKPP/vnLtv+oGzcI9tAgux3RrAsxtogwwq1o44fM3Wk0NQivo7xhis5dJA
xfgrmoKu8kK7JypYvP9Qq8GZus6MN04Q2YgwhUqd9PModZAmk13jSVkZ7OKzMdKMV7p5ZYBHJFQT
yMOf75espiruwjXm4tTWSlPbGlDosU6DS6WfTCUuXIt2RW7gHimTIbUMOKf1Qud3Jx16FyfATnNl
OmK34r+Ae2Kfq7+gi4uNWO6ncS3pPzrwzOoSpih5/CYxdSGfN07OtZvgu3S6O7z682Bh/d3XP4hd
ksfX384oVakE/twJljWjHA8DeRAL8PU0GLXtvt3GrZdmQy/we+x+3DxzH8yCyw1fMgCCWBH5EM0w
LH6R9yh2DxkXO0ySj/Ed1kd9iIAZkTGpAKbLnyybjUAQ8qoUq/yDy+aSoMSALOOxUFKLvrK02at7
dSQhRr8GjO9lTntmF3/rmE4OUM6gNxR/wWo27JYWhtwlqRZ2lxc0b0TNb6625/b+d0HbVEdolHDo
09hkayl1aI8PbImBIxwFwMVu32oiDxW4aCtmpFZF7kaR6XpeHpvoQm+4ExcZtxbnW5v/lu9OMrb6
9NkhWQp2xdvLEphwvoaK6WqaMHRMvmc2P16AJdRJpLB8wST+MqZ5UCvBgCHr+Q9P+R4XNmnYgL3W
zmK2qGOWvJeLcdWbt8yvFoK/JM997jYjXUvH27ae6vBDwMm/C3Sulnv3Z2f3tqY+pUyurizeKAN2
FX0a4F9VZIX/dhw6ziyGqBlepseji97KU1XorQkV5gmJDeQ5dkCJkPhpUTyxKXXo/apy6S6EbnZN
DIqs9GpNRHSQcX10+MI9bE5eldvu+dbPB4cco4TmqSFwQ3Kgivj5h/HJHcArXn7myLseoEV9CvQ/
hWnWxGOd+NL/NFJ0Esb4w+uY7x27sOiH5fFQgaiw6cEG8K5OdzwgWC9iUj8+YfplRGVtunSXIiLV
HBJgxNmVwFsjcJQWtpwCbkVNqm3v4YJG06C9v9T/AveoKlNqx60JLTpE2Y0TH2QDG/gT6evgqLrY
LzUm08WbV9oehNn608YX/YViImyU7r1ft69I8rQqpqjCz8gFxBqbZOsuDgPb8rVdLN6YAw4vEyqD
9oUR8jQmQ2rSZEmGs4K96PPywPwct+ccQbfb0FwHoUJCWEeAoBNo4OUklIm+mdtiCg7a3IsV/GQ+
Y5Ie4FnPnxA/Yczl5dZQ0NvvQpJBrTOV5S6RJpmhtt9ngRjAhfX2RYkelWwqmmYVrVIpqQEXYGAJ
bp4kXlwC+/M8AFghPuWVZDoGRnqU7BOY2vkDw+nysOrBTU85MnyJbNUfnown3pnsoygszP3ni+0p
uYe1Diqmd3xj4nwZx/KAzVxWK4QShPfX82eph+xLUWNcmRHYZuNj8B7bUf4QxeUTiEk/YTpklYwn
1qTebJWgYDQujWCOEswV4+bg/OgGnLgbZVgzNHuG8YOtyHUTBPtZpTn+kwycZq8CH7PNEQbTlVfm
aUj1yiSi4WUE+edyTq6CnCyQZjHHj87EKVgmwArsFCVW6dA8kPf56WxZPslv8tjBqMQZqqAz9POt
TzDy4MkyPzVpCopgCU4LZBzI9IHTyG2mzlClWHCZtuSyaHMa2yM3dScrWL2AAHK/mF/xErEN09EW
OxYeJwGlczoFeRnosYCOFwGJ3nur5knoo+pUDhZ5A/tYJivicgqPXNPKrrYHomgF8ZWXYZ9nH11Q
HujbCMPnaRyAjOQYkC7qk23LdC4mk3C1BYYt/1uLeOD9+W00wz9LfOIHJaNUcO9bHFuo8lOD0C2c
gboYAo/F7gEfd+oAAMGsYjkRIIhBJGlywGFLW0fLmdkqBbq8PsqSHbhV0TW2Wj+p30ApRSowzQtn
k1NXWLVI/k/UrkrisIRDR+tGEOW182z6dOYkBfPm0jwH+key7rr+rhnz3LshXndDu06W9uSN8qJh
kJBst0k/ALukyN86fmSw/I8kqFhc5hauYnXEyr/0ICR+oVYnCyp8tk0k6FrJ6gFMZJHCvenTKKx7
8oukSlD7C/J30TUP+JeYgA68c1fl0gvI07nJm7N87n6R86nxYvFp/gc0QCdZFVFTjLwBB0Q17KnM
ZBTiqXxkYxhwTXJY
`protect end_protected
