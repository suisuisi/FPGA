`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LidfS+Ir2q2ks5gVe0rvcBo62Xql8G78EZOOsgdf7WedAZFg4NPhJrZwiv+XISBKCMSlQvrsmvaS
PLiwBEN2/w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aRmWNsckoHsFozB+1r+Tp7sCGwM64BEvhPZL3P8FFOPkG2fUd3A+fYiNc7f6+VY+yRY9Et9/Www3
bi7fDuveMEwmMcat81vdra4/xnnsZWCtBYfZl7tTCYqUftG4xS7Ru76yxNUhZWxKOmNzQUhPGt65
R7HAmB+0HMF3SarZIlM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
r8S3wU4slN6TZD5PFmr3sjxEbCf/VqBKg6oxkYFalIMwMkZSuaF0u5171R/yIwfvdqjecF3ZJPUs
HAn5/DJH1XkDnWWDej2IMmQnXqizCx090uI/PenoEAejSEBNDTMgF3V7IEYZyQC3AdizGTu3Lu1k
fCZLd0vUdSsKSC3xrjW0orDOVNs/lhDaZ2b2O25fMw5+CKbk1RzWXilQlUJTkRxOI6p/R23k/8A/
/zdBTq9CEk83Z/ksYPPBaljALsZ7j0X+IQon7fqgao0kuR90mXxrQmDSsPCJRPkLIM1Iw1zT5ZXF
R1JK0tZ03tMTbzzakgy0EBcNZBUg39xzklGp+w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EDm7VL5RTPdPuZ4fRoLJyLsQMwnNZ1v+I5aRtPOcIVqZJg9/RHJLd5utUqOCMdccgYNXYqoEYBNM
dj8D/Fc51Sam4m8APGgT6MPZQm6Hh+jYbGvuEmutC1miS2Cm+140EFL7UHaCKM21KShK/KHOA+i0
9sicgqB0sMbSNdJAA9WvRDb+pHElsVV0PAsCklVbCVlamfSlpRlAwmQHp+R+q6bkot+TyHWM8oWi
XDKQ2GHM6mXhIjGORNxoqMTUCtqasTh4q/IoVUuHNlZiSSyb2WErrtIhb6wFpqBqzkT860NIsUwy
HNFF5NytTH+Egg8S7cHeizUiiijuzDv27AD3KA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U88LaUq0gE4SvRYG4IiDvHnXD62Q6horN8wuJtFHu+RWnx0kodtGTQIZDxXCroay23QLb2jg5QHf
Ti8sJv8OGKIrRcPjwhPy8f7NAmXSFJzMBxLEmAeNZMLLGbGTcGGDh6KQHPO/WrbpXRdDRUDn6ZaN
cwKUEO02cXdQaFSagd07Er43sQb9jwBloBYu57zxSlweaVd0utIPZ5XP3WePNGbiYBqKUmGeVkzJ
3uqc0U+ZKBAqUdy403TjTlyyQBMfgfffDtyvYSndOScOxBbxDklmPh7FrvigRa0V1FkjTptW25oP
lKKyZJYrJQsR+4BGrsGdPrh4J2xEhp7VDc3Vww==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GusyF95ZmKtQuC5uTLzHCLs2PQGyKsciRCV+m88AgHM0KD0LZ+txdfnCPT8wJ8y93Ra02tge36m+
oyJz0EyuWRxZ7tjJ8IEIHpJsMnX1XuZ8/RGc5VBQDnsZpT1CtWBvedMg14tn2c0TIKkxMo6uq7ut
nq9Zleh9A3/5fqbDjwM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OcMMQhgaBmkAQf5RIMetA1RdgiDYGS+e9FIklvlemWcBqsNjnjmEj7ZvEWTsAosXwATf5zOBFBKo
R2WR/FCMtbD4ZvW5XUNxOvDcH+u4GtvlxOm6rpxgUhAyVfECz+p4c+wxHcIL/JX/jQPmhhc4o0KF
SHsHgArZ6RZ3kGoxktYyF7xkc2NvJrZp57v+zrHy0EekwPaNqdCZVXk4aQmDbaTPa9AqxQ35dkft
3XRJM+5VxFQb3NEQE8JE2E2hF24MTuC/FRq62Nd3f/BsozBtFVsEzkKRTbM+xQR9dqZ6tkbu9OdD
w7fkcfYf0RutzC2zGel2iJaCvu+54Swn1UrAHg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
828edt0fd+wcAkdmOATIYKz2TJPyo4CrJVf6HVNFp0qQ3oQt07L0RaK5+DXiY+ymxStZ2/6D+W4+
FLw1d4UTT8k/YHg//GDagD61N3klMQCMPabCZtEOLVleizI56gQ33TA6mTKK8SNHLyUeSOsI27FV
BNV/iemYTNQd1d2Z+vCMZnWd9M4O1SPe/XloC1Uk7AK0FohTFfDmZYhyPuuBbWap68e3bQksxPOo
hECxsStkyI1e+Wwpc+FHmW8SO8muRYphJzLsS17xrpAAO2h72ZGMySpPpsRpz4Jcfhq5Y4GhGIMX
nX6Cx0KOrFhh/WF0j1kbFT+2fa0yX6EXGMxrdyt2LPbbT3qn/QtF/vpK8+O7pbjYi6FHeiMjSS7N
6+EsCQDWMogDeWP5SjM9B/M9D9wkadQJ/oVDZ6aMxX+EXXD4Z8HSdB13tynLVe9HYTlR/pAGc3HF
3wVNYXrVU6AqKlp6NCvdHjrux2iTbFY2kTEcnIA+BHBTwyo2r31KtchnDXpk1pyQAXChkXlU4N8O
Kh4ZS/6Zsxr4lRxDLmNHIt+wbofBQcO6D2YMmHjYzeZc6YOQ4plQ7ZCr0VqQaSY6hd7LJukRTJ9s
1p9FVxazYzWFR25SVdd37Oohn+DX3HF3Py/iMUjQKpLIlyKDC5c58SrqZKFF3F6vpccFqVa/+V+g
qiS+Tc85r1bqxZTygiF6PMXpt4Tf1fqF1wOCWhwnp5i3xhbzfQ3YVNnnim4wqxgMW3OqhWXz6hlr
J+WHpogr8Sc6WV27r6PKu/HDchCajQ8+DzM4E9jIwqRKtHf4+74ZsUpG5pddcI5fOlP8R0pKZxUC
PRQiiQHOlehF3dz1VbneFCqDN6yJIw6mafunCElf2ZI/j7DH22nPAYqF+RY7xqQMoMKRLqEE2uI5
zdULgApAMGACLRQLYi/carWhhI81TPfAxJ5PCTEU6tSkQS7OtdYAC4eZ8IXpIJl5pxFbd+OHg9Mr
iAIAUsPsPrh1B2g+KvvjuMUponf/oQWXe77CPri8RTTO92J55FnemLQm1PDG4oWjNVpHrwlimczQ
JgKcg47unnCLLOrqPN0ZtVEVZOigLvPx01OWYpEIlF8CSh3EfTfR+6U7yIbcloWP2oCRsd6enZ5Y
nh1YB3PwLrSIUR0QgIoHkqB2CXz5CCfhUHzMzNGbPYr6xEI24DPattp0dBny1LjQ6CoQ3cMqBOUT
9+LIsCr6Jc7wL1TO4kc1OC4nrllw/WdIrmPN1/y+pXxeOWQaP9rR3Fw31zPQ32C6Ywa5C/s9LXqM
OiXc6Yl6aFWLkQcWNrc7KV4WwYtbxLUEtMcP+SxxQQz/t2C6x/jzj96O3G6lNlMTAQEfEwJQhQcK
lkVnHdMNI6OqfyCjL4jGV42Ow1O0MvT9hOQj1gLBm1PqJfLiUc04g3T02lNxZJ8AFlG1U7m/gJxz
TtJBCpuNgNRlZwOy9qRhWvdo3JJTvbPNrg8qsfsmbyW5zqZeIppzBoidHAckQDXJLzmOP8nr0moL
inbLkr1F9DUBJ0LCOYKrijel0dukxy89N6L8o+djtwQcKxzQhR8hNnprbS7oxUSaI8Ic+Z4mdneL
qdVtw7ewkZXGu7ZLWL5dMFwI5alezfGgziW1MRUOVHFUay5WsyT3ynlYlQS+F0xiLfuvgr+bv8Ur
L4S92b3L+5v/GRto1qsOVlVSco+4Xn193SRyvfNAo2xaukrzNEc/RFOwkj07zq1r8xxnFXEbecxx
W9sD4TQbLOTxT8oggrpSEKZYJS/rzQOjEn536K9dK3ZEklTUrQi/Py8IFCnYEB/o1mNXsjns2JRj
fe0r7N8r/L5sDG5bIsnlT7rVnyk0hULQ2BvOZmJ5RUClx52WoTXEWASotNJJTokYl8PhzGoBQsLL
iXqIeRwosRnuXWugJVVwZW7jZPO+p6VkQZFrlLl6yXpxPD7X3Y8REvYFLM2SHJTECu/jcaljjEdU
TjWtkwp0GRzavUawngarXOpFQISQWrSH89X+VKv/4yHfQSQmAYLeQXIDmbU96e+g5RlMX+UcoAB0
OYlDFHkRyKh/wr9s1L4JFidDHk1sG5YRni3K5XNrl6pfrZ6QELKRXC7Tpdh2EL0sYemLAMw1zlLC
QXVzSpywvp2UxLbR/DysXeNIRNhM7xE6rjw6vHxZOcVrjYlTkjJIVptYhYvHwMSB5EUQ6HkM4Psf
al74kQHhcNBh4L+B7/MLPB3vdjulzrjJTxKOBDSnrQDHesZ50W9Uk9CRjz7c4fQsDKMjCE/bzWMv
2vrOhvfJRrKZbAGTvbYBPfTbXWRInSJfn2xibhWXWLyMNrVhPQjK6CUguWTVu0jtOPrRCvc7RAxF
usw+Ci7XQ9z+u+GqiAF/mQqgHha09IqemLNUBG3fTOAKoNx7rYkWO6owmw+RrP1fUGiLQelf+Jeu
ESLar/l4cvMc4jsLI4NGrqVDgwnq1cUWPpysnGxUbp4qilAlSkUlrJl+zuM1rHQwQ6QxEDpDcEkN
BhRHUIYqZ/SuMaoSprPHmEv1QbGVO8chZT/4gNILNbxzf468QV1h3agVz9llSqDbnUHtWgk4nM4s
vycnC1/NCylaqhZxcV4lTDoX1m/3MqsvFPPqXbuNwtkcdOX2xQs9+O/cNYweT2iVtzdAX+/JZFsA
vY5UL+tbV4O2b72pzqxAfa/U7uNigaTck0ADBabXnT2CFybo6QoTIWg1upO3BtIW3mlMNDHK8XgI
66WUF75cnSXWOYh0+RxzjGGTdWFsbYYHzScgoZcb4ihWxNEh82rLaXGgoE04AnwgL69M9NiG/fpx
oV3VEmjSzvmioUMuvlnen3KiDaa4oEM+rz3lbewR+CSPpwykOg61+/E6ioGvOMSte5GzNYfLVPf9
DtJbCUAYaqTAQRpgF2c+C6rRwzWEjLBW8L4TS/7xrJM+BzgGqSwl9VmuCqjePoO4H2eCE/xmx3WJ
Qbg0Ve2Qv6QQMcczjcQeZkGZwWArbz1w+tFJwOmZqAeyhYCSdQirGwWrN4h0e6W38gytsRMp6yRm
JFsIcDAKKg1ode1aYQjaRNeo6E21YElwcVKWG0M84wovpZcwY2ahysdcJ5vut9t0PUxCwJmw3QGe
uKKUhgbeU4AWGxgGcDYjwWqF2Qwt1ey2HA3v+Q0/jVXHHFXoacAQnYrKhzugCt5mdLuNqckjwhg8
8ZDV4gNKs+BX4AkI0rnZKUqIzQy/NolDQS+5krxFi9s9RYvcJWjNwWbh3QzA4Po04eqvfdVyiugc
v5MSuWa+vd/MtGMEvWS43n6vGlsmf/m3vDaLo1xoFjRa1QqYleowCP1SsamShmmRWeovo4X1DSwu
WGC1ZPIH+ZV3QQOw+4mkrTisMuOvEeSocUB6TWEBG0t84mexcUOj9J7bEYLKSZhS2JhclgOHitLM
P8/p6pevVG5i8wcY/tcQwpypMCZuacv2sNdT7q+nYSxv4rcFtqefMmWc7G+4uViDT5s5X/xx3FdY
PietUdjI8aWSNjuUPJbDO00EkDJD2WI1wWy1YNGwx7znY5pMF0VMh8aD+j4bDZVF3LjCENcl1T/i
sdaSUlRYKMKFPN27HrXT65z291posa9mv/uQ6fOpvbmgf2xFUzgdCFtv3jNUGSpoqmeqb0GM/mVs
cgrfP6BcGUG8b2T1fDk2tQYnGgMnY5M+tWEAsJA1cteftBmKNWDc225T3xHqJEp2S3Vx+vTfswjc
NuDbyjTTWQvpTU0OW3H31VVP1Z7hM3gJaEDUcw+/Wr52pFTgp24Mjuubc4FsC7Azehw5P72ye7ww
Q1KRYtlZHFKN0gLQpIZeOSFmg6ebXBf975W1UdRdFU+mkaAC3cO8TJLx3ePag0acHSjPm6i7TNj8
p5cbQiWZewhtC/DWDtl+E2/yDusBCICOzg0GSxFRs8tb0/xTjJ6uIdsecdzt8N2dSDdSZX9EmtmE
4ecDKAaNayeNFJNDI26MoVs8+WJ+Wbu0QFuhq9yvsy2dINVUHKFPVnC6LV4HkHU77C9KKocOPOEq
qfusnn/yxec8A1xniwJ0DEb3X1AU6wbHUD6T2oNtOjiBKApDy1eA1NwT0nDQzr6Z6Xzj7S/wp7Ht
4cdLAuHHFSqWti8g3VHfh5EJ2pO06fFKedWhVHJcNYnwPnfdyA7MD4kkCqqtvFkotnmV7C1r+Je2
ov5l7KK1ae8yvvvKjHzYdLkQY1gy2/Z86uWT4/VaYP+xw5IGe2/9DcKtN4MuaP0ilLTQzL7IM5bm
agbznM2qolBBlvZFfccX6zZn+R4YmizscenpsMFps5V8RyDvzRy1zHLOjuF5knKKkSrrZJBWFTRw
tZA+uf40nW783gK0ah4EzgzvCRPBzLn/f08m4NF9kMEx7KjWit+nP5vlGpmxPzqK5rEOQH/fu52j
U+ezOCJnkEW7OIzVK1kJH4TnWwTebWxgaGUqwe8VpMthTJh1IgO8ApKtoV2O5jjsvZDflwJzVxEJ
o7RRGBilPIExeu3c2GnJ+MZrgDmS+8KNVov0Yx+toF9XlQotMO3NWrHMcWnsnQnR31VKJ64K+FRM
QnTVz6DhjdDRkspEtxbhXvTN+b8hncNcxa1dvVk0Rw1YCfKkoJXt80Nfinx9B1AIwPu9sBpLieIS
riX25MzB8CFQr88/BhnhYcmfMgV9/sloGjAW3++GVgxU+fwPP5AAcVtFxZuG/jglye+YFKfU5Hfl
I4rV1dnAg3iQVOQwp+S6H9qbg+6zvbkWXFyxonu1fiTXI1QGYc5D7rTKZUwge9w5rg9T7lscGLB9
2NeW5MLLMCBLjTwz0zATwJu3Ajpk4ZLo5YRvJOjy9Slx8+DbfwS1kGsRw4JVj36ao2jCChStYcl7
++Fe7JMpRu+tc8QnbBs0VgjGvik7Ih5///vGxvU7eGVwGhpP7FDyWv2VRwTkAFinI7IMETa/DCs5
WDp8W4XxjxnryQjmFrYDQe/j8HQs/M4hZ476PWUQv3o99g2X38RvAhQ0YFEaJVC0Xj/+YtDJwBJm
yuw5K5UbFF07GKcPAym+aOIk8zOJXNh9UfHzlvBRgn8bVhiZ4J01BOuOqnxJVsd60gpOWRRClb2A
WRprWA1YwDCUKU3L1oOCNnWV+p8Hsb1dqZflzxBmCFTcab/Zovkd1lU70c5CV6Nn4kdDATU9uzTD
MWGBhv5DhuS1YcIJA0jPN1l/DSFIpjZ+966Drj7cMLYbsUGjKfH+y2fVxr5q1tMDwLERJlZEYEAg
bwm1aETXUeFKcdsYXFW3xIJynk1Z37J3zJXxr8LsT9iQNQGHzXuVn5CBNwUt+yVgRmLJeaP2FGAd
9F/8n6nDFkuarzQD3pIliJcbsSl1TEDo5DNmaaozzgyjaLb5c+Zac22+54pvQDvQG6D47FRjzMws
IIiKG3FmL3/943RXvgju0C5EoPh35UZp4hlK7DabkvevPXSWOnUOeJCaR6nKMEMrqbCJ8USJuksK
tTk5IqAxn30LNZfPnR/6CzIC3ffo/v4P9grjKVTvW01jiQrLumlmwe2BeYlOKYEBKqtOOvK9ExKw
UP1R5+35aBj76nBWdhDfi25OQMnLEGFMJ6LD9o8shdWlSoWjc4MGFQox3hMbW1nx6PyPBgG0IyXr
XSOaD9Wq+bHJc3tfrZOnbaYtjez5KtFluKor94vOphgwu1zeXl5gYadjlNqEOw1nz8Bt79yBi7eB
ezpCd77XyddRLCn8d7h2ddsZJvwCSfmnuoz+VHCT7Q1Qi9zZAuj4Ql1D8JTtWjWQhU1CEAScKhfc
aAvejBl0KLlhp1RhiHIZE6yoaq+z8/WnNKcbT0f1ZATXcDdhGOWef5gyLAVtzUX2WgvgkHFEiQX2
R8CInDDvDUXdiPzzxMiJk4fMAZAGX6HY/99zieVY4l96MToCsqGT3f4BwBCzcpYUE12rxfrY2Tkq
uvAfCGdqifmxqRiMc+d59gsLjeFMJOFPllzF0wBNvC9o0dV2tV0O/7tHLb8bwMvcyJaBOujXoowr
vxMGqNtCjucLted6NVLi1nuKJcVr7pzOefGmUm8IlvuiVR8eSSbn6bq54SQG2q3V4rcPMiQfgikK
1s54bU05c7OIHSSB1gKXW+z8qXk084OqxMCk6ibqto5t0yZglDVkn6EGupOqgW8Ao13V8IfaU28R
dWFjtTb6AETpt7Phjgq5Wwl3JfWv510YEQW4n0K7q1R8uGkDP9HwLqAVz138Q1FObfbHCYkYNf6a
CSGXpnrlwVpj6NoXiZ04VcCsQqhruBMuxMs9ATobuH8O7rOkiSBkO5cCT+aMEoHMdRmvbQXiK+YV
i1A2xYQenMfbktPfZfPl6Elf7+ifWPYvdX2xKxY3lVXqz3+8sxyGW5MrLai2iZ3Wy6hIzTDQeDi5
lXqVkVg+EgkXL2lsuY9CrTdxdKr9CjabeWawSEM8tiibIdKNVOT74IeO9jTD+MsTXPYbw/eZ6jdP
h6xfjfHcoe0fjpu0t/s7SZsZUlZUMM+tDHCsLpu5H1Fwr9V6boi1ohMgtcloUjQtR4m4vtuGWUkO
I8O6TBkjwYVi6wKG+pHduDCYCoXERM5/2drsvW/FeuHefcObqRk+EvSSod6O4R4Er0tHhPZR5aj1
Z98PNQ8+FICCobWU406x+A5wLOlYBgi9MFIw6y92mYIsVaJwYUIr6vRJsru7Y5eh6/YUgbrs8HVN
nAHtUfMNH7FIgDoMo8lbrDxm9wrMzf7TInbBYMhaitifkuIwsc36S9gjzZ+ZUcHwE57AhX8Eqoju
1VX5dgTGhH9XJ1ujY8atpczZLVX/cMH8xY7onRpq7JU669znz5tTcwEIrk2wCJd0SWYs3ID5Xurw
OfCM2FppqMFN59bcCjrgtZnv7ot5CsxkyB2mCjTd+KeNkGHukfCXhp2Okcm0ukz/WXXKkUyQ9TyM
5wFrMA5XUSzbkDcM8daEFTIxnZGyxLM9QExx15+YvMsY0MS2t8vqvp4nKiQa1NBDP6CFArifoSpH
J14mh3E1MLZE6+Y4s2hZt38Sp2MBPV7SwJQ2BRkxeH9q+QzMFHQ441BAs+rvD5P6m8aJKhBV6vd0
ni25Orp8sjkVTHiI44svjol6kMFksWqsE68LtydDoj1gn6CwRoxNFHVE1tN3FBvsWI1h7vMsw0+O
xakrKp5alZGx7QI8WIBKJYUh1LBX2e920FXkeBTbVxMicmZJq/fvaplUJHm5204hxMF927WDE8N3
TLSAmmRdKKdqM1kURwzNUuHWnPgcMDFA1PmYgaNXedqnl1hpJRrwS5t7MMXVXUuNoabiR+o3iJYI
4/Cd/gWfV/93KeHOr8IGTw4wa9hEbbT+8+kDMe/n9oNr/IQad+ba4ArNfBcIky9+hCFw5oFMP4tb
cEmPyS1LbybKdcPAQk1oHHvABWMhE8Yxy8ZYE3Wz2w/q2FYBCZVafNal+0wZKWqLPYr5w37CjkWU
4+gPga03UtVgfM2O74OyWy3fIJhdch8wr66prgs04z8BKV1JofbrBabxe8QgoHHpbr+7MMQMSDvH
m+d0k4Wh70U47XD5wbdpIeSAJSlqgPn2NP16phhgXJeB4dCuAKZN4dzV9WLh3v70xncQEXiSv+Ng
A3E4j0yzRZKqkTjBKKhKo3cILPeSxMvIH2Y7NNgvSXMRWH6+vgJeEouI6CmuLHyvccKDGxYJu+vk
JkqnLTu3y+IcAn0JRFECu7QYDwftZavJDjPbyXMdF2UM+2k2aNUbSSOs8k3KY3BPH1ubkYephZuY
q/pTFdj/yiw4INRqPJyGZ9Vec8+q5YEcAdYCpRk1aCqSw5r8CxLr9X2vuc6psI1nKnxtBig7zTus
mjsJfPlCiAlrcmMztscgG3jBs1OthPKnjGL4Mr0BwZWdf1GeHGw2k1BmkWyWg3/ugXuFfj3z/Wql
/PTnZC8QjyTZ04lO68/p7G+mo902d8zmxncJFvc+SZW3w5A1N/ns8Xdw4U1UgLn0IAqgavCQ6Rrh
ERg+/zu8pPhigoBoskHD7kVQMxckynfqAs/oFNmBUV0QT0UOcfDxtkCwxK3w9Mq/3yMDP2vag9Zd
ypStS9CfpIrh/WbI2p8ts5wT0qdHkwZR2FR64pC+oJ63d8hFTn3Pov0kW2qBuHH30huOHwqGm81O
qNqjhm4fQ0mSUwJspQb1vpnIeDpNhMaG2oCHv696wSbXHdn6X2PsC8SL9LyHh3FRRkpaZjFERvj2
uPUYKUUvoQzYlZN63RdAJ3JpJFoPidi6OGSCCu0l4+qWpzHhky6T4CL2+KJ1tMIvJCCV707/GVxe
RWImXU82La/161Hu7i8upmE6+VeH85gjKQPcKsY70XWSeNLR3d68DN3wACXoY7KvJyhmxaviqHPf
sGah1zliQuTfNDsTUaQSkkYRivf5y4B6ZeiRuQYQAIiIcf1y8W5+5gVOjDexHJKsU1R5UFGK7auJ
g4Ebdpl5I7L+lDAeFDiCLt+cz7ll8qz/SOhZZJ5cKEJd9oFxD9tmjHYvdaDEhvEoM8WyRfrMFzeu
w+Z+Px9Y7oFa7vIToGYtH5Aw4UcvuLOjRLJ1qNbf1lOeZsNvfhs79vHr/ki7v4LYbjsxInmOkT+5
2nKAN8RBmBrNydbb7u8/m6Vq/Ul+xddiq3UATRSG6GzG9Cw2wEu2u8cxngdP43Q5oPm9ibGLKDPw
Sbs1caphkM64qy+c/GYNdSdd5FBjIIZ1S+dgisFQtcvN5nkCHHGWuVgcRnDp3CTJlb/rXQykl8rG
U2lAQOHquMk6kp0rVP9rgLkX5GJHTiZrXeaTKTRY10NG+aD0FQlZIk6AAg6J7o5gj3o0APJAL+gY
iZivjDCSjMTkvy9oGP1ggdFRdoyiZuXUz1SX059gpcEnXXxXMoql8JGElG+ez78S8AOpKQX2Bm2y
OyTrgU5mwUtwJ9QMOfwuFIkJ3pdJE+XhMaAvATbGOip7j9l9vgRjlURq8tdHJu3k7gjW2o2M6N4Y
seF8G3fWP5rTV6TLL6bGo99IDtEkHR7LFtgOWJmmEaZys4CkbOdlvwSKpjG5IEOr0MG5VyjTHRU8
4EHCZqj5P4j5RoXjIaFliRfp9bJ6eWBPbB+WvM6trFCPL8O7v1SPXOamE9xAVr0OhnHKtVt4qJT4
EvHUhsc1fUAbHImF7nybbKBtWfbEhxRwderjsPfTre98VBEbffgGhY1OD5fJtW/guG7W5iaIkcIC
2x0Mzm+dFz5ZmdiRZZHi/cFi3R3xlypbET4a8SqysxZaV3AjMT5ziVIiFk6H2g8b5zxv263LNkdC
1zxOMl4e5Kximxhgk0wNn/3luFJs35mJ8rvE/nFMWumKD5EMuYOXasqEW2aRulMLL58QkflRkv47
y03dX+WIPGNR4QFeBndndYVQ2REY/TBC9xFabWT8qeA1MeHHUhoL94cN2LOgQ0yDrKdIAQFr+TS1
bgC2JaQV8TrPJM9rERpPS7d2+o4/gHlxG1/ahy9bwrLs3YTzIW8e93Cljtx/i6I1F1StqEXG3HLe
EG1ETM8zOZ5uOEwgG9DZq/oVg+CcK+u9G76O4ioM5yRBp6toCgKu4PI8jNhYGRlCJ5PB0YYI3S5h
MC+0hiUhVY44mFtv2XXsq0QqmqPNnOdu94R+iCcwQDNxd6xIRZq9jh/zKSBIwMZc7aUOuWPb7LgA
Uv+wvkp56MNVu9Q3OAyhTA4RWuwn5Aa8LHVHIr9ENLPPCAo9CVJf8gagyVNUc+q0RF065BmeerBY
DWPeute9syqoKpWafwmwY84hNN5574MXlgvEK+KY38pAEpXK7w+EYS9op/bL/ci5M6qpnfkGHT7Z
+3ZyT6EP03xdRcedDXkxccyRENmidiLZQzZU3L1dFnRLmQBUqveaAqDm0DS8ZtiM9VbJYKjpwr9F
Vwj9xC/wy2UM6zbth7OdoIBAt2J3szPyYmPwbr56+Fy05DrFU8I1J5s3uughMBZHXrQqI8X3o4ki
PMv1REGdhkMZJXHdM3Ra9z4t3IOKCp90ReHqp71Lw17G905ho9u3wsIMKBBsybMvfSuyA60c18pt
afMkugtIgHpojHpzLYqbH5iKuygvPSKFS99RKZD3nQEzlS9YYe8ajR5vC3VyAFT2bNr2RX0oHcO1
GzhDGFv4Yx/dNvf2mQ14MK4ACbgH7ikPG8Ed9RAkBXCHp6bqQFHkmhdGbsGMeWIS0kXpDMpclChC
JCBVgW/lje2WLTTiVCYp4SCdc+6FCsxP2nO9DRnA4549LoKxsPrJHK7R4MBzPCtVWXIYjpQckAhw
8hJbC/AIuLngazpdckRb5gyngW+ZGJYkcQzLSHfohMgq5hTmu2aPPrwEMfDUFlpHKUtc/2g8wNJS
MPvP9nYJS0dC/Ez/Bl7jzzUbcPq+NPTkSph4LEU+k297x2XeWUgP4XHBEawP+OAtbZbTmDl4Sb7r
a0NAhJFUz70KQJkrcHxOyWswCcXbo/SLWlcE4mVkKErzcaSnLLSt3imHHtEDZkRpSXNBPnMzqGRC
P5m2eF+pUFC/RNWfgs73wm5oZYRc1X8uGPAfn6VswFRxW8VqgMjqf9bvSNFxZcQClXolbMdf5x0K
LeXB1kv9qJ3yLuYABpQLM1PosSZwYW4o3Qu8i+zZLHF9C6XL0bmxcrdKdLc+Xa3OvpHAuVfeAQsD
H1iZksF3LRbq1AeEq3YtDS0CshOgfOxn40XsHTZcc8S+VE13HbNQp2TjFUKY1JN5C2FyBZGxzMor
l3oGjo/+X+F8U7xIXiOVtXpRq5Heg0II90hVK/bVfTTHZaPRM0soySrrFkaamJPbAzB+aWbVq4mu
uZkOhJyf+RA87ojqUvvPd5gmKi76F7GxZgMGiENOoq58YgKkgcV44ZYcbxMiVpEa5bvOmThnPdLX
V2RJmTANBSqy3L9Fh+2QVAN/tftF4h0vlTLii/39qoH6nUU+ICAskbaqGxC36jPCp6rMvI527bY0
owda8EO4c7jb5GQ08xZikouCgzxwiI7qYBq7g4sc8rpkZtvpYJz6C40NOeEszEiYrJkmgLBz27a8
mpaUPT6cEg55SNkzVVU8BKc5nmfljVeHMdt4kY0DR6cvlcvf9HWo2xJ4eLe2hOP6zIWnJ9fF1yVk
6KJNZj2+KFEBOkMVzgSkr5qjJpPjg7szHlC10LoWCriumJY3eKEZJ936krdsdEC+WuFYZzpnQ2vF
rLQxgdpxmTGG5ewfIEZPuI4nUTngMrBvsyqYCKmPKsuP1XCA8Mp+XnylIQZSYUCu1TgtIwZCJqNi
JCLiV9lGQbXFYKdP9RwyLowQgg/QU3rn6y15AzWHTyE1fW7WCTYI0GfWrLeWsZycrqC8C+jT6+nP
y3lrRH1wOSqz8SpCc3CNTdAkjzYHUozNOjp3M1DQBpT0h/iFwmxgDnK4vjlorVzmSlJy7ToZslB6
jcR+lFlNoGTVrVl4Zz1sPl7QyyQbtUukU+50kFXOTrsxofEaWMpREHq5K/a2tI/jMudGzINNdI7x
1Zck4J5PYgrFL+MQ/qGr/rKcPHpkLeq5EWkHX/E2lJPFaZTpyZly1ft98dAuwQvBteHWtvpdp13l
CJh7iKtLiIztSHL9b2foQz/VohCrl6nD9Lok1sygnQxl08GT0mvx/8D792wKTT5z+L6fO4UpJ8H5
CGwsjLJrWXZrTnNjGLBWguxfKTLjaZpsh7CEfrVzDYMMyODuAuLY4bFHR8I/NXftGYFsvxrNJz1Z
jTy43PYPv5Bc5v/y6oxJqQpXv0JqO/fszRt9s5xI9X6A605WOz5uid2v/hm07PedUcG2neaFNMsH
nzEy/whbzg/d3s6HrurW3sL3+QBfpLn0sgayhc92YnBByag4V3NymedhLKl08zeMP16HPNlTkH/o
yDK5pGY3M+MhKbe1kDj2oUL2Z6cEY+dLch13iaiTUEoQo1gisOsc99BFivY+DUUwYmTlInq5dfUt
qZGJqsCeIP0iI1IAoQaTuBII+ofUK8g7AmpwebHzurbGqgUzXs6XXkOa5O4ZbN28ixFy7Gcw+rHt
/5mctY4Ulb2uN/5nuJUO8tK++/ffZoLx86QJ9YZgS8Bv8yETuNHGMVv1g2RYR/2LIbqu2H+N5+7t
/PUd8Lxn4plinQ2xcKfCnT/0g1IcY46czybuh7y90/TxB+qtMtH1jBL9RprzqavE75TnPJltD3Vc
1BekKFX4fhSjCMM1dov2BQ7ww/dmbjjOw552KSzA201UGdNPDOCR0NrIHBmTEnnWAtH1mIUEK4E9
WXzoRYtp58AwdwMfpeYGRVLqcYTQTEwCz3Dh6LzjpI0+vuLJpr9CQszQBWqcga5Tr8wuBK2cvcNQ
QLcVOMdIlLV1faHaA1BeJDW4J7xpTfjg9qgY45He2EZy2RVmKPk1c6sm+M0qVAPSclN8XbFKnAgC
Qec814F0IWNmx8TYMZ91LGvzlWNa57Nq9PbFGM2H0cnS/sJKp2OSfO20+9sSHW9mR2/cFSI/rmjz
TlhLCoIkXrPuToA307wjuRvm7WcRejpkzNIF+C4oGFoGhUFTchnxCkBIXz+xDx1AIMsWQsNX4Sj7
PfqQdXiO6yBpUXsGeakZQUH/Ywrlfu1q0hdu2uiGsvxCkSLCENNfQQdT+FkYb8oZqa3l2lBgh591
Pc+eOG7NXuPANmPhU6lALpw4njbC6ZaHAi/vJzs5a13G5L3GSSa31bMx0NW7n9M+Y/tCiWeKX1qZ
aRsaJcpSfv6DTVZdMcDupHaBZ/Bn35/xYHs7d1GaKxFATq+w7N7idrleiBv55XahUHw/ygidv+rv
DCpf7NqNlvL/Ca8eDygby5HLAw5SygFCaNHaBQA/D+mEszgcM960xR65/pAQap23LiEOytg2rd0K
PJvoF2uASB2EX9/YO6JzHTkdZodTg6Sd3TnrSgXU3aV8XRL4K0k/owq+eESt1uc7Z7EPgH0+r92g
L4j/uDYIn5rlzVQETzhsRJlpEwvUe/UxY4oLf5EP2DrVvQ8SnYrw4SwbTuttJOXR05vNJnYZVAPC
9JJVa9wSU6VBEewcWJ16/aEDXU/pk9Q7e9pnmmvp5zqMh8EsPMVwEPDB2FA8QUUvE/HSmePaKRKh
OseZ3AUcNGZXeBnNtWPTY/L6wHF3eC4+taA5ERbC7fz4eBDt60kFOsO0TtMxRtoFXHYwizNwXRwo
ETUBawv88VgtgpjELLImJEZlb1DsRI5gFzb6pcrEVP9JKSuyrvZi7LAckG1jdgaogBMZjboORrOq
5EroXTdOxu9jc89WQ/uRt5ohWA6Uj42JA4T4wWDoMfbVRZ9PARGdbCIwz2LdUenSxWYcLrnOofZO
prh/e12Qedu98bW3odsh9qKJdHFaqK/eOCBwoVc3KPiRw042lWg+2qvxkpJDu9dhRdeUuj0vRbLR
u7HkU6yy/B6Kbuux2d/geb9DC0ESr8H5OWxVKFkC1+7iDfLwkSd1EOwWhwj+N+aItu8/kSltgQeT
qkvshq8kQ/VGQb7Mt6s2H+tXPjYK+Jbco5QtIpkVTOz9A5mmtC0/bpZNCac7abHzzzQ5b9n6LfQ5
Ojj+4DmsWBnshXAyIjCcq0AcqExvMTROp8IRIE+fU0BB24hPXWVxrPb7OX2ZE0+iMh2in0PprN5q
GpSWDjEkhN+wGDm3CpxVQwolpqHwPaeAPI7zwAVR1xDnNz882OlXkFHooBQ89xUfQhMnHWAxREj+
+ZcUDw7yb+gIQHc/4asqITKqrbsb9ewtoAAduvCKh1HBH+b8DjAGFK9W+3EWFx0HJwI1uOFRusNr
nHdf+eurjrRe2gZs0pJ0ogaEfPAVy/Ozwumt3T+YJCKy+BiCt55YmcIrPyftZts49AUIGO0NU42U
xgEK42SjdTUPecv+2BFPO98Gdkuqi1o5Nh8YEm9PMBGxUP+bWBhrKkNLbjj1VvoOGr8ugf+1Mb6f
03+9mQAgxcDw3zedGRQrKEwG7Frhb6mV/wB6bDwvgd+lMNlvzpz4i28JwPYoIUTWz9UIKuZ8zZFg
al5IszVT6VWxP8JkeKjdKXCpjXtb9LK/SH/4pCPykVHXNnM1UZS8XRECXo3fRiqkbUv8Lf5YmlfI
g5Qh2TUzV67ir+yZ6fmnCulo3ilrz2uAYzD2BY7IgKGVSHkaI9V0KpVOVw9Pzr514ls7dEzw0AZj
gdXBO26oCf7O1r1LlmLcMYqGn72Tn4BNt4ur2VrbohZPTOFrp+LVEUWAvJtWLWPF6CSjMZHf2h5C
uG1pkKUBkMpzesIqOhUBFUEpGO8l0VLjqLimOO+jkuO11sAcPKPDEr4uTF4IELixZQI3FyeEJkvw
Z1rb/VaszcsAlZiQ65u1aP/LDMZocy/AFlZzDqPBrrbznKba+DpZWTZSbtEXz3A/QKldyhoMPMdp
qnliEsk7v27PMq++CsxN4DmhLyHxdhQKhLX2ydbq6Pwv6Fv6mePTRLNAp2XL+IeisnrfRtg0GNEg
3vu0brwXcdK8unZVshqUkz/555mIFhFQSp86B4vcxTeGzU6QtYt/7KLcKvwZSLs2RAXPeShOuarX
vlHJ4utYBdXY0R6CmJSWwtboMuvfjjTB1dibWyWcTYHui0IkcVFozmjpGihauPSevObxW59sraMB
TpFr2SQay54AkCNAKK6fMmt9p2FB3UEA7iAG/CB26307KLtDKo+TP/Jpgyg8FDL7uVks4/LX2jMm
BK/dJ/d8ADfocw9NQtLZskKMhLJYDg67dsdblP5EPQ1C8JFiqbdO7ZL3OByW342NsGrv5amHu/Lc
VvZGpRFJz8qImTHrQ5vULNg8GoeVlqy2PEfmFtYMthVGIvIqnpRf2GfoznzXoSfjqeIFCeQl5CmN
UxJUeBbCnbF7g8G5aTr2r5+VJ4nYXQqkHRTwDzbq7jm4gGEgI0ZVfQKFX7f8BoJFH4NkMdHPM+AV
Zz+laqOSHJ35ZrfWw+6ucATmVa0NUihR5XIsk9RY4ZFuLxDIR2dYHmSfOg/PqH2xZdfdce7SPRJS
4T5QqK3D0kJSvKzHBw/xxnbYQDYYjZV2xQq9IglRBVQkXLJN9Q7QXsfBvsEN0smuLe42ZLHbrjBf
zssC2OkL8BOG2le5ydivCzHmb8PuBVNiyZ1n/DFfpz97SzZNF3Z/1CiRZUKobG6oJC7zkYqwEvri
hH0+RmUWJrVQCm3SmIUxs/aXOqCOm3XiK7I8cNi8VzxN/DwHkCIVTXPY9z+aCI3OpZ+2sbM9vHT+
2P60VLn1AdusrShABJmyeorLlSQc4eHcC/nCyHoEaLHf8jeBLUSiDVWybYHYnZKRyXkgcGCS2hJP
Eq2Zqk5HlH66LKu+57TqFVjubj/DrajdkhuNbhxR/tx4LOtMBibnhCKzQHa4EtYMo4hCliBnCKRs
zbZw6lEaEP05qdZo+SIxF0jPIRGlHwDfp3U/snP5+Xs/lmDFeGBmAepAIvlHUJQZYPM402Vjz8xz
LjZMYlQI/WGgVO+I0xDewK0PB3Xevxf2rjsSGfhOTiXFpjuS4xbzPgUfTsjBsSOx6NvH9+bKbV8z
wWJYu6XTBR684r3wNi8rnL3qTNPgTbkXJAUByxZ866eXaB+hICwxGrwy/CWifrlEJwbWQtd3+MiB
g0SSPuvSkAGJsZ12Ls2vDYylojbHZH0AjRVX/dY53wYIjdPA3RU3OBJwHP7b0pn9ABAUMjiAoZvE
hb8vFDapYaKWm7YHy6fWPMgFu+x01JUTAmAr0RE9WlA4u/jQOxD+/PKz9PG4YtSM6Mj/U5brN9OF
o9TMP7pq5bOBpjMnPpqHm9qGqZgzIhIQDcfctiyGpxvLV+9SVIOa/DfsATiMBfmLLwO3TGvtSoxu
P9dotbGLZAtiUejrI6XCHKeY66CwTLE8oBpYA91yoLSzpyxDw2TZFBZ00PU3CQmqOBOth0V69mn5
ioG32Y03goCTknqXFtvPPXA9bz05uGUNlZWFPrRBqnaUR7szTlBWYlxmBpsrOBAil4uM3YRBapKQ
BbTxT44tQVVb5OsVIiTRAg2z/CU1FSey6mAjSALv3NgCqWbE+GGTh9jTbhS4VzfufsBtKpgM8xJK
9pNyMgfgcNBzhg78qBHIk5YUQ+wR2+27NgibUiL7wkyPp8aWyV+vaOhhkgkJcUDmak4ll0GBz6YL
VoPWYXjir4/BBnRpNxBpbxqGy/IUr3hrCd9qleV965M22UHjaGYx8UZzF3qGWRzSFU4ldMAdmumT
zdOmdZglQExai1kfP56kFJs3orlzCEMuHhIcXJo2uN0O1NCbuALFNb0X9f6eQ9OGJ4ZvWcD6BMvs
dLG8G9YiuqAo7NJ9vwvX/QGUL0cVcgh/N99ED+ytwFu2L59MluhmOO8N9GAhORZcVLdT7aQjjcom
KfCbKHBW/WR06aTdD49lmSwKjiihEWjFpKly1mVxdW0Q+60CbNVnnjbxxZhOQ7KBbScLsv84Frnp
rQZpDpW5X02bKe6uFWjCbve5Q+wogL6H5htPp16edjMhcstw2opMoTFqm9cY65K4hG8RBpAFCLi3
vpiT7pAraw3Fwmaf0riTSSPn6CsISuTy1bRLl23oDMpr7+zBy7JYbfBvFTm4I3ZpdRHu+JKamBjy
V5IEmqjampCTAovnh3O4vt7VOHXVb3lE2WsrpshdYv1k0/Mzix3vD7KVLkFFvDVq8m5tCgfSrjHY
oHHL0yu5jvhBVvvuv5LXPoB/wpQHmfXB5bzGB3W58w5sNsmL2X5uqYOiGm1Dtxumn6eKc6mJ0jXY
bqNlqKV3trHKEzzuozIAUHG3M36SYX2kbs9xaEenXbCBf7ATtNRI5qX+zyNDg1TPf1w9MUm1MPJn
FxSZhA+WGfpfgAqJQR+lxrEPjA7ZmtB4MFyRr4101GUQnRUsC6vx5FM0+1I80FwYfHTYrFXbysZK
j3YcliFDGCDGg0Aug5liIaPzZSE2q+L11l3RPkpMp/UAjXGbGFMxI0IETso4GTT8OLLw7By1v/86
E2pS0gzjZms/AKXQbt/b1WfwarA7Nwrmk7QxMP6wMwaf13UwRePBcj2GQfdTMjHNfAuykAS67dfu
YWRK59mlo97EY/gJp/78nOl2phQ93tJqnqYXDzFH9ezPYyO8zA0+kXh9WhXv/yYDI8TV2ifBJwPS
PZdbimfieFnWZSUM2l6HohBlMPSHfXnw6nj4mTLF4498bNLIt9W1AzBgN0wFbzAH6eSh+ZxIKziM
9uaDkO/4D/1/Qodn25zWizH8oHxO/A5Mie128bCyJCN8A/S7vM1J+/ryO81gb2yJ6N0bIhqHonId
q/lno5QjplFZksh2Ep4eavcKVcsWlFg54itqVw4JDnGenkbPjSCjgP4b3kbghwbscPQih+0+CUMR
R0kTzbA2kYi9JTBRmEJKVMyFlLfRBEI+wHcXZwejzIUydzzCNJgzZl4Zdux91Gy3SbX8yQimLkmq
WaqrREPn/mkvghBslsGBtI0XiUsTgbbtnY9DsKWWmFvOWVcv7c0nr20epojfDHEOyAlmLQ1wllUM
DVaR/VaazioSi+7+3GO4e61gpoVVVisiG5XV1cKFKA2OY77CfLxVCxwZPbCoVxq4DiFN3SEmH3n9
Dl6ThCbGj/wx1zufKARuxNcZ/Zlf9x8Rm3eOhCij3sW+i6XTTwLs1InMMwYx9RnI+2wMMn4HR0xq
3hLNeSrN0vp+k+gaa5qisPe6dXolcZc/wAX4aZhkIgM0AV+TT/0DmZ4Ohicl0OB1e8Z2rSoT0nbb
RcuSlN1nsImIk4fhjlqniZcql3SPrapRa+bGtpp1A6p21wQ4L1RY+O3Iz5epAmlXMcAf6/fRuoiT
1cQMXNTj8/PCAPX/P5dNoRU/cbQ5WRjfIKGA8++rOn9rjZd0kPmIBWio4dMkAjmoNyNpY5dM6cDT
1D34hGAXQmJ687pWalWRGFbkzRjQXZveDSrR2Hl5PaYe1DxLEyX+QcwhL4hFohLEJj8rGgaLsaBH
Eizj69I/nTK8BkOoNxVYLz/GqDYtutgTPvmffD3vAn6h/fDMOdliH2CZDgaGeDEGkqellf4eiHQA
rJ/r6ItYpokqX//5TJLAMZZ256PPaL81F22EqpVqw7L7hf/Zd76y/rw8VD8qj2NIoKjGPOZmTZyw
J3tV5pQpgp5lrLWJvagBI6SXOeffuKQUTyfNc87DEHP2rMrwkypoSr270NUjwdUcUC25o3zpoqZd
jzseGFCm6Wj3bjuicbaJ68UlBK//N7LCwIOSPYstUqkCJentpP3coWo14FW4l5scehZ137ZS0nR2
pLvl0D432Lvuz0rzT1npPz+iy0YK/T6WB8TcYhg8wrVIT4Y9YTvI9LYsBdQq02EQ4culn0sljqDW
kRsdwQxHXpK3Nhha/rE5u+SfU+VQLMB9IvGlzMSu17X1wS3GPi6iUCJkdNduPVfHeKLkXv1vH1kR
F1tLnBXPUl1tx7zAsmlejNILQ7eAnZHtaE/RUmNDfdD4mtO8g6zgblds7aSPVA3GbP08oZALgJj1
qyomlhyliZvKaYVAd5+lKsFkG3FdmhHm3XY+piCGj0kp5+GehDHuVeB9EJkb1+mwwDZsohJ6u/uY
SQYOmveHf2YPMN/fwkZXkdumq//JYaEZx0uaCcOZV/W7HWQGQcEdb2VA0DFk4j1KV9SQQB3lPnp/
ehk6Orbn0CYIFIytBEIUoggy/wrrwHaGdVsnxeg+K2bVOa9ZsKYIUQTT/z9++5U4/uFn1Zt8Dtv4
PeXbIg3ogFgJOsMoXhOXRVEGWV5j0KVbqTpBgzYOcFRtRp6QGs+Ye0UUjtXhQnzamecQ+QI1y6V6
QLf3jRYJzbRKGmfA1PUO8eYCAvH/KhVBnS9L4399ukkEU03DW7nHfWL8VUfOWgmC6/Xyf8ctLNzh
u/4oOXB+Nr3SW54fJBi/rSYJKwhttf0tRDzTP8BxrTUIIUVo3iXFm+4Ev9bHIttegNbpLyY5TBc5
vmhiUXZ6Ffi5SR8pcSnJubGCpXlnVmv+YMQva6RXg3sKJlQ0s1hbKKeGc/za6B2OefRZTs1z22l0
azBgcsDb/b0CN0jZOEfIbhVY1Sc9TbrrxQhFr+Bq5nHW17B0EXhUyrTHa3flnycG1pZitwoqeb5G
KW+pAyebKoQ68rxwKGsE88wH8wz2AHpjyiSeoHpJQ0rknnxUXwuV7LizX5VHn/JXu+kyOpL5DhW1
/S7DLmUxyREh7cfDk9UuSmp88ex1Jv3OLWD0CE0NomLk1uPiOF6oQxbdpWS4krFUhD05s1erX6Uv
JTvrlJGfyQNwC1raBNsamnmpc93h5xPJesZd6u3vmM9g9mE90IFl46ElUAyVI3ubf+xA+Vv9kGju
pSJO/r7LiAHaAkaOzUKxlrpT7X6wBRfBKrgjl88ns7h3nUW8bPzMcEegBjcaKp3fsFRgPY0kawU1
pwcffEd4CnvQfP4hfx+er/DZRvstQzCwZP+0t8SeVQV7nkPz7+fOwbq3bjkJRG6avnpqlICDzxgg
XIhlwzfcUiDg8NmwiiXkLVTl2K2Kxk1pO2hw7njSfixeClc5iPWAqW10ydj7Phspz88HAOrXKVM7
Z3iY3bcN7/QirThOizc1DSEkFu5Ka/yPW+VRROHwuV2Qg1zn5moxCTBkZbdXDiohyaiJMnMK3LOE
Zm6WJdNtNlOwJoHPofAQOHA9Vt9m2eyxZYdC2my4btAYxE3TiYqhiFBr9RWy9yNq9t86WGnSjGz5
zqkUnhv2IN7k+A2npP0EyVX2VR4za8TFYqaxyyH09ImvQFMgHXLa8kqhp2Kl3QGes0SckYJyysfY
NRncAd+vPOZnFooi9l9jbIKRXB6fKucMAu85eayD5GM7tYEIJQvVTkhYm3wRI6TKt+cib1lsD+NG
xcjvbJjPGNdtIwHQsr+pkY270RTDrQhrPfW4Rrw2sr4pF0xIk2II3/203WDXqeBg8rLwvnQa2d1Q
OiQRqZBwvf2mp4FASe1BcgGa1ceqIMeFPP+NrWspx2hnZ++YJb/RDyHETRk90A81tSvldnfP+rQx
pW49A3BdXagrNmt/InEVwNWSCOUU8U7GbKVAdDDgAVxflU3fEHw97DNOY7gcG0IBARGQ2WZP6oVp
KLlvwavIFlEFrmdg3FfWDlQtGXbBDOSeCeIU3N8fOGyLwZSWDPxnLn9rbXApinu/tWTCNN6Wt6DH
Nl9yVwo4NMdDpMQc8+fyflN1t90m4k6INBK2jbmHuRQBcR0xKWGjbYkp+5pzAiLwEmQ2X5eNTh25
39KMKMCDCUPeTX2U/V9YTLBpeneouJKmkRLkbySCgEvl79mVgKvZ8gT81fSBDwdH3cyOMqFovy8g
xJF+B3LrhvRFSiVdjO1xRr7+e/b7oafFfLWwdZYzZarH6u9Fp89MWHz2qfo+yfbC0QZWz5y0quZW
AzK92/YP28sPUavyndx3uyXpAFL2IirVw1OgvJWH/zMFJWDAfb4g43nY/03mosuFLu7XFOmEAULZ
PB2beHQ+yrFsysG98GeDCjJnyZlTy4MwztF5GD9W0N+nq1vygZ/fKSQZqHz5zf9BSwg23CdJt2rK
72xnOA1hPh+swD3mDltxchDyt3wjEKmhO+A93410INDOIfgw2zmda8tcYQDsyFBgAbmkZD5M/FgG
N+GvDX2Rb3pP/KeoDBKu3PPuo74EkUtecpc4exEo0yMmChoRGRWBO9rBag6i1ds2o0K6ldfkQPWg
j71Yel3GZBE6+3QW7q4L0Z0+K0JttTMHWoH43Bj6R9Nuobu+bXtcI1XL6UZeDF248Mlua25fewbm
8lbv1ymm6pF3S7qpauZjBTVwTeUHdemV9vGRO1tz332dvdph84HnEQt1x/cPy8qBeFWEqgBQ+QNg
ywPfE2D86KScTfeGk7+EfoS3Pr9t8dgKYI8+TgfIdPsh39uC0tPxh+SRRM3QAzD8K9sMVTzh0J9x
UZKIz6K9/rE0nwI4gynywDhQopsrdg7O9WkgvQUVWqOetRVasLCqYET2TMt9SWs6oHp12ThwGObL
8q/LRzOuA1l4LGN8ZsqQxTc4pg+FoYvCW4n5ZUWakzUyXO/5/47gMV33HXeGeiH0e57U3zCNfgIn
uy06bKdS/tB3ec3Z24/oeCTrM5RMv0iX/2lk0GuXVtrUsIuSJBDariXKHAwnPF4t/3GnxjcH9H3j
dbSG6G1rnAwBm1rAaH2XOJFSpHk37PgQGUdPnshxSzTDBCoFurpD+GvfkRf3FMuQZoBKkT66q4J0
H0KLflcozyXDlfsEky5zi+mei8gA52x9cufNCTqqPnDnfUgIoTwNAHVz04r0+h4lirn5uvekArcW
UJ7BTxqUgWlMTbRlHVnQzSk/D1I+2pZ6hmypNeXVEupRA18Jm0VyZmqzp3amwUBKFq9N0ZKQ5sVp
FJyYeP6dvXTXYeL3KkJdamdC9alC/XCuTf9ueIwEDgQo/S5gqu6QnQBrqhtZIrj8Va8VRqCdUNtL
CjAC1+iDziqYzlXiL6jc1rDv0VfsrNgCpcJzFWrX8E/xu045/D8rPu45Ua6opEl8GDYLdzN1oHDy
9SReYqUvPfrxQ30S17gBcnujoIhaaAg47kDTdxRU+5qe2qQ6PmXpSC4zYz1g+4tdZcNGO9DXBr15
SPOJPcrgy1QClNtRUq3UrHihGiKrvvL31LXbY7o7rIokMGn9jtmYO9gDNku2ow3c85/RAFMXK2Of
MbR9EEAVZx/t4Tdi3ZRx/ASFFB7Yt3jgPHxKD0Pkx6Fe+CQ0BEDREowO8LbRGfKOH2uYjkbtJaxD
LL/iuxqjqvKYpviYIesAoR370UAzgrdxbW+ZC9Qulm4bb5ah0DZEovM57QSXgfCxmajV73Gcldo8
pb43M7DpVs6Vz1HSfFPj8klYB/yO/4uhrYe0iEtus7kob4EIo7xdsAE+RxPOvCUPjrPHHWqd2bwU
jOcPyzlYrNDoH+OarUYBOsBy7PCzydcopyWTIVLVSWBBQWt1XPBixv/CgueBOH6vIXVTCk/cFSAt
P+xTOInL6+HIq00KX0JyJiFBEYccE4SC5YfPmF24LYy0fe9FKJQFIpvqjB53d0Z6Q7Aygimzilqc
0Lkz7h7XJLokcV9V6puvf58n3TjFz08tEpp1lh2wor5y3mLWiwXhFAAbne/MMhnkFC0x3nc8oh4A
MzACH6IChYzPhpDabcpEvU57l3Pdkq8usuuXF2yhVrIX9GBiwj9099TJPgc7Fa4+D9htxsC0pQN7
vYB73hO3xIa10lhYIp73RuC7zJEdcbuh4jmu0OVmOE3NaYeJgYrH92TiHC62/0R8rRpksr6kBG5D
82iGTuSnAevUCGieFreQIIJK7KNmu41n4DO62JOtETQCYwuFftPymoAsZ5lihsQg9ZrBXvH2is/9
cMvsiw01Mf8sJcoiswCl1czfECwns+pFCH/4zzQP+LCFWIAOOR0OElaxX7v2blOmpcAZRjpUqNh7
CtuW4jGJNq5AQCpjhsE8IySAIEJsupFMPyum9P8hJRAa9bB9MkkaOcxjMAT/949lzjOubt2+ngz/
3kB+wYkILVuG2wBGXQgYsb+Ts2MaVswpbPpDPinhiH4h+JxaHJh2drgNqw+p4y6Ki88P83H6SvhJ
IjU0AKDZPMzu6/EINyoT/nR/2HeK2YUbQwjemWXQ2OzTWyf0xf9IqpVzX4kyq3hzedwlYQjzmGV8
D5SeqgBwC+EeLxK6Kbl3lwLc26NKq1XgLcMzr++SJJu0vgJ4I2pXAK7/wa7GOY8ntTQt2TDf8W6Z
leLyxZT6PJe9Tm2nIXPa9YhFYFIjPl/yrYfPyb0tMgHC8nuR+DCBkQRqhMnkKT7R7OfOv0MDe1fo
jSowe3KiorKCcElUrPa8MbIpmvFrM52vBPJF7bgifz7NyRN/IKTRM7JaGC/fO1Rx195QzfDgW3uP
d/28nBgFDZ/oywQ/JMHsbR1wmoNbzzkJ/kBZnQOPWTG3z1UpCnhOorvbSOqp/vsgp2tIl2vEIMbM
b8eRYB25j9nlaRiaX46q3nNJW42sM0C1xyuz8iYtxEvylL5xiIfD/H9GddLDFbDuPO/KW++sO/MS
JnuGbKtEngRkqRvzKhsLqs9X5aXZrJqS4QRBd55D40qOQEAbEbtYD95eth7GTPQ4cIOilnptmwgb
TycffU9gOZYs6EFYwXV4esdj4XhLcHxyEY6xvBaqw29UBkocPRauRQQSXEiBusOAg0E1SNKL4yv8
NqS5XpiUOZoWp+1eJqEQUwgBHSTXm4h3LQ04MYDXMyXTfRFfVpqDX2V9g3x7ozJCaw/HKSShUOfy
oK7l828WbG7SiDO7bR5vGDYD16NWl8gwxw5+FAq8MXAM3gxcHKbBzmmXvDzehQd5gZv7TTytXR1g
mE2ANsgCbmSotwqiCRr8yjri+h7gf5aVC2A+0raI1zQisBl4TxhdZ/50gpw9XaR0n5MYxbn7N3V/
P/Ko0x9Y3QYmDhDBpT8HUfEJyoukRmRfNt+lKDP4IajpV8SkmYAnJMQ+s0Pg7rYECa5shUK3dXc3
EcVM2R82lanTbNcU+ghWmLmqteQrkTF49CiSNfgMq3i8vxC0cUWz4urhOrC14GuBrYv+Gxj6MY3P
WX4zsBuA0PBKjooIzVWE28Q8Ib1xHvdFLYRuCZ/ctAPWj7SNr2LyXngfceJRxaQov6jLzEGXVjLV
UmWlltn8ksO524aP7L9uHwgFAAf36D3B4hrYV9H8SFvJqnr6OJjTQvfhy9HlIDRBbDKk2wqU6ti2
ne/K4kE+xSCJ2xvlUS13Kzluko7TPiBYL+xgv/8Rx2UhQKcBv4u9EYx7GtnDHrfIwO/Fr/xT+P7Z
fQaniqrvL/YbxgNSvjf/LQTJHw/cl+MnyAac/7OHqw1qDUE0lrkEHvcbs/dpU2Z1Ux+8QlZPxceW
9QvGl2U1jpPz9KxIl+LHVZWtx+1QH5LGf4Wd3v0djIfFOYe/c1yuzith5IenoMgwB6xbIKMO6P6w
L1sugWELtJ6l9eR0gQIaVD3hOmqbJZAZDqEtnzmngWErzBnGCmzTZLQwJsB/HsqGFhwSMbbahnMS
Fdg5FB27cRfxlcPHtDh/cP9l1f9dvx72a+qjdq+WsNr/DZdWcTTfiI0jfbLB4nLgqhbKbWgG9tVE
D7rgcxQTN5XWD0EFtPBVOpBkOBrTnJ6s6azO0MJiQOMrXJ/CDBuQD6rma9GN5hnYfNj7skxVsq3B
6fZVuIJhty1A/s5kOvM39fquy0fWpQvJopJihHdcWxdDY1TZ4Bas7txNLSoVg784rHEEm5MG4V2M
7/7VG0cxuHZCxVKI8jzl8Wrf3TgPsTMN5o0jxbcgZu/sijJTaZX0ihbUO59/39FhPdapf5T+chPJ
5cCAIG8PqSh5sPAPH1TumaeIqg54fxwP6p2GgS1sapdQWguZU/KcPhn9nHwOl6oS9WjjVEiemYrS
jLqm33ZeuTZ6Fom/C/2OYwqedPpPOwPJAEczqpNuboTmNbMDh4G3KoszjY6W46M06eUKhP0mlr5p
uxw/i5tBXzQrOgek4SrAVLJBrs9GJPPstT9ABbtKJ6Ij2vY5+ptF7Np48ZbEKDlVhPX38hyP6Xfd
KCChOPr3PvTIADczG+UuSDGz1K6sJliuW05sGEkGlmipQgVi0qO+uiTr8PCneM0++WvdQue0lv5i
amo6ObLeubX8Ma9/JR/Mz9OddC4OJNiw4MIQMhyKFXOM7lcgiuDlBv4giulPJdSa9+vFeGKQt/+e
K3X4IdurxfSrpdVJ5cuuF/jmudf+MebvVzleQIuZfizsr383mg0eOmxndUEBIWeRYFNSJ5fbVdo5
zkvP+wCDTNuvJX6K9y8a7y/nS29CDwpxdJL8CuQWIuEwNmrcquvE+EijET3bygDrToamth0Zr4XQ
bL0UcpcgVGlH9cB1jCjh3XluZtuGnL8VT1Q6Ic7oOF8BCrnP/Vs82R9tQ5grp0ROCX2T9a6J7Bbz
exQLTJNF1DOE9yhkXVvz1DAJg1//OnOJsqXEHibS3w16xk5V+156GMblraNoLzBPahOXpkGwm8SB
467KZKln0R74np+EieFtj0gKjCcgEKDUIO7qOiZaiSCA6YzRRXWqkMZ6Vh78YKibU1bU5r52PK8P
9XdgyXy/EvkE+I74FLFyT3Up1Bw74YKVKkf+2zoUPOzROVQvVfJ6ps8ewDImZ9rRG6TpmA+JNjd2
MSboy6QnU0wVjcZmGIqKYpKUVClaha8yWoHthnOv1iuXp9VdD00weKMIMA7Rg5vdtSZWiTDfAl0v
xyWlKTMt/VOiBEuRMsOT00R9eHFY5w6O0FiWMhL95q9NL73ld2wJOq1VFHM0GYHvJPQuzHRXLcJc
/Q7HEtJnVjcANujQ69DHWsa57Opnzca3liyirN0/wSitaYS8mxdX+avtISPlHPtygL1wRU8xo05G
moZo5e2wLtQ61Y1z6VYQGRX5v21GLTLRmgqOoTCnlyLGqJZKMTCu+nxvDHJyZ3WcpBU0St9v7GFD
SxRIGQpmcg+dYs4AEwomhG4KV/J859HC0Dw/NbaRHSwARha975gFIvsqpIEBndT8wYmtjth6cG2b
FXGTspTCO/rE/slKWxH0CxGmgCU9UQ3mULvjhy0xQWeqSARXTr1Hcn6H+j2q3iAGEr/u+YQkIik8
2XtuoAZxFkFq4+VCRUOH1LS6ZAB+dj0ukgCI/6y2ow3Reo+FSPdpxdlkPo0IHnJni930e37IIgOh
Y+c8Nu43iTUKjCOd04cOrix0I3NfvrXN4iKYsegHGbJdHshGWRLywDM/gkqxhnlHXldPMuJ352Q/
rozYDg9NHLpDfjbwf0AUrMGEqxKEbtXvd9Y4OoGN5l6oAKLka9ZzzSw/K4CCBkZANf8wYQ1iHW3k
3vp6rbdPzFPCnqMzD3RzW3XBu46Vn77wwAsKh7R5WncabgQiOjGuVEqlODZ3cbmx+Na58i3dFATg
Y9kqc1cpiIt1VZeJS16BXf36G2A22XBVd6VnRYPy2gbLq9BHex6QkISU6B3zpJCMd7JUOUJ7KpeV
4a7m5+TTVQ404yPxpqNB4GJZ8mPphpzzrbwuZ48s/QaoCKEl+G4r6l7EDD+ORrbf5Z672lc45kFX
afEvptjyaoWX/e2p98agZlh7XhESM+/iUMSL9q2Ngayo0UnIpXIyv2+68TzP3Xk7+JTXH6Hiv/Kw
uGb6b/M+nuctf/uqYdnyIy9tUS8sQxcuFBP9/c876axIfRneXSAiW8Gb9FgYL4ueR+tvTnxq4rTR
o9a5C0Nonb5X8VppxoM+eryivxuIeX8kI0wjbcuy3RUIOXdRkjIQkXnbxrdfkEJZ2gcd/dG7hao/
rOPtSkgOC07+/LCsktkhZQc6zUaGqQnLtoCiWB58gjKHy28vGNwsDBMD06v6JQAzsde5pMydx/sc
KmthZqLqXTVUkhJFpQbAp3oY76yFPnGj5JCz1OYBg+vN2Y0lccBytV4gMZqTu3fYJMl2nJ4Gt9sk
XM2KWgtIAtcKIvrkWyLORDRBvYWVRwtvCVzoBYLeJ+1j6moYQMyO/qc5qs3nY7Zka3DZ4d+8R4Kq
oqBrYwQ6apJyIzNCfA1vbAeKTdOoyg4vMkXLeKOcD8uQR8GqhTq/AbRNKF4fAj1OAgOUzDQIv/Rf
kFukhBGqPVFZD0wARqGPPAMgR496GZLcEGHTg3kIG/awVBf997e4oYW2Tv4CYlGiqrA/TSsUOW0D
mkFNTDIRd0ibhP6D8DFlo1a1Eh47ATSHgc2Zx58+FrJtyjnQLKNxIJhbjs4cI9IlPjJXMFPe6ZC7
XYiIIYmhQlRqqle7bgAQ69+hH948RsOOpktOnTjq0metZsk9kk1zqTfNloBolcNSFiIJ4Bn5vMOI
GfEoRXwsoLeIT8rUlMq7V5Bsz/rDeZQHqCtYM7BIva5CP6ZpDtnWSK142n/eShUVlci0nuZlkq9K
G4pzLJK9o4i0cWnD/uPjWACLjnpRqpKoxZ/kB5IjDTzl7XpoLg+C8sJKLhYoiBgVKL0BpOAIqQZM
Q3YDxHhwYEdswq1sHAzoiMbFJmNBxUQdw7OjcvnGUTDAmh6hYeDMDC3XuqA0qyO2xeYMocbrD1N0
ZbBDK0Bq2WZ95U0hddlRLf34AJJtJ+AhaJQHCIuIaDZwRk0nmdZ9fOw/7fbipMCn6ysNSts5XPGu
DfvHC5OmNnPjZ5eq/01Spbfy1korT1DU6BHVRzpUqwXwej8DjPlX07TGay5aal/byIIep2GKmnGU
sVX61ZNAvdlc8avnoZ3uqYPm8b0f6c6050aOXyPYTPcbBmvzC1h723axmuZViMkQiklG6Lg05qsL
M9IgaOKXvcxFoDXP4rVbSfCqlS6nxIJTI8WQOTLqvhQy604paAAtUs3vhRQr8u+HTXF21EDr7dMO
qX50IHVGcBv699++hkp9PrnMcUgQAbn10clKTaD8n7Jb52Wpzz3uHqhkDLEPBc5rcfVMS0J/b9JK
XxlK95ptZe8nRf471FiZADosCRYZgM/waMJwaxe7splR/3B82/eI5Up6L9ZAwnQu3oBIEuZJ6Gek
QcJs3dHO1b3sMgbvdUTRKEea9I6IKEBzGO7XI+sSGKfv41mjAVuAsFi7cVp5pbcN/22c2KGq645W
QIikvW2ArLzh9p0qlAkDg2fOQDA2WpVEKS1XTTIyrPdqBbw1llzYxdH3zcq4Gq7Zemm/tDOTgLWj
MKjmBydtEDidnKM9zvS1Ot2hoKKXm8gaItuBt7Owy+evjfGPoheYl7kt4sQBHZXweWcBHldDWWHP
w38gVks6id0Fg4qflxKlfeGWMJuJrZ/PbxSoLi7f9DeTB1rOe9E94cmXjErVfob6mWLfdWVwMuhk
4tSFAd0VPfheXz0yRoyvt1tOxTSanPHgbjd7X/JonFcWOTFmAevjUsuF1pw4OPOACGgmeZXGiMHc
zJswQMP1lWKrdpIsOBJMHqpywtKKiNdnhS4248/40N3+XdPPu8nuTm1JE4edY5MsGOD7WFT1Z69h
yDFKfmmMtnxxVO1fUsl2UBomvrcimmGHb8PI5w5QylB+n6g5jjJaelC5GgL6fpxT6r8zynWhgwfz
lPBYNu7ihCTY77YpJ1DzJaBpzHvdTbQIODGzWwZlyokWBi3A8xxeZKUJLK76PmyI1GifImU0Oa31
89dL08ks6pFIhR60wZSmDemEcAYS59vat/n5RBbZBdigkIDjT1dJOwE7S7gc9lqsqb13MTH1lEaa
6urSnQDhzJ1isBHirdUu8eNNnWDsTmInkHjx+6MwKsijrP5Pl1aoaSsmoltY36douj+I2DIe98Dz
Q7pjIisA9+LMpw6gZgw2uK8rdJWdQFq6+SakdHfde+1bWVYLedc9wQqpkglyTabnEW82SZ0Rxcgt
tbqZ9C5vCGlBTjRWOY+2ssYFrOn/BfplNJ/Bm/LewV/DnuCtgAOrlcPFD4903sc3Pq5KKMzbGyRb
Twq2LPrCurZjEsRH75WKnCkBKNd/K28mhkuB1cls+EQkF/ttbw9a5UihAudMfKq4/GHCtxj9pV68
AOGj1qqpxeG2Y/McB56Ic/rCvSZWLUk1s8SF8tkKqry4QZ6LGfaVuVSklW0R7ELaaavfCscM4ytI
hKVNc9d2pfCkhXdK4BERvWKyWGgO36v2zBxbAXF8VzDYn1dNm0Spi7e7UQVUnmdCDnBqB/mUOghR
RfMTU6RJ4HcpD0f41qLMDPmaQRv8v+dESTdxGBrW+4Uz61WCdl3/4V28qH2kZhy6q0GOHFVeLVVN
Jv55lLp/QzBnpOrMLa+nNFf867c5avywteczs89AOw9lUdmaeSkClFvCRWMVaxX83yui7FZrrWsS
MTnHzOOrFaI3CwKofVAq4xhShLAeGos/UGtOQEe3tQMbMuiexaHzeOiWcLDmBia2LmRo8w/jL9us
vqqED7W5kDJvM6GaIWQLNoOQDR/MS7DbZ7mOFSnumxEvfyeuOhgb1vP+SNo+0ps6jSALMtbexurC
TxFV3/1yCEE81k9QGL1S1QtaWwHxHWAOD/96x6j+cY/abH22pbQmVe9jQhLm2LFGbfVN2y33o6qL
krmYwYonNc5VLu8kNSSfbKY4qTNPk42H4nb5/e6FNgPNAn3ekmz+x+gChQHXbISGRNFMeBRgOCF4
KB3dCxg0WuWRI/CYDR9bvQoeXB883T+T39V5xaCBhdZu164qRN7DlCBGlDs3Ng2R9TZBoTs9l5g5
KXpmY3yinxmVqTHL2NpV2Bc5jaeH7f/SFWEqW5Gg9Ia628Z2feFPWt+V0iZp0H/vQfBL8idASc82
0olD++Kx+nfpGgzFB2++omlgDQ4DT2++VVgwDogqzPw0u2Q0FCjbYuhOzd561SWovL5Db4gkzc/q
BellG599jTfuECqEgkQxR8B9IbaJ5mE124X4lsXObhw38Pw4PNjIn38S/eQgbE9Jp1sg7xW7BOpN
2bK1SZzQT2pLz2YoytKeqY4Vb1cjA1fpJK3nwllF9rnkDbTFi8XyOUciPCTAuRXR6t+8oe7Mx6Vk
sTBAVy/y+vKi+5lOCtzkWAzgqTyYa0K9kL2pKVY9YneaQeQx7k+93Dsy2jPdGHruhY8Rd82Q7Bnv
on0OEp/6ylB5VScf7DBGhyr7XzB2E9sDthLgkA1Tj4j0J/hg+xxTwGa/tGqBFEcOCko4+EQFQSbV
ugCBuMvrQoCqWEooQDBZ6QLMtN6o0xDF47SFCuWEHjK0mCWTJpw1iWhCeOR5rPyJPMTBFOP6B4AZ
/D6AA41Py6HN6CI51xvFUbxhoSf2dOeC1y4EbzvHu4sZqNrMIvFOlOCUgUCkeUUuo0iljBG7WQPl
nzmtWXnYnpYGUxinVj8SNskguET9JB49C4dEcymo1+hSTz2PkAgeIQXr2sjzdalEeSXfw/5M6QMJ
/r7U304hI5diR/FvgeRIXCT6oWqtmk7ukqxsPnx213Fw5+3J/AJZYUvNKmdmKa99FB2wEWlT1bg8
TFjgG/5o4HAfdbBmj2GDalHDn558JctRsoueRKrgvrmpyzR96ToCzi3v0XWvB+pxGifagHzX7u4y
iYxJI6kH4fa8Q8HzsBdUteg+8yVB4bjr1yhQu7fXQ5KT10Dxxm/ixJ7ZdUdvk3MuUBnamJ22o2Wy
uBa5W5iqbSu97UGb32Q0y38upvWxPVleYStHaMzui2+X8puXOyQgX0krUrUU5oTUNR5klZU1foZZ
tpEGog1A3f3Qj8G0JPgpX7rH2SQjkrdkF0nBzWV6Ky+jjefz8nWLHYZT+oboODwacmH6nC2Wi1v1
Wc9E7RWvajdq2NWhLzR8ghKc0YKLfC34K6GkMlWHS1qRo1ZOUwgtcHoejdVvJ8IiK6ACYB/PM0z0
TxAfFw3psn15kcq49jAPsn0w58rmr6O94kosfuUzN2zFnAGmys71vtQiO0F/eeojdGRMPj/GLuio
++fjlLyZ8VLItODRahvcAO6UOJJgl62vvA736SYriZd4CT3qPbv0t7KtOeYTly1HC17Oguxz0DNs
W3nQ4cjjz4gpgPrn4sJycIw2rcKauomvpwMqoxPUx9pZZRFvgXhKhsm2VUpIatIRCnFkVgfuoOiJ
bIR3sBfwd3YpdkP2GqPTdNOSE8LV89bsuTQeQjC2
`protect end_protected
